
module mult_N1024_CC128 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [7:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2039]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U11 ( .A(n42018), .B(n42017), .Z(n41999) );
  XOR U12 ( .A(n42000), .B(n41999), .Z(n42001) );
  NANDN U13 ( .A(n4065), .B(n41890), .Z(n1) );
  NANDN U14 ( .A(n41848), .B(n42115), .Z(n2) );
  AND U15 ( .A(n1), .B(n2), .Z(n41894) );
  XOR U16 ( .A(n41923), .B(n41922), .Z(n41925) );
  XOR U17 ( .A(n41969), .B(n41968), .Z(n41970) );
  XOR U18 ( .A(n41986), .B(n41985), .Z(n41987) );
  XOR U19 ( .A(n42002), .B(n42001), .Z(n42021) );
  XOR U20 ( .A(n42109), .B(n42108), .Z(n42111) );
  XOR U21 ( .A(n42164), .B(n42163), .Z(n42165) );
  NANDN U22 ( .A(n4437), .B(n4068), .Z(n3) );
  NANDN U23 ( .A(n4403), .B(n42115), .Z(n4) );
  AND U24 ( .A(n3), .B(n4), .Z(n4439) );
  NANDN U25 ( .A(n4433), .B(n42047), .Z(n5) );
  NANDN U26 ( .A(n4481), .B(n4067), .Z(n6) );
  NAND U27 ( .A(n5), .B(n6), .Z(n4492) );
  NANDN U28 ( .A(n4514), .B(n4068), .Z(n7) );
  NANDN U29 ( .A(n4485), .B(n42115), .Z(n8) );
  AND U30 ( .A(n7), .B(n8), .Z(n4519) );
  NANDN U31 ( .A(n4513), .B(n42047), .Z(n9) );
  NANDN U32 ( .A(n4550), .B(n4067), .Z(n10) );
  NAND U33 ( .A(n9), .B(n10), .Z(n4561) );
  NANDN U34 ( .A(n4588), .B(n4068), .Z(n11) );
  NANDN U35 ( .A(n4554), .B(n42115), .Z(n12) );
  AND U36 ( .A(n11), .B(n12), .Z(n4593) );
  NANDN U37 ( .A(n4587), .B(n42047), .Z(n13) );
  NANDN U38 ( .A(n4624), .B(n4067), .Z(n14) );
  NAND U39 ( .A(n13), .B(n14), .Z(n4635) );
  NANDN U40 ( .A(n4665), .B(n4068), .Z(n15) );
  NANDN U41 ( .A(n4628), .B(n42115), .Z(n16) );
  AND U42 ( .A(n15), .B(n16), .Z(n4667) );
  NANDN U43 ( .A(n4661), .B(n42047), .Z(n17) );
  NANDN U44 ( .A(n4698), .B(n4067), .Z(n18) );
  NAND U45 ( .A(n17), .B(n18), .Z(n4709) );
  NANDN U46 ( .A(n4736), .B(n4068), .Z(n19) );
  NANDN U47 ( .A(n4702), .B(n42115), .Z(n20) );
  AND U48 ( .A(n19), .B(n20), .Z(n4741) );
  NANDN U49 ( .A(n4735), .B(n42047), .Z(n21) );
  NANDN U50 ( .A(n4772), .B(n4067), .Z(n22) );
  NAND U51 ( .A(n21), .B(n22), .Z(n4783) );
  NANDN U52 ( .A(n4813), .B(n4068), .Z(n23) );
  NANDN U53 ( .A(n4776), .B(n42115), .Z(n24) );
  AND U54 ( .A(n23), .B(n24), .Z(n4815) );
  NANDN U55 ( .A(n4809), .B(n42047), .Z(n25) );
  NANDN U56 ( .A(n4846), .B(n4067), .Z(n26) );
  NAND U57 ( .A(n25), .B(n26), .Z(n4857) );
  NANDN U58 ( .A(n4884), .B(n4068), .Z(n27) );
  NANDN U59 ( .A(n4847), .B(n42115), .Z(n28) );
  AND U60 ( .A(n27), .B(n28), .Z(n4889) );
  NANDN U61 ( .A(n4883), .B(n42047), .Z(n29) );
  NANDN U62 ( .A(n4920), .B(n4067), .Z(n30) );
  NAND U63 ( .A(n29), .B(n30), .Z(n4931) );
  NANDN U64 ( .A(n4958), .B(n4068), .Z(n31) );
  NANDN U65 ( .A(n4924), .B(n42115), .Z(n32) );
  AND U66 ( .A(n31), .B(n32), .Z(n4963) );
  NANDN U67 ( .A(n4957), .B(n42047), .Z(n33) );
  NANDN U68 ( .A(n4994), .B(n4067), .Z(n34) );
  NAND U69 ( .A(n33), .B(n34), .Z(n5005) );
  NANDN U70 ( .A(n5035), .B(n4068), .Z(n35) );
  NANDN U71 ( .A(n4998), .B(n42115), .Z(n36) );
  AND U72 ( .A(n35), .B(n36), .Z(n5037) );
  NANDN U73 ( .A(n5031), .B(n42047), .Z(n37) );
  NANDN U74 ( .A(n5068), .B(n4067), .Z(n38) );
  NAND U75 ( .A(n37), .B(n38), .Z(n5079) );
  NANDN U76 ( .A(n5106), .B(n4068), .Z(n39) );
  NANDN U77 ( .A(n5069), .B(n42115), .Z(n40) );
  AND U78 ( .A(n39), .B(n40), .Z(n5111) );
  NANDN U79 ( .A(n5105), .B(n42047), .Z(n41) );
  NANDN U80 ( .A(n5142), .B(n4067), .Z(n42) );
  NAND U81 ( .A(n41), .B(n42), .Z(n5153) );
  NANDN U82 ( .A(n5183), .B(n4068), .Z(n43) );
  NANDN U83 ( .A(n5146), .B(n42115), .Z(n44) );
  AND U84 ( .A(n43), .B(n44), .Z(n5185) );
  NANDN U85 ( .A(n5179), .B(n42047), .Z(n45) );
  NANDN U86 ( .A(n5216), .B(n4067), .Z(n46) );
  NAND U87 ( .A(n45), .B(n46), .Z(n5227) );
  NANDN U88 ( .A(n5254), .B(n4068), .Z(n47) );
  NANDN U89 ( .A(n5220), .B(n42115), .Z(n48) );
  AND U90 ( .A(n47), .B(n48), .Z(n5259) );
  NANDN U91 ( .A(n5253), .B(n42047), .Z(n49) );
  NANDN U92 ( .A(n5290), .B(n4067), .Z(n50) );
  NAND U93 ( .A(n49), .B(n50), .Z(n5301) );
  NANDN U94 ( .A(n5331), .B(n4068), .Z(n51) );
  NANDN U95 ( .A(n5294), .B(n42115), .Z(n52) );
  AND U96 ( .A(n51), .B(n52), .Z(n5333) );
  NANDN U97 ( .A(n5327), .B(n42047), .Z(n53) );
  NANDN U98 ( .A(n5364), .B(n4067), .Z(n54) );
  NAND U99 ( .A(n53), .B(n54), .Z(n5375) );
  NANDN U100 ( .A(n5405), .B(n4068), .Z(n55) );
  NANDN U101 ( .A(n5365), .B(n42115), .Z(n56) );
  AND U102 ( .A(n55), .B(n56), .Z(n5407) );
  NANDN U103 ( .A(n5401), .B(n42047), .Z(n57) );
  NANDN U104 ( .A(n5438), .B(n4067), .Z(n58) );
  NAND U105 ( .A(n57), .B(n58), .Z(n5449) );
  NANDN U106 ( .A(n5476), .B(n4068), .Z(n59) );
  NANDN U107 ( .A(n5442), .B(n42115), .Z(n60) );
  AND U108 ( .A(n59), .B(n60), .Z(n5481) );
  NANDN U109 ( .A(n5475), .B(n42047), .Z(n61) );
  NANDN U110 ( .A(n5512), .B(n4067), .Z(n62) );
  NAND U111 ( .A(n61), .B(n62), .Z(n5523) );
  NANDN U112 ( .A(n5553), .B(n4068), .Z(n63) );
  NANDN U113 ( .A(n5516), .B(n42115), .Z(n64) );
  AND U114 ( .A(n63), .B(n64), .Z(n5555) );
  NANDN U115 ( .A(n5549), .B(n42047), .Z(n65) );
  NANDN U116 ( .A(n5586), .B(n4067), .Z(n66) );
  NAND U117 ( .A(n65), .B(n66), .Z(n5597) );
  NANDN U118 ( .A(n5627), .B(n4068), .Z(n67) );
  NANDN U119 ( .A(n5590), .B(n42115), .Z(n68) );
  AND U120 ( .A(n67), .B(n68), .Z(n5629) );
  NANDN U121 ( .A(n5623), .B(n42047), .Z(n69) );
  NANDN U122 ( .A(n5660), .B(n4067), .Z(n70) );
  NAND U123 ( .A(n69), .B(n70), .Z(n5671) );
  NANDN U124 ( .A(n5701), .B(n4068), .Z(n71) );
  NANDN U125 ( .A(n5661), .B(n42115), .Z(n72) );
  AND U126 ( .A(n71), .B(n72), .Z(n5703) );
  NANDN U127 ( .A(n5697), .B(n42047), .Z(n73) );
  NANDN U128 ( .A(n5734), .B(n4067), .Z(n74) );
  NAND U129 ( .A(n73), .B(n74), .Z(n5745) );
  NANDN U130 ( .A(n5775), .B(n4068), .Z(n75) );
  NANDN U131 ( .A(n5735), .B(n42115), .Z(n76) );
  AND U132 ( .A(n75), .B(n76), .Z(n5777) );
  NANDN U133 ( .A(n5771), .B(n42047), .Z(n77) );
  NANDN U134 ( .A(n5808), .B(n4067), .Z(n78) );
  NAND U135 ( .A(n77), .B(n78), .Z(n5819) );
  NANDN U136 ( .A(n5849), .B(n4068), .Z(n79) );
  NANDN U137 ( .A(n5812), .B(n42115), .Z(n80) );
  AND U138 ( .A(n79), .B(n80), .Z(n5851) );
  NANDN U139 ( .A(n5845), .B(n42047), .Z(n81) );
  NANDN U140 ( .A(n5882), .B(n4067), .Z(n82) );
  NAND U141 ( .A(n81), .B(n82), .Z(n5893) );
  NANDN U142 ( .A(n5923), .B(n4068), .Z(n83) );
  NANDN U143 ( .A(n5886), .B(n42115), .Z(n84) );
  AND U144 ( .A(n83), .B(n84), .Z(n5925) );
  NANDN U145 ( .A(n5919), .B(n42047), .Z(n85) );
  NANDN U146 ( .A(n5956), .B(n4067), .Z(n86) );
  NAND U147 ( .A(n85), .B(n86), .Z(n5967) );
  NANDN U148 ( .A(n5997), .B(n4068), .Z(n87) );
  NANDN U149 ( .A(n5957), .B(n42115), .Z(n88) );
  AND U150 ( .A(n87), .B(n88), .Z(n5999) );
  NANDN U151 ( .A(n5993), .B(n42047), .Z(n89) );
  NANDN U152 ( .A(n6030), .B(n4067), .Z(n90) );
  NAND U153 ( .A(n89), .B(n90), .Z(n6041) );
  NANDN U154 ( .A(n6071), .B(n4068), .Z(n91) );
  NANDN U155 ( .A(n6034), .B(n42115), .Z(n92) );
  AND U156 ( .A(n91), .B(n92), .Z(n6073) );
  NANDN U157 ( .A(n6067), .B(n42047), .Z(n93) );
  NANDN U158 ( .A(n6104), .B(n4067), .Z(n94) );
  NAND U159 ( .A(n93), .B(n94), .Z(n6115) );
  NANDN U160 ( .A(n6142), .B(n4068), .Z(n95) );
  NANDN U161 ( .A(n6108), .B(n42115), .Z(n96) );
  AND U162 ( .A(n95), .B(n96), .Z(n6147) );
  NANDN U163 ( .A(n6141), .B(n42047), .Z(n97) );
  NANDN U164 ( .A(n6178), .B(n4067), .Z(n98) );
  NAND U165 ( .A(n97), .B(n98), .Z(n6189) );
  NANDN U166 ( .A(n6216), .B(n4068), .Z(n99) );
  NANDN U167 ( .A(n6182), .B(n42115), .Z(n100) );
  AND U168 ( .A(n99), .B(n100), .Z(n6221) );
  NANDN U169 ( .A(n6215), .B(n42047), .Z(n101) );
  NANDN U170 ( .A(n6252), .B(n4067), .Z(n102) );
  NAND U171 ( .A(n101), .B(n102), .Z(n6263) );
  NANDN U172 ( .A(n6293), .B(n4068), .Z(n103) );
  NANDN U173 ( .A(n6256), .B(n42115), .Z(n104) );
  AND U174 ( .A(n103), .B(n104), .Z(n6295) );
  NANDN U175 ( .A(n6289), .B(n42047), .Z(n105) );
  NANDN U176 ( .A(n6326), .B(n4067), .Z(n106) );
  NAND U177 ( .A(n105), .B(n106), .Z(n6337) );
  NANDN U178 ( .A(n6367), .B(n4068), .Z(n107) );
  NANDN U179 ( .A(n6330), .B(n42115), .Z(n108) );
  AND U180 ( .A(n107), .B(n108), .Z(n6369) );
  NANDN U181 ( .A(n6363), .B(n42047), .Z(n109) );
  NANDN U182 ( .A(n6400), .B(n4067), .Z(n110) );
  NAND U183 ( .A(n109), .B(n110), .Z(n6411) );
  NANDN U184 ( .A(n6438), .B(n4068), .Z(n111) );
  NANDN U185 ( .A(n6404), .B(n42115), .Z(n112) );
  AND U186 ( .A(n111), .B(n112), .Z(n6443) );
  NANDN U187 ( .A(n6437), .B(n42047), .Z(n113) );
  NANDN U188 ( .A(n6474), .B(n4067), .Z(n114) );
  NAND U189 ( .A(n113), .B(n114), .Z(n6485) );
  NANDN U190 ( .A(n6515), .B(n4068), .Z(n115) );
  NANDN U191 ( .A(n6478), .B(n42115), .Z(n116) );
  AND U192 ( .A(n115), .B(n116), .Z(n6517) );
  NANDN U193 ( .A(n6511), .B(n42047), .Z(n117) );
  NANDN U194 ( .A(n6548), .B(n4067), .Z(n118) );
  NAND U195 ( .A(n117), .B(n118), .Z(n6559) );
  NANDN U196 ( .A(n6589), .B(n4068), .Z(n119) );
  NANDN U197 ( .A(n6552), .B(n42115), .Z(n120) );
  AND U198 ( .A(n119), .B(n120), .Z(n6591) );
  NANDN U199 ( .A(n6585), .B(n42047), .Z(n121) );
  NANDN U200 ( .A(n6622), .B(n4067), .Z(n122) );
  NAND U201 ( .A(n121), .B(n122), .Z(n6633) );
  NANDN U202 ( .A(n6663), .B(n4068), .Z(n123) );
  NANDN U203 ( .A(n6626), .B(n42115), .Z(n124) );
  AND U204 ( .A(n123), .B(n124), .Z(n6665) );
  NANDN U205 ( .A(n6659), .B(n42047), .Z(n125) );
  NANDN U206 ( .A(n6696), .B(n4067), .Z(n126) );
  NAND U207 ( .A(n125), .B(n126), .Z(n6707) );
  NANDN U208 ( .A(n6734), .B(n4068), .Z(n127) );
  NANDN U209 ( .A(n6700), .B(n42115), .Z(n128) );
  AND U210 ( .A(n127), .B(n128), .Z(n6739) );
  NANDN U211 ( .A(n6733), .B(n42047), .Z(n129) );
  NANDN U212 ( .A(n6770), .B(n4067), .Z(n130) );
  NAND U213 ( .A(n129), .B(n130), .Z(n6781) );
  NANDN U214 ( .A(n6811), .B(n4068), .Z(n131) );
  NANDN U215 ( .A(n6774), .B(n42115), .Z(n132) );
  AND U216 ( .A(n131), .B(n132), .Z(n6813) );
  NANDN U217 ( .A(n6807), .B(n42047), .Z(n133) );
  NANDN U218 ( .A(n6844), .B(n4067), .Z(n134) );
  NAND U219 ( .A(n133), .B(n134), .Z(n6855) );
  NANDN U220 ( .A(n6885), .B(n4068), .Z(n135) );
  NANDN U221 ( .A(n6845), .B(n42115), .Z(n136) );
  AND U222 ( .A(n135), .B(n136), .Z(n6887) );
  NANDN U223 ( .A(n6881), .B(n42047), .Z(n137) );
  NANDN U224 ( .A(n6923), .B(n4067), .Z(n138) );
  NAND U225 ( .A(n137), .B(n138), .Z(n6934) );
  NANDN U226 ( .A(n6959), .B(n4068), .Z(n139) );
  NANDN U227 ( .A(n6924), .B(n42115), .Z(n140) );
  AND U228 ( .A(n139), .B(n140), .Z(n6961) );
  NANDN U229 ( .A(n6955), .B(n42047), .Z(n141) );
  NANDN U230 ( .A(n6992), .B(n4067), .Z(n142) );
  NAND U231 ( .A(n141), .B(n142), .Z(n7003) );
  NANDN U232 ( .A(n7035), .B(n4068), .Z(n143) );
  NANDN U233 ( .A(n6996), .B(n42115), .Z(n144) );
  AND U234 ( .A(n143), .B(n144), .Z(n7040) );
  NANDN U235 ( .A(n7034), .B(n42047), .Z(n145) );
  NANDN U236 ( .A(n7066), .B(n4067), .Z(n146) );
  NAND U237 ( .A(n145), .B(n146), .Z(n7077) );
  NANDN U238 ( .A(n7104), .B(n4068), .Z(n147) );
  NANDN U239 ( .A(n7067), .B(n42115), .Z(n148) );
  AND U240 ( .A(n147), .B(n148), .Z(n7109) );
  NANDN U241 ( .A(n7103), .B(n42047), .Z(n149) );
  NANDN U242 ( .A(n7140), .B(n4067), .Z(n150) );
  NAND U243 ( .A(n149), .B(n150), .Z(n7151) );
  NANDN U244 ( .A(n7178), .B(n4068), .Z(n151) );
  NANDN U245 ( .A(n7144), .B(n42115), .Z(n152) );
  AND U246 ( .A(n151), .B(n152), .Z(n7183) );
  NANDN U247 ( .A(n7177), .B(n42047), .Z(n153) );
  NANDN U248 ( .A(n7214), .B(n4067), .Z(n154) );
  NAND U249 ( .A(n153), .B(n154), .Z(n7225) );
  NANDN U250 ( .A(n7255), .B(n4068), .Z(n155) );
  NANDN U251 ( .A(n7218), .B(n42115), .Z(n156) );
  AND U252 ( .A(n155), .B(n156), .Z(n7257) );
  NANDN U253 ( .A(n7251), .B(n42047), .Z(n157) );
  NANDN U254 ( .A(n7288), .B(n4067), .Z(n158) );
  NAND U255 ( .A(n157), .B(n158), .Z(n7299) );
  NANDN U256 ( .A(n7329), .B(n4068), .Z(n159) );
  NANDN U257 ( .A(n7292), .B(n42115), .Z(n160) );
  AND U258 ( .A(n159), .B(n160), .Z(n7331) );
  NANDN U259 ( .A(n7325), .B(n42047), .Z(n161) );
  NANDN U260 ( .A(n7362), .B(n4067), .Z(n162) );
  NAND U261 ( .A(n161), .B(n162), .Z(n7373) );
  NANDN U262 ( .A(n7403), .B(n4068), .Z(n163) );
  NANDN U263 ( .A(n7363), .B(n42115), .Z(n164) );
  AND U264 ( .A(n163), .B(n164), .Z(n7405) );
  NANDN U265 ( .A(n7399), .B(n42047), .Z(n165) );
  NANDN U266 ( .A(n7436), .B(n4067), .Z(n166) );
  NAND U267 ( .A(n165), .B(n166), .Z(n7447) );
  NANDN U268 ( .A(n7477), .B(n4068), .Z(n167) );
  NANDN U269 ( .A(n7440), .B(n42115), .Z(n168) );
  AND U270 ( .A(n167), .B(n168), .Z(n7479) );
  NANDN U271 ( .A(n7473), .B(n42047), .Z(n169) );
  NANDN U272 ( .A(n7510), .B(n4067), .Z(n170) );
  NAND U273 ( .A(n169), .B(n170), .Z(n7521) );
  NANDN U274 ( .A(n7551), .B(n4068), .Z(n171) );
  NANDN U275 ( .A(n7514), .B(n42115), .Z(n172) );
  AND U276 ( .A(n171), .B(n172), .Z(n7553) );
  NANDN U277 ( .A(n7547), .B(n42047), .Z(n173) );
  NANDN U278 ( .A(n7584), .B(n4067), .Z(n174) );
  NAND U279 ( .A(n173), .B(n174), .Z(n7595) );
  NANDN U280 ( .A(n7625), .B(n4068), .Z(n175) );
  NANDN U281 ( .A(n7588), .B(n42115), .Z(n176) );
  AND U282 ( .A(n175), .B(n176), .Z(n7627) );
  NANDN U283 ( .A(n7621), .B(n42047), .Z(n177) );
  NANDN U284 ( .A(n7658), .B(n4067), .Z(n178) );
  NAND U285 ( .A(n177), .B(n178), .Z(n7669) );
  NANDN U286 ( .A(n7699), .B(n4068), .Z(n179) );
  NANDN U287 ( .A(n7662), .B(n42115), .Z(n180) );
  AND U288 ( .A(n179), .B(n180), .Z(n7701) );
  NANDN U289 ( .A(n7695), .B(n42047), .Z(n181) );
  NANDN U290 ( .A(n7732), .B(n4067), .Z(n182) );
  NAND U291 ( .A(n181), .B(n182), .Z(n7743) );
  NANDN U292 ( .A(n7773), .B(n4068), .Z(n183) );
  NANDN U293 ( .A(n7736), .B(n42115), .Z(n184) );
  AND U294 ( .A(n183), .B(n184), .Z(n7775) );
  NANDN U295 ( .A(n7769), .B(n42047), .Z(n185) );
  NANDN U296 ( .A(n7806), .B(n4067), .Z(n186) );
  NAND U297 ( .A(n185), .B(n186), .Z(n7817) );
  NANDN U298 ( .A(n7847), .B(n4068), .Z(n187) );
  NANDN U299 ( .A(n7810), .B(n42115), .Z(n188) );
  AND U300 ( .A(n187), .B(n188), .Z(n7849) );
  NANDN U301 ( .A(n7843), .B(n42047), .Z(n189) );
  NANDN U302 ( .A(n7880), .B(n4067), .Z(n190) );
  NAND U303 ( .A(n189), .B(n190), .Z(n7891) );
  NANDN U304 ( .A(n7921), .B(n4068), .Z(n191) );
  NANDN U305 ( .A(n7881), .B(n42115), .Z(n192) );
  AND U306 ( .A(n191), .B(n192), .Z(n7923) );
  NANDN U307 ( .A(n7917), .B(n42047), .Z(n193) );
  NANDN U308 ( .A(n7954), .B(n4067), .Z(n194) );
  NAND U309 ( .A(n193), .B(n194), .Z(n7965) );
  NANDN U310 ( .A(n7995), .B(n4068), .Z(n195) );
  NANDN U311 ( .A(n7958), .B(n42115), .Z(n196) );
  AND U312 ( .A(n195), .B(n196), .Z(n7997) );
  NANDN U313 ( .A(n7991), .B(n42047), .Z(n197) );
  NANDN U314 ( .A(n8028), .B(n4067), .Z(n198) );
  NAND U315 ( .A(n197), .B(n198), .Z(n8039) );
  NANDN U316 ( .A(n8069), .B(n4068), .Z(n199) );
  NANDN U317 ( .A(n8032), .B(n42115), .Z(n200) );
  AND U318 ( .A(n199), .B(n200), .Z(n8071) );
  NANDN U319 ( .A(n8065), .B(n42047), .Z(n201) );
  NANDN U320 ( .A(n8102), .B(n4067), .Z(n202) );
  NAND U321 ( .A(n201), .B(n202), .Z(n8113) );
  NANDN U322 ( .A(n8140), .B(n4068), .Z(n203) );
  NANDN U323 ( .A(n8103), .B(n42115), .Z(n204) );
  AND U324 ( .A(n203), .B(n204), .Z(n8145) );
  NANDN U325 ( .A(n8139), .B(n42047), .Z(n205) );
  NANDN U326 ( .A(n8176), .B(n4067), .Z(n206) );
  NAND U327 ( .A(n205), .B(n206), .Z(n8187) );
  NANDN U328 ( .A(n8217), .B(n4068), .Z(n207) );
  NANDN U329 ( .A(n8177), .B(n42115), .Z(n208) );
  AND U330 ( .A(n207), .B(n208), .Z(n8219) );
  NANDN U331 ( .A(n8213), .B(n42047), .Z(n209) );
  NANDN U332 ( .A(n8250), .B(n4067), .Z(n210) );
  NAND U333 ( .A(n209), .B(n210), .Z(n8261) );
  NANDN U334 ( .A(n8291), .B(n4068), .Z(n211) );
  NANDN U335 ( .A(n8251), .B(n42115), .Z(n212) );
  AND U336 ( .A(n211), .B(n212), .Z(n8293) );
  NANDN U337 ( .A(n8287), .B(n42047), .Z(n213) );
  NANDN U338 ( .A(n8324), .B(n4067), .Z(n214) );
  NAND U339 ( .A(n213), .B(n214), .Z(n8335) );
  NANDN U340 ( .A(n8365), .B(n4068), .Z(n215) );
  NANDN U341 ( .A(n8328), .B(n42115), .Z(n216) );
  AND U342 ( .A(n215), .B(n216), .Z(n8367) );
  NANDN U343 ( .A(n8361), .B(n42047), .Z(n217) );
  NANDN U344 ( .A(n8398), .B(n4067), .Z(n218) );
  NAND U345 ( .A(n217), .B(n218), .Z(n8409) );
  NANDN U346 ( .A(n8439), .B(n4068), .Z(n219) );
  NANDN U347 ( .A(n8402), .B(n42115), .Z(n220) );
  AND U348 ( .A(n219), .B(n220), .Z(n8441) );
  NANDN U349 ( .A(n8435), .B(n42047), .Z(n221) );
  NANDN U350 ( .A(n8472), .B(n4067), .Z(n222) );
  NAND U351 ( .A(n221), .B(n222), .Z(n8483) );
  NANDN U352 ( .A(n8513), .B(n4068), .Z(n223) );
  NANDN U353 ( .A(n8476), .B(n42115), .Z(n224) );
  AND U354 ( .A(n223), .B(n224), .Z(n8515) );
  NANDN U355 ( .A(n8509), .B(n42047), .Z(n225) );
  NANDN U356 ( .A(n8546), .B(n4067), .Z(n226) );
  NAND U357 ( .A(n225), .B(n226), .Z(n8557) );
  NANDN U358 ( .A(n8587), .B(n4068), .Z(n227) );
  NANDN U359 ( .A(n8547), .B(n42115), .Z(n228) );
  AND U360 ( .A(n227), .B(n228), .Z(n8589) );
  NANDN U361 ( .A(n8583), .B(n42047), .Z(n229) );
  NANDN U362 ( .A(n8620), .B(n4067), .Z(n230) );
  NAND U363 ( .A(n229), .B(n230), .Z(n8631) );
  NANDN U364 ( .A(n8661), .B(n4068), .Z(n231) );
  NANDN U365 ( .A(n8624), .B(n42115), .Z(n232) );
  AND U366 ( .A(n231), .B(n232), .Z(n8663) );
  NANDN U367 ( .A(n8657), .B(n42047), .Z(n233) );
  NANDN U368 ( .A(n8694), .B(n4067), .Z(n234) );
  NAND U369 ( .A(n233), .B(n234), .Z(n8705) );
  NANDN U370 ( .A(n8732), .B(n4068), .Z(n235) );
  NANDN U371 ( .A(n8695), .B(n42115), .Z(n236) );
  AND U372 ( .A(n235), .B(n236), .Z(n8737) );
  NANDN U373 ( .A(n8731), .B(n42047), .Z(n237) );
  NANDN U374 ( .A(n8768), .B(n4067), .Z(n238) );
  NAND U375 ( .A(n237), .B(n238), .Z(n8779) );
  NANDN U376 ( .A(n8806), .B(n4068), .Z(n239) );
  NANDN U377 ( .A(n8772), .B(n42115), .Z(n240) );
  AND U378 ( .A(n239), .B(n240), .Z(n8811) );
  NANDN U379 ( .A(n8805), .B(n42047), .Z(n241) );
  NANDN U380 ( .A(n8842), .B(n4067), .Z(n242) );
  NAND U381 ( .A(n241), .B(n242), .Z(n8853) );
  NANDN U382 ( .A(n8883), .B(n4068), .Z(n243) );
  NANDN U383 ( .A(n8843), .B(n42115), .Z(n244) );
  AND U384 ( .A(n243), .B(n244), .Z(n8885) );
  NANDN U385 ( .A(n8879), .B(n42047), .Z(n245) );
  NANDN U386 ( .A(n8916), .B(n4067), .Z(n246) );
  NAND U387 ( .A(n245), .B(n246), .Z(n8927) );
  NANDN U388 ( .A(n8957), .B(n4068), .Z(n247) );
  NANDN U389 ( .A(n8920), .B(n42115), .Z(n248) );
  AND U390 ( .A(n247), .B(n248), .Z(n8959) );
  NANDN U391 ( .A(n8953), .B(n42047), .Z(n249) );
  NANDN U392 ( .A(n8990), .B(n4067), .Z(n250) );
  NAND U393 ( .A(n249), .B(n250), .Z(n9001) );
  NANDN U394 ( .A(n9033), .B(n4068), .Z(n251) );
  NANDN U395 ( .A(n8994), .B(n42115), .Z(n252) );
  AND U396 ( .A(n251), .B(n252), .Z(n9038) );
  NANDN U397 ( .A(n9032), .B(n42047), .Z(n253) );
  NANDN U398 ( .A(n9064), .B(n4067), .Z(n254) );
  NAND U399 ( .A(n253), .B(n254), .Z(n9075) );
  NANDN U400 ( .A(n9105), .B(n4068), .Z(n255) );
  NANDN U401 ( .A(n9068), .B(n42115), .Z(n256) );
  AND U402 ( .A(n255), .B(n256), .Z(n9107) );
  NANDN U403 ( .A(n9101), .B(n42047), .Z(n257) );
  NANDN U404 ( .A(n9138), .B(n4067), .Z(n258) );
  NAND U405 ( .A(n257), .B(n258), .Z(n9149) );
  NANDN U406 ( .A(n9179), .B(n4068), .Z(n259) );
  NANDN U407 ( .A(n9142), .B(n42115), .Z(n260) );
  AND U408 ( .A(n259), .B(n260), .Z(n9181) );
  NANDN U409 ( .A(n9175), .B(n42047), .Z(n261) );
  NANDN U410 ( .A(n9212), .B(n4067), .Z(n262) );
  NAND U411 ( .A(n261), .B(n262), .Z(n9223) );
  NANDN U412 ( .A(n9253), .B(n4068), .Z(n263) );
  NANDN U413 ( .A(n9216), .B(n42115), .Z(n264) );
  AND U414 ( .A(n263), .B(n264), .Z(n9255) );
  NANDN U415 ( .A(n9249), .B(n42047), .Z(n265) );
  NANDN U416 ( .A(n9286), .B(n4067), .Z(n266) );
  NAND U417 ( .A(n265), .B(n266), .Z(n9297) );
  NANDN U418 ( .A(n9327), .B(n4068), .Z(n267) );
  NANDN U419 ( .A(n9290), .B(n42115), .Z(n268) );
  AND U420 ( .A(n267), .B(n268), .Z(n9329) );
  NANDN U421 ( .A(n9323), .B(n42047), .Z(n269) );
  NANDN U422 ( .A(n9360), .B(n4067), .Z(n270) );
  NAND U423 ( .A(n269), .B(n270), .Z(n9371) );
  NANDN U424 ( .A(n9398), .B(n4068), .Z(n271) );
  NANDN U425 ( .A(n9364), .B(n42115), .Z(n272) );
  AND U426 ( .A(n271), .B(n272), .Z(n9403) );
  NANDN U427 ( .A(n9397), .B(n42047), .Z(n273) );
  NANDN U428 ( .A(n9434), .B(n4067), .Z(n274) );
  NAND U429 ( .A(n273), .B(n274), .Z(n9445) );
  NANDN U430 ( .A(n9475), .B(n4068), .Z(n275) );
  NANDN U431 ( .A(n9435), .B(n42115), .Z(n276) );
  AND U432 ( .A(n275), .B(n276), .Z(n9477) );
  NANDN U433 ( .A(n9471), .B(n42047), .Z(n277) );
  NANDN U434 ( .A(n9508), .B(n4067), .Z(n278) );
  NAND U435 ( .A(n277), .B(n278), .Z(n9519) );
  NANDN U436 ( .A(n9546), .B(n4068), .Z(n279) );
  NANDN U437 ( .A(n9509), .B(n42115), .Z(n280) );
  AND U438 ( .A(n279), .B(n280), .Z(n9551) );
  NANDN U439 ( .A(n9545), .B(n42047), .Z(n281) );
  NANDN U440 ( .A(n9582), .B(n4067), .Z(n282) );
  NAND U441 ( .A(n281), .B(n282), .Z(n9593) );
  NANDN U442 ( .A(n9623), .B(n4068), .Z(n283) );
  NANDN U443 ( .A(n9586), .B(n42115), .Z(n284) );
  AND U444 ( .A(n283), .B(n284), .Z(n9625) );
  NANDN U445 ( .A(n9619), .B(n42047), .Z(n285) );
  NANDN U446 ( .A(n9656), .B(n4067), .Z(n286) );
  NAND U447 ( .A(n285), .B(n286), .Z(n9667) );
  NANDN U448 ( .A(n9702), .B(n4068), .Z(n287) );
  NANDN U449 ( .A(n9657), .B(n42115), .Z(n288) );
  AND U450 ( .A(n287), .B(n288), .Z(n9704) );
  NANDN U451 ( .A(n9698), .B(n42047), .Z(n289) );
  NANDN U452 ( .A(n9730), .B(n4067), .Z(n290) );
  NAND U453 ( .A(n289), .B(n290), .Z(n9741) );
  NANDN U454 ( .A(n9771), .B(n4068), .Z(n291) );
  NANDN U455 ( .A(n9734), .B(n42115), .Z(n292) );
  AND U456 ( .A(n291), .B(n292), .Z(n9773) );
  NANDN U457 ( .A(n9767), .B(n42047), .Z(n293) );
  NANDN U458 ( .A(n9804), .B(n4067), .Z(n294) );
  NAND U459 ( .A(n293), .B(n294), .Z(n9815) );
  NANDN U460 ( .A(n9842), .B(n4068), .Z(n295) );
  NANDN U461 ( .A(n9808), .B(n42115), .Z(n296) );
  AND U462 ( .A(n295), .B(n296), .Z(n9847) );
  NANDN U463 ( .A(n9841), .B(n42047), .Z(n297) );
  NANDN U464 ( .A(n9878), .B(n4067), .Z(n298) );
  NAND U465 ( .A(n297), .B(n298), .Z(n9889) );
  NANDN U466 ( .A(n9919), .B(n4068), .Z(n299) );
  NANDN U467 ( .A(n9882), .B(n42115), .Z(n300) );
  AND U468 ( .A(n299), .B(n300), .Z(n9921) );
  NANDN U469 ( .A(n9915), .B(n42047), .Z(n301) );
  NANDN U470 ( .A(n9952), .B(n4067), .Z(n302) );
  NAND U471 ( .A(n301), .B(n302), .Z(n9963) );
  NANDN U472 ( .A(n9993), .B(n4068), .Z(n303) );
  NANDN U473 ( .A(n9956), .B(n42115), .Z(n304) );
  AND U474 ( .A(n303), .B(n304), .Z(n9995) );
  NANDN U475 ( .A(n9989), .B(n42047), .Z(n305) );
  NANDN U476 ( .A(n10026), .B(n4067), .Z(n306) );
  NAND U477 ( .A(n305), .B(n306), .Z(n10037) );
  NANDN U478 ( .A(n10067), .B(n4068), .Z(n307) );
  NANDN U479 ( .A(n10030), .B(n42115), .Z(n308) );
  AND U480 ( .A(n307), .B(n308), .Z(n10069) );
  NANDN U481 ( .A(n10063), .B(n42047), .Z(n309) );
  NANDN U482 ( .A(n10100), .B(n4067), .Z(n310) );
  NAND U483 ( .A(n309), .B(n310), .Z(n10111) );
  NANDN U484 ( .A(n10138), .B(n4068), .Z(n311) );
  NANDN U485 ( .A(n10104), .B(n42115), .Z(n312) );
  AND U486 ( .A(n311), .B(n312), .Z(n10143) );
  NANDN U487 ( .A(n10137), .B(n42047), .Z(n313) );
  NANDN U488 ( .A(n10174), .B(n4067), .Z(n314) );
  NAND U489 ( .A(n313), .B(n314), .Z(n10185) );
  NANDN U490 ( .A(n10215), .B(n4068), .Z(n315) );
  NANDN U491 ( .A(n10175), .B(n42115), .Z(n316) );
  AND U492 ( .A(n315), .B(n316), .Z(n10217) );
  NANDN U493 ( .A(n10211), .B(n42047), .Z(n317) );
  NANDN U494 ( .A(n10248), .B(n4067), .Z(n318) );
  NAND U495 ( .A(n317), .B(n318), .Z(n10259) );
  NANDN U496 ( .A(n10289), .B(n4068), .Z(n319) );
  NANDN U497 ( .A(n10252), .B(n42115), .Z(n320) );
  AND U498 ( .A(n319), .B(n320), .Z(n10291) );
  NANDN U499 ( .A(n10285), .B(n42047), .Z(n321) );
  NANDN U500 ( .A(n10322), .B(n4067), .Z(n322) );
  NAND U501 ( .A(n321), .B(n322), .Z(n10333) );
  NANDN U502 ( .A(n10363), .B(n4068), .Z(n323) );
  NANDN U503 ( .A(n10326), .B(n42115), .Z(n324) );
  AND U504 ( .A(n323), .B(n324), .Z(n10365) );
  NANDN U505 ( .A(n10359), .B(n42047), .Z(n325) );
  NANDN U506 ( .A(n10396), .B(n4067), .Z(n326) );
  NAND U507 ( .A(n325), .B(n326), .Z(n10407) );
  NANDN U508 ( .A(n10437), .B(n4068), .Z(n327) );
  NANDN U509 ( .A(n10400), .B(n42115), .Z(n328) );
  AND U510 ( .A(n327), .B(n328), .Z(n10439) );
  NANDN U511 ( .A(n10433), .B(n42047), .Z(n329) );
  NANDN U512 ( .A(n10470), .B(n4067), .Z(n330) );
  NAND U513 ( .A(n329), .B(n330), .Z(n10481) );
  NANDN U514 ( .A(n10511), .B(n4068), .Z(n331) );
  NANDN U515 ( .A(n10474), .B(n42115), .Z(n332) );
  AND U516 ( .A(n331), .B(n332), .Z(n10513) );
  NANDN U517 ( .A(n10507), .B(n42047), .Z(n333) );
  NANDN U518 ( .A(n10544), .B(n4067), .Z(n334) );
  NAND U519 ( .A(n333), .B(n334), .Z(n10555) );
  NANDN U520 ( .A(n10585), .B(n4068), .Z(n335) );
  NANDN U521 ( .A(n10548), .B(n42115), .Z(n336) );
  AND U522 ( .A(n335), .B(n336), .Z(n10587) );
  NANDN U523 ( .A(n10581), .B(n42047), .Z(n337) );
  NANDN U524 ( .A(n10618), .B(n4067), .Z(n338) );
  NAND U525 ( .A(n337), .B(n338), .Z(n10629) );
  NANDN U526 ( .A(n10656), .B(n4068), .Z(n339) );
  NANDN U527 ( .A(n10619), .B(n42115), .Z(n340) );
  AND U528 ( .A(n339), .B(n340), .Z(n10661) );
  NANDN U529 ( .A(n10655), .B(n42047), .Z(n341) );
  NANDN U530 ( .A(n10692), .B(n4067), .Z(n342) );
  NAND U531 ( .A(n341), .B(n342), .Z(n10703) );
  NANDN U532 ( .A(n10730), .B(n4068), .Z(n343) );
  NANDN U533 ( .A(n10696), .B(n42115), .Z(n344) );
  AND U534 ( .A(n343), .B(n344), .Z(n10735) );
  NANDN U535 ( .A(n10729), .B(n42047), .Z(n345) );
  NANDN U536 ( .A(n10766), .B(n4067), .Z(n346) );
  NAND U537 ( .A(n345), .B(n346), .Z(n10777) );
  NANDN U538 ( .A(n10807), .B(n4068), .Z(n347) );
  NANDN U539 ( .A(n10770), .B(n42115), .Z(n348) );
  AND U540 ( .A(n347), .B(n348), .Z(n10809) );
  NANDN U541 ( .A(n10803), .B(n42047), .Z(n349) );
  NANDN U542 ( .A(n10840), .B(n4067), .Z(n350) );
  NAND U543 ( .A(n349), .B(n350), .Z(n10851) );
  NANDN U544 ( .A(n10881), .B(n4068), .Z(n351) );
  NANDN U545 ( .A(n10844), .B(n42115), .Z(n352) );
  AND U546 ( .A(n351), .B(n352), .Z(n10883) );
  NANDN U547 ( .A(n10877), .B(n42047), .Z(n353) );
  NANDN U548 ( .A(n10914), .B(n4067), .Z(n354) );
  NAND U549 ( .A(n353), .B(n354), .Z(n10925) );
  NANDN U550 ( .A(n10955), .B(n4068), .Z(n355) );
  NANDN U551 ( .A(n10918), .B(n42115), .Z(n356) );
  AND U552 ( .A(n355), .B(n356), .Z(n10957) );
  NANDN U553 ( .A(n10951), .B(n42047), .Z(n357) );
  NANDN U554 ( .A(n10988), .B(n4067), .Z(n358) );
  NAND U555 ( .A(n357), .B(n358), .Z(n10999) );
  NANDN U556 ( .A(n11026), .B(n4068), .Z(n359) );
  NANDN U557 ( .A(n10992), .B(n42115), .Z(n360) );
  AND U558 ( .A(n359), .B(n360), .Z(n11031) );
  NANDN U559 ( .A(n11025), .B(n42047), .Z(n361) );
  NANDN U560 ( .A(n11062), .B(n4067), .Z(n362) );
  NAND U561 ( .A(n361), .B(n362), .Z(n11073) );
  NANDN U562 ( .A(n11100), .B(n4068), .Z(n363) );
  NANDN U563 ( .A(n11066), .B(n42115), .Z(n364) );
  AND U564 ( .A(n363), .B(n364), .Z(n11105) );
  NANDN U565 ( .A(n11099), .B(n42047), .Z(n365) );
  NANDN U566 ( .A(n11136), .B(n4067), .Z(n366) );
  NAND U567 ( .A(n365), .B(n366), .Z(n11147) );
  NANDN U568 ( .A(n11177), .B(n4068), .Z(n367) );
  NANDN U569 ( .A(n11137), .B(n42115), .Z(n368) );
  AND U570 ( .A(n367), .B(n368), .Z(n11179) );
  NANDN U571 ( .A(n11173), .B(n42047), .Z(n369) );
  NANDN U572 ( .A(n11210), .B(n4067), .Z(n370) );
  NAND U573 ( .A(n369), .B(n370), .Z(n11221) );
  NANDN U574 ( .A(n11251), .B(n4068), .Z(n371) );
  NANDN U575 ( .A(n11214), .B(n42115), .Z(n372) );
  AND U576 ( .A(n371), .B(n372), .Z(n11253) );
  NANDN U577 ( .A(n11247), .B(n42047), .Z(n373) );
  NANDN U578 ( .A(n11284), .B(n4067), .Z(n374) );
  NAND U579 ( .A(n373), .B(n374), .Z(n11295) );
  NANDN U580 ( .A(n11322), .B(n4068), .Z(n375) );
  NANDN U581 ( .A(n11285), .B(n42115), .Z(n376) );
  AND U582 ( .A(n375), .B(n376), .Z(n11327) );
  NANDN U583 ( .A(n11321), .B(n42047), .Z(n377) );
  NANDN U584 ( .A(n11358), .B(n4067), .Z(n378) );
  NAND U585 ( .A(n377), .B(n378), .Z(n11369) );
  NANDN U586 ( .A(n11396), .B(n4068), .Z(n379) );
  NANDN U587 ( .A(n11362), .B(n42115), .Z(n380) );
  AND U588 ( .A(n379), .B(n380), .Z(n11401) );
  NANDN U589 ( .A(n11395), .B(n42047), .Z(n381) );
  NANDN U590 ( .A(n11432), .B(n4067), .Z(n382) );
  NAND U591 ( .A(n381), .B(n382), .Z(n11443) );
  NANDN U592 ( .A(n11473), .B(n4068), .Z(n383) );
  NANDN U593 ( .A(n11433), .B(n42115), .Z(n384) );
  AND U594 ( .A(n383), .B(n384), .Z(n11475) );
  NANDN U595 ( .A(n11469), .B(n42047), .Z(n385) );
  NANDN U596 ( .A(n11506), .B(n4067), .Z(n386) );
  NAND U597 ( .A(n385), .B(n386), .Z(n11517) );
  NANDN U598 ( .A(n11547), .B(n4068), .Z(n387) );
  NANDN U599 ( .A(n11510), .B(n42115), .Z(n388) );
  AND U600 ( .A(n387), .B(n388), .Z(n11549) );
  NANDN U601 ( .A(n11543), .B(n42047), .Z(n389) );
  NANDN U602 ( .A(n11580), .B(n4067), .Z(n390) );
  NAND U603 ( .A(n389), .B(n390), .Z(n11591) );
  NANDN U604 ( .A(n11621), .B(n4068), .Z(n391) );
  NANDN U605 ( .A(n11581), .B(n42115), .Z(n392) );
  AND U606 ( .A(n391), .B(n392), .Z(n11623) );
  NANDN U607 ( .A(n11617), .B(n42047), .Z(n393) );
  NANDN U608 ( .A(n11654), .B(n4067), .Z(n394) );
  NAND U609 ( .A(n393), .B(n394), .Z(n11665) );
  NANDN U610 ( .A(n11695), .B(n4068), .Z(n395) );
  NANDN U611 ( .A(n11655), .B(n42115), .Z(n396) );
  AND U612 ( .A(n395), .B(n396), .Z(n11697) );
  NANDN U613 ( .A(n11691), .B(n42047), .Z(n397) );
  NANDN U614 ( .A(n11728), .B(n4067), .Z(n398) );
  NAND U615 ( .A(n397), .B(n398), .Z(n11739) );
  NANDN U616 ( .A(n11769), .B(n4068), .Z(n399) );
  NANDN U617 ( .A(n11732), .B(n42115), .Z(n400) );
  AND U618 ( .A(n399), .B(n400), .Z(n11771) );
  NANDN U619 ( .A(n11765), .B(n42047), .Z(n401) );
  NANDN U620 ( .A(n11802), .B(n4067), .Z(n402) );
  NAND U621 ( .A(n401), .B(n402), .Z(n11813) );
  NANDN U622 ( .A(n11843), .B(n4068), .Z(n403) );
  NANDN U623 ( .A(n11803), .B(n42115), .Z(n404) );
  AND U624 ( .A(n403), .B(n404), .Z(n11845) );
  NANDN U625 ( .A(n11839), .B(n42047), .Z(n405) );
  NANDN U626 ( .A(n11876), .B(n4067), .Z(n406) );
  NAND U627 ( .A(n405), .B(n406), .Z(n11887) );
  NANDN U628 ( .A(n11917), .B(n4068), .Z(n407) );
  NANDN U629 ( .A(n11880), .B(n42115), .Z(n408) );
  AND U630 ( .A(n407), .B(n408), .Z(n11919) );
  NANDN U631 ( .A(n11913), .B(n42047), .Z(n409) );
  NANDN U632 ( .A(n11950), .B(n4067), .Z(n410) );
  NAND U633 ( .A(n409), .B(n410), .Z(n11961) );
  NANDN U634 ( .A(n11991), .B(n4068), .Z(n411) );
  NANDN U635 ( .A(n11954), .B(n42115), .Z(n412) );
  AND U636 ( .A(n411), .B(n412), .Z(n11993) );
  NANDN U637 ( .A(n11987), .B(n42047), .Z(n413) );
  NANDN U638 ( .A(n12024), .B(n4067), .Z(n414) );
  NAND U639 ( .A(n413), .B(n414), .Z(n12035) );
  NANDN U640 ( .A(n12065), .B(n4068), .Z(n415) );
  NANDN U641 ( .A(n12025), .B(n42115), .Z(n416) );
  AND U642 ( .A(n415), .B(n416), .Z(n12067) );
  NANDN U643 ( .A(n12061), .B(n42047), .Z(n417) );
  NANDN U644 ( .A(n12098), .B(n4067), .Z(n418) );
  NAND U645 ( .A(n417), .B(n418), .Z(n12109) );
  NANDN U646 ( .A(n12139), .B(n4068), .Z(n419) );
  NANDN U647 ( .A(n12099), .B(n42115), .Z(n420) );
  AND U648 ( .A(n419), .B(n420), .Z(n12141) );
  NANDN U649 ( .A(n12135), .B(n42047), .Z(n421) );
  NANDN U650 ( .A(n12172), .B(n4067), .Z(n422) );
  NAND U651 ( .A(n421), .B(n422), .Z(n12183) );
  NANDN U652 ( .A(n12213), .B(n4068), .Z(n423) );
  NANDN U653 ( .A(n12176), .B(n42115), .Z(n424) );
  AND U654 ( .A(n423), .B(n424), .Z(n12215) );
  NANDN U655 ( .A(n12209), .B(n42047), .Z(n425) );
  NANDN U656 ( .A(n12246), .B(n4067), .Z(n426) );
  NAND U657 ( .A(n425), .B(n426), .Z(n12257) );
  NANDN U658 ( .A(n12284), .B(n4068), .Z(n427) );
  NANDN U659 ( .A(n12250), .B(n42115), .Z(n428) );
  AND U660 ( .A(n427), .B(n428), .Z(n12289) );
  NANDN U661 ( .A(n12283), .B(n42047), .Z(n429) );
  NANDN U662 ( .A(n12320), .B(n4067), .Z(n430) );
  NAND U663 ( .A(n429), .B(n430), .Z(n12331) );
  NANDN U664 ( .A(n12361), .B(n4068), .Z(n431) );
  NANDN U665 ( .A(n12324), .B(n42115), .Z(n432) );
  AND U666 ( .A(n431), .B(n432), .Z(n12363) );
  NANDN U667 ( .A(n12357), .B(n42047), .Z(n433) );
  NANDN U668 ( .A(n12394), .B(n4067), .Z(n434) );
  NAND U669 ( .A(n433), .B(n434), .Z(n12405) );
  NANDN U670 ( .A(n12435), .B(n4068), .Z(n435) );
  NANDN U671 ( .A(n12395), .B(n42115), .Z(n436) );
  AND U672 ( .A(n435), .B(n436), .Z(n12437) );
  NANDN U673 ( .A(n12431), .B(n42047), .Z(n437) );
  NANDN U674 ( .A(n12468), .B(n4067), .Z(n438) );
  NAND U675 ( .A(n437), .B(n438), .Z(n12479) );
  NANDN U676 ( .A(n12506), .B(n4068), .Z(n439) );
  NANDN U677 ( .A(n12472), .B(n42115), .Z(n440) );
  AND U678 ( .A(n439), .B(n440), .Z(n12511) );
  NANDN U679 ( .A(n12505), .B(n42047), .Z(n441) );
  NANDN U680 ( .A(n12542), .B(n4067), .Z(n442) );
  NAND U681 ( .A(n441), .B(n442), .Z(n12553) );
  NANDN U682 ( .A(n12580), .B(n4068), .Z(n443) );
  NANDN U683 ( .A(n12546), .B(n42115), .Z(n444) );
  AND U684 ( .A(n443), .B(n444), .Z(n12585) );
  NANDN U685 ( .A(n12579), .B(n42047), .Z(n445) );
  NANDN U686 ( .A(n12616), .B(n4067), .Z(n446) );
  NAND U687 ( .A(n445), .B(n446), .Z(n12627) );
  NANDN U688 ( .A(n12657), .B(n4068), .Z(n447) );
  NANDN U689 ( .A(n12620), .B(n42115), .Z(n448) );
  AND U690 ( .A(n447), .B(n448), .Z(n12659) );
  NANDN U691 ( .A(n12653), .B(n42047), .Z(n449) );
  NANDN U692 ( .A(n12690), .B(n4067), .Z(n450) );
  NAND U693 ( .A(n449), .B(n450), .Z(n12701) );
  NANDN U694 ( .A(n12731), .B(n4068), .Z(n451) );
  NANDN U695 ( .A(n12694), .B(n42115), .Z(n452) );
  AND U696 ( .A(n451), .B(n452), .Z(n12733) );
  NANDN U697 ( .A(n12727), .B(n42047), .Z(n453) );
  NANDN U698 ( .A(n12764), .B(n4067), .Z(n454) );
  NAND U699 ( .A(n453), .B(n454), .Z(n12775) );
  NANDN U700 ( .A(n12805), .B(n4068), .Z(n455) );
  NANDN U701 ( .A(n12768), .B(n42115), .Z(n456) );
  AND U702 ( .A(n455), .B(n456), .Z(n12807) );
  NANDN U703 ( .A(n12801), .B(n42047), .Z(n457) );
  NANDN U704 ( .A(n12838), .B(n4067), .Z(n458) );
  NAND U705 ( .A(n457), .B(n458), .Z(n12849) );
  NANDN U706 ( .A(n12879), .B(n4068), .Z(n459) );
  NANDN U707 ( .A(n12842), .B(n42115), .Z(n460) );
  AND U708 ( .A(n459), .B(n460), .Z(n12881) );
  NANDN U709 ( .A(n12875), .B(n42047), .Z(n461) );
  NANDN U710 ( .A(n12912), .B(n4067), .Z(n462) );
  NAND U711 ( .A(n461), .B(n462), .Z(n12923) );
  NANDN U712 ( .A(n12950), .B(n4068), .Z(n463) );
  NANDN U713 ( .A(n12916), .B(n42115), .Z(n464) );
  AND U714 ( .A(n463), .B(n464), .Z(n12955) );
  NANDN U715 ( .A(n12949), .B(n42047), .Z(n465) );
  NANDN U716 ( .A(n12986), .B(n4067), .Z(n466) );
  NAND U717 ( .A(n465), .B(n466), .Z(n12997) );
  NANDN U718 ( .A(n13024), .B(n4068), .Z(n467) );
  NANDN U719 ( .A(n12990), .B(n42115), .Z(n468) );
  AND U720 ( .A(n467), .B(n468), .Z(n13029) );
  NANDN U721 ( .A(n13023), .B(n42047), .Z(n469) );
  NANDN U722 ( .A(n13060), .B(n4067), .Z(n470) );
  NAND U723 ( .A(n469), .B(n470), .Z(n13071) );
  NANDN U724 ( .A(n13101), .B(n4068), .Z(n471) );
  NANDN U725 ( .A(n13064), .B(n42115), .Z(n472) );
  AND U726 ( .A(n471), .B(n472), .Z(n13103) );
  NANDN U727 ( .A(n13097), .B(n42047), .Z(n473) );
  NANDN U728 ( .A(n13134), .B(n4067), .Z(n474) );
  NAND U729 ( .A(n473), .B(n474), .Z(n13145) );
  NANDN U730 ( .A(n13175), .B(n4068), .Z(n475) );
  NANDN U731 ( .A(n13138), .B(n42115), .Z(n476) );
  AND U732 ( .A(n475), .B(n476), .Z(n13177) );
  NANDN U733 ( .A(n13171), .B(n42047), .Z(n477) );
  NANDN U734 ( .A(n13208), .B(n4067), .Z(n478) );
  NAND U735 ( .A(n477), .B(n478), .Z(n13219) );
  NANDN U736 ( .A(n13249), .B(n4068), .Z(n479) );
  NANDN U737 ( .A(n13212), .B(n42115), .Z(n480) );
  AND U738 ( .A(n479), .B(n480), .Z(n13251) );
  NANDN U739 ( .A(n13245), .B(n42047), .Z(n481) );
  NANDN U740 ( .A(n13282), .B(n4067), .Z(n482) );
  NAND U741 ( .A(n481), .B(n482), .Z(n13293) );
  NANDN U742 ( .A(n13320), .B(n4068), .Z(n483) );
  NANDN U743 ( .A(n13286), .B(n42115), .Z(n484) );
  AND U744 ( .A(n483), .B(n484), .Z(n13325) );
  NANDN U745 ( .A(n13319), .B(n42047), .Z(n485) );
  NANDN U746 ( .A(n13356), .B(n4067), .Z(n486) );
  NAND U747 ( .A(n485), .B(n486), .Z(n13367) );
  NANDN U748 ( .A(n13397), .B(n4068), .Z(n487) );
  NANDN U749 ( .A(n13360), .B(n42115), .Z(n488) );
  AND U750 ( .A(n487), .B(n488), .Z(n13399) );
  NANDN U751 ( .A(n13393), .B(n42047), .Z(n489) );
  NANDN U752 ( .A(n13430), .B(n4067), .Z(n490) );
  NAND U753 ( .A(n489), .B(n490), .Z(n13441) );
  NANDN U754 ( .A(n13471), .B(n4068), .Z(n491) );
  NANDN U755 ( .A(n13431), .B(n42115), .Z(n492) );
  AND U756 ( .A(n491), .B(n492), .Z(n13473) );
  NANDN U757 ( .A(n13467), .B(n42047), .Z(n493) );
  NANDN U758 ( .A(n13504), .B(n4067), .Z(n494) );
  NAND U759 ( .A(n493), .B(n494), .Z(n13515) );
  NANDN U760 ( .A(n13545), .B(n4068), .Z(n495) );
  NANDN U761 ( .A(n13505), .B(n42115), .Z(n496) );
  AND U762 ( .A(n495), .B(n496), .Z(n13547) );
  NANDN U763 ( .A(n13541), .B(n42047), .Z(n497) );
  NANDN U764 ( .A(n13578), .B(n4067), .Z(n498) );
  NAND U765 ( .A(n497), .B(n498), .Z(n13589) );
  NANDN U766 ( .A(n13619), .B(n4068), .Z(n499) );
  NANDN U767 ( .A(n13582), .B(n42115), .Z(n500) );
  AND U768 ( .A(n499), .B(n500), .Z(n13621) );
  NANDN U769 ( .A(n13615), .B(n42047), .Z(n501) );
  NANDN U770 ( .A(n13652), .B(n4067), .Z(n502) );
  NAND U771 ( .A(n501), .B(n502), .Z(n13663) );
  NANDN U772 ( .A(n13693), .B(n4068), .Z(n503) );
  NANDN U773 ( .A(n13656), .B(n42115), .Z(n504) );
  AND U774 ( .A(n503), .B(n504), .Z(n13695) );
  NANDN U775 ( .A(n13689), .B(n42047), .Z(n505) );
  NANDN U776 ( .A(n13726), .B(n4067), .Z(n506) );
  NAND U777 ( .A(n505), .B(n506), .Z(n13737) );
  NANDN U778 ( .A(n13767), .B(n4068), .Z(n507) );
  NANDN U779 ( .A(n13727), .B(n42115), .Z(n508) );
  AND U780 ( .A(n507), .B(n508), .Z(n13769) );
  NANDN U781 ( .A(n13763), .B(n42047), .Z(n509) );
  NANDN U782 ( .A(n13800), .B(n4067), .Z(n510) );
  NAND U783 ( .A(n509), .B(n510), .Z(n13811) );
  NANDN U784 ( .A(n13841), .B(n4068), .Z(n511) );
  NANDN U785 ( .A(n13804), .B(n42115), .Z(n512) );
  AND U786 ( .A(n511), .B(n512), .Z(n13843) );
  NANDN U787 ( .A(n13837), .B(n42047), .Z(n513) );
  NANDN U788 ( .A(n13874), .B(n4067), .Z(n514) );
  NAND U789 ( .A(n513), .B(n514), .Z(n13885) );
  NANDN U790 ( .A(n13915), .B(n4068), .Z(n515) );
  NANDN U791 ( .A(n13878), .B(n42115), .Z(n516) );
  AND U792 ( .A(n515), .B(n516), .Z(n13917) );
  NANDN U793 ( .A(n13911), .B(n42047), .Z(n517) );
  NANDN U794 ( .A(n13948), .B(n4067), .Z(n518) );
  NAND U795 ( .A(n517), .B(n518), .Z(n13959) );
  NANDN U796 ( .A(n13986), .B(n4068), .Z(n519) );
  NANDN U797 ( .A(n13952), .B(n42115), .Z(n520) );
  AND U798 ( .A(n519), .B(n520), .Z(n13991) );
  NANDN U799 ( .A(n13985), .B(n42047), .Z(n521) );
  NANDN U800 ( .A(n14022), .B(n4067), .Z(n522) );
  NAND U801 ( .A(n521), .B(n522), .Z(n14033) );
  NANDN U802 ( .A(n14063), .B(n4068), .Z(n523) );
  NANDN U803 ( .A(n14026), .B(n42115), .Z(n524) );
  AND U804 ( .A(n523), .B(n524), .Z(n14065) );
  NANDN U805 ( .A(n14059), .B(n42047), .Z(n525) );
  NANDN U806 ( .A(n14101), .B(n4067), .Z(n526) );
  NAND U807 ( .A(n525), .B(n526), .Z(n14112) );
  NANDN U808 ( .A(n14139), .B(n4068), .Z(n527) );
  NANDN U809 ( .A(n14105), .B(n42115), .Z(n528) );
  AND U810 ( .A(n527), .B(n528), .Z(n14144) );
  NANDN U811 ( .A(n14138), .B(n42047), .Z(n529) );
  NANDN U812 ( .A(n14170), .B(n4067), .Z(n530) );
  NAND U813 ( .A(n529), .B(n530), .Z(n14181) );
  NANDN U814 ( .A(n14211), .B(n4068), .Z(n531) );
  NANDN U815 ( .A(n14174), .B(n42115), .Z(n532) );
  AND U816 ( .A(n531), .B(n532), .Z(n14213) );
  NANDN U817 ( .A(n14207), .B(n42047), .Z(n533) );
  NANDN U818 ( .A(n14249), .B(n4067), .Z(n534) );
  NAND U819 ( .A(n533), .B(n534), .Z(n14260) );
  NANDN U820 ( .A(n14285), .B(n4068), .Z(n535) );
  NANDN U821 ( .A(n14253), .B(n42115), .Z(n536) );
  AND U822 ( .A(n535), .B(n536), .Z(n14287) );
  NANDN U823 ( .A(n14281), .B(n42047), .Z(n537) );
  NANDN U824 ( .A(n14318), .B(n4067), .Z(n538) );
  NAND U825 ( .A(n537), .B(n538), .Z(n14329) );
  NANDN U826 ( .A(n14359), .B(n4068), .Z(n539) );
  NANDN U827 ( .A(n14319), .B(n42115), .Z(n540) );
  AND U828 ( .A(n539), .B(n540), .Z(n14361) );
  NANDN U829 ( .A(n14355), .B(n42047), .Z(n541) );
  NANDN U830 ( .A(n14392), .B(n4067), .Z(n542) );
  NAND U831 ( .A(n541), .B(n542), .Z(n14403) );
  NANDN U832 ( .A(n14433), .B(n4068), .Z(n543) );
  NANDN U833 ( .A(n14396), .B(n42115), .Z(n544) );
  AND U834 ( .A(n543), .B(n544), .Z(n14435) );
  NANDN U835 ( .A(n14429), .B(n42047), .Z(n545) );
  NANDN U836 ( .A(n14466), .B(n4067), .Z(n546) );
  NAND U837 ( .A(n545), .B(n546), .Z(n14477) );
  NANDN U838 ( .A(n14504), .B(n4068), .Z(n547) );
  NANDN U839 ( .A(n14470), .B(n42115), .Z(n548) );
  AND U840 ( .A(n547), .B(n548), .Z(n14509) );
  NANDN U841 ( .A(n14503), .B(n42047), .Z(n549) );
  NANDN U842 ( .A(n14540), .B(n4067), .Z(n550) );
  NAND U843 ( .A(n549), .B(n550), .Z(n14551) );
  NANDN U844 ( .A(n14581), .B(n4068), .Z(n551) );
  NANDN U845 ( .A(n14541), .B(n42115), .Z(n552) );
  AND U846 ( .A(n551), .B(n552), .Z(n14583) );
  NANDN U847 ( .A(n14577), .B(n42047), .Z(n553) );
  NANDN U848 ( .A(n14614), .B(n4067), .Z(n554) );
  NAND U849 ( .A(n553), .B(n554), .Z(n14625) );
  NANDN U850 ( .A(n14655), .B(n4068), .Z(n555) );
  NANDN U851 ( .A(n14618), .B(n42115), .Z(n556) );
  AND U852 ( .A(n555), .B(n556), .Z(n14657) );
  NANDN U853 ( .A(n14651), .B(n42047), .Z(n557) );
  NANDN U854 ( .A(n14688), .B(n4067), .Z(n558) );
  NAND U855 ( .A(n557), .B(n558), .Z(n14699) );
  NANDN U856 ( .A(n14729), .B(n4068), .Z(n559) );
  NANDN U857 ( .A(n14692), .B(n42115), .Z(n560) );
  AND U858 ( .A(n559), .B(n560), .Z(n14731) );
  NANDN U859 ( .A(n14725), .B(n42047), .Z(n561) );
  NANDN U860 ( .A(n14762), .B(n4067), .Z(n562) );
  NAND U861 ( .A(n561), .B(n562), .Z(n14773) );
  NANDN U862 ( .A(n14800), .B(n4068), .Z(n563) );
  NANDN U863 ( .A(n14766), .B(n42115), .Z(n564) );
  AND U864 ( .A(n563), .B(n564), .Z(n14805) );
  NANDN U865 ( .A(n14799), .B(n42047), .Z(n565) );
  NANDN U866 ( .A(n14836), .B(n4067), .Z(n566) );
  NAND U867 ( .A(n565), .B(n566), .Z(n14847) );
  NANDN U868 ( .A(n14877), .B(n4068), .Z(n567) );
  NANDN U869 ( .A(n14837), .B(n42115), .Z(n568) );
  AND U870 ( .A(n567), .B(n568), .Z(n14879) );
  NANDN U871 ( .A(n14873), .B(n42047), .Z(n569) );
  NANDN U872 ( .A(n14910), .B(n4067), .Z(n570) );
  NAND U873 ( .A(n569), .B(n570), .Z(n14921) );
  NANDN U874 ( .A(n14951), .B(n4068), .Z(n571) );
  NANDN U875 ( .A(n14914), .B(n42115), .Z(n572) );
  AND U876 ( .A(n571), .B(n572), .Z(n14953) );
  NANDN U877 ( .A(n14947), .B(n42047), .Z(n573) );
  NANDN U878 ( .A(n14984), .B(n4067), .Z(n574) );
  NAND U879 ( .A(n573), .B(n574), .Z(n14995) );
  NANDN U880 ( .A(n15025), .B(n4068), .Z(n575) );
  NANDN U881 ( .A(n14985), .B(n42115), .Z(n576) );
  AND U882 ( .A(n575), .B(n576), .Z(n15027) );
  NANDN U883 ( .A(n15021), .B(n42047), .Z(n577) );
  NANDN U884 ( .A(n15058), .B(n4067), .Z(n578) );
  NAND U885 ( .A(n577), .B(n578), .Z(n15069) );
  NANDN U886 ( .A(n15099), .B(n4068), .Z(n579) );
  NANDN U887 ( .A(n15062), .B(n42115), .Z(n580) );
  AND U888 ( .A(n579), .B(n580), .Z(n15101) );
  NANDN U889 ( .A(n15095), .B(n42047), .Z(n581) );
  NANDN U890 ( .A(n15132), .B(n4067), .Z(n582) );
  NAND U891 ( .A(n581), .B(n582), .Z(n15143) );
  NANDN U892 ( .A(n15170), .B(n4068), .Z(n583) );
  NANDN U893 ( .A(n15136), .B(n42115), .Z(n584) );
  AND U894 ( .A(n583), .B(n584), .Z(n15175) );
  NANDN U895 ( .A(n15169), .B(n42047), .Z(n585) );
  NANDN U896 ( .A(n15206), .B(n4067), .Z(n586) );
  NAND U897 ( .A(n585), .B(n586), .Z(n15217) );
  NANDN U898 ( .A(n15244), .B(n4068), .Z(n587) );
  NANDN U899 ( .A(n15210), .B(n42115), .Z(n588) );
  AND U900 ( .A(n587), .B(n588), .Z(n15249) );
  NANDN U901 ( .A(n15243), .B(n42047), .Z(n589) );
  NANDN U902 ( .A(n15280), .B(n4067), .Z(n590) );
  NAND U903 ( .A(n589), .B(n590), .Z(n15291) );
  NANDN U904 ( .A(n15318), .B(n4068), .Z(n591) );
  NANDN U905 ( .A(n15284), .B(n42115), .Z(n592) );
  AND U906 ( .A(n591), .B(n592), .Z(n15323) );
  NANDN U907 ( .A(n15317), .B(n42047), .Z(n593) );
  NANDN U908 ( .A(n15354), .B(n4067), .Z(n594) );
  NAND U909 ( .A(n593), .B(n594), .Z(n15365) );
  NANDN U910 ( .A(n15395), .B(n4068), .Z(n595) );
  NANDN U911 ( .A(n15355), .B(n42115), .Z(n596) );
  AND U912 ( .A(n595), .B(n596), .Z(n15397) );
  NANDN U913 ( .A(n15391), .B(n42047), .Z(n597) );
  NANDN U914 ( .A(n15428), .B(n4067), .Z(n598) );
  NAND U915 ( .A(n597), .B(n598), .Z(n15439) );
  NANDN U916 ( .A(n15469), .B(n4068), .Z(n599) );
  NANDN U917 ( .A(n15429), .B(n42115), .Z(n600) );
  AND U918 ( .A(n599), .B(n600), .Z(n15471) );
  NANDN U919 ( .A(n15465), .B(n42047), .Z(n601) );
  NANDN U920 ( .A(n15502), .B(n4067), .Z(n602) );
  NAND U921 ( .A(n601), .B(n602), .Z(n15513) );
  NANDN U922 ( .A(n15543), .B(n4068), .Z(n603) );
  NANDN U923 ( .A(n15503), .B(n42115), .Z(n604) );
  AND U924 ( .A(n603), .B(n604), .Z(n15545) );
  NANDN U925 ( .A(n15539), .B(n42047), .Z(n605) );
  NANDN U926 ( .A(n15576), .B(n4067), .Z(n606) );
  NAND U927 ( .A(n605), .B(n606), .Z(n15587) );
  NANDN U928 ( .A(n15617), .B(n4068), .Z(n607) );
  NANDN U929 ( .A(n15580), .B(n42115), .Z(n608) );
  AND U930 ( .A(n607), .B(n608), .Z(n15619) );
  NANDN U931 ( .A(n15613), .B(n42047), .Z(n609) );
  NANDN U932 ( .A(n15650), .B(n4067), .Z(n610) );
  NAND U933 ( .A(n609), .B(n610), .Z(n15661) );
  NANDN U934 ( .A(n15691), .B(n4068), .Z(n611) );
  NANDN U935 ( .A(n15651), .B(n42115), .Z(n612) );
  AND U936 ( .A(n611), .B(n612), .Z(n15693) );
  NANDN U937 ( .A(n15687), .B(n42047), .Z(n613) );
  NANDN U938 ( .A(n15724), .B(n4067), .Z(n614) );
  NAND U939 ( .A(n613), .B(n614), .Z(n15735) );
  NANDN U940 ( .A(n15762), .B(n4068), .Z(n615) );
  NANDN U941 ( .A(n15728), .B(n42115), .Z(n616) );
  AND U942 ( .A(n615), .B(n616), .Z(n15767) );
  NANDN U943 ( .A(n15761), .B(n42047), .Z(n617) );
  NANDN U944 ( .A(n15798), .B(n4067), .Z(n618) );
  NAND U945 ( .A(n617), .B(n618), .Z(n15809) );
  NANDN U946 ( .A(n15836), .B(n4068), .Z(n619) );
  NANDN U947 ( .A(n15802), .B(n42115), .Z(n620) );
  AND U948 ( .A(n619), .B(n620), .Z(n15841) );
  NANDN U949 ( .A(n15835), .B(n42047), .Z(n621) );
  NANDN U950 ( .A(n15872), .B(n4067), .Z(n622) );
  NAND U951 ( .A(n621), .B(n622), .Z(n15883) );
  NANDN U952 ( .A(n15913), .B(n4068), .Z(n623) );
  NANDN U953 ( .A(n15876), .B(n42115), .Z(n624) );
  AND U954 ( .A(n623), .B(n624), .Z(n15915) );
  NANDN U955 ( .A(n15909), .B(n42047), .Z(n625) );
  NANDN U956 ( .A(n15946), .B(n4067), .Z(n626) );
  NAND U957 ( .A(n625), .B(n626), .Z(n15957) );
  NANDN U958 ( .A(n15984), .B(n4068), .Z(n627) );
  NANDN U959 ( .A(n15950), .B(n42115), .Z(n628) );
  AND U960 ( .A(n627), .B(n628), .Z(n15989) );
  NANDN U961 ( .A(n15983), .B(n42047), .Z(n629) );
  NANDN U962 ( .A(n16020), .B(n4067), .Z(n630) );
  NAND U963 ( .A(n629), .B(n630), .Z(n16031) );
  NANDN U964 ( .A(n16058), .B(n4068), .Z(n631) );
  NANDN U965 ( .A(n16024), .B(n42115), .Z(n632) );
  AND U966 ( .A(n631), .B(n632), .Z(n16063) );
  NANDN U967 ( .A(n16057), .B(n42047), .Z(n633) );
  NANDN U968 ( .A(n16094), .B(n4067), .Z(n634) );
  NAND U969 ( .A(n633), .B(n634), .Z(n16105) );
  NANDN U970 ( .A(n16135), .B(n4068), .Z(n635) );
  NANDN U971 ( .A(n16098), .B(n42115), .Z(n636) );
  AND U972 ( .A(n635), .B(n636), .Z(n16137) );
  NANDN U973 ( .A(n16131), .B(n42047), .Z(n637) );
  NANDN U974 ( .A(n16168), .B(n4067), .Z(n638) );
  NAND U975 ( .A(n637), .B(n638), .Z(n16179) );
  NANDN U976 ( .A(n16209), .B(n4068), .Z(n639) );
  NANDN U977 ( .A(n16172), .B(n42115), .Z(n640) );
  AND U978 ( .A(n639), .B(n640), .Z(n16211) );
  NANDN U979 ( .A(n16205), .B(n42047), .Z(n641) );
  NANDN U980 ( .A(n16242), .B(n4067), .Z(n642) );
  NAND U981 ( .A(n641), .B(n642), .Z(n16253) );
  NANDN U982 ( .A(n16283), .B(n4068), .Z(n643) );
  NANDN U983 ( .A(n16243), .B(n42115), .Z(n644) );
  AND U984 ( .A(n643), .B(n644), .Z(n16285) );
  NANDN U985 ( .A(n16279), .B(n42047), .Z(n645) );
  NANDN U986 ( .A(n16316), .B(n4067), .Z(n646) );
  NAND U987 ( .A(n645), .B(n646), .Z(n16327) );
  NANDN U988 ( .A(n16357), .B(n4068), .Z(n647) );
  NANDN U989 ( .A(n16320), .B(n42115), .Z(n648) );
  AND U990 ( .A(n647), .B(n648), .Z(n16359) );
  NANDN U991 ( .A(n16353), .B(n42047), .Z(n649) );
  NANDN U992 ( .A(n16390), .B(n4067), .Z(n650) );
  NAND U993 ( .A(n649), .B(n650), .Z(n16401) );
  NANDN U994 ( .A(n16431), .B(n4068), .Z(n651) );
  NANDN U995 ( .A(n16391), .B(n42115), .Z(n652) );
  AND U996 ( .A(n651), .B(n652), .Z(n16433) );
  NANDN U997 ( .A(n16427), .B(n42047), .Z(n653) );
  NANDN U998 ( .A(n16464), .B(n4067), .Z(n654) );
  NAND U999 ( .A(n653), .B(n654), .Z(n16475) );
  NANDN U1000 ( .A(n16505), .B(n4068), .Z(n655) );
  NANDN U1001 ( .A(n16465), .B(n42115), .Z(n656) );
  AND U1002 ( .A(n655), .B(n656), .Z(n16507) );
  NANDN U1003 ( .A(n16501), .B(n42047), .Z(n657) );
  NANDN U1004 ( .A(n16538), .B(n4067), .Z(n658) );
  NAND U1005 ( .A(n657), .B(n658), .Z(n16549) );
  NANDN U1006 ( .A(n16579), .B(n4068), .Z(n659) );
  NANDN U1007 ( .A(n16539), .B(n42115), .Z(n660) );
  AND U1008 ( .A(n659), .B(n660), .Z(n16581) );
  NANDN U1009 ( .A(n16575), .B(n42047), .Z(n661) );
  NANDN U1010 ( .A(n16612), .B(n4067), .Z(n662) );
  NAND U1011 ( .A(n661), .B(n662), .Z(n16623) );
  NANDN U1012 ( .A(n16653), .B(n4068), .Z(n663) );
  NANDN U1013 ( .A(n16616), .B(n42115), .Z(n664) );
  AND U1014 ( .A(n663), .B(n664), .Z(n16655) );
  NANDN U1015 ( .A(n16649), .B(n42047), .Z(n665) );
  NANDN U1016 ( .A(n16686), .B(n4067), .Z(n666) );
  NAND U1017 ( .A(n665), .B(n666), .Z(n16697) );
  NANDN U1018 ( .A(n16727), .B(n4068), .Z(n667) );
  NANDN U1019 ( .A(n16690), .B(n42115), .Z(n668) );
  AND U1020 ( .A(n667), .B(n668), .Z(n16729) );
  NANDN U1021 ( .A(n16723), .B(n42047), .Z(n669) );
  NANDN U1022 ( .A(n16760), .B(n4067), .Z(n670) );
  NAND U1023 ( .A(n669), .B(n670), .Z(n16771) );
  NANDN U1024 ( .A(n16801), .B(n4068), .Z(n671) );
  NANDN U1025 ( .A(n16764), .B(n42115), .Z(n672) );
  AND U1026 ( .A(n671), .B(n672), .Z(n16803) );
  NANDN U1027 ( .A(n16797), .B(n42047), .Z(n673) );
  NANDN U1028 ( .A(n16834), .B(n4067), .Z(n674) );
  NAND U1029 ( .A(n673), .B(n674), .Z(n16845) );
  NANDN U1030 ( .A(n16872), .B(n4068), .Z(n675) );
  NANDN U1031 ( .A(n16838), .B(n42115), .Z(n676) );
  AND U1032 ( .A(n675), .B(n676), .Z(n16877) );
  NANDN U1033 ( .A(n16871), .B(n42047), .Z(n677) );
  NANDN U1034 ( .A(n16908), .B(n4067), .Z(n678) );
  NAND U1035 ( .A(n677), .B(n678), .Z(n16919) );
  NANDN U1036 ( .A(n16949), .B(n4068), .Z(n679) );
  NANDN U1037 ( .A(n16912), .B(n42115), .Z(n680) );
  AND U1038 ( .A(n679), .B(n680), .Z(n16951) );
  NANDN U1039 ( .A(n16945), .B(n42047), .Z(n681) );
  NANDN U1040 ( .A(n16982), .B(n4067), .Z(n682) );
  NAND U1041 ( .A(n681), .B(n682), .Z(n16993) );
  NANDN U1042 ( .A(n17023), .B(n4068), .Z(n683) );
  NANDN U1043 ( .A(n16986), .B(n42115), .Z(n684) );
  AND U1044 ( .A(n683), .B(n684), .Z(n17025) );
  NANDN U1045 ( .A(n17019), .B(n42047), .Z(n685) );
  NANDN U1046 ( .A(n17056), .B(n4067), .Z(n686) );
  NAND U1047 ( .A(n685), .B(n686), .Z(n17067) );
  NANDN U1048 ( .A(n17094), .B(n4068), .Z(n687) );
  NANDN U1049 ( .A(n17060), .B(n42115), .Z(n688) );
  AND U1050 ( .A(n687), .B(n688), .Z(n17099) );
  NANDN U1051 ( .A(n17093), .B(n42047), .Z(n689) );
  NANDN U1052 ( .A(n17130), .B(n4067), .Z(n690) );
  NAND U1053 ( .A(n689), .B(n690), .Z(n17141) );
  NANDN U1054 ( .A(n17168), .B(n4068), .Z(n691) );
  NANDN U1055 ( .A(n17134), .B(n42115), .Z(n692) );
  AND U1056 ( .A(n691), .B(n692), .Z(n17173) );
  NANDN U1057 ( .A(n17167), .B(n42047), .Z(n693) );
  NANDN U1058 ( .A(n17204), .B(n4067), .Z(n694) );
  NAND U1059 ( .A(n693), .B(n694), .Z(n17215) );
  NANDN U1060 ( .A(n17242), .B(n4068), .Z(n695) );
  NANDN U1061 ( .A(n17208), .B(n42115), .Z(n696) );
  AND U1062 ( .A(n695), .B(n696), .Z(n17247) );
  NANDN U1063 ( .A(n17241), .B(n42047), .Z(n697) );
  NANDN U1064 ( .A(n17278), .B(n4067), .Z(n698) );
  NAND U1065 ( .A(n697), .B(n698), .Z(n17289) );
  NANDN U1066 ( .A(n17319), .B(n4068), .Z(n699) );
  NANDN U1067 ( .A(n17282), .B(n42115), .Z(n700) );
  AND U1068 ( .A(n699), .B(n700), .Z(n17321) );
  NANDN U1069 ( .A(n17315), .B(n42047), .Z(n701) );
  NANDN U1070 ( .A(n17352), .B(n4067), .Z(n702) );
  NAND U1071 ( .A(n701), .B(n702), .Z(n17363) );
  NANDN U1072 ( .A(n17390), .B(n4068), .Z(n703) );
  NANDN U1073 ( .A(n17356), .B(n42115), .Z(n704) );
  AND U1074 ( .A(n703), .B(n704), .Z(n17395) );
  NANDN U1075 ( .A(n17389), .B(n42047), .Z(n705) );
  NANDN U1076 ( .A(n17426), .B(n4067), .Z(n706) );
  NAND U1077 ( .A(n705), .B(n706), .Z(n17437) );
  NANDN U1078 ( .A(n17467), .B(n4068), .Z(n707) );
  NANDN U1079 ( .A(n17430), .B(n42115), .Z(n708) );
  AND U1080 ( .A(n707), .B(n708), .Z(n17469) );
  NANDN U1081 ( .A(n17463), .B(n42047), .Z(n709) );
  NANDN U1082 ( .A(n17500), .B(n4067), .Z(n710) );
  NAND U1083 ( .A(n709), .B(n710), .Z(n17511) );
  NANDN U1084 ( .A(n17541), .B(n4068), .Z(n711) );
  NANDN U1085 ( .A(n17504), .B(n42115), .Z(n712) );
  AND U1086 ( .A(n711), .B(n712), .Z(n17543) );
  NANDN U1087 ( .A(n17537), .B(n42047), .Z(n713) );
  NANDN U1088 ( .A(n17574), .B(n4067), .Z(n714) );
  NAND U1089 ( .A(n713), .B(n714), .Z(n17585) );
  NANDN U1090 ( .A(n17615), .B(n4068), .Z(n715) );
  NANDN U1091 ( .A(n17578), .B(n42115), .Z(n716) );
  AND U1092 ( .A(n715), .B(n716), .Z(n17617) );
  NANDN U1093 ( .A(n17611), .B(n42047), .Z(n717) );
  NANDN U1094 ( .A(n17648), .B(n4067), .Z(n718) );
  NAND U1095 ( .A(n717), .B(n718), .Z(n17659) );
  NANDN U1096 ( .A(n17689), .B(n4068), .Z(n719) );
  NANDN U1097 ( .A(n17649), .B(n42115), .Z(n720) );
  AND U1098 ( .A(n719), .B(n720), .Z(n17691) );
  NANDN U1099 ( .A(n17685), .B(n42047), .Z(n721) );
  NANDN U1100 ( .A(n17722), .B(n4067), .Z(n722) );
  NAND U1101 ( .A(n721), .B(n722), .Z(n17733) );
  NANDN U1102 ( .A(n17763), .B(n4068), .Z(n723) );
  NANDN U1103 ( .A(n17726), .B(n42115), .Z(n724) );
  AND U1104 ( .A(n723), .B(n724), .Z(n17765) );
  NANDN U1105 ( .A(n17759), .B(n42047), .Z(n725) );
  NANDN U1106 ( .A(n17796), .B(n4067), .Z(n726) );
  NAND U1107 ( .A(n725), .B(n726), .Z(n17807) );
  NANDN U1108 ( .A(n17837), .B(n4068), .Z(n727) );
  NANDN U1109 ( .A(n17797), .B(n42115), .Z(n728) );
  AND U1110 ( .A(n727), .B(n728), .Z(n17839) );
  NANDN U1111 ( .A(n17833), .B(n42047), .Z(n729) );
  NANDN U1112 ( .A(n17870), .B(n4067), .Z(n730) );
  NAND U1113 ( .A(n729), .B(n730), .Z(n17881) );
  NANDN U1114 ( .A(n17911), .B(n4068), .Z(n731) );
  NANDN U1115 ( .A(n17874), .B(n42115), .Z(n732) );
  AND U1116 ( .A(n731), .B(n732), .Z(n17913) );
  NANDN U1117 ( .A(n17907), .B(n42047), .Z(n733) );
  NANDN U1118 ( .A(n17944), .B(n4067), .Z(n734) );
  NAND U1119 ( .A(n733), .B(n734), .Z(n17955) );
  NANDN U1120 ( .A(n17985), .B(n4068), .Z(n735) );
  NANDN U1121 ( .A(n17948), .B(n42115), .Z(n736) );
  AND U1122 ( .A(n735), .B(n736), .Z(n17987) );
  NANDN U1123 ( .A(n17981), .B(n42047), .Z(n737) );
  NANDN U1124 ( .A(n18018), .B(n4067), .Z(n738) );
  NAND U1125 ( .A(n737), .B(n738), .Z(n18029) );
  NANDN U1126 ( .A(n18059), .B(n4068), .Z(n739) );
  NANDN U1127 ( .A(n18022), .B(n42115), .Z(n740) );
  AND U1128 ( .A(n739), .B(n740), .Z(n18061) );
  NANDN U1129 ( .A(n18055), .B(n42047), .Z(n741) );
  NANDN U1130 ( .A(n18092), .B(n4067), .Z(n742) );
  NAND U1131 ( .A(n741), .B(n742), .Z(n18103) );
  NANDN U1132 ( .A(n18133), .B(n4068), .Z(n743) );
  NANDN U1133 ( .A(n18096), .B(n42115), .Z(n744) );
  AND U1134 ( .A(n743), .B(n744), .Z(n18135) );
  NANDN U1135 ( .A(n18129), .B(n42047), .Z(n745) );
  NANDN U1136 ( .A(n18166), .B(n4067), .Z(n746) );
  NAND U1137 ( .A(n745), .B(n746), .Z(n18177) );
  NANDN U1138 ( .A(n18207), .B(n4068), .Z(n747) );
  NANDN U1139 ( .A(n18167), .B(n42115), .Z(n748) );
  AND U1140 ( .A(n747), .B(n748), .Z(n18209) );
  NANDN U1141 ( .A(n18203), .B(n42047), .Z(n749) );
  NANDN U1142 ( .A(n18240), .B(n4067), .Z(n750) );
  NAND U1143 ( .A(n749), .B(n750), .Z(n18251) );
  NANDN U1144 ( .A(n18281), .B(n4068), .Z(n751) );
  NANDN U1145 ( .A(n18244), .B(n42115), .Z(n752) );
  AND U1146 ( .A(n751), .B(n752), .Z(n18283) );
  NANDN U1147 ( .A(n18277), .B(n42047), .Z(n753) );
  NANDN U1148 ( .A(n18314), .B(n4067), .Z(n754) );
  NAND U1149 ( .A(n753), .B(n754), .Z(n18325) );
  NANDN U1150 ( .A(n18355), .B(n4068), .Z(n755) );
  NANDN U1151 ( .A(n18318), .B(n42115), .Z(n756) );
  AND U1152 ( .A(n755), .B(n756), .Z(n18357) );
  NANDN U1153 ( .A(n18351), .B(n42047), .Z(n757) );
  NANDN U1154 ( .A(n18388), .B(n4067), .Z(n758) );
  NAND U1155 ( .A(n757), .B(n758), .Z(n18399) );
  NANDN U1156 ( .A(n18429), .B(n4068), .Z(n759) );
  NANDN U1157 ( .A(n18392), .B(n42115), .Z(n760) );
  AND U1158 ( .A(n759), .B(n760), .Z(n18431) );
  NANDN U1159 ( .A(n18425), .B(n42047), .Z(n761) );
  NANDN U1160 ( .A(n18462), .B(n4067), .Z(n762) );
  NAND U1161 ( .A(n761), .B(n762), .Z(n18473) );
  NANDN U1162 ( .A(n18503), .B(n4068), .Z(n763) );
  NANDN U1163 ( .A(n18463), .B(n42115), .Z(n764) );
  AND U1164 ( .A(n763), .B(n764), .Z(n18505) );
  NANDN U1165 ( .A(n18499), .B(n42047), .Z(n765) );
  NANDN U1166 ( .A(n18536), .B(n4067), .Z(n766) );
  NAND U1167 ( .A(n765), .B(n766), .Z(n18547) );
  NANDN U1168 ( .A(n18577), .B(n4068), .Z(n767) );
  NANDN U1169 ( .A(n18540), .B(n42115), .Z(n768) );
  AND U1170 ( .A(n767), .B(n768), .Z(n18579) );
  NANDN U1171 ( .A(n18573), .B(n42047), .Z(n769) );
  NANDN U1172 ( .A(n18610), .B(n4067), .Z(n770) );
  NAND U1173 ( .A(n769), .B(n770), .Z(n18621) );
  NANDN U1174 ( .A(n18648), .B(n4068), .Z(n771) );
  NANDN U1175 ( .A(n18611), .B(n42115), .Z(n772) );
  AND U1176 ( .A(n771), .B(n772), .Z(n18653) );
  NANDN U1177 ( .A(n18647), .B(n42047), .Z(n773) );
  NANDN U1178 ( .A(n18684), .B(n4067), .Z(n774) );
  NAND U1179 ( .A(n773), .B(n774), .Z(n18695) );
  NANDN U1180 ( .A(n18725), .B(n4068), .Z(n775) );
  NANDN U1181 ( .A(n18688), .B(n42115), .Z(n776) );
  AND U1182 ( .A(n775), .B(n776), .Z(n18727) );
  NANDN U1183 ( .A(n18721), .B(n42047), .Z(n777) );
  NANDN U1184 ( .A(n18758), .B(n4067), .Z(n778) );
  NAND U1185 ( .A(n777), .B(n778), .Z(n18769) );
  NANDN U1186 ( .A(n18796), .B(n4068), .Z(n779) );
  NANDN U1187 ( .A(n18759), .B(n42115), .Z(n780) );
  AND U1188 ( .A(n779), .B(n780), .Z(n18801) );
  NANDN U1189 ( .A(n18795), .B(n42047), .Z(n781) );
  NANDN U1190 ( .A(n18832), .B(n4067), .Z(n782) );
  NAND U1191 ( .A(n781), .B(n782), .Z(n18843) );
  NANDN U1192 ( .A(n18873), .B(n4068), .Z(n783) );
  NANDN U1193 ( .A(n18833), .B(n42115), .Z(n784) );
  AND U1194 ( .A(n783), .B(n784), .Z(n18875) );
  NANDN U1195 ( .A(n18869), .B(n42047), .Z(n785) );
  NANDN U1196 ( .A(n18906), .B(n4067), .Z(n786) );
  NAND U1197 ( .A(n785), .B(n786), .Z(n18917) );
  NANDN U1198 ( .A(n18944), .B(n4068), .Z(n787) );
  NANDN U1199 ( .A(n18907), .B(n42115), .Z(n788) );
  AND U1200 ( .A(n787), .B(n788), .Z(n18949) );
  NANDN U1201 ( .A(n18943), .B(n42047), .Z(n789) );
  NANDN U1202 ( .A(n18980), .B(n4067), .Z(n790) );
  NAND U1203 ( .A(n789), .B(n790), .Z(n18991) );
  NANDN U1204 ( .A(n19018), .B(n4068), .Z(n791) );
  NANDN U1205 ( .A(n18984), .B(n42115), .Z(n792) );
  AND U1206 ( .A(n791), .B(n792), .Z(n19023) );
  NANDN U1207 ( .A(n19017), .B(n42047), .Z(n793) );
  NANDN U1208 ( .A(n19054), .B(n4067), .Z(n794) );
  NAND U1209 ( .A(n793), .B(n794), .Z(n19065) );
  NANDN U1210 ( .A(n19092), .B(n4068), .Z(n795) );
  NANDN U1211 ( .A(n19058), .B(n42115), .Z(n796) );
  AND U1212 ( .A(n795), .B(n796), .Z(n19097) );
  NANDN U1213 ( .A(n19091), .B(n42047), .Z(n797) );
  NANDN U1214 ( .A(n19128), .B(n4067), .Z(n798) );
  NAND U1215 ( .A(n797), .B(n798), .Z(n19139) );
  NANDN U1216 ( .A(n19166), .B(n4068), .Z(n799) );
  NANDN U1217 ( .A(n19132), .B(n42115), .Z(n800) );
  AND U1218 ( .A(n799), .B(n800), .Z(n19171) );
  NANDN U1219 ( .A(n19165), .B(n42047), .Z(n801) );
  NANDN U1220 ( .A(n19202), .B(n4067), .Z(n802) );
  NAND U1221 ( .A(n801), .B(n802), .Z(n19213) );
  NANDN U1222 ( .A(n19243), .B(n4068), .Z(n803) );
  NANDN U1223 ( .A(n19206), .B(n42115), .Z(n804) );
  AND U1224 ( .A(n803), .B(n804), .Z(n19245) );
  NANDN U1225 ( .A(n19239), .B(n42047), .Z(n805) );
  NANDN U1226 ( .A(n19276), .B(n4067), .Z(n806) );
  NAND U1227 ( .A(n805), .B(n806), .Z(n19287) );
  NANDN U1228 ( .A(n19317), .B(n4068), .Z(n807) );
  NANDN U1229 ( .A(n19280), .B(n42115), .Z(n808) );
  AND U1230 ( .A(n807), .B(n808), .Z(n19319) );
  NANDN U1231 ( .A(n19313), .B(n42047), .Z(n809) );
  NANDN U1232 ( .A(n19350), .B(n4067), .Z(n810) );
  NAND U1233 ( .A(n809), .B(n810), .Z(n19361) );
  NANDN U1234 ( .A(n19391), .B(n4068), .Z(n811) );
  NANDN U1235 ( .A(n19354), .B(n42115), .Z(n812) );
  AND U1236 ( .A(n811), .B(n812), .Z(n19393) );
  NANDN U1237 ( .A(n19387), .B(n42047), .Z(n813) );
  NANDN U1238 ( .A(n19424), .B(n4067), .Z(n814) );
  NAND U1239 ( .A(n813), .B(n814), .Z(n19435) );
  NANDN U1240 ( .A(n19465), .B(n4068), .Z(n815) );
  NANDN U1241 ( .A(n19425), .B(n42115), .Z(n816) );
  AND U1242 ( .A(n815), .B(n816), .Z(n19467) );
  NANDN U1243 ( .A(n19461), .B(n42047), .Z(n817) );
  NANDN U1244 ( .A(n19498), .B(n4067), .Z(n818) );
  NAND U1245 ( .A(n817), .B(n818), .Z(n19509) );
  NANDN U1246 ( .A(n19539), .B(n4068), .Z(n819) );
  NANDN U1247 ( .A(n19502), .B(n42115), .Z(n820) );
  AND U1248 ( .A(n819), .B(n820), .Z(n19541) );
  NANDN U1249 ( .A(n19535), .B(n42047), .Z(n821) );
  NANDN U1250 ( .A(n19572), .B(n4067), .Z(n822) );
  NAND U1251 ( .A(n821), .B(n822), .Z(n19583) );
  NANDN U1252 ( .A(n19613), .B(n4068), .Z(n823) );
  NANDN U1253 ( .A(n19576), .B(n42115), .Z(n824) );
  AND U1254 ( .A(n823), .B(n824), .Z(n19615) );
  NANDN U1255 ( .A(n19609), .B(n42047), .Z(n825) );
  NANDN U1256 ( .A(n19646), .B(n4067), .Z(n826) );
  NAND U1257 ( .A(n825), .B(n826), .Z(n19657) );
  NANDN U1258 ( .A(n19687), .B(n4068), .Z(n827) );
  NANDN U1259 ( .A(n19650), .B(n42115), .Z(n828) );
  AND U1260 ( .A(n827), .B(n828), .Z(n19689) );
  NANDN U1261 ( .A(n19683), .B(n42047), .Z(n829) );
  NANDN U1262 ( .A(n19720), .B(n4067), .Z(n830) );
  NAND U1263 ( .A(n829), .B(n830), .Z(n19731) );
  NANDN U1264 ( .A(n19761), .B(n4068), .Z(n831) );
  NANDN U1265 ( .A(n19721), .B(n42115), .Z(n832) );
  AND U1266 ( .A(n831), .B(n832), .Z(n19763) );
  NANDN U1267 ( .A(n19757), .B(n42047), .Z(n833) );
  NANDN U1268 ( .A(n19794), .B(n4067), .Z(n834) );
  NAND U1269 ( .A(n833), .B(n834), .Z(n19805) );
  NANDN U1270 ( .A(n19832), .B(n4068), .Z(n835) );
  NANDN U1271 ( .A(n19798), .B(n42115), .Z(n836) );
  AND U1272 ( .A(n835), .B(n836), .Z(n19837) );
  NANDN U1273 ( .A(n19831), .B(n42047), .Z(n837) );
  NANDN U1274 ( .A(n19868), .B(n4067), .Z(n838) );
  NAND U1275 ( .A(n837), .B(n838), .Z(n19879) );
  NANDN U1276 ( .A(n19909), .B(n4068), .Z(n839) );
  NANDN U1277 ( .A(n19872), .B(n42115), .Z(n840) );
  AND U1278 ( .A(n839), .B(n840), .Z(n19911) );
  NANDN U1279 ( .A(n19905), .B(n42047), .Z(n841) );
  NANDN U1280 ( .A(n19942), .B(n4067), .Z(n842) );
  NAND U1281 ( .A(n841), .B(n842), .Z(n19953) );
  NANDN U1282 ( .A(n19980), .B(n4068), .Z(n843) );
  NANDN U1283 ( .A(n19946), .B(n42115), .Z(n844) );
  AND U1284 ( .A(n843), .B(n844), .Z(n19985) );
  NANDN U1285 ( .A(n19979), .B(n42047), .Z(n845) );
  NANDN U1286 ( .A(n20016), .B(n4067), .Z(n846) );
  NAND U1287 ( .A(n845), .B(n846), .Z(n20027) );
  NANDN U1288 ( .A(n20057), .B(n4068), .Z(n847) );
  NANDN U1289 ( .A(n20020), .B(n42115), .Z(n848) );
  AND U1290 ( .A(n847), .B(n848), .Z(n20059) );
  NANDN U1291 ( .A(n20053), .B(n42047), .Z(n849) );
  NANDN U1292 ( .A(n20090), .B(n4067), .Z(n850) );
  NAND U1293 ( .A(n849), .B(n850), .Z(n20101) );
  NANDN U1294 ( .A(n20131), .B(n4068), .Z(n851) );
  NANDN U1295 ( .A(n20094), .B(n42115), .Z(n852) );
  AND U1296 ( .A(n851), .B(n852), .Z(n20133) );
  NANDN U1297 ( .A(n20127), .B(n42047), .Z(n853) );
  NANDN U1298 ( .A(n20164), .B(n4067), .Z(n854) );
  NAND U1299 ( .A(n853), .B(n854), .Z(n20175) );
  NANDN U1300 ( .A(n20205), .B(n4068), .Z(n855) );
  NANDN U1301 ( .A(n20165), .B(n42115), .Z(n856) );
  AND U1302 ( .A(n855), .B(n856), .Z(n20207) );
  NANDN U1303 ( .A(n20201), .B(n42047), .Z(n857) );
  NANDN U1304 ( .A(n20238), .B(n4067), .Z(n858) );
  NAND U1305 ( .A(n857), .B(n858), .Z(n20249) );
  NANDN U1306 ( .A(n20279), .B(n4068), .Z(n859) );
  NANDN U1307 ( .A(n20242), .B(n42115), .Z(n860) );
  AND U1308 ( .A(n859), .B(n860), .Z(n20281) );
  NANDN U1309 ( .A(n20275), .B(n42047), .Z(n861) );
  NANDN U1310 ( .A(n20312), .B(n4067), .Z(n862) );
  NAND U1311 ( .A(n861), .B(n862), .Z(n20323) );
  NANDN U1312 ( .A(n20353), .B(n4068), .Z(n863) );
  NANDN U1313 ( .A(n20316), .B(n42115), .Z(n864) );
  AND U1314 ( .A(n863), .B(n864), .Z(n20355) );
  NANDN U1315 ( .A(n20349), .B(n42047), .Z(n865) );
  NANDN U1316 ( .A(n20386), .B(n4067), .Z(n866) );
  NAND U1317 ( .A(n865), .B(n866), .Z(n20397) );
  NANDN U1318 ( .A(n20424), .B(n4068), .Z(n867) );
  NANDN U1319 ( .A(n20390), .B(n42115), .Z(n868) );
  AND U1320 ( .A(n867), .B(n868), .Z(n20429) );
  NANDN U1321 ( .A(n20423), .B(n42047), .Z(n869) );
  NANDN U1322 ( .A(n20460), .B(n4067), .Z(n870) );
  NAND U1323 ( .A(n869), .B(n870), .Z(n20471) );
  NANDN U1324 ( .A(n20501), .B(n4068), .Z(n871) );
  NANDN U1325 ( .A(n20464), .B(n42115), .Z(n872) );
  AND U1326 ( .A(n871), .B(n872), .Z(n20503) );
  NANDN U1327 ( .A(n20497), .B(n42047), .Z(n873) );
  NANDN U1328 ( .A(n20534), .B(n4067), .Z(n874) );
  NAND U1329 ( .A(n873), .B(n874), .Z(n20545) );
  NANDN U1330 ( .A(n20572), .B(n4068), .Z(n875) );
  NANDN U1331 ( .A(n20538), .B(n42115), .Z(n876) );
  AND U1332 ( .A(n875), .B(n876), .Z(n20577) );
  NANDN U1333 ( .A(n20571), .B(n42047), .Z(n877) );
  NANDN U1334 ( .A(n20608), .B(n4067), .Z(n878) );
  NAND U1335 ( .A(n877), .B(n878), .Z(n20619) );
  NANDN U1336 ( .A(n20649), .B(n4068), .Z(n879) );
  NANDN U1337 ( .A(n20612), .B(n42115), .Z(n880) );
  AND U1338 ( .A(n879), .B(n880), .Z(n20651) );
  NANDN U1339 ( .A(n20645), .B(n42047), .Z(n881) );
  NANDN U1340 ( .A(n20682), .B(n4067), .Z(n882) );
  NAND U1341 ( .A(n881), .B(n882), .Z(n20693) );
  NANDN U1342 ( .A(n20723), .B(n4068), .Z(n883) );
  NANDN U1343 ( .A(n20686), .B(n42115), .Z(n884) );
  AND U1344 ( .A(n883), .B(n884), .Z(n20725) );
  NANDN U1345 ( .A(n20719), .B(n42047), .Z(n885) );
  NANDN U1346 ( .A(n20756), .B(n4067), .Z(n886) );
  NAND U1347 ( .A(n885), .B(n886), .Z(n20767) );
  NANDN U1348 ( .A(n20797), .B(n4068), .Z(n887) );
  NANDN U1349 ( .A(n20760), .B(n42115), .Z(n888) );
  AND U1350 ( .A(n887), .B(n888), .Z(n20799) );
  NANDN U1351 ( .A(n20793), .B(n42047), .Z(n889) );
  NANDN U1352 ( .A(n20830), .B(n4067), .Z(n890) );
  NAND U1353 ( .A(n889), .B(n890), .Z(n20841) );
  NANDN U1354 ( .A(n20871), .B(n4068), .Z(n891) );
  NANDN U1355 ( .A(n20834), .B(n42115), .Z(n892) );
  AND U1356 ( .A(n891), .B(n892), .Z(n20873) );
  NANDN U1357 ( .A(n20867), .B(n42047), .Z(n893) );
  NANDN U1358 ( .A(n20904), .B(n4067), .Z(n894) );
  NAND U1359 ( .A(n893), .B(n894), .Z(n20915) );
  NANDN U1360 ( .A(n20945), .B(n4068), .Z(n895) );
  NANDN U1361 ( .A(n20908), .B(n42115), .Z(n896) );
  AND U1362 ( .A(n895), .B(n896), .Z(n20947) );
  NANDN U1363 ( .A(n20941), .B(n42047), .Z(n897) );
  NANDN U1364 ( .A(n20978), .B(n4067), .Z(n898) );
  NAND U1365 ( .A(n897), .B(n898), .Z(n20989) );
  NANDN U1366 ( .A(n21019), .B(n4068), .Z(n899) );
  NANDN U1367 ( .A(n20982), .B(n42115), .Z(n900) );
  AND U1368 ( .A(n899), .B(n900), .Z(n21021) );
  NANDN U1369 ( .A(n21015), .B(n42047), .Z(n901) );
  NANDN U1370 ( .A(n21052), .B(n4067), .Z(n902) );
  NAND U1371 ( .A(n901), .B(n902), .Z(n21063) );
  NANDN U1372 ( .A(n21093), .B(n4068), .Z(n903) );
  NANDN U1373 ( .A(n21053), .B(n42115), .Z(n904) );
  AND U1374 ( .A(n903), .B(n904), .Z(n21095) );
  NANDN U1375 ( .A(n21089), .B(n42047), .Z(n905) );
  NANDN U1376 ( .A(n21126), .B(n4067), .Z(n906) );
  NAND U1377 ( .A(n905), .B(n906), .Z(n21137) );
  NANDN U1378 ( .A(n21167), .B(n4068), .Z(n907) );
  NANDN U1379 ( .A(n21130), .B(n42115), .Z(n908) );
  AND U1380 ( .A(n907), .B(n908), .Z(n21169) );
  NANDN U1381 ( .A(n21163), .B(n42047), .Z(n909) );
  NANDN U1382 ( .A(n21200), .B(n4067), .Z(n910) );
  NAND U1383 ( .A(n909), .B(n910), .Z(n21211) );
  NANDN U1384 ( .A(n21238), .B(n4068), .Z(n911) );
  NANDN U1385 ( .A(n21201), .B(n42115), .Z(n912) );
  AND U1386 ( .A(n911), .B(n912), .Z(n21243) );
  NANDN U1387 ( .A(n21237), .B(n42047), .Z(n913) );
  NANDN U1388 ( .A(n21274), .B(n4067), .Z(n914) );
  NAND U1389 ( .A(n913), .B(n914), .Z(n21285) );
  NANDN U1390 ( .A(n21312), .B(n4068), .Z(n915) );
  NANDN U1391 ( .A(n21278), .B(n42115), .Z(n916) );
  AND U1392 ( .A(n915), .B(n916), .Z(n21317) );
  NANDN U1393 ( .A(n21311), .B(n42047), .Z(n917) );
  NANDN U1394 ( .A(n21348), .B(n4067), .Z(n918) );
  NAND U1395 ( .A(n917), .B(n918), .Z(n21359) );
  NANDN U1396 ( .A(n21389), .B(n4068), .Z(n919) );
  NANDN U1397 ( .A(n21352), .B(n42115), .Z(n920) );
  AND U1398 ( .A(n919), .B(n920), .Z(n21391) );
  NANDN U1399 ( .A(n21385), .B(n42047), .Z(n921) );
  NANDN U1400 ( .A(n21422), .B(n4067), .Z(n922) );
  NAND U1401 ( .A(n921), .B(n922), .Z(n21433) );
  NANDN U1402 ( .A(n21463), .B(n4068), .Z(n923) );
  NANDN U1403 ( .A(n21423), .B(n42115), .Z(n924) );
  AND U1404 ( .A(n923), .B(n924), .Z(n21465) );
  NANDN U1405 ( .A(n21459), .B(n42047), .Z(n925) );
  NANDN U1406 ( .A(n21496), .B(n4067), .Z(n926) );
  NAND U1407 ( .A(n925), .B(n926), .Z(n21507) );
  NANDN U1408 ( .A(n21537), .B(n4068), .Z(n927) );
  NANDN U1409 ( .A(n21500), .B(n42115), .Z(n928) );
  AND U1410 ( .A(n927), .B(n928), .Z(n21539) );
  NANDN U1411 ( .A(n21533), .B(n42047), .Z(n929) );
  NANDN U1412 ( .A(n21570), .B(n4067), .Z(n930) );
  NAND U1413 ( .A(n929), .B(n930), .Z(n21581) );
  NANDN U1414 ( .A(n21611), .B(n4068), .Z(n931) );
  NANDN U1415 ( .A(n21571), .B(n42115), .Z(n932) );
  AND U1416 ( .A(n931), .B(n932), .Z(n21613) );
  NANDN U1417 ( .A(n21607), .B(n42047), .Z(n933) );
  NANDN U1418 ( .A(n21644), .B(n4067), .Z(n934) );
  NAND U1419 ( .A(n933), .B(n934), .Z(n21655) );
  NANDN U1420 ( .A(n21685), .B(n4068), .Z(n935) );
  NANDN U1421 ( .A(n21645), .B(n42115), .Z(n936) );
  AND U1422 ( .A(n935), .B(n936), .Z(n21687) );
  NANDN U1423 ( .A(n21681), .B(n42047), .Z(n937) );
  NANDN U1424 ( .A(n21718), .B(n4067), .Z(n938) );
  NAND U1425 ( .A(n937), .B(n938), .Z(n21729) );
  NANDN U1426 ( .A(n21759), .B(n4068), .Z(n939) );
  NANDN U1427 ( .A(n21722), .B(n42115), .Z(n940) );
  AND U1428 ( .A(n939), .B(n940), .Z(n21761) );
  NANDN U1429 ( .A(n21755), .B(n42047), .Z(n941) );
  NANDN U1430 ( .A(n21792), .B(n4067), .Z(n942) );
  NAND U1431 ( .A(n941), .B(n942), .Z(n21803) );
  NANDN U1432 ( .A(n21833), .B(n4068), .Z(n943) );
  NANDN U1433 ( .A(n21793), .B(n42115), .Z(n944) );
  AND U1434 ( .A(n943), .B(n944), .Z(n21835) );
  NANDN U1435 ( .A(n21829), .B(n42047), .Z(n945) );
  NANDN U1436 ( .A(n21866), .B(n4067), .Z(n946) );
  NAND U1437 ( .A(n945), .B(n946), .Z(n21877) );
  NANDN U1438 ( .A(n21907), .B(n4068), .Z(n947) );
  NANDN U1439 ( .A(n21870), .B(n42115), .Z(n948) );
  AND U1440 ( .A(n947), .B(n948), .Z(n21909) );
  NANDN U1441 ( .A(n21903), .B(n42047), .Z(n949) );
  NANDN U1442 ( .A(n21940), .B(n4067), .Z(n950) );
  NAND U1443 ( .A(n949), .B(n950), .Z(n21951) );
  NANDN U1444 ( .A(n21981), .B(n4068), .Z(n951) );
  NANDN U1445 ( .A(n21941), .B(n42115), .Z(n952) );
  AND U1446 ( .A(n951), .B(n952), .Z(n21983) );
  NANDN U1447 ( .A(n21977), .B(n42047), .Z(n953) );
  NANDN U1448 ( .A(n22014), .B(n4067), .Z(n954) );
  NAND U1449 ( .A(n953), .B(n954), .Z(n22025) );
  NANDN U1450 ( .A(n22052), .B(n4068), .Z(n955) );
  NANDN U1451 ( .A(n22018), .B(n42115), .Z(n956) );
  AND U1452 ( .A(n955), .B(n956), .Z(n22057) );
  NANDN U1453 ( .A(n22051), .B(n42047), .Z(n957) );
  NANDN U1454 ( .A(n22088), .B(n4067), .Z(n958) );
  NAND U1455 ( .A(n957), .B(n958), .Z(n22099) );
  NANDN U1456 ( .A(n22126), .B(n4068), .Z(n959) );
  NANDN U1457 ( .A(n22092), .B(n42115), .Z(n960) );
  AND U1458 ( .A(n959), .B(n960), .Z(n22131) );
  NANDN U1459 ( .A(n22125), .B(n42047), .Z(n961) );
  NANDN U1460 ( .A(n22162), .B(n4067), .Z(n962) );
  NAND U1461 ( .A(n961), .B(n962), .Z(n22173) );
  NANDN U1462 ( .A(n22203), .B(n4068), .Z(n963) );
  NANDN U1463 ( .A(n22166), .B(n42115), .Z(n964) );
  AND U1464 ( .A(n963), .B(n964), .Z(n22205) );
  NANDN U1465 ( .A(n22199), .B(n42047), .Z(n965) );
  NANDN U1466 ( .A(n22236), .B(n4067), .Z(n966) );
  NAND U1467 ( .A(n965), .B(n966), .Z(n22247) );
  NANDN U1468 ( .A(n22277), .B(n4068), .Z(n967) );
  NANDN U1469 ( .A(n22237), .B(n42115), .Z(n968) );
  AND U1470 ( .A(n967), .B(n968), .Z(n22279) );
  NANDN U1471 ( .A(n22273), .B(n42047), .Z(n969) );
  NANDN U1472 ( .A(n22310), .B(n4067), .Z(n970) );
  NAND U1473 ( .A(n969), .B(n970), .Z(n22321) );
  NANDN U1474 ( .A(n22351), .B(n4068), .Z(n971) );
  NANDN U1475 ( .A(n22314), .B(n42115), .Z(n972) );
  AND U1476 ( .A(n971), .B(n972), .Z(n22353) );
  NANDN U1477 ( .A(n22347), .B(n42047), .Z(n973) );
  NANDN U1478 ( .A(n22384), .B(n4067), .Z(n974) );
  NAND U1479 ( .A(n973), .B(n974), .Z(n22395) );
  NANDN U1480 ( .A(n22425), .B(n4068), .Z(n975) );
  NANDN U1481 ( .A(n22388), .B(n42115), .Z(n976) );
  AND U1482 ( .A(n975), .B(n976), .Z(n22427) );
  NANDN U1483 ( .A(n22421), .B(n42047), .Z(n977) );
  NANDN U1484 ( .A(n22458), .B(n4067), .Z(n978) );
  NAND U1485 ( .A(n977), .B(n978), .Z(n22469) );
  NANDN U1486 ( .A(n22496), .B(n4068), .Z(n979) );
  NANDN U1487 ( .A(n22462), .B(n42115), .Z(n980) );
  AND U1488 ( .A(n979), .B(n980), .Z(n22501) );
  NANDN U1489 ( .A(n22495), .B(n42047), .Z(n981) );
  NANDN U1490 ( .A(n22532), .B(n4067), .Z(n982) );
  NAND U1491 ( .A(n981), .B(n982), .Z(n22543) );
  NANDN U1492 ( .A(n22573), .B(n4068), .Z(n983) );
  NANDN U1493 ( .A(n22536), .B(n42115), .Z(n984) );
  AND U1494 ( .A(n983), .B(n984), .Z(n22575) );
  NANDN U1495 ( .A(n22569), .B(n42047), .Z(n985) );
  NANDN U1496 ( .A(n22606), .B(n4067), .Z(n986) );
  NAND U1497 ( .A(n985), .B(n986), .Z(n22617) );
  NANDN U1498 ( .A(n22647), .B(n4068), .Z(n987) );
  NANDN U1499 ( .A(n22610), .B(n42115), .Z(n988) );
  AND U1500 ( .A(n987), .B(n988), .Z(n22649) );
  NANDN U1501 ( .A(n22643), .B(n42047), .Z(n989) );
  NANDN U1502 ( .A(n22680), .B(n4067), .Z(n990) );
  NAND U1503 ( .A(n989), .B(n990), .Z(n22691) );
  NANDN U1504 ( .A(n22718), .B(n4068), .Z(n991) );
  NANDN U1505 ( .A(n22684), .B(n42115), .Z(n992) );
  AND U1506 ( .A(n991), .B(n992), .Z(n22723) );
  NANDN U1507 ( .A(n22717), .B(n42047), .Z(n993) );
  NANDN U1508 ( .A(n22759), .B(n4067), .Z(n994) );
  NAND U1509 ( .A(n993), .B(n994), .Z(n22770) );
  NANDN U1510 ( .A(n22792), .B(n4068), .Z(n995) );
  NANDN U1511 ( .A(n22763), .B(n42115), .Z(n996) );
  AND U1512 ( .A(n995), .B(n996), .Z(n22797) );
  NANDN U1513 ( .A(n22791), .B(n42047), .Z(n997) );
  NANDN U1514 ( .A(n22828), .B(n4067), .Z(n998) );
  NAND U1515 ( .A(n997), .B(n998), .Z(n22839) );
  NANDN U1516 ( .A(n22869), .B(n4068), .Z(n999) );
  NANDN U1517 ( .A(n22829), .B(n42115), .Z(n1000) );
  AND U1518 ( .A(n999), .B(n1000), .Z(n22871) );
  NANDN U1519 ( .A(n22865), .B(n42047), .Z(n1001) );
  NANDN U1520 ( .A(n22902), .B(n4067), .Z(n1002) );
  NAND U1521 ( .A(n1001), .B(n1002), .Z(n22913) );
  NANDN U1522 ( .A(n22943), .B(n4068), .Z(n1003) );
  NANDN U1523 ( .A(n22903), .B(n42115), .Z(n1004) );
  AND U1524 ( .A(n1003), .B(n1004), .Z(n22945) );
  NANDN U1525 ( .A(n22939), .B(n42047), .Z(n1005) );
  NANDN U1526 ( .A(n22976), .B(n4067), .Z(n1006) );
  NAND U1527 ( .A(n1005), .B(n1006), .Z(n22987) );
  NANDN U1528 ( .A(n23017), .B(n4068), .Z(n1007) );
  NANDN U1529 ( .A(n22980), .B(n42115), .Z(n1008) );
  AND U1530 ( .A(n1007), .B(n1008), .Z(n23019) );
  NANDN U1531 ( .A(n23013), .B(n42047), .Z(n1009) );
  NANDN U1532 ( .A(n23050), .B(n4067), .Z(n1010) );
  NAND U1533 ( .A(n1009), .B(n1010), .Z(n23061) );
  NANDN U1534 ( .A(n23088), .B(n4068), .Z(n1011) );
  NANDN U1535 ( .A(n23054), .B(n42115), .Z(n1012) );
  AND U1536 ( .A(n1011), .B(n1012), .Z(n23093) );
  NANDN U1537 ( .A(n23087), .B(n42047), .Z(n1013) );
  NANDN U1538 ( .A(n23124), .B(n4067), .Z(n1014) );
  NAND U1539 ( .A(n1013), .B(n1014), .Z(n23135) );
  NANDN U1540 ( .A(n23165), .B(n4068), .Z(n1015) );
  NANDN U1541 ( .A(n23128), .B(n42115), .Z(n1016) );
  AND U1542 ( .A(n1015), .B(n1016), .Z(n23167) );
  NANDN U1543 ( .A(n23161), .B(n42047), .Z(n1017) );
  NANDN U1544 ( .A(n23198), .B(n4067), .Z(n1018) );
  NAND U1545 ( .A(n1017), .B(n1018), .Z(n23209) );
  NANDN U1546 ( .A(n23239), .B(n4068), .Z(n1019) );
  NANDN U1547 ( .A(n23199), .B(n42115), .Z(n1020) );
  AND U1548 ( .A(n1019), .B(n1020), .Z(n23241) );
  NANDN U1549 ( .A(n23235), .B(n42047), .Z(n1021) );
  NANDN U1550 ( .A(n23272), .B(n4067), .Z(n1022) );
  NAND U1551 ( .A(n1021), .B(n1022), .Z(n23283) );
  NANDN U1552 ( .A(n23313), .B(n4068), .Z(n1023) );
  NANDN U1553 ( .A(n23273), .B(n42115), .Z(n1024) );
  AND U1554 ( .A(n1023), .B(n1024), .Z(n23315) );
  NANDN U1555 ( .A(n23309), .B(n42047), .Z(n1025) );
  NANDN U1556 ( .A(n23346), .B(n4067), .Z(n1026) );
  NAND U1557 ( .A(n1025), .B(n1026), .Z(n23357) );
  NANDN U1558 ( .A(n23384), .B(n4068), .Z(n1027) );
  NANDN U1559 ( .A(n23350), .B(n42115), .Z(n1028) );
  AND U1560 ( .A(n1027), .B(n1028), .Z(n23389) );
  NANDN U1561 ( .A(n23383), .B(n42047), .Z(n1029) );
  NANDN U1562 ( .A(n23420), .B(n4067), .Z(n1030) );
  NAND U1563 ( .A(n1029), .B(n1030), .Z(n23431) );
  NANDN U1564 ( .A(n23458), .B(n4068), .Z(n1031) );
  NANDN U1565 ( .A(n23421), .B(n42115), .Z(n1032) );
  AND U1566 ( .A(n1031), .B(n1032), .Z(n23463) );
  NANDN U1567 ( .A(n23457), .B(n42047), .Z(n1033) );
  NANDN U1568 ( .A(n23494), .B(n4067), .Z(n1034) );
  NAND U1569 ( .A(n1033), .B(n1034), .Z(n23505) );
  NANDN U1570 ( .A(n23535), .B(n4068), .Z(n1035) );
  NANDN U1571 ( .A(n23498), .B(n42115), .Z(n1036) );
  AND U1572 ( .A(n1035), .B(n1036), .Z(n23537) );
  NANDN U1573 ( .A(n23531), .B(n42047), .Z(n1037) );
  NANDN U1574 ( .A(n23568), .B(n4067), .Z(n1038) );
  NAND U1575 ( .A(n1037), .B(n1038), .Z(n23579) );
  NANDN U1576 ( .A(n23606), .B(n4068), .Z(n1039) );
  NANDN U1577 ( .A(n23572), .B(n42115), .Z(n1040) );
  AND U1578 ( .A(n1039), .B(n1040), .Z(n23611) );
  NANDN U1579 ( .A(n23605), .B(n42047), .Z(n1041) );
  NANDN U1580 ( .A(n23642), .B(n4067), .Z(n1042) );
  NAND U1581 ( .A(n1041), .B(n1042), .Z(n23653) );
  NANDN U1582 ( .A(n23683), .B(n4068), .Z(n1043) );
  NANDN U1583 ( .A(n23646), .B(n42115), .Z(n1044) );
  AND U1584 ( .A(n1043), .B(n1044), .Z(n23685) );
  NANDN U1585 ( .A(n23679), .B(n42047), .Z(n1045) );
  NANDN U1586 ( .A(n23716), .B(n4067), .Z(n1046) );
  NAND U1587 ( .A(n1045), .B(n1046), .Z(n23727) );
  NANDN U1588 ( .A(n23757), .B(n4068), .Z(n1047) );
  NANDN U1589 ( .A(n23717), .B(n42115), .Z(n1048) );
  AND U1590 ( .A(n1047), .B(n1048), .Z(n23759) );
  NANDN U1591 ( .A(n23753), .B(n42047), .Z(n1049) );
  NANDN U1592 ( .A(n23790), .B(n4067), .Z(n1050) );
  NAND U1593 ( .A(n1049), .B(n1050), .Z(n23801) );
  NANDN U1594 ( .A(n23828), .B(n4068), .Z(n1051) );
  NANDN U1595 ( .A(n23794), .B(n42115), .Z(n1052) );
  AND U1596 ( .A(n1051), .B(n1052), .Z(n23833) );
  NANDN U1597 ( .A(n23827), .B(n42047), .Z(n1053) );
  NANDN U1598 ( .A(n23864), .B(n4067), .Z(n1054) );
  NAND U1599 ( .A(n1053), .B(n1054), .Z(n23875) );
  NANDN U1600 ( .A(n23905), .B(n4068), .Z(n1055) );
  NANDN U1601 ( .A(n23868), .B(n42115), .Z(n1056) );
  AND U1602 ( .A(n1055), .B(n1056), .Z(n23907) );
  NANDN U1603 ( .A(n23901), .B(n42047), .Z(n1057) );
  NANDN U1604 ( .A(n23938), .B(n4067), .Z(n1058) );
  NAND U1605 ( .A(n1057), .B(n1058), .Z(n23949) );
  NANDN U1606 ( .A(n23979), .B(n4068), .Z(n1059) );
  NANDN U1607 ( .A(n23939), .B(n42115), .Z(n1060) );
  AND U1608 ( .A(n1059), .B(n1060), .Z(n23981) );
  NANDN U1609 ( .A(n23975), .B(n42047), .Z(n1061) );
  NANDN U1610 ( .A(n24012), .B(n4067), .Z(n1062) );
  NAND U1611 ( .A(n1061), .B(n1062), .Z(n24023) );
  NANDN U1612 ( .A(n24053), .B(n4068), .Z(n1063) );
  NANDN U1613 ( .A(n24016), .B(n42115), .Z(n1064) );
  AND U1614 ( .A(n1063), .B(n1064), .Z(n24055) );
  NANDN U1615 ( .A(n24049), .B(n42047), .Z(n1065) );
  NANDN U1616 ( .A(n24086), .B(n4067), .Z(n1066) );
  NAND U1617 ( .A(n1065), .B(n1066), .Z(n24097) );
  NANDN U1618 ( .A(n24124), .B(n4068), .Z(n1067) );
  NANDN U1619 ( .A(n24087), .B(n42115), .Z(n1068) );
  AND U1620 ( .A(n1067), .B(n1068), .Z(n24129) );
  NANDN U1621 ( .A(n24123), .B(n42047), .Z(n1069) );
  NANDN U1622 ( .A(n24160), .B(n4067), .Z(n1070) );
  NAND U1623 ( .A(n1069), .B(n1070), .Z(n24171) );
  NANDN U1624 ( .A(n24201), .B(n4068), .Z(n1071) );
  NANDN U1625 ( .A(n24164), .B(n42115), .Z(n1072) );
  AND U1626 ( .A(n1071), .B(n1072), .Z(n24203) );
  NANDN U1627 ( .A(n24197), .B(n42047), .Z(n1073) );
  NANDN U1628 ( .A(n24234), .B(n4067), .Z(n1074) );
  NAND U1629 ( .A(n1073), .B(n1074), .Z(n24245) );
  NANDN U1630 ( .A(n24275), .B(n4068), .Z(n1075) );
  NANDN U1631 ( .A(n24238), .B(n42115), .Z(n1076) );
  AND U1632 ( .A(n1075), .B(n1076), .Z(n24277) );
  NANDN U1633 ( .A(n24271), .B(n42047), .Z(n1077) );
  NANDN U1634 ( .A(n24308), .B(n4067), .Z(n1078) );
  NAND U1635 ( .A(n1077), .B(n1078), .Z(n24319) );
  NANDN U1636 ( .A(n24349), .B(n4068), .Z(n1079) );
  NANDN U1637 ( .A(n24312), .B(n42115), .Z(n1080) );
  AND U1638 ( .A(n1079), .B(n1080), .Z(n24351) );
  NANDN U1639 ( .A(n24345), .B(n42047), .Z(n1081) );
  NANDN U1640 ( .A(n24382), .B(n4067), .Z(n1082) );
  NAND U1641 ( .A(n1081), .B(n1082), .Z(n24393) );
  NANDN U1642 ( .A(n24423), .B(n4068), .Z(n1083) );
  NANDN U1643 ( .A(n24386), .B(n42115), .Z(n1084) );
  AND U1644 ( .A(n1083), .B(n1084), .Z(n24425) );
  NANDN U1645 ( .A(n24419), .B(n42047), .Z(n1085) );
  NANDN U1646 ( .A(n24456), .B(n4067), .Z(n1086) );
  NAND U1647 ( .A(n1085), .B(n1086), .Z(n24467) );
  NANDN U1648 ( .A(n24497), .B(n4068), .Z(n1087) );
  NANDN U1649 ( .A(n24460), .B(n42115), .Z(n1088) );
  AND U1650 ( .A(n1087), .B(n1088), .Z(n24499) );
  NANDN U1651 ( .A(n24493), .B(n42047), .Z(n1089) );
  NANDN U1652 ( .A(n24530), .B(n4067), .Z(n1090) );
  NAND U1653 ( .A(n1089), .B(n1090), .Z(n24541) );
  NANDN U1654 ( .A(n24571), .B(n4068), .Z(n1091) );
  NANDN U1655 ( .A(n24531), .B(n42115), .Z(n1092) );
  AND U1656 ( .A(n1091), .B(n1092), .Z(n24573) );
  NANDN U1657 ( .A(n24567), .B(n42047), .Z(n1093) );
  NANDN U1658 ( .A(n24604), .B(n4067), .Z(n1094) );
  NAND U1659 ( .A(n1093), .B(n1094), .Z(n24615) );
  NANDN U1660 ( .A(n24645), .B(n4068), .Z(n1095) );
  NANDN U1661 ( .A(n24605), .B(n42115), .Z(n1096) );
  AND U1662 ( .A(n1095), .B(n1096), .Z(n24647) );
  NANDN U1663 ( .A(n24641), .B(n42047), .Z(n1097) );
  NANDN U1664 ( .A(n24678), .B(n4067), .Z(n1098) );
  NAND U1665 ( .A(n1097), .B(n1098), .Z(n24689) );
  NANDN U1666 ( .A(n24716), .B(n4068), .Z(n1099) );
  NANDN U1667 ( .A(n24682), .B(n42115), .Z(n1100) );
  AND U1668 ( .A(n1099), .B(n1100), .Z(n24721) );
  NANDN U1669 ( .A(n24715), .B(n42047), .Z(n1101) );
  NANDN U1670 ( .A(n24752), .B(n4067), .Z(n1102) );
  NAND U1671 ( .A(n1101), .B(n1102), .Z(n24763) );
  NANDN U1672 ( .A(n24790), .B(n4068), .Z(n1103) );
  NANDN U1673 ( .A(n24756), .B(n42115), .Z(n1104) );
  AND U1674 ( .A(n1103), .B(n1104), .Z(n24795) );
  NANDN U1675 ( .A(n24789), .B(n42047), .Z(n1105) );
  NANDN U1676 ( .A(n24826), .B(n4067), .Z(n1106) );
  NAND U1677 ( .A(n1105), .B(n1106), .Z(n24837) );
  NANDN U1678 ( .A(n24867), .B(n4068), .Z(n1107) );
  NANDN U1679 ( .A(n24830), .B(n42115), .Z(n1108) );
  AND U1680 ( .A(n1107), .B(n1108), .Z(n24869) );
  NANDN U1681 ( .A(n24863), .B(n42047), .Z(n1109) );
  NANDN U1682 ( .A(n24900), .B(n4067), .Z(n1110) );
  NAND U1683 ( .A(n1109), .B(n1110), .Z(n24911) );
  NANDN U1684 ( .A(n24941), .B(n4068), .Z(n1111) );
  NANDN U1685 ( .A(n24901), .B(n42115), .Z(n1112) );
  AND U1686 ( .A(n1111), .B(n1112), .Z(n24943) );
  NANDN U1687 ( .A(n24937), .B(n42047), .Z(n1113) );
  NANDN U1688 ( .A(n24974), .B(n4067), .Z(n1114) );
  NAND U1689 ( .A(n1113), .B(n1114), .Z(n24985) );
  NANDN U1690 ( .A(n25015), .B(n4068), .Z(n1115) );
  NANDN U1691 ( .A(n24978), .B(n42115), .Z(n1116) );
  AND U1692 ( .A(n1115), .B(n1116), .Z(n25017) );
  NANDN U1693 ( .A(n25011), .B(n42047), .Z(n1117) );
  NANDN U1694 ( .A(n25048), .B(n4067), .Z(n1118) );
  NAND U1695 ( .A(n1117), .B(n1118), .Z(n25059) );
  NANDN U1696 ( .A(n25089), .B(n4068), .Z(n1119) );
  NANDN U1697 ( .A(n25052), .B(n42115), .Z(n1120) );
  AND U1698 ( .A(n1119), .B(n1120), .Z(n25091) );
  NANDN U1699 ( .A(n25085), .B(n42047), .Z(n1121) );
  NANDN U1700 ( .A(n25122), .B(n4067), .Z(n1122) );
  NAND U1701 ( .A(n1121), .B(n1122), .Z(n25133) );
  NANDN U1702 ( .A(n25163), .B(n4068), .Z(n1123) );
  NANDN U1703 ( .A(n25126), .B(n42115), .Z(n1124) );
  AND U1704 ( .A(n1123), .B(n1124), .Z(n25165) );
  NANDN U1705 ( .A(n25159), .B(n42047), .Z(n1125) );
  NANDN U1706 ( .A(n25196), .B(n4067), .Z(n1126) );
  NAND U1707 ( .A(n1125), .B(n1126), .Z(n25207) );
  NANDN U1708 ( .A(n25234), .B(n4068), .Z(n1127) );
  NANDN U1709 ( .A(n25200), .B(n42115), .Z(n1128) );
  AND U1710 ( .A(n1127), .B(n1128), .Z(n25239) );
  NANDN U1711 ( .A(n25233), .B(n42047), .Z(n1129) );
  NANDN U1712 ( .A(n25270), .B(n4067), .Z(n1130) );
  NAND U1713 ( .A(n1129), .B(n1130), .Z(n25281) );
  NANDN U1714 ( .A(n25311), .B(n4068), .Z(n1131) );
  NANDN U1715 ( .A(n25271), .B(n42115), .Z(n1132) );
  AND U1716 ( .A(n1131), .B(n1132), .Z(n25313) );
  NANDN U1717 ( .A(n25307), .B(n42047), .Z(n1133) );
  NANDN U1718 ( .A(n25344), .B(n4067), .Z(n1134) );
  NAND U1719 ( .A(n1133), .B(n1134), .Z(n25355) );
  NANDN U1720 ( .A(n25382), .B(n4068), .Z(n1135) );
  NANDN U1721 ( .A(n25348), .B(n42115), .Z(n1136) );
  AND U1722 ( .A(n1135), .B(n1136), .Z(n25387) );
  NANDN U1723 ( .A(n25381), .B(n42047), .Z(n1137) );
  NANDN U1724 ( .A(n25418), .B(n4067), .Z(n1138) );
  NAND U1725 ( .A(n1137), .B(n1138), .Z(n25429) );
  NANDN U1726 ( .A(n25459), .B(n4068), .Z(n1139) );
  NANDN U1727 ( .A(n25422), .B(n42115), .Z(n1140) );
  AND U1728 ( .A(n1139), .B(n1140), .Z(n25461) );
  NANDN U1729 ( .A(n25455), .B(n42047), .Z(n1141) );
  NANDN U1730 ( .A(n25492), .B(n4067), .Z(n1142) );
  NAND U1731 ( .A(n1141), .B(n1142), .Z(n25503) );
  NANDN U1732 ( .A(n25530), .B(n4068), .Z(n1143) );
  NANDN U1733 ( .A(n25493), .B(n42115), .Z(n1144) );
  AND U1734 ( .A(n1143), .B(n1144), .Z(n25535) );
  NANDN U1735 ( .A(n25529), .B(n42047), .Z(n1145) );
  NANDN U1736 ( .A(n25566), .B(n4067), .Z(n1146) );
  NAND U1737 ( .A(n1145), .B(n1146), .Z(n25577) );
  NANDN U1738 ( .A(n25604), .B(n4068), .Z(n1147) );
  NANDN U1739 ( .A(n25567), .B(n42115), .Z(n1148) );
  AND U1740 ( .A(n1147), .B(n1148), .Z(n25609) );
  NANDN U1741 ( .A(n25603), .B(n42047), .Z(n1149) );
  NANDN U1742 ( .A(n25640), .B(n4067), .Z(n1150) );
  NAND U1743 ( .A(n1149), .B(n1150), .Z(n25651) );
  NANDN U1744 ( .A(n25681), .B(n4068), .Z(n1151) );
  NANDN U1745 ( .A(n25644), .B(n42115), .Z(n1152) );
  AND U1746 ( .A(n1151), .B(n1152), .Z(n25683) );
  NANDN U1747 ( .A(n25677), .B(n42047), .Z(n1153) );
  NANDN U1748 ( .A(n25714), .B(n4067), .Z(n1154) );
  NAND U1749 ( .A(n1153), .B(n1154), .Z(n25725) );
  NANDN U1750 ( .A(n25755), .B(n4068), .Z(n1155) );
  NANDN U1751 ( .A(n25718), .B(n42115), .Z(n1156) );
  AND U1752 ( .A(n1155), .B(n1156), .Z(n25757) );
  NANDN U1753 ( .A(n25751), .B(n42047), .Z(n1157) );
  NANDN U1754 ( .A(n25788), .B(n4067), .Z(n1158) );
  NAND U1755 ( .A(n1157), .B(n1158), .Z(n25799) );
  NANDN U1756 ( .A(n25829), .B(n4068), .Z(n1159) );
  NANDN U1757 ( .A(n25789), .B(n42115), .Z(n1160) );
  AND U1758 ( .A(n1159), .B(n1160), .Z(n25831) );
  NANDN U1759 ( .A(n25825), .B(n42047), .Z(n1161) );
  NANDN U1760 ( .A(n25862), .B(n4067), .Z(n1162) );
  NAND U1761 ( .A(n1161), .B(n1162), .Z(n25873) );
  NANDN U1762 ( .A(n25900), .B(n4068), .Z(n1163) );
  NANDN U1763 ( .A(n25866), .B(n42115), .Z(n1164) );
  AND U1764 ( .A(n1163), .B(n1164), .Z(n25905) );
  NANDN U1765 ( .A(n25899), .B(n42047), .Z(n1165) );
  NANDN U1766 ( .A(n25936), .B(n4067), .Z(n1166) );
  NAND U1767 ( .A(n1165), .B(n1166), .Z(n25947) );
  NANDN U1768 ( .A(n25974), .B(n4068), .Z(n1167) );
  NANDN U1769 ( .A(n25940), .B(n42115), .Z(n1168) );
  AND U1770 ( .A(n1167), .B(n1168), .Z(n25979) );
  NANDN U1771 ( .A(n25973), .B(n42047), .Z(n1169) );
  NANDN U1772 ( .A(n26010), .B(n4067), .Z(n1170) );
  NAND U1773 ( .A(n1169), .B(n1170), .Z(n26021) );
  NANDN U1774 ( .A(n26051), .B(n4068), .Z(n1171) );
  NANDN U1775 ( .A(n26014), .B(n42115), .Z(n1172) );
  AND U1776 ( .A(n1171), .B(n1172), .Z(n26053) );
  NANDN U1777 ( .A(n26047), .B(n42047), .Z(n1173) );
  NANDN U1778 ( .A(n26084), .B(n4067), .Z(n1174) );
  NAND U1779 ( .A(n1173), .B(n1174), .Z(n26095) );
  NANDN U1780 ( .A(n26125), .B(n4068), .Z(n1175) );
  NANDN U1781 ( .A(n26088), .B(n42115), .Z(n1176) );
  AND U1782 ( .A(n1175), .B(n1176), .Z(n26127) );
  NANDN U1783 ( .A(n26121), .B(n42047), .Z(n1177) );
  NANDN U1784 ( .A(n26158), .B(n4067), .Z(n1178) );
  NAND U1785 ( .A(n1177), .B(n1178), .Z(n26169) );
  NANDN U1786 ( .A(n26199), .B(n4068), .Z(n1179) );
  NANDN U1787 ( .A(n26159), .B(n42115), .Z(n1180) );
  AND U1788 ( .A(n1179), .B(n1180), .Z(n26201) );
  NANDN U1789 ( .A(n26195), .B(n42047), .Z(n1181) );
  NANDN U1790 ( .A(n26232), .B(n4067), .Z(n1182) );
  NAND U1791 ( .A(n1181), .B(n1182), .Z(n26243) );
  NANDN U1792 ( .A(n26273), .B(n4068), .Z(n1183) );
  NANDN U1793 ( .A(n26233), .B(n42115), .Z(n1184) );
  AND U1794 ( .A(n1183), .B(n1184), .Z(n26275) );
  NANDN U1795 ( .A(n26269), .B(n42047), .Z(n1185) );
  NANDN U1796 ( .A(n26306), .B(n4067), .Z(n1186) );
  NAND U1797 ( .A(n1185), .B(n1186), .Z(n26317) );
  NANDN U1798 ( .A(n26347), .B(n4068), .Z(n1187) );
  NANDN U1799 ( .A(n26310), .B(n42115), .Z(n1188) );
  AND U1800 ( .A(n1187), .B(n1188), .Z(n26349) );
  NANDN U1801 ( .A(n26343), .B(n42047), .Z(n1189) );
  NANDN U1802 ( .A(n26380), .B(n4067), .Z(n1190) );
  NAND U1803 ( .A(n1189), .B(n1190), .Z(n26391) );
  NANDN U1804 ( .A(n26421), .B(n4068), .Z(n1191) );
  NANDN U1805 ( .A(n26381), .B(n42115), .Z(n1192) );
  AND U1806 ( .A(n1191), .B(n1192), .Z(n26423) );
  NANDN U1807 ( .A(n26417), .B(n42047), .Z(n1193) );
  NANDN U1808 ( .A(n26454), .B(n4067), .Z(n1194) );
  NAND U1809 ( .A(n1193), .B(n1194), .Z(n26465) );
  NANDN U1810 ( .A(n26495), .B(n4068), .Z(n1195) );
  NANDN U1811 ( .A(n26455), .B(n42115), .Z(n1196) );
  AND U1812 ( .A(n1195), .B(n1196), .Z(n26497) );
  NANDN U1813 ( .A(n26491), .B(n42047), .Z(n1197) );
  NANDN U1814 ( .A(n26528), .B(n4067), .Z(n1198) );
  NAND U1815 ( .A(n1197), .B(n1198), .Z(n26539) );
  NANDN U1816 ( .A(n26569), .B(n4068), .Z(n1199) );
  NANDN U1817 ( .A(n26532), .B(n42115), .Z(n1200) );
  AND U1818 ( .A(n1199), .B(n1200), .Z(n26571) );
  NANDN U1819 ( .A(n26565), .B(n42047), .Z(n1201) );
  NANDN U1820 ( .A(n26602), .B(n4067), .Z(n1202) );
  NAND U1821 ( .A(n1201), .B(n1202), .Z(n26613) );
  NANDN U1822 ( .A(n26640), .B(n4068), .Z(n1203) );
  NANDN U1823 ( .A(n26603), .B(n42115), .Z(n1204) );
  AND U1824 ( .A(n1203), .B(n1204), .Z(n26645) );
  NANDN U1825 ( .A(n26639), .B(n42047), .Z(n1205) );
  NANDN U1826 ( .A(n26676), .B(n4067), .Z(n1206) );
  NAND U1827 ( .A(n1205), .B(n1206), .Z(n26687) );
  NANDN U1828 ( .A(n26717), .B(n4068), .Z(n1207) );
  NANDN U1829 ( .A(n26680), .B(n42115), .Z(n1208) );
  AND U1830 ( .A(n1207), .B(n1208), .Z(n26719) );
  NANDN U1831 ( .A(n26713), .B(n42047), .Z(n1209) );
  NANDN U1832 ( .A(n26750), .B(n4067), .Z(n1210) );
  NAND U1833 ( .A(n1209), .B(n1210), .Z(n26761) );
  NANDN U1834 ( .A(n26788), .B(n4068), .Z(n1211) );
  NANDN U1835 ( .A(n26751), .B(n42115), .Z(n1212) );
  AND U1836 ( .A(n1211), .B(n1212), .Z(n26793) );
  NANDN U1837 ( .A(n26787), .B(n42047), .Z(n1213) );
  NANDN U1838 ( .A(n26824), .B(n4067), .Z(n1214) );
  NAND U1839 ( .A(n1213), .B(n1214), .Z(n26835) );
  NANDN U1840 ( .A(n26865), .B(n4068), .Z(n1215) );
  NANDN U1841 ( .A(n26828), .B(n42115), .Z(n1216) );
  AND U1842 ( .A(n1215), .B(n1216), .Z(n26867) );
  NANDN U1843 ( .A(n26861), .B(n42047), .Z(n1217) );
  NANDN U1844 ( .A(n26898), .B(n4067), .Z(n1218) );
  NAND U1845 ( .A(n1217), .B(n1218), .Z(n26909) );
  NANDN U1846 ( .A(n26939), .B(n4068), .Z(n1219) );
  NANDN U1847 ( .A(n26902), .B(n42115), .Z(n1220) );
  AND U1848 ( .A(n1219), .B(n1220), .Z(n26941) );
  NANDN U1849 ( .A(n26935), .B(n42047), .Z(n1221) );
  NANDN U1850 ( .A(n26972), .B(n4067), .Z(n1222) );
  NAND U1851 ( .A(n1221), .B(n1222), .Z(n26983) );
  NANDN U1852 ( .A(n27010), .B(n4068), .Z(n1223) );
  NANDN U1853 ( .A(n26976), .B(n42115), .Z(n1224) );
  AND U1854 ( .A(n1223), .B(n1224), .Z(n27015) );
  NANDN U1855 ( .A(n27009), .B(n42047), .Z(n1225) );
  NANDN U1856 ( .A(n27046), .B(n4067), .Z(n1226) );
  NAND U1857 ( .A(n1225), .B(n1226), .Z(n27057) );
  NANDN U1858 ( .A(n27084), .B(n4068), .Z(n1227) );
  NANDN U1859 ( .A(n27050), .B(n42115), .Z(n1228) );
  AND U1860 ( .A(n1227), .B(n1228), .Z(n27089) );
  NANDN U1861 ( .A(n27083), .B(n42047), .Z(n1229) );
  NANDN U1862 ( .A(n27120), .B(n4067), .Z(n1230) );
  NAND U1863 ( .A(n1229), .B(n1230), .Z(n27131) );
  NANDN U1864 ( .A(n27158), .B(n4068), .Z(n1231) );
  NANDN U1865 ( .A(n27124), .B(n42115), .Z(n1232) );
  AND U1866 ( .A(n1231), .B(n1232), .Z(n27163) );
  NANDN U1867 ( .A(n27157), .B(n42047), .Z(n1233) );
  NANDN U1868 ( .A(n27194), .B(n4067), .Z(n1234) );
  NAND U1869 ( .A(n1233), .B(n1234), .Z(n27205) );
  NANDN U1870 ( .A(n27235), .B(n4068), .Z(n1235) );
  NANDN U1871 ( .A(n27198), .B(n42115), .Z(n1236) );
  AND U1872 ( .A(n1235), .B(n1236), .Z(n27237) );
  NANDN U1873 ( .A(n27231), .B(n42047), .Z(n1237) );
  NANDN U1874 ( .A(n27268), .B(n4067), .Z(n1238) );
  NAND U1875 ( .A(n1237), .B(n1238), .Z(n27279) );
  NANDN U1876 ( .A(n27306), .B(n4068), .Z(n1239) );
  NANDN U1877 ( .A(n27272), .B(n42115), .Z(n1240) );
  AND U1878 ( .A(n1239), .B(n1240), .Z(n27311) );
  NANDN U1879 ( .A(n27305), .B(n42047), .Z(n1241) );
  NANDN U1880 ( .A(n27342), .B(n4067), .Z(n1242) );
  NAND U1881 ( .A(n1241), .B(n1242), .Z(n27353) );
  NANDN U1882 ( .A(n27383), .B(n4068), .Z(n1243) );
  NANDN U1883 ( .A(n27346), .B(n42115), .Z(n1244) );
  AND U1884 ( .A(n1243), .B(n1244), .Z(n27385) );
  NANDN U1885 ( .A(n27379), .B(n42047), .Z(n1245) );
  NANDN U1886 ( .A(n27416), .B(n4067), .Z(n1246) );
  NAND U1887 ( .A(n1245), .B(n1246), .Z(n27427) );
  NANDN U1888 ( .A(n27457), .B(n4068), .Z(n1247) );
  NANDN U1889 ( .A(n27420), .B(n42115), .Z(n1248) );
  AND U1890 ( .A(n1247), .B(n1248), .Z(n27459) );
  NANDN U1891 ( .A(n27453), .B(n42047), .Z(n1249) );
  NANDN U1892 ( .A(n27490), .B(n4067), .Z(n1250) );
  NAND U1893 ( .A(n1249), .B(n1250), .Z(n27501) );
  NANDN U1894 ( .A(n27531), .B(n4068), .Z(n1251) );
  NANDN U1895 ( .A(n27494), .B(n42115), .Z(n1252) );
  AND U1896 ( .A(n1251), .B(n1252), .Z(n27533) );
  NANDN U1897 ( .A(n27527), .B(n42047), .Z(n1253) );
  NANDN U1898 ( .A(n27564), .B(n4067), .Z(n1254) );
  NAND U1899 ( .A(n1253), .B(n1254), .Z(n27575) );
  NANDN U1900 ( .A(n27605), .B(n4068), .Z(n1255) );
  NANDN U1901 ( .A(n27568), .B(n42115), .Z(n1256) );
  AND U1902 ( .A(n1255), .B(n1256), .Z(n27607) );
  NANDN U1903 ( .A(n27601), .B(n42047), .Z(n1257) );
  NANDN U1904 ( .A(n27638), .B(n4067), .Z(n1258) );
  NAND U1905 ( .A(n1257), .B(n1258), .Z(n27649) );
  NANDN U1906 ( .A(n27676), .B(n4068), .Z(n1259) );
  NANDN U1907 ( .A(n27642), .B(n42115), .Z(n1260) );
  AND U1908 ( .A(n1259), .B(n1260), .Z(n27681) );
  NANDN U1909 ( .A(n27675), .B(n42047), .Z(n1261) );
  NANDN U1910 ( .A(n27712), .B(n4067), .Z(n1262) );
  NAND U1911 ( .A(n1261), .B(n1262), .Z(n27723) );
  NANDN U1912 ( .A(n27750), .B(n4068), .Z(n1263) );
  NANDN U1913 ( .A(n27716), .B(n42115), .Z(n1264) );
  AND U1914 ( .A(n1263), .B(n1264), .Z(n27755) );
  NANDN U1915 ( .A(n27749), .B(n42047), .Z(n1265) );
  NANDN U1916 ( .A(n27786), .B(n4067), .Z(n1266) );
  NAND U1917 ( .A(n1265), .B(n1266), .Z(n27797) );
  NANDN U1918 ( .A(n27827), .B(n4068), .Z(n1267) );
  NANDN U1919 ( .A(n27790), .B(n42115), .Z(n1268) );
  AND U1920 ( .A(n1267), .B(n1268), .Z(n27829) );
  NANDN U1921 ( .A(n27823), .B(n42047), .Z(n1269) );
  NANDN U1922 ( .A(n27860), .B(n4067), .Z(n1270) );
  NAND U1923 ( .A(n1269), .B(n1270), .Z(n27871) );
  NANDN U1924 ( .A(n27898), .B(n4068), .Z(n1271) );
  NANDN U1925 ( .A(n27864), .B(n42115), .Z(n1272) );
  AND U1926 ( .A(n1271), .B(n1272), .Z(n27903) );
  NANDN U1927 ( .A(n27897), .B(n42047), .Z(n1273) );
  NANDN U1928 ( .A(n27934), .B(n4067), .Z(n1274) );
  NAND U1929 ( .A(n1273), .B(n1274), .Z(n27945) );
  NANDN U1930 ( .A(n27972), .B(n4068), .Z(n1275) );
  NANDN U1931 ( .A(n27935), .B(n42115), .Z(n1276) );
  AND U1932 ( .A(n1275), .B(n1276), .Z(n27977) );
  NANDN U1933 ( .A(n27971), .B(n42047), .Z(n1277) );
  NANDN U1934 ( .A(n28008), .B(n4067), .Z(n1278) );
  NAND U1935 ( .A(n1277), .B(n1278), .Z(n28019) );
  NANDN U1936 ( .A(n28046), .B(n4068), .Z(n1279) );
  NANDN U1937 ( .A(n28012), .B(n42115), .Z(n1280) );
  AND U1938 ( .A(n1279), .B(n1280), .Z(n28051) );
  NANDN U1939 ( .A(n28045), .B(n42047), .Z(n1281) );
  NANDN U1940 ( .A(n28082), .B(n4067), .Z(n1282) );
  NAND U1941 ( .A(n1281), .B(n1282), .Z(n28093) );
  NANDN U1942 ( .A(n28123), .B(n4068), .Z(n1283) );
  NANDN U1943 ( .A(n28086), .B(n42115), .Z(n1284) );
  AND U1944 ( .A(n1283), .B(n1284), .Z(n28125) );
  NANDN U1945 ( .A(n28119), .B(n42047), .Z(n1285) );
  NANDN U1946 ( .A(n28156), .B(n4067), .Z(n1286) );
  NAND U1947 ( .A(n1285), .B(n1286), .Z(n28167) );
  NANDN U1948 ( .A(n28197), .B(n4068), .Z(n1287) );
  NANDN U1949 ( .A(n28160), .B(n42115), .Z(n1288) );
  AND U1950 ( .A(n1287), .B(n1288), .Z(n28199) );
  NANDN U1951 ( .A(n28193), .B(n42047), .Z(n1289) );
  NANDN U1952 ( .A(n28230), .B(n4067), .Z(n1290) );
  NAND U1953 ( .A(n1289), .B(n1290), .Z(n28241) );
  NANDN U1954 ( .A(n28271), .B(n4068), .Z(n1291) );
  NANDN U1955 ( .A(n28234), .B(n42115), .Z(n1292) );
  AND U1956 ( .A(n1291), .B(n1292), .Z(n28273) );
  NANDN U1957 ( .A(n28267), .B(n42047), .Z(n1293) );
  NANDN U1958 ( .A(n28304), .B(n4067), .Z(n1294) );
  NAND U1959 ( .A(n1293), .B(n1294), .Z(n28315) );
  NANDN U1960 ( .A(n28345), .B(n4068), .Z(n1295) );
  NANDN U1961 ( .A(n28308), .B(n42115), .Z(n1296) );
  AND U1962 ( .A(n1295), .B(n1296), .Z(n28347) );
  NANDN U1963 ( .A(n28341), .B(n42047), .Z(n1297) );
  NANDN U1964 ( .A(n28378), .B(n4067), .Z(n1298) );
  NAND U1965 ( .A(n1297), .B(n1298), .Z(n28389) );
  NANDN U1966 ( .A(n28416), .B(n4068), .Z(n1299) );
  NANDN U1967 ( .A(n28382), .B(n42115), .Z(n1300) );
  AND U1968 ( .A(n1299), .B(n1300), .Z(n28421) );
  NANDN U1969 ( .A(n28415), .B(n42047), .Z(n1301) );
  NANDN U1970 ( .A(n28452), .B(n4067), .Z(n1302) );
  NAND U1971 ( .A(n1301), .B(n1302), .Z(n28463) );
  NANDN U1972 ( .A(n28493), .B(n4068), .Z(n1303) );
  NANDN U1973 ( .A(n28453), .B(n42115), .Z(n1304) );
  AND U1974 ( .A(n1303), .B(n1304), .Z(n28495) );
  NANDN U1975 ( .A(n28489), .B(n42047), .Z(n1305) );
  NANDN U1976 ( .A(n28526), .B(n4067), .Z(n1306) );
  NAND U1977 ( .A(n1305), .B(n1306), .Z(n28537) );
  NANDN U1978 ( .A(n28564), .B(n4068), .Z(n1307) );
  NANDN U1979 ( .A(n28530), .B(n42115), .Z(n1308) );
  AND U1980 ( .A(n1307), .B(n1308), .Z(n28569) );
  NANDN U1981 ( .A(n28563), .B(n42047), .Z(n1309) );
  NANDN U1982 ( .A(n28600), .B(n4067), .Z(n1310) );
  NAND U1983 ( .A(n1309), .B(n1310), .Z(n28611) );
  NANDN U1984 ( .A(n28641), .B(n4068), .Z(n1311) );
  NANDN U1985 ( .A(n28604), .B(n42115), .Z(n1312) );
  AND U1986 ( .A(n1311), .B(n1312), .Z(n28643) );
  NANDN U1987 ( .A(n28637), .B(n42047), .Z(n1313) );
  NANDN U1988 ( .A(n28674), .B(n4067), .Z(n1314) );
  NAND U1989 ( .A(n1313), .B(n1314), .Z(n28685) );
  NANDN U1990 ( .A(n28715), .B(n4068), .Z(n1315) );
  NANDN U1991 ( .A(n28678), .B(n42115), .Z(n1316) );
  AND U1992 ( .A(n1315), .B(n1316), .Z(n28717) );
  NANDN U1993 ( .A(n28711), .B(n42047), .Z(n1317) );
  NANDN U1994 ( .A(n28748), .B(n4067), .Z(n1318) );
  NAND U1995 ( .A(n1317), .B(n1318), .Z(n28759) );
  NANDN U1996 ( .A(n28789), .B(n4068), .Z(n1319) );
  NANDN U1997 ( .A(n28752), .B(n42115), .Z(n1320) );
  AND U1998 ( .A(n1319), .B(n1320), .Z(n28791) );
  NANDN U1999 ( .A(n28785), .B(n42047), .Z(n1321) );
  NANDN U2000 ( .A(n28822), .B(n4067), .Z(n1322) );
  NAND U2001 ( .A(n1321), .B(n1322), .Z(n28833) );
  NANDN U2002 ( .A(n28860), .B(n4068), .Z(n1323) );
  NANDN U2003 ( .A(n28823), .B(n42115), .Z(n1324) );
  AND U2004 ( .A(n1323), .B(n1324), .Z(n28865) );
  NANDN U2005 ( .A(n28859), .B(n42047), .Z(n1325) );
  NANDN U2006 ( .A(n28896), .B(n4067), .Z(n1326) );
  NAND U2007 ( .A(n1325), .B(n1326), .Z(n28907) );
  NANDN U2008 ( .A(n28934), .B(n4068), .Z(n1327) );
  NANDN U2009 ( .A(n28900), .B(n42115), .Z(n1328) );
  AND U2010 ( .A(n1327), .B(n1328), .Z(n28939) );
  NANDN U2011 ( .A(n28933), .B(n42047), .Z(n1329) );
  NANDN U2012 ( .A(n28970), .B(n4067), .Z(n1330) );
  NAND U2013 ( .A(n1329), .B(n1330), .Z(n28981) );
  NANDN U2014 ( .A(n29011), .B(n4068), .Z(n1331) );
  NANDN U2015 ( .A(n28974), .B(n42115), .Z(n1332) );
  AND U2016 ( .A(n1331), .B(n1332), .Z(n29013) );
  NANDN U2017 ( .A(n29007), .B(n42047), .Z(n1333) );
  NANDN U2018 ( .A(n29044), .B(n4067), .Z(n1334) );
  NAND U2019 ( .A(n1333), .B(n1334), .Z(n29055) );
  NANDN U2020 ( .A(n29082), .B(n4068), .Z(n1335) );
  NANDN U2021 ( .A(n29045), .B(n42115), .Z(n1336) );
  AND U2022 ( .A(n1335), .B(n1336), .Z(n29087) );
  NANDN U2023 ( .A(n29081), .B(n42047), .Z(n1337) );
  NANDN U2024 ( .A(n29118), .B(n4067), .Z(n1338) );
  NAND U2025 ( .A(n1337), .B(n1338), .Z(n29129) );
  NANDN U2026 ( .A(n29159), .B(n4068), .Z(n1339) );
  NANDN U2027 ( .A(n29122), .B(n42115), .Z(n1340) );
  AND U2028 ( .A(n1339), .B(n1340), .Z(n29161) );
  NANDN U2029 ( .A(n29155), .B(n42047), .Z(n1341) );
  NANDN U2030 ( .A(n29192), .B(n4067), .Z(n1342) );
  NAND U2031 ( .A(n1341), .B(n1342), .Z(n29203) );
  NANDN U2032 ( .A(n29230), .B(n4068), .Z(n1343) );
  NANDN U2033 ( .A(n29196), .B(n42115), .Z(n1344) );
  AND U2034 ( .A(n1343), .B(n1344), .Z(n29235) );
  NANDN U2035 ( .A(n29229), .B(n42047), .Z(n1345) );
  NANDN U2036 ( .A(n29266), .B(n4067), .Z(n1346) );
  NAND U2037 ( .A(n1345), .B(n1346), .Z(n29277) );
  NANDN U2038 ( .A(n29307), .B(n4068), .Z(n1347) );
  NANDN U2039 ( .A(n29270), .B(n42115), .Z(n1348) );
  AND U2040 ( .A(n1347), .B(n1348), .Z(n29309) );
  NANDN U2041 ( .A(n29303), .B(n42047), .Z(n1349) );
  NANDN U2042 ( .A(n29340), .B(n4067), .Z(n1350) );
  NAND U2043 ( .A(n1349), .B(n1350), .Z(n29351) );
  NANDN U2044 ( .A(n29381), .B(n4068), .Z(n1351) );
  NANDN U2045 ( .A(n29344), .B(n42115), .Z(n1352) );
  AND U2046 ( .A(n1351), .B(n1352), .Z(n29383) );
  NANDN U2047 ( .A(n29377), .B(n42047), .Z(n1353) );
  NANDN U2048 ( .A(n29414), .B(n4067), .Z(n1354) );
  NAND U2049 ( .A(n1353), .B(n1354), .Z(n29425) );
  NANDN U2050 ( .A(n29455), .B(n4068), .Z(n1355) );
  NANDN U2051 ( .A(n29418), .B(n42115), .Z(n1356) );
  AND U2052 ( .A(n1355), .B(n1356), .Z(n29457) );
  NANDN U2053 ( .A(n29451), .B(n42047), .Z(n1357) );
  NANDN U2054 ( .A(n29488), .B(n4067), .Z(n1358) );
  NAND U2055 ( .A(n1357), .B(n1358), .Z(n29499) );
  NANDN U2056 ( .A(n29526), .B(n4068), .Z(n1359) );
  NANDN U2057 ( .A(n29489), .B(n42115), .Z(n1360) );
  AND U2058 ( .A(n1359), .B(n1360), .Z(n29531) );
  NANDN U2059 ( .A(n29525), .B(n42047), .Z(n1361) );
  NANDN U2060 ( .A(n29562), .B(n4067), .Z(n1362) );
  NAND U2061 ( .A(n1361), .B(n1362), .Z(n29574) );
  NANDN U2062 ( .A(n29604), .B(n4068), .Z(n1363) );
  NANDN U2063 ( .A(n29567), .B(n42115), .Z(n1364) );
  AND U2064 ( .A(n1363), .B(n1364), .Z(n29606) );
  NANDN U2065 ( .A(n29600), .B(n42047), .Z(n1365) );
  NANDN U2066 ( .A(n29637), .B(n4067), .Z(n1366) );
  NAND U2067 ( .A(n1365), .B(n1366), .Z(n29648) );
  NANDN U2068 ( .A(n29678), .B(n4068), .Z(n1367) );
  NANDN U2069 ( .A(n29641), .B(n42115), .Z(n1368) );
  AND U2070 ( .A(n1367), .B(n1368), .Z(n29680) );
  NANDN U2071 ( .A(n29674), .B(n42047), .Z(n1369) );
  NANDN U2072 ( .A(n29711), .B(n4067), .Z(n1370) );
  NAND U2073 ( .A(n1369), .B(n1370), .Z(n29722) );
  NANDN U2074 ( .A(n29752), .B(n4068), .Z(n1371) );
  NANDN U2075 ( .A(n29712), .B(n42115), .Z(n1372) );
  AND U2076 ( .A(n1371), .B(n1372), .Z(n29754) );
  NANDN U2077 ( .A(n29748), .B(n42047), .Z(n1373) );
  NANDN U2078 ( .A(n29785), .B(n4067), .Z(n1374) );
  NAND U2079 ( .A(n1373), .B(n1374), .Z(n29796) );
  NANDN U2080 ( .A(n29826), .B(n4068), .Z(n1375) );
  NANDN U2081 ( .A(n29786), .B(n42115), .Z(n1376) );
  AND U2082 ( .A(n1375), .B(n1376), .Z(n29828) );
  NANDN U2083 ( .A(n29822), .B(n42047), .Z(n1377) );
  NANDN U2084 ( .A(n29859), .B(n4067), .Z(n1378) );
  NAND U2085 ( .A(n1377), .B(n1378), .Z(n29870) );
  NANDN U2086 ( .A(n29897), .B(n4068), .Z(n1379) );
  NANDN U2087 ( .A(n29863), .B(n42115), .Z(n1380) );
  AND U2088 ( .A(n1379), .B(n1380), .Z(n29902) );
  NANDN U2089 ( .A(n29896), .B(n42047), .Z(n1381) );
  NANDN U2090 ( .A(n29933), .B(n4067), .Z(n1382) );
  NAND U2091 ( .A(n1381), .B(n1382), .Z(n29944) );
  NANDN U2092 ( .A(n29974), .B(n4068), .Z(n1383) );
  NANDN U2093 ( .A(n29934), .B(n42115), .Z(n1384) );
  AND U2094 ( .A(n1383), .B(n1384), .Z(n29976) );
  NANDN U2095 ( .A(n29970), .B(n42047), .Z(n1385) );
  NANDN U2096 ( .A(n30007), .B(n4067), .Z(n1386) );
  NAND U2097 ( .A(n1385), .B(n1386), .Z(n30018) );
  NANDN U2098 ( .A(n30045), .B(n4068), .Z(n1387) );
  NANDN U2099 ( .A(n30011), .B(n42115), .Z(n1388) );
  AND U2100 ( .A(n1387), .B(n1388), .Z(n30050) );
  NANDN U2101 ( .A(n30044), .B(n42047), .Z(n1389) );
  NANDN U2102 ( .A(n30081), .B(n4067), .Z(n1390) );
  NAND U2103 ( .A(n1389), .B(n1390), .Z(n30092) );
  NANDN U2104 ( .A(n30122), .B(n4068), .Z(n1391) );
  NANDN U2105 ( .A(n30085), .B(n42115), .Z(n1392) );
  AND U2106 ( .A(n1391), .B(n1392), .Z(n30124) );
  NANDN U2107 ( .A(n30118), .B(n42047), .Z(n1393) );
  NANDN U2108 ( .A(n30155), .B(n4067), .Z(n1394) );
  NAND U2109 ( .A(n1393), .B(n1394), .Z(n30166) );
  NANDN U2110 ( .A(n30193), .B(n4068), .Z(n1395) );
  NANDN U2111 ( .A(n30159), .B(n42115), .Z(n1396) );
  AND U2112 ( .A(n1395), .B(n1396), .Z(n30198) );
  NANDN U2113 ( .A(n30192), .B(n42047), .Z(n1397) );
  NANDN U2114 ( .A(n30229), .B(n4067), .Z(n1398) );
  NAND U2115 ( .A(n1397), .B(n1398), .Z(n30240) );
  NANDN U2116 ( .A(n30270), .B(n4068), .Z(n1399) );
  NANDN U2117 ( .A(n30230), .B(n42115), .Z(n1400) );
  AND U2118 ( .A(n1399), .B(n1400), .Z(n30272) );
  NANDN U2119 ( .A(n30266), .B(n42047), .Z(n1401) );
  NANDN U2120 ( .A(n30303), .B(n4067), .Z(n1402) );
  NAND U2121 ( .A(n1401), .B(n1402), .Z(n30314) );
  NANDN U2122 ( .A(n30344), .B(n4068), .Z(n1403) );
  NANDN U2123 ( .A(n30304), .B(n42115), .Z(n1404) );
  AND U2124 ( .A(n1403), .B(n1404), .Z(n30346) );
  NANDN U2125 ( .A(n30340), .B(n42047), .Z(n1405) );
  NANDN U2126 ( .A(n30377), .B(n4067), .Z(n1406) );
  NAND U2127 ( .A(n1405), .B(n1406), .Z(n30388) );
  NANDN U2128 ( .A(n30418), .B(n4068), .Z(n1407) );
  NANDN U2129 ( .A(n30381), .B(n42115), .Z(n1408) );
  AND U2130 ( .A(n1407), .B(n1408), .Z(n30420) );
  NANDN U2131 ( .A(n30414), .B(n42047), .Z(n1409) );
  NANDN U2132 ( .A(n30451), .B(n4067), .Z(n1410) );
  NAND U2133 ( .A(n1409), .B(n1410), .Z(n30462) );
  NANDN U2134 ( .A(n30492), .B(n4068), .Z(n1411) );
  NANDN U2135 ( .A(n30452), .B(n42115), .Z(n1412) );
  AND U2136 ( .A(n1411), .B(n1412), .Z(n30494) );
  NANDN U2137 ( .A(n30488), .B(n42047), .Z(n1413) );
  NANDN U2138 ( .A(n30525), .B(n4067), .Z(n1414) );
  NAND U2139 ( .A(n1413), .B(n1414), .Z(n30536) );
  NANDN U2140 ( .A(n30563), .B(n4068), .Z(n1415) );
  NANDN U2141 ( .A(n30529), .B(n42115), .Z(n1416) );
  AND U2142 ( .A(n1415), .B(n1416), .Z(n30568) );
  NANDN U2143 ( .A(n30562), .B(n42047), .Z(n1417) );
  NANDN U2144 ( .A(n30599), .B(n4067), .Z(n1418) );
  NAND U2145 ( .A(n1417), .B(n1418), .Z(n30610) );
  NANDN U2146 ( .A(n30640), .B(n4068), .Z(n1419) );
  NANDN U2147 ( .A(n30603), .B(n42115), .Z(n1420) );
  AND U2148 ( .A(n1419), .B(n1420), .Z(n30642) );
  NANDN U2149 ( .A(n30636), .B(n42047), .Z(n1421) );
  NANDN U2150 ( .A(n30673), .B(n4067), .Z(n1422) );
  NAND U2151 ( .A(n1421), .B(n1422), .Z(n30684) );
  NANDN U2152 ( .A(n30711), .B(n4068), .Z(n1423) );
  NANDN U2153 ( .A(n30677), .B(n42115), .Z(n1424) );
  AND U2154 ( .A(n1423), .B(n1424), .Z(n30716) );
  NANDN U2155 ( .A(n30710), .B(n42047), .Z(n1425) );
  NANDN U2156 ( .A(n30747), .B(n4067), .Z(n1426) );
  NAND U2157 ( .A(n1425), .B(n1426), .Z(n30758) );
  NANDN U2158 ( .A(n30788), .B(n4068), .Z(n1427) );
  NANDN U2159 ( .A(n30748), .B(n42115), .Z(n1428) );
  AND U2160 ( .A(n1427), .B(n1428), .Z(n30790) );
  NANDN U2161 ( .A(n30784), .B(n42047), .Z(n1429) );
  NANDN U2162 ( .A(n30821), .B(n4067), .Z(n1430) );
  NAND U2163 ( .A(n1429), .B(n1430), .Z(n30832) );
  NANDN U2164 ( .A(n30862), .B(n4068), .Z(n1431) );
  NANDN U2165 ( .A(n30822), .B(n42115), .Z(n1432) );
  AND U2166 ( .A(n1431), .B(n1432), .Z(n30864) );
  NANDN U2167 ( .A(n30858), .B(n42047), .Z(n1433) );
  NANDN U2168 ( .A(n30895), .B(n4067), .Z(n1434) );
  NAND U2169 ( .A(n1433), .B(n1434), .Z(n30906) );
  NANDN U2170 ( .A(n30936), .B(n4068), .Z(n1435) );
  NANDN U2171 ( .A(n30899), .B(n42115), .Z(n1436) );
  AND U2172 ( .A(n1435), .B(n1436), .Z(n30938) );
  NANDN U2173 ( .A(n30932), .B(n42047), .Z(n1437) );
  NANDN U2174 ( .A(n30969), .B(n4067), .Z(n1438) );
  NAND U2175 ( .A(n1437), .B(n1438), .Z(n30980) );
  NANDN U2176 ( .A(n31010), .B(n4068), .Z(n1439) );
  NANDN U2177 ( .A(n30970), .B(n42115), .Z(n1440) );
  AND U2178 ( .A(n1439), .B(n1440), .Z(n31012) );
  NANDN U2179 ( .A(n31006), .B(n42047), .Z(n1441) );
  NANDN U2180 ( .A(n31043), .B(n4067), .Z(n1442) );
  NAND U2181 ( .A(n1441), .B(n1442), .Z(n31054) );
  NANDN U2182 ( .A(n31084), .B(n4068), .Z(n1443) );
  NANDN U2183 ( .A(n31047), .B(n42115), .Z(n1444) );
  AND U2184 ( .A(n1443), .B(n1444), .Z(n31086) );
  NANDN U2185 ( .A(n31080), .B(n42047), .Z(n1445) );
  NANDN U2186 ( .A(n31117), .B(n4067), .Z(n1446) );
  NAND U2187 ( .A(n1445), .B(n1446), .Z(n31128) );
  NANDN U2188 ( .A(n31155), .B(n4068), .Z(n1447) );
  NANDN U2189 ( .A(n31121), .B(n42115), .Z(n1448) );
  AND U2190 ( .A(n1447), .B(n1448), .Z(n31160) );
  NANDN U2191 ( .A(n31154), .B(n42047), .Z(n1449) );
  NANDN U2192 ( .A(n31191), .B(n4067), .Z(n1450) );
  NAND U2193 ( .A(n1449), .B(n1450), .Z(n31202) );
  NANDN U2194 ( .A(n31232), .B(n4068), .Z(n1451) );
  NANDN U2195 ( .A(n31195), .B(n42115), .Z(n1452) );
  AND U2196 ( .A(n1451), .B(n1452), .Z(n31234) );
  NANDN U2197 ( .A(n31228), .B(n42047), .Z(n1453) );
  NANDN U2198 ( .A(n31265), .B(n4067), .Z(n1454) );
  NAND U2199 ( .A(n1453), .B(n1454), .Z(n31276) );
  NANDN U2200 ( .A(n31306), .B(n4068), .Z(n1455) );
  NANDN U2201 ( .A(n31269), .B(n42115), .Z(n1456) );
  AND U2202 ( .A(n1455), .B(n1456), .Z(n31308) );
  NANDN U2203 ( .A(n31302), .B(n42047), .Z(n1457) );
  NANDN U2204 ( .A(n31339), .B(n4067), .Z(n1458) );
  NAND U2205 ( .A(n1457), .B(n1458), .Z(n31350) );
  NANDN U2206 ( .A(n31380), .B(n4068), .Z(n1459) );
  NANDN U2207 ( .A(n31340), .B(n42115), .Z(n1460) );
  AND U2208 ( .A(n1459), .B(n1460), .Z(n31382) );
  NANDN U2209 ( .A(n31376), .B(n42047), .Z(n1461) );
  NANDN U2210 ( .A(n31413), .B(n4067), .Z(n1462) );
  NAND U2211 ( .A(n1461), .B(n1462), .Z(n31424) );
  NANDN U2212 ( .A(n31454), .B(n4068), .Z(n1463) );
  NANDN U2213 ( .A(n31417), .B(n42115), .Z(n1464) );
  AND U2214 ( .A(n1463), .B(n1464), .Z(n31456) );
  NANDN U2215 ( .A(n31450), .B(n42047), .Z(n1465) );
  NANDN U2216 ( .A(n31487), .B(n4067), .Z(n1466) );
  NAND U2217 ( .A(n1465), .B(n1466), .Z(n31498) );
  NANDN U2218 ( .A(n31525), .B(n4068), .Z(n1467) );
  NANDN U2219 ( .A(n31491), .B(n42115), .Z(n1468) );
  AND U2220 ( .A(n1467), .B(n1468), .Z(n31530) );
  NANDN U2221 ( .A(n31524), .B(n42047), .Z(n1469) );
  NANDN U2222 ( .A(n31561), .B(n4067), .Z(n1470) );
  NAND U2223 ( .A(n1469), .B(n1470), .Z(n31572) );
  NANDN U2224 ( .A(n31602), .B(n4068), .Z(n1471) );
  NANDN U2225 ( .A(n31562), .B(n42115), .Z(n1472) );
  AND U2226 ( .A(n1471), .B(n1472), .Z(n31604) );
  NANDN U2227 ( .A(n31598), .B(n42047), .Z(n1473) );
  NANDN U2228 ( .A(n31635), .B(n4067), .Z(n1474) );
  NAND U2229 ( .A(n1473), .B(n1474), .Z(n31646) );
  NANDN U2230 ( .A(n31673), .B(n4068), .Z(n1475) );
  NANDN U2231 ( .A(n31639), .B(n42115), .Z(n1476) );
  AND U2232 ( .A(n1475), .B(n1476), .Z(n31678) );
  NANDN U2233 ( .A(n31672), .B(n42047), .Z(n1477) );
  NANDN U2234 ( .A(n31709), .B(n4067), .Z(n1478) );
  NAND U2235 ( .A(n1477), .B(n1478), .Z(n31720) );
  NANDN U2236 ( .A(n31747), .B(n4068), .Z(n1479) );
  NANDN U2237 ( .A(n31713), .B(n42115), .Z(n1480) );
  AND U2238 ( .A(n1479), .B(n1480), .Z(n31752) );
  NANDN U2239 ( .A(n31746), .B(n42047), .Z(n1481) );
  NANDN U2240 ( .A(n31783), .B(n4067), .Z(n1482) );
  NAND U2241 ( .A(n1481), .B(n1482), .Z(n31794) );
  NANDN U2242 ( .A(n31824), .B(n4068), .Z(n1483) );
  NANDN U2243 ( .A(n31787), .B(n42115), .Z(n1484) );
  AND U2244 ( .A(n1483), .B(n1484), .Z(n31826) );
  NANDN U2245 ( .A(n31820), .B(n42047), .Z(n1485) );
  NANDN U2246 ( .A(n31857), .B(n4067), .Z(n1486) );
  NAND U2247 ( .A(n1485), .B(n1486), .Z(n31868) );
  NANDN U2248 ( .A(n31898), .B(n4068), .Z(n1487) );
  NANDN U2249 ( .A(n31858), .B(n42115), .Z(n1488) );
  AND U2250 ( .A(n1487), .B(n1488), .Z(n31900) );
  NANDN U2251 ( .A(n31894), .B(n42047), .Z(n1489) );
  NANDN U2252 ( .A(n31931), .B(n4067), .Z(n1490) );
  NAND U2253 ( .A(n1489), .B(n1490), .Z(n31942) );
  NANDN U2254 ( .A(n31972), .B(n4068), .Z(n1491) );
  NANDN U2255 ( .A(n31935), .B(n42115), .Z(n1492) );
  AND U2256 ( .A(n1491), .B(n1492), .Z(n31974) );
  NANDN U2257 ( .A(n31968), .B(n42047), .Z(n1493) );
  NANDN U2258 ( .A(n32005), .B(n4067), .Z(n1494) );
  NAND U2259 ( .A(n1493), .B(n1494), .Z(n32016) );
  NANDN U2260 ( .A(n32046), .B(n4068), .Z(n1495) );
  NANDN U2261 ( .A(n32006), .B(n42115), .Z(n1496) );
  AND U2262 ( .A(n1495), .B(n1496), .Z(n32048) );
  NANDN U2263 ( .A(n32042), .B(n42047), .Z(n1497) );
  NANDN U2264 ( .A(n32079), .B(n4067), .Z(n1498) );
  NAND U2265 ( .A(n1497), .B(n1498), .Z(n32090) );
  NANDN U2266 ( .A(n32120), .B(n4068), .Z(n1499) );
  NANDN U2267 ( .A(n32083), .B(n42115), .Z(n1500) );
  AND U2268 ( .A(n1499), .B(n1500), .Z(n32122) );
  NANDN U2269 ( .A(n32116), .B(n42047), .Z(n1501) );
  NANDN U2270 ( .A(n32153), .B(n4067), .Z(n1502) );
  NAND U2271 ( .A(n1501), .B(n1502), .Z(n32164) );
  NANDN U2272 ( .A(n32194), .B(n4068), .Z(n1503) );
  NANDN U2273 ( .A(n32157), .B(n42115), .Z(n1504) );
  AND U2274 ( .A(n1503), .B(n1504), .Z(n32196) );
  NANDN U2275 ( .A(n32190), .B(n42047), .Z(n1505) );
  NANDN U2276 ( .A(n32227), .B(n4067), .Z(n1506) );
  NAND U2277 ( .A(n1505), .B(n1506), .Z(n32238) );
  NANDN U2278 ( .A(n32268), .B(n4068), .Z(n1507) );
  NANDN U2279 ( .A(n32231), .B(n42115), .Z(n1508) );
  AND U2280 ( .A(n1507), .B(n1508), .Z(n32270) );
  NANDN U2281 ( .A(n32264), .B(n42047), .Z(n1509) );
  NANDN U2282 ( .A(n32301), .B(n4067), .Z(n1510) );
  NAND U2283 ( .A(n1509), .B(n1510), .Z(n32312) );
  NANDN U2284 ( .A(n32339), .B(n4068), .Z(n1511) );
  NANDN U2285 ( .A(n32302), .B(n42115), .Z(n1512) );
  AND U2286 ( .A(n1511), .B(n1512), .Z(n32344) );
  NANDN U2287 ( .A(n32338), .B(n42047), .Z(n1513) );
  NANDN U2288 ( .A(n32375), .B(n4067), .Z(n1514) );
  NAND U2289 ( .A(n1513), .B(n1514), .Z(n32386) );
  NANDN U2290 ( .A(n32416), .B(n4068), .Z(n1515) );
  NANDN U2291 ( .A(n32376), .B(n42115), .Z(n1516) );
  AND U2292 ( .A(n1515), .B(n1516), .Z(n32418) );
  NANDN U2293 ( .A(n32412), .B(n42047), .Z(n1517) );
  NANDN U2294 ( .A(n32449), .B(n4067), .Z(n1518) );
  NAND U2295 ( .A(n1517), .B(n1518), .Z(n32460) );
  NANDN U2296 ( .A(n32490), .B(n4068), .Z(n1519) );
  NANDN U2297 ( .A(n32453), .B(n42115), .Z(n1520) );
  AND U2298 ( .A(n1519), .B(n1520), .Z(n32492) );
  NANDN U2299 ( .A(n32486), .B(n42047), .Z(n1521) );
  NANDN U2300 ( .A(n32523), .B(n4067), .Z(n1522) );
  NAND U2301 ( .A(n1521), .B(n1522), .Z(n32534) );
  NANDN U2302 ( .A(n32564), .B(n4068), .Z(n1523) );
  NANDN U2303 ( .A(n32527), .B(n42115), .Z(n1524) );
  AND U2304 ( .A(n1523), .B(n1524), .Z(n32566) );
  NANDN U2305 ( .A(n32560), .B(n42047), .Z(n1525) );
  NANDN U2306 ( .A(n32597), .B(n4067), .Z(n1526) );
  NAND U2307 ( .A(n1525), .B(n1526), .Z(n32608) );
  NANDN U2308 ( .A(n32635), .B(n4068), .Z(n1527) );
  NANDN U2309 ( .A(n32598), .B(n42115), .Z(n1528) );
  AND U2310 ( .A(n1527), .B(n1528), .Z(n32640) );
  NANDN U2311 ( .A(n32634), .B(n42047), .Z(n1529) );
  NANDN U2312 ( .A(n32671), .B(n4067), .Z(n1530) );
  NAND U2313 ( .A(n1529), .B(n1530), .Z(n32682) );
  NANDN U2314 ( .A(n32709), .B(n4068), .Z(n1531) );
  NANDN U2315 ( .A(n32672), .B(n42115), .Z(n1532) );
  AND U2316 ( .A(n1531), .B(n1532), .Z(n32714) );
  NANDN U2317 ( .A(n32708), .B(n42047), .Z(n1533) );
  NANDN U2318 ( .A(n32745), .B(n4067), .Z(n1534) );
  NAND U2319 ( .A(n1533), .B(n1534), .Z(n32756) );
  NANDN U2320 ( .A(n32783), .B(n4068), .Z(n1535) );
  NANDN U2321 ( .A(n32746), .B(n42115), .Z(n1536) );
  AND U2322 ( .A(n1535), .B(n1536), .Z(n32788) );
  NANDN U2323 ( .A(n32782), .B(n42047), .Z(n1537) );
  NANDN U2324 ( .A(n32819), .B(n4067), .Z(n1538) );
  NAND U2325 ( .A(n1537), .B(n1538), .Z(n32830) );
  NANDN U2326 ( .A(n32857), .B(n4068), .Z(n1539) );
  NANDN U2327 ( .A(n32820), .B(n42115), .Z(n1540) );
  AND U2328 ( .A(n1539), .B(n1540), .Z(n32862) );
  NANDN U2329 ( .A(n32856), .B(n42047), .Z(n1541) );
  NANDN U2330 ( .A(n32893), .B(n4067), .Z(n1542) );
  NAND U2331 ( .A(n1541), .B(n1542), .Z(n32904) );
  NANDN U2332 ( .A(n32934), .B(n4068), .Z(n1543) );
  NANDN U2333 ( .A(n32897), .B(n42115), .Z(n1544) );
  AND U2334 ( .A(n1543), .B(n1544), .Z(n32936) );
  NANDN U2335 ( .A(n32930), .B(n42047), .Z(n1545) );
  NANDN U2336 ( .A(n32967), .B(n4067), .Z(n1546) );
  NAND U2337 ( .A(n1545), .B(n1546), .Z(n32978) );
  NANDN U2338 ( .A(n33008), .B(n4068), .Z(n1547) );
  NANDN U2339 ( .A(n32971), .B(n42115), .Z(n1548) );
  AND U2340 ( .A(n1547), .B(n1548), .Z(n33010) );
  NANDN U2341 ( .A(n33004), .B(n42047), .Z(n1549) );
  NANDN U2342 ( .A(n33041), .B(n4067), .Z(n1550) );
  NAND U2343 ( .A(n1549), .B(n1550), .Z(n33052) );
  NANDN U2344 ( .A(n33082), .B(n4068), .Z(n1551) );
  NANDN U2345 ( .A(n33045), .B(n42115), .Z(n1552) );
  AND U2346 ( .A(n1551), .B(n1552), .Z(n33084) );
  NANDN U2347 ( .A(n33078), .B(n42047), .Z(n1553) );
  NANDN U2348 ( .A(n33115), .B(n4067), .Z(n1554) );
  NAND U2349 ( .A(n1553), .B(n1554), .Z(n33126) );
  NANDN U2350 ( .A(n33156), .B(n4068), .Z(n1555) );
  NANDN U2351 ( .A(n33116), .B(n42115), .Z(n1556) );
  AND U2352 ( .A(n1555), .B(n1556), .Z(n33158) );
  NANDN U2353 ( .A(n33152), .B(n42047), .Z(n1557) );
  NANDN U2354 ( .A(n33189), .B(n4067), .Z(n1558) );
  NAND U2355 ( .A(n1557), .B(n1558), .Z(n33200) );
  NANDN U2356 ( .A(n33227), .B(n4068), .Z(n1559) );
  NANDN U2357 ( .A(n33190), .B(n42115), .Z(n1560) );
  AND U2358 ( .A(n1559), .B(n1560), .Z(n33232) );
  NANDN U2359 ( .A(n33226), .B(n42047), .Z(n1561) );
  NANDN U2360 ( .A(n33263), .B(n4067), .Z(n1562) );
  NAND U2361 ( .A(n1561), .B(n1562), .Z(n33274) );
  NANDN U2362 ( .A(n33301), .B(n4068), .Z(n1563) );
  NANDN U2363 ( .A(n33267), .B(n42115), .Z(n1564) );
  AND U2364 ( .A(n1563), .B(n1564), .Z(n33306) );
  NANDN U2365 ( .A(n33300), .B(n42047), .Z(n1565) );
  NANDN U2366 ( .A(n33337), .B(n4067), .Z(n1566) );
  NAND U2367 ( .A(n1565), .B(n1566), .Z(n33348) );
  NANDN U2368 ( .A(n33378), .B(n4068), .Z(n1567) );
  NANDN U2369 ( .A(n33341), .B(n42115), .Z(n1568) );
  AND U2370 ( .A(n1567), .B(n1568), .Z(n33380) );
  NANDN U2371 ( .A(n33374), .B(n42047), .Z(n1569) );
  NANDN U2372 ( .A(n33411), .B(n4067), .Z(n1570) );
  NAND U2373 ( .A(n1569), .B(n1570), .Z(n33422) );
  NANDN U2374 ( .A(n33449), .B(n4068), .Z(n1571) );
  NANDN U2375 ( .A(n33415), .B(n42115), .Z(n1572) );
  AND U2376 ( .A(n1571), .B(n1572), .Z(n33454) );
  NANDN U2377 ( .A(n33448), .B(n42047), .Z(n1573) );
  NANDN U2378 ( .A(n33485), .B(n4067), .Z(n1574) );
  NAND U2379 ( .A(n1573), .B(n1574), .Z(n33496) );
  NANDN U2380 ( .A(n33523), .B(n4068), .Z(n1575) );
  NANDN U2381 ( .A(n33489), .B(n42115), .Z(n1576) );
  AND U2382 ( .A(n1575), .B(n1576), .Z(n33528) );
  NANDN U2383 ( .A(n33522), .B(n42047), .Z(n1577) );
  NANDN U2384 ( .A(n33559), .B(n4067), .Z(n1578) );
  NAND U2385 ( .A(n1577), .B(n1578), .Z(n33570) );
  NANDN U2386 ( .A(n33600), .B(n4068), .Z(n1579) );
  NANDN U2387 ( .A(n33563), .B(n42115), .Z(n1580) );
  AND U2388 ( .A(n1579), .B(n1580), .Z(n33602) );
  NANDN U2389 ( .A(n33596), .B(n42047), .Z(n1581) );
  NANDN U2390 ( .A(n33633), .B(n4067), .Z(n1582) );
  NAND U2391 ( .A(n1581), .B(n1582), .Z(n33644) );
  NANDN U2392 ( .A(n33674), .B(n4068), .Z(n1583) );
  NANDN U2393 ( .A(n33634), .B(n42115), .Z(n1584) );
  AND U2394 ( .A(n1583), .B(n1584), .Z(n33676) );
  NANDN U2395 ( .A(n33670), .B(n42047), .Z(n1585) );
  NANDN U2396 ( .A(n33707), .B(n4067), .Z(n1586) );
  NAND U2397 ( .A(n1585), .B(n1586), .Z(n33718) );
  NANDN U2398 ( .A(n33748), .B(n4068), .Z(n1587) );
  NANDN U2399 ( .A(n33711), .B(n42115), .Z(n1588) );
  AND U2400 ( .A(n1587), .B(n1588), .Z(n33750) );
  NANDN U2401 ( .A(n33744), .B(n42047), .Z(n1589) );
  NANDN U2402 ( .A(n33781), .B(n4067), .Z(n1590) );
  NAND U2403 ( .A(n1589), .B(n1590), .Z(n33792) );
  NANDN U2404 ( .A(n33822), .B(n4068), .Z(n1591) );
  NANDN U2405 ( .A(n33782), .B(n42115), .Z(n1592) );
  AND U2406 ( .A(n1591), .B(n1592), .Z(n33824) );
  NANDN U2407 ( .A(n33818), .B(n42047), .Z(n1593) );
  NANDN U2408 ( .A(n33855), .B(n4067), .Z(n1594) );
  NAND U2409 ( .A(n1593), .B(n1594), .Z(n33866) );
  NANDN U2410 ( .A(n33893), .B(n4068), .Z(n1595) );
  NANDN U2411 ( .A(n33859), .B(n42115), .Z(n1596) );
  AND U2412 ( .A(n1595), .B(n1596), .Z(n33898) );
  NANDN U2413 ( .A(n33892), .B(n42047), .Z(n1597) );
  NANDN U2414 ( .A(n33929), .B(n4067), .Z(n1598) );
  NAND U2415 ( .A(n1597), .B(n1598), .Z(n33940) );
  NANDN U2416 ( .A(n33967), .B(n4068), .Z(n1599) );
  NANDN U2417 ( .A(n33933), .B(n42115), .Z(n1600) );
  AND U2418 ( .A(n1599), .B(n1600), .Z(n33972) );
  NANDN U2419 ( .A(n33966), .B(n42047), .Z(n1601) );
  NANDN U2420 ( .A(n34003), .B(n4067), .Z(n1602) );
  NAND U2421 ( .A(n1601), .B(n1602), .Z(n34014) );
  NANDN U2422 ( .A(n34044), .B(n4068), .Z(n1603) );
  NANDN U2423 ( .A(n34007), .B(n42115), .Z(n1604) );
  AND U2424 ( .A(n1603), .B(n1604), .Z(n34046) );
  NANDN U2425 ( .A(n34040), .B(n42047), .Z(n1605) );
  NANDN U2426 ( .A(n34077), .B(n4067), .Z(n1606) );
  NAND U2427 ( .A(n1605), .B(n1606), .Z(n34088) );
  NANDN U2428 ( .A(n34115), .B(n4068), .Z(n1607) );
  NANDN U2429 ( .A(n34078), .B(n42115), .Z(n1608) );
  AND U2430 ( .A(n1607), .B(n1608), .Z(n34120) );
  NANDN U2431 ( .A(n34114), .B(n42047), .Z(n1609) );
  NANDN U2432 ( .A(n34151), .B(n4067), .Z(n1610) );
  NAND U2433 ( .A(n1609), .B(n1610), .Z(n34162) );
  NANDN U2434 ( .A(n34189), .B(n4068), .Z(n1611) );
  NANDN U2435 ( .A(n34155), .B(n42115), .Z(n1612) );
  AND U2436 ( .A(n1611), .B(n1612), .Z(n34194) );
  NANDN U2437 ( .A(n34188), .B(n42047), .Z(n1613) );
  NANDN U2438 ( .A(n34225), .B(n4067), .Z(n1614) );
  NAND U2439 ( .A(n1613), .B(n1614), .Z(n34236) );
  NANDN U2440 ( .A(n34266), .B(n4068), .Z(n1615) );
  NANDN U2441 ( .A(n34229), .B(n42115), .Z(n1616) );
  AND U2442 ( .A(n1615), .B(n1616), .Z(n34268) );
  NANDN U2443 ( .A(n34262), .B(n42047), .Z(n1617) );
  NANDN U2444 ( .A(n34299), .B(n4067), .Z(n1618) );
  NAND U2445 ( .A(n1617), .B(n1618), .Z(n34310) );
  NANDN U2446 ( .A(n34340), .B(n4068), .Z(n1619) );
  NANDN U2447 ( .A(n34300), .B(n42115), .Z(n1620) );
  AND U2448 ( .A(n1619), .B(n1620), .Z(n34342) );
  NANDN U2449 ( .A(n34336), .B(n42047), .Z(n1621) );
  NANDN U2450 ( .A(n34373), .B(n4067), .Z(n1622) );
  NAND U2451 ( .A(n1621), .B(n1622), .Z(n34384) );
  NANDN U2452 ( .A(n34411), .B(n4068), .Z(n1623) );
  NANDN U2453 ( .A(n34374), .B(n42115), .Z(n1624) );
  AND U2454 ( .A(n1623), .B(n1624), .Z(n34416) );
  NANDN U2455 ( .A(n34410), .B(n42047), .Z(n1625) );
  NANDN U2456 ( .A(n34447), .B(n4067), .Z(n1626) );
  NAND U2457 ( .A(n1625), .B(n1626), .Z(n34458) );
  NANDN U2458 ( .A(n34485), .B(n4068), .Z(n1627) );
  NANDN U2459 ( .A(n34448), .B(n42115), .Z(n1628) );
  AND U2460 ( .A(n1627), .B(n1628), .Z(n34490) );
  NANDN U2461 ( .A(n34484), .B(n42047), .Z(n1629) );
  NANDN U2462 ( .A(n34521), .B(n4067), .Z(n1630) );
  NAND U2463 ( .A(n1629), .B(n1630), .Z(n34532) );
  NANDN U2464 ( .A(n34562), .B(n4068), .Z(n1631) );
  NANDN U2465 ( .A(n34525), .B(n42115), .Z(n1632) );
  AND U2466 ( .A(n1631), .B(n1632), .Z(n34564) );
  NANDN U2467 ( .A(n34558), .B(n42047), .Z(n1633) );
  NANDN U2468 ( .A(n34595), .B(n4067), .Z(n1634) );
  NAND U2469 ( .A(n1633), .B(n1634), .Z(n34606) );
  NANDN U2470 ( .A(n34636), .B(n4068), .Z(n1635) );
  NANDN U2471 ( .A(n34596), .B(n42115), .Z(n1636) );
  AND U2472 ( .A(n1635), .B(n1636), .Z(n34638) );
  NANDN U2473 ( .A(n34632), .B(n42047), .Z(n1637) );
  NANDN U2474 ( .A(n34669), .B(n4067), .Z(n1638) );
  NAND U2475 ( .A(n1637), .B(n1638), .Z(n34680) );
  NANDN U2476 ( .A(n34707), .B(n4068), .Z(n1639) );
  NANDN U2477 ( .A(n34670), .B(n42115), .Z(n1640) );
  AND U2478 ( .A(n1639), .B(n1640), .Z(n34712) );
  NANDN U2479 ( .A(n34706), .B(n42047), .Z(n1641) );
  NANDN U2480 ( .A(n34743), .B(n4067), .Z(n1642) );
  NAND U2481 ( .A(n1641), .B(n1642), .Z(n34754) );
  NANDN U2482 ( .A(n34781), .B(n4068), .Z(n1643) );
  NANDN U2483 ( .A(n34744), .B(n42115), .Z(n1644) );
  AND U2484 ( .A(n1643), .B(n1644), .Z(n34786) );
  NANDN U2485 ( .A(n34780), .B(n42047), .Z(n1645) );
  NANDN U2486 ( .A(n34817), .B(n4067), .Z(n1646) );
  NAND U2487 ( .A(n1645), .B(n1646), .Z(n34828) );
  NANDN U2488 ( .A(n34855), .B(n4068), .Z(n1647) );
  NANDN U2489 ( .A(n34818), .B(n42115), .Z(n1648) );
  AND U2490 ( .A(n1647), .B(n1648), .Z(n34860) );
  NANDN U2491 ( .A(n34854), .B(n42047), .Z(n1649) );
  NANDN U2492 ( .A(n34891), .B(n4067), .Z(n1650) );
  NAND U2493 ( .A(n1649), .B(n1650), .Z(n34902) );
  NANDN U2494 ( .A(n34929), .B(n4068), .Z(n1651) );
  NANDN U2495 ( .A(n34892), .B(n42115), .Z(n1652) );
  AND U2496 ( .A(n1651), .B(n1652), .Z(n34934) );
  NANDN U2497 ( .A(n34928), .B(n42047), .Z(n1653) );
  NANDN U2498 ( .A(n34965), .B(n4067), .Z(n1654) );
  NAND U2499 ( .A(n1653), .B(n1654), .Z(n34976) );
  NANDN U2500 ( .A(n35006), .B(n4068), .Z(n1655) );
  NANDN U2501 ( .A(n34969), .B(n42115), .Z(n1656) );
  AND U2502 ( .A(n1655), .B(n1656), .Z(n35008) );
  NANDN U2503 ( .A(n35002), .B(n42047), .Z(n1657) );
  NANDN U2504 ( .A(n35039), .B(n4067), .Z(n1658) );
  NAND U2505 ( .A(n1657), .B(n1658), .Z(n35050) );
  NANDN U2506 ( .A(n35077), .B(n4068), .Z(n1659) );
  NANDN U2507 ( .A(n35043), .B(n42115), .Z(n1660) );
  AND U2508 ( .A(n1659), .B(n1660), .Z(n35082) );
  NANDN U2509 ( .A(n35076), .B(n42047), .Z(n1661) );
  NANDN U2510 ( .A(n35113), .B(n4067), .Z(n1662) );
  NAND U2511 ( .A(n1661), .B(n1662), .Z(n35124) );
  NANDN U2512 ( .A(n35154), .B(n4068), .Z(n1663) );
  NANDN U2513 ( .A(n35114), .B(n42115), .Z(n1664) );
  AND U2514 ( .A(n1663), .B(n1664), .Z(n35156) );
  NANDN U2515 ( .A(n35150), .B(n42047), .Z(n1665) );
  NANDN U2516 ( .A(n35187), .B(n4067), .Z(n1666) );
  NAND U2517 ( .A(n1665), .B(n1666), .Z(n35198) );
  NANDN U2518 ( .A(n35228), .B(n4068), .Z(n1667) );
  NANDN U2519 ( .A(n35191), .B(n42115), .Z(n1668) );
  AND U2520 ( .A(n1667), .B(n1668), .Z(n35230) );
  NANDN U2521 ( .A(n35224), .B(n42047), .Z(n1669) );
  NANDN U2522 ( .A(n35261), .B(n4067), .Z(n1670) );
  NAND U2523 ( .A(n1669), .B(n1670), .Z(n35272) );
  NANDN U2524 ( .A(n35299), .B(n4068), .Z(n1671) );
  NANDN U2525 ( .A(n35265), .B(n42115), .Z(n1672) );
  AND U2526 ( .A(n1671), .B(n1672), .Z(n35304) );
  NANDN U2527 ( .A(n35298), .B(n42047), .Z(n1673) );
  NANDN U2528 ( .A(n35335), .B(n4067), .Z(n1674) );
  NAND U2529 ( .A(n1673), .B(n1674), .Z(n35346) );
  NANDN U2530 ( .A(n35373), .B(n4068), .Z(n1675) );
  NANDN U2531 ( .A(n35336), .B(n42115), .Z(n1676) );
  AND U2532 ( .A(n1675), .B(n1676), .Z(n35378) );
  NANDN U2533 ( .A(n35372), .B(n42047), .Z(n1677) );
  NANDN U2534 ( .A(n35409), .B(n4067), .Z(n1678) );
  NAND U2535 ( .A(n1677), .B(n1678), .Z(n35420) );
  NANDN U2536 ( .A(n35447), .B(n4068), .Z(n1679) );
  NANDN U2537 ( .A(n35410), .B(n42115), .Z(n1680) );
  AND U2538 ( .A(n1679), .B(n1680), .Z(n35452) );
  NANDN U2539 ( .A(n35446), .B(n42047), .Z(n1681) );
  NANDN U2540 ( .A(n35483), .B(n4067), .Z(n1682) );
  NAND U2541 ( .A(n1681), .B(n1682), .Z(n35494) );
  NANDN U2542 ( .A(n35521), .B(n4068), .Z(n1683) );
  NANDN U2543 ( .A(n35484), .B(n42115), .Z(n1684) );
  AND U2544 ( .A(n1683), .B(n1684), .Z(n35526) );
  NANDN U2545 ( .A(n35520), .B(n42047), .Z(n1685) );
  NANDN U2546 ( .A(n35557), .B(n4067), .Z(n1686) );
  NAND U2547 ( .A(n1685), .B(n1686), .Z(n35568) );
  NANDN U2548 ( .A(n35598), .B(n4068), .Z(n1687) );
  NANDN U2549 ( .A(n35558), .B(n42115), .Z(n1688) );
  AND U2550 ( .A(n1687), .B(n1688), .Z(n35600) );
  NANDN U2551 ( .A(n35594), .B(n42047), .Z(n1689) );
  NANDN U2552 ( .A(n35631), .B(n4067), .Z(n1690) );
  NAND U2553 ( .A(n1689), .B(n1690), .Z(n35642) );
  NANDN U2554 ( .A(n35669), .B(n4068), .Z(n1691) );
  NANDN U2555 ( .A(n35635), .B(n42115), .Z(n1692) );
  AND U2556 ( .A(n1691), .B(n1692), .Z(n35674) );
  NANDN U2557 ( .A(n35668), .B(n42047), .Z(n1693) );
  NANDN U2558 ( .A(n35705), .B(n4067), .Z(n1694) );
  NAND U2559 ( .A(n1693), .B(n1694), .Z(n35716) );
  NANDN U2560 ( .A(n35743), .B(n4068), .Z(n1695) );
  NANDN U2561 ( .A(n35706), .B(n42115), .Z(n1696) );
  AND U2562 ( .A(n1695), .B(n1696), .Z(n35748) );
  NANDN U2563 ( .A(n35742), .B(n42047), .Z(n1697) );
  NANDN U2564 ( .A(n35779), .B(n4067), .Z(n1698) );
  NAND U2565 ( .A(n1697), .B(n1698), .Z(n35790) );
  NANDN U2566 ( .A(n35820), .B(n4068), .Z(n1699) );
  NANDN U2567 ( .A(n35780), .B(n42115), .Z(n1700) );
  AND U2568 ( .A(n1699), .B(n1700), .Z(n35822) );
  NANDN U2569 ( .A(n35816), .B(n42047), .Z(n1701) );
  NANDN U2570 ( .A(n35853), .B(n4067), .Z(n1702) );
  NAND U2571 ( .A(n1701), .B(n1702), .Z(n35864) );
  NANDN U2572 ( .A(n35894), .B(n4068), .Z(n1703) );
  NANDN U2573 ( .A(n35857), .B(n42115), .Z(n1704) );
  AND U2574 ( .A(n1703), .B(n1704), .Z(n35896) );
  NANDN U2575 ( .A(n35890), .B(n42047), .Z(n1705) );
  NANDN U2576 ( .A(n35927), .B(n4067), .Z(n1706) );
  NAND U2577 ( .A(n1705), .B(n1706), .Z(n35938) );
  NANDN U2578 ( .A(n35968), .B(n4068), .Z(n1707) );
  NANDN U2579 ( .A(n35928), .B(n42115), .Z(n1708) );
  AND U2580 ( .A(n1707), .B(n1708), .Z(n35970) );
  NANDN U2581 ( .A(n35964), .B(n42047), .Z(n1709) );
  NANDN U2582 ( .A(n36001), .B(n4067), .Z(n1710) );
  NAND U2583 ( .A(n1709), .B(n1710), .Z(n36012) );
  NANDN U2584 ( .A(n36042), .B(n4068), .Z(n1711) );
  NANDN U2585 ( .A(n36002), .B(n42115), .Z(n1712) );
  AND U2586 ( .A(n1711), .B(n1712), .Z(n36044) );
  NANDN U2587 ( .A(n36038), .B(n42047), .Z(n1713) );
  NANDN U2588 ( .A(n36075), .B(n4067), .Z(n1714) );
  NAND U2589 ( .A(n1713), .B(n1714), .Z(n36086) );
  NANDN U2590 ( .A(n36113), .B(n4068), .Z(n1715) );
  NANDN U2591 ( .A(n36079), .B(n42115), .Z(n1716) );
  AND U2592 ( .A(n1715), .B(n1716), .Z(n36118) );
  NANDN U2593 ( .A(n36112), .B(n42047), .Z(n1717) );
  NANDN U2594 ( .A(n36149), .B(n4067), .Z(n1718) );
  NAND U2595 ( .A(n1717), .B(n1718), .Z(n36160) );
  NANDN U2596 ( .A(n36190), .B(n4068), .Z(n1719) );
  NANDN U2597 ( .A(n36153), .B(n42115), .Z(n1720) );
  AND U2598 ( .A(n1719), .B(n1720), .Z(n36192) );
  NANDN U2599 ( .A(n36186), .B(n42047), .Z(n1721) );
  NANDN U2600 ( .A(n36223), .B(n4067), .Z(n1722) );
  NAND U2601 ( .A(n1721), .B(n1722), .Z(n36234) );
  NANDN U2602 ( .A(n36261), .B(n4068), .Z(n1723) );
  NANDN U2603 ( .A(n36224), .B(n42115), .Z(n1724) );
  AND U2604 ( .A(n1723), .B(n1724), .Z(n36266) );
  NANDN U2605 ( .A(n36260), .B(n42047), .Z(n1725) );
  NANDN U2606 ( .A(n36302), .B(n4067), .Z(n1726) );
  NAND U2607 ( .A(n1725), .B(n1726), .Z(n36313) );
  NANDN U2608 ( .A(n36335), .B(n4068), .Z(n1727) );
  NANDN U2609 ( .A(n36306), .B(n42115), .Z(n1728) );
  AND U2610 ( .A(n1727), .B(n1728), .Z(n36340) );
  NANDN U2611 ( .A(n36334), .B(n42047), .Z(n1729) );
  NANDN U2612 ( .A(n36371), .B(n4067), .Z(n1730) );
  NAND U2613 ( .A(n1729), .B(n1730), .Z(n36382) );
  NANDN U2614 ( .A(n36412), .B(n4068), .Z(n1731) );
  NANDN U2615 ( .A(n36372), .B(n42115), .Z(n1732) );
  AND U2616 ( .A(n1731), .B(n1732), .Z(n36414) );
  NANDN U2617 ( .A(n36408), .B(n42047), .Z(n1733) );
  NANDN U2618 ( .A(n36445), .B(n4067), .Z(n1734) );
  NAND U2619 ( .A(n1733), .B(n1734), .Z(n36456) );
  NANDN U2620 ( .A(n36486), .B(n4068), .Z(n1735) );
  NANDN U2621 ( .A(n36449), .B(n42115), .Z(n1736) );
  AND U2622 ( .A(n1735), .B(n1736), .Z(n36488) );
  NANDN U2623 ( .A(n36482), .B(n42047), .Z(n1737) );
  NANDN U2624 ( .A(n36519), .B(n4067), .Z(n1738) );
  NAND U2625 ( .A(n1737), .B(n1738), .Z(n36530) );
  NANDN U2626 ( .A(n36560), .B(n4068), .Z(n1739) );
  NANDN U2627 ( .A(n36523), .B(n42115), .Z(n1740) );
  AND U2628 ( .A(n1739), .B(n1740), .Z(n36562) );
  NANDN U2629 ( .A(n36556), .B(n42047), .Z(n1741) );
  NANDN U2630 ( .A(n36593), .B(n4067), .Z(n1742) );
  NAND U2631 ( .A(n1741), .B(n1742), .Z(n36604) );
  NANDN U2632 ( .A(n36631), .B(n4068), .Z(n1743) );
  NANDN U2633 ( .A(n36597), .B(n42115), .Z(n1744) );
  AND U2634 ( .A(n1743), .B(n1744), .Z(n36636) );
  NANDN U2635 ( .A(n36630), .B(n42047), .Z(n1745) );
  NANDN U2636 ( .A(n36667), .B(n4067), .Z(n1746) );
  NAND U2637 ( .A(n1745), .B(n1746), .Z(n36678) );
  NANDN U2638 ( .A(n36708), .B(n4068), .Z(n1747) );
  NANDN U2639 ( .A(n36671), .B(n42115), .Z(n1748) );
  AND U2640 ( .A(n1747), .B(n1748), .Z(n36710) );
  NANDN U2641 ( .A(n36704), .B(n42047), .Z(n1749) );
  NANDN U2642 ( .A(n36741), .B(n4067), .Z(n1750) );
  NAND U2643 ( .A(n1749), .B(n1750), .Z(n36752) );
  NANDN U2644 ( .A(n36782), .B(n4068), .Z(n1751) );
  NANDN U2645 ( .A(n36742), .B(n42115), .Z(n1752) );
  AND U2646 ( .A(n1751), .B(n1752), .Z(n36784) );
  NANDN U2647 ( .A(n36778), .B(n42047), .Z(n1753) );
  NANDN U2648 ( .A(n36815), .B(n4067), .Z(n1754) );
  NAND U2649 ( .A(n1753), .B(n1754), .Z(n36826) );
  NANDN U2650 ( .A(n36856), .B(n4068), .Z(n1755) );
  NANDN U2651 ( .A(n36816), .B(n42115), .Z(n1756) );
  AND U2652 ( .A(n1755), .B(n1756), .Z(n36858) );
  NANDN U2653 ( .A(n36852), .B(n42047), .Z(n1757) );
  NANDN U2654 ( .A(n36889), .B(n4067), .Z(n1758) );
  NAND U2655 ( .A(n1757), .B(n1758), .Z(n36900) );
  NANDN U2656 ( .A(n36927), .B(n4068), .Z(n1759) );
  NANDN U2657 ( .A(n36893), .B(n42115), .Z(n1760) );
  AND U2658 ( .A(n1759), .B(n1760), .Z(n36932) );
  NANDN U2659 ( .A(n36926), .B(n42047), .Z(n1761) );
  NANDN U2660 ( .A(n36963), .B(n4067), .Z(n1762) );
  NAND U2661 ( .A(n1761), .B(n1762), .Z(n36974) );
  NANDN U2662 ( .A(n37001), .B(n4068), .Z(n1763) );
  NANDN U2663 ( .A(n36967), .B(n42115), .Z(n1764) );
  AND U2664 ( .A(n1763), .B(n1764), .Z(n37006) );
  NANDN U2665 ( .A(n37000), .B(n42047), .Z(n1765) );
  NANDN U2666 ( .A(n37037), .B(n4067), .Z(n1766) );
  NAND U2667 ( .A(n1765), .B(n1766), .Z(n37048) );
  NANDN U2668 ( .A(n37078), .B(n4068), .Z(n1767) );
  NANDN U2669 ( .A(n37041), .B(n42115), .Z(n1768) );
  AND U2670 ( .A(n1767), .B(n1768), .Z(n37080) );
  NANDN U2671 ( .A(n37074), .B(n42047), .Z(n1769) );
  NANDN U2672 ( .A(n37111), .B(n4067), .Z(n1770) );
  NAND U2673 ( .A(n1769), .B(n1770), .Z(n37122) );
  NANDN U2674 ( .A(n37152), .B(n4068), .Z(n1771) );
  NANDN U2675 ( .A(n37112), .B(n42115), .Z(n1772) );
  AND U2676 ( .A(n1771), .B(n1772), .Z(n37154) );
  NANDN U2677 ( .A(n37148), .B(n42047), .Z(n1773) );
  NANDN U2678 ( .A(n37185), .B(n4067), .Z(n1774) );
  NAND U2679 ( .A(n1773), .B(n1774), .Z(n37196) );
  NANDN U2680 ( .A(n37226), .B(n4068), .Z(n1775) );
  NANDN U2681 ( .A(n37189), .B(n42115), .Z(n1776) );
  AND U2682 ( .A(n1775), .B(n1776), .Z(n37228) );
  NANDN U2683 ( .A(n37222), .B(n42047), .Z(n1777) );
  NANDN U2684 ( .A(n37259), .B(n4067), .Z(n1778) );
  NAND U2685 ( .A(n1777), .B(n1778), .Z(n37270) );
  NANDN U2686 ( .A(n37297), .B(n4068), .Z(n1779) );
  NANDN U2687 ( .A(n37263), .B(n42115), .Z(n1780) );
  AND U2688 ( .A(n1779), .B(n1780), .Z(n37302) );
  NANDN U2689 ( .A(n37296), .B(n42047), .Z(n1781) );
  NANDN U2690 ( .A(n37333), .B(n4067), .Z(n1782) );
  NAND U2691 ( .A(n1781), .B(n1782), .Z(n37344) );
  NANDN U2692 ( .A(n37371), .B(n4068), .Z(n1783) );
  NANDN U2693 ( .A(n37334), .B(n42115), .Z(n1784) );
  AND U2694 ( .A(n1783), .B(n1784), .Z(n37376) );
  NANDN U2695 ( .A(n37370), .B(n42047), .Z(n1785) );
  NANDN U2696 ( .A(n37407), .B(n4067), .Z(n1786) );
  NAND U2697 ( .A(n1785), .B(n1786), .Z(n37418) );
  NANDN U2698 ( .A(n37445), .B(n4068), .Z(n1787) );
  NANDN U2699 ( .A(n37411), .B(n42115), .Z(n1788) );
  AND U2700 ( .A(n1787), .B(n1788), .Z(n37450) );
  NANDN U2701 ( .A(n37444), .B(n42047), .Z(n1789) );
  NANDN U2702 ( .A(n37481), .B(n4067), .Z(n1790) );
  NAND U2703 ( .A(n1789), .B(n1790), .Z(n37492) );
  NANDN U2704 ( .A(n37519), .B(n4068), .Z(n1791) );
  NANDN U2705 ( .A(n37482), .B(n42115), .Z(n1792) );
  AND U2706 ( .A(n1791), .B(n1792), .Z(n37524) );
  NANDN U2707 ( .A(n37518), .B(n42047), .Z(n1793) );
  NANDN U2708 ( .A(n37555), .B(n4067), .Z(n1794) );
  NAND U2709 ( .A(n1793), .B(n1794), .Z(n37566) );
  NANDN U2710 ( .A(n37596), .B(n4068), .Z(n1795) );
  NANDN U2711 ( .A(n37559), .B(n42115), .Z(n1796) );
  AND U2712 ( .A(n1795), .B(n1796), .Z(n37598) );
  NANDN U2713 ( .A(n37592), .B(n42047), .Z(n1797) );
  NANDN U2714 ( .A(n37629), .B(n4067), .Z(n1798) );
  NAND U2715 ( .A(n1797), .B(n1798), .Z(n37640) );
  NANDN U2716 ( .A(n37670), .B(n4068), .Z(n1799) );
  NANDN U2717 ( .A(n37630), .B(n42115), .Z(n1800) );
  AND U2718 ( .A(n1799), .B(n1800), .Z(n37672) );
  NANDN U2719 ( .A(n37666), .B(n42047), .Z(n1801) );
  NANDN U2720 ( .A(n37703), .B(n4067), .Z(n1802) );
  NAND U2721 ( .A(n1801), .B(n1802), .Z(n37714) );
  NANDN U2722 ( .A(n37744), .B(n4068), .Z(n1803) );
  NANDN U2723 ( .A(n37707), .B(n42115), .Z(n1804) );
  AND U2724 ( .A(n1803), .B(n1804), .Z(n37746) );
  NANDN U2725 ( .A(n37740), .B(n42047), .Z(n1805) );
  NANDN U2726 ( .A(n37777), .B(n4067), .Z(n1806) );
  NAND U2727 ( .A(n1805), .B(n1806), .Z(n37788) );
  NANDN U2728 ( .A(n37818), .B(n4068), .Z(n1807) );
  NANDN U2729 ( .A(n37778), .B(n42115), .Z(n1808) );
  AND U2730 ( .A(n1807), .B(n1808), .Z(n37820) );
  NANDN U2731 ( .A(n37814), .B(n42047), .Z(n1809) );
  NANDN U2732 ( .A(n37851), .B(n4067), .Z(n1810) );
  NAND U2733 ( .A(n1809), .B(n1810), .Z(n37862) );
  NANDN U2734 ( .A(n37889), .B(n4068), .Z(n1811) );
  NANDN U2735 ( .A(n37855), .B(n42115), .Z(n1812) );
  AND U2736 ( .A(n1811), .B(n1812), .Z(n37894) );
  NANDN U2737 ( .A(n37888), .B(n42047), .Z(n1813) );
  NANDN U2738 ( .A(n37925), .B(n4067), .Z(n1814) );
  NAND U2739 ( .A(n1813), .B(n1814), .Z(n37936) );
  NANDN U2740 ( .A(n37963), .B(n4068), .Z(n1815) );
  NANDN U2741 ( .A(n37929), .B(n42115), .Z(n1816) );
  AND U2742 ( .A(n1815), .B(n1816), .Z(n37968) );
  NANDN U2743 ( .A(n37962), .B(n42047), .Z(n1817) );
  NANDN U2744 ( .A(n37999), .B(n4067), .Z(n1818) );
  NAND U2745 ( .A(n1817), .B(n1818), .Z(n38010) );
  NANDN U2746 ( .A(n38040), .B(n4068), .Z(n1819) );
  NANDN U2747 ( .A(n38003), .B(n42115), .Z(n1820) );
  AND U2748 ( .A(n1819), .B(n1820), .Z(n38042) );
  NANDN U2749 ( .A(n38036), .B(n42047), .Z(n1821) );
  NANDN U2750 ( .A(n38073), .B(n4067), .Z(n1822) );
  NAND U2751 ( .A(n1821), .B(n1822), .Z(n38084) );
  NANDN U2752 ( .A(n38114), .B(n4068), .Z(n1823) );
  NANDN U2753 ( .A(n38077), .B(n42115), .Z(n1824) );
  AND U2754 ( .A(n1823), .B(n1824), .Z(n38116) );
  NANDN U2755 ( .A(n38110), .B(n42047), .Z(n1825) );
  NANDN U2756 ( .A(n38147), .B(n4067), .Z(n1826) );
  NAND U2757 ( .A(n1825), .B(n1826), .Z(n38158) );
  NANDN U2758 ( .A(n38188), .B(n4068), .Z(n1827) );
  NANDN U2759 ( .A(n38151), .B(n42115), .Z(n1828) );
  AND U2760 ( .A(n1827), .B(n1828), .Z(n38190) );
  NANDN U2761 ( .A(n38184), .B(n42047), .Z(n1829) );
  NANDN U2762 ( .A(n38221), .B(n4067), .Z(n1830) );
  NAND U2763 ( .A(n1829), .B(n1830), .Z(n38232) );
  NANDN U2764 ( .A(n38262), .B(n4068), .Z(n1831) );
  NANDN U2765 ( .A(n38225), .B(n42115), .Z(n1832) );
  AND U2766 ( .A(n1831), .B(n1832), .Z(n38264) );
  NANDN U2767 ( .A(n38258), .B(n42047), .Z(n1833) );
  NANDN U2768 ( .A(n38295), .B(n4067), .Z(n1834) );
  NAND U2769 ( .A(n1833), .B(n1834), .Z(n38306) );
  NANDN U2770 ( .A(n38333), .B(n4068), .Z(n1835) );
  NANDN U2771 ( .A(n38296), .B(n42115), .Z(n1836) );
  AND U2772 ( .A(n1835), .B(n1836), .Z(n38338) );
  NANDN U2773 ( .A(n38332), .B(n42047), .Z(n1837) );
  NANDN U2774 ( .A(n38369), .B(n4067), .Z(n1838) );
  NAND U2775 ( .A(n1837), .B(n1838), .Z(n38380) );
  NANDN U2776 ( .A(n38407), .B(n4068), .Z(n1839) );
  NANDN U2777 ( .A(n38373), .B(n42115), .Z(n1840) );
  AND U2778 ( .A(n1839), .B(n1840), .Z(n38412) );
  NANDN U2779 ( .A(n38406), .B(n42047), .Z(n1841) );
  NANDN U2780 ( .A(n38443), .B(n4067), .Z(n1842) );
  NAND U2781 ( .A(n1841), .B(n1842), .Z(n38454) );
  NANDN U2782 ( .A(n38481), .B(n4068), .Z(n1843) );
  NANDN U2783 ( .A(n38447), .B(n42115), .Z(n1844) );
  AND U2784 ( .A(n1843), .B(n1844), .Z(n38486) );
  NANDN U2785 ( .A(n38480), .B(n42047), .Z(n1845) );
  NANDN U2786 ( .A(n38517), .B(n4067), .Z(n1846) );
  NAND U2787 ( .A(n1845), .B(n1846), .Z(n38528) );
  NANDN U2788 ( .A(n38558), .B(n4068), .Z(n1847) );
  NANDN U2789 ( .A(n38518), .B(n42115), .Z(n1848) );
  AND U2790 ( .A(n1847), .B(n1848), .Z(n38560) );
  NANDN U2791 ( .A(n38554), .B(n42047), .Z(n1849) );
  NANDN U2792 ( .A(n38591), .B(n4067), .Z(n1850) );
  NAND U2793 ( .A(n1849), .B(n1850), .Z(n38602) );
  NANDN U2794 ( .A(n38629), .B(n4068), .Z(n1851) );
  NANDN U2795 ( .A(n38595), .B(n42115), .Z(n1852) );
  AND U2796 ( .A(n1851), .B(n1852), .Z(n38634) );
  NANDN U2797 ( .A(n38628), .B(n42047), .Z(n1853) );
  NANDN U2798 ( .A(n38665), .B(n4067), .Z(n1854) );
  NAND U2799 ( .A(n1853), .B(n1854), .Z(n38676) );
  NANDN U2800 ( .A(n38706), .B(n4068), .Z(n1855) );
  NANDN U2801 ( .A(n38669), .B(n42115), .Z(n1856) );
  AND U2802 ( .A(n1855), .B(n1856), .Z(n38708) );
  NANDN U2803 ( .A(n38702), .B(n42047), .Z(n1857) );
  NANDN U2804 ( .A(n38739), .B(n4067), .Z(n1858) );
  NAND U2805 ( .A(n1857), .B(n1858), .Z(n38750) );
  NANDN U2806 ( .A(n38780), .B(n4068), .Z(n1859) );
  NANDN U2807 ( .A(n38743), .B(n42115), .Z(n1860) );
  AND U2808 ( .A(n1859), .B(n1860), .Z(n38782) );
  NANDN U2809 ( .A(n38776), .B(n42047), .Z(n1861) );
  NANDN U2810 ( .A(n38813), .B(n4067), .Z(n1862) );
  NAND U2811 ( .A(n1861), .B(n1862), .Z(n38824) );
  NANDN U2812 ( .A(n38854), .B(n4068), .Z(n1863) );
  NANDN U2813 ( .A(n38817), .B(n42115), .Z(n1864) );
  AND U2814 ( .A(n1863), .B(n1864), .Z(n38856) );
  NANDN U2815 ( .A(n38850), .B(n42047), .Z(n1865) );
  NANDN U2816 ( .A(n38887), .B(n4067), .Z(n1866) );
  NAND U2817 ( .A(n1865), .B(n1866), .Z(n38898) );
  NANDN U2818 ( .A(n38928), .B(n4068), .Z(n1867) );
  NANDN U2819 ( .A(n38891), .B(n42115), .Z(n1868) );
  AND U2820 ( .A(n1867), .B(n1868), .Z(n38930) );
  NANDN U2821 ( .A(n38924), .B(n42047), .Z(n1869) );
  NANDN U2822 ( .A(n38961), .B(n4067), .Z(n1870) );
  NAND U2823 ( .A(n1869), .B(n1870), .Z(n38972) );
  NANDN U2824 ( .A(n39002), .B(n4068), .Z(n1871) );
  NANDN U2825 ( .A(n38962), .B(n42115), .Z(n1872) );
  AND U2826 ( .A(n1871), .B(n1872), .Z(n39004) );
  NANDN U2827 ( .A(n38998), .B(n42047), .Z(n1873) );
  NANDN U2828 ( .A(n39035), .B(n4067), .Z(n1874) );
  NAND U2829 ( .A(n1873), .B(n1874), .Z(n39046) );
  NANDN U2830 ( .A(n39076), .B(n4068), .Z(n1875) );
  NANDN U2831 ( .A(n39039), .B(n42115), .Z(n1876) );
  AND U2832 ( .A(n1875), .B(n1876), .Z(n39078) );
  NANDN U2833 ( .A(n39072), .B(n42047), .Z(n1877) );
  NANDN U2834 ( .A(n39109), .B(n4067), .Z(n1878) );
  NAND U2835 ( .A(n1877), .B(n1878), .Z(n39120) );
  NANDN U2836 ( .A(n39147), .B(n4068), .Z(n1879) );
  NANDN U2837 ( .A(n39110), .B(n42115), .Z(n1880) );
  AND U2838 ( .A(n1879), .B(n1880), .Z(n39152) );
  NANDN U2839 ( .A(n39146), .B(n42047), .Z(n1881) );
  NANDN U2840 ( .A(n39183), .B(n4067), .Z(n1882) );
  NAND U2841 ( .A(n1881), .B(n1882), .Z(n39194) );
  NANDN U2842 ( .A(n39224), .B(n4068), .Z(n1883) );
  NANDN U2843 ( .A(n39184), .B(n42115), .Z(n1884) );
  AND U2844 ( .A(n1883), .B(n1884), .Z(n39226) );
  NANDN U2845 ( .A(n39220), .B(n42047), .Z(n1885) );
  NANDN U2846 ( .A(n39257), .B(n4067), .Z(n1886) );
  NAND U2847 ( .A(n1885), .B(n1886), .Z(n39268) );
  NANDN U2848 ( .A(n39298), .B(n4068), .Z(n1887) );
  NANDN U2849 ( .A(n39258), .B(n42115), .Z(n1888) );
  AND U2850 ( .A(n1887), .B(n1888), .Z(n39300) );
  NANDN U2851 ( .A(n39294), .B(n42047), .Z(n1889) );
  NANDN U2852 ( .A(n39331), .B(n4067), .Z(n1890) );
  NAND U2853 ( .A(n1889), .B(n1890), .Z(n39342) );
  NANDN U2854 ( .A(n39372), .B(n4068), .Z(n1891) );
  NANDN U2855 ( .A(n39332), .B(n42115), .Z(n1892) );
  AND U2856 ( .A(n1891), .B(n1892), .Z(n39374) );
  NANDN U2857 ( .A(n39368), .B(n42047), .Z(n1893) );
  NANDN U2858 ( .A(n39405), .B(n4067), .Z(n1894) );
  NAND U2859 ( .A(n1893), .B(n1894), .Z(n39416) );
  NANDN U2860 ( .A(n39446), .B(n4068), .Z(n1895) );
  NANDN U2861 ( .A(n39409), .B(n42115), .Z(n1896) );
  AND U2862 ( .A(n1895), .B(n1896), .Z(n39448) );
  NANDN U2863 ( .A(n39442), .B(n42047), .Z(n1897) );
  NANDN U2864 ( .A(n39479), .B(n4067), .Z(n1898) );
  NAND U2865 ( .A(n1897), .B(n1898), .Z(n39490) );
  NANDN U2866 ( .A(n39520), .B(n4068), .Z(n1899) );
  NANDN U2867 ( .A(n39483), .B(n42115), .Z(n1900) );
  AND U2868 ( .A(n1899), .B(n1900), .Z(n39522) );
  NANDN U2869 ( .A(n39516), .B(n42047), .Z(n1901) );
  NANDN U2870 ( .A(n39553), .B(n4067), .Z(n1902) );
  NAND U2871 ( .A(n1901), .B(n1902), .Z(n39564) );
  NANDN U2872 ( .A(n39594), .B(n4068), .Z(n1903) );
  NANDN U2873 ( .A(n39557), .B(n42115), .Z(n1904) );
  AND U2874 ( .A(n1903), .B(n1904), .Z(n39596) );
  NANDN U2875 ( .A(n39590), .B(n42047), .Z(n1905) );
  NANDN U2876 ( .A(n39627), .B(n4067), .Z(n1906) );
  NAND U2877 ( .A(n1905), .B(n1906), .Z(n39638) );
  NANDN U2878 ( .A(n39665), .B(n4068), .Z(n1907) );
  NANDN U2879 ( .A(n39631), .B(n42115), .Z(n1908) );
  AND U2880 ( .A(n1907), .B(n1908), .Z(n39670) );
  NANDN U2881 ( .A(n39664), .B(n42047), .Z(n1909) );
  NANDN U2882 ( .A(n39701), .B(n4067), .Z(n1910) );
  NAND U2883 ( .A(n1909), .B(n1910), .Z(n39712) );
  NANDN U2884 ( .A(n39742), .B(n4068), .Z(n1911) );
  NANDN U2885 ( .A(n39705), .B(n42115), .Z(n1912) );
  AND U2886 ( .A(n1911), .B(n1912), .Z(n39744) );
  NANDN U2887 ( .A(n39738), .B(n42047), .Z(n1913) );
  NANDN U2888 ( .A(n39775), .B(n4067), .Z(n1914) );
  NAND U2889 ( .A(n1913), .B(n1914), .Z(n39786) );
  NANDN U2890 ( .A(n39813), .B(n4068), .Z(n1915) );
  NANDN U2891 ( .A(n39779), .B(n42115), .Z(n1916) );
  AND U2892 ( .A(n1915), .B(n1916), .Z(n39818) );
  NANDN U2893 ( .A(n39812), .B(n42047), .Z(n1917) );
  NANDN U2894 ( .A(n39849), .B(n4067), .Z(n1918) );
  NAND U2895 ( .A(n1917), .B(n1918), .Z(n39860) );
  NANDN U2896 ( .A(n39890), .B(n4068), .Z(n1919) );
  NANDN U2897 ( .A(n39853), .B(n42115), .Z(n1920) );
  AND U2898 ( .A(n1919), .B(n1920), .Z(n39892) );
  NANDN U2899 ( .A(n39886), .B(n42047), .Z(n1921) );
  NANDN U2900 ( .A(n39923), .B(n4067), .Z(n1922) );
  NAND U2901 ( .A(n1921), .B(n1922), .Z(n39934) );
  NANDN U2902 ( .A(n39964), .B(n4068), .Z(n1923) );
  NANDN U2903 ( .A(n39924), .B(n42115), .Z(n1924) );
  AND U2904 ( .A(n1923), .B(n1924), .Z(n39966) );
  NANDN U2905 ( .A(n39960), .B(n42047), .Z(n1925) );
  NANDN U2906 ( .A(n39997), .B(n4067), .Z(n1926) );
  NAND U2907 ( .A(n1925), .B(n1926), .Z(n40008) );
  NANDN U2908 ( .A(n40035), .B(n4068), .Z(n1927) );
  NANDN U2909 ( .A(n39998), .B(n42115), .Z(n1928) );
  AND U2910 ( .A(n1927), .B(n1928), .Z(n40040) );
  NANDN U2911 ( .A(n40034), .B(n42047), .Z(n1929) );
  NANDN U2912 ( .A(n40071), .B(n4067), .Z(n1930) );
  NAND U2913 ( .A(n1929), .B(n1930), .Z(n40082) );
  NANDN U2914 ( .A(n40112), .B(n4068), .Z(n1931) );
  NANDN U2915 ( .A(n40072), .B(n42115), .Z(n1932) );
  AND U2916 ( .A(n1931), .B(n1932), .Z(n40114) );
  NANDN U2917 ( .A(n40108), .B(n42047), .Z(n1933) );
  NANDN U2918 ( .A(n40145), .B(n4067), .Z(n1934) );
  NAND U2919 ( .A(n1933), .B(n1934), .Z(n40156) );
  NANDN U2920 ( .A(n40186), .B(n4068), .Z(n1935) );
  NANDN U2921 ( .A(n40149), .B(n42115), .Z(n1936) );
  AND U2922 ( .A(n1935), .B(n1936), .Z(n40188) );
  NANDN U2923 ( .A(n40182), .B(n42047), .Z(n1937) );
  NANDN U2924 ( .A(n40219), .B(n4067), .Z(n1938) );
  NAND U2925 ( .A(n1937), .B(n1938), .Z(n40230) );
  NANDN U2926 ( .A(n40260), .B(n4068), .Z(n1939) );
  NANDN U2927 ( .A(n40223), .B(n42115), .Z(n1940) );
  AND U2928 ( .A(n1939), .B(n1940), .Z(n40262) );
  NANDN U2929 ( .A(n40256), .B(n42047), .Z(n1941) );
  NANDN U2930 ( .A(n40293), .B(n4067), .Z(n1942) );
  NAND U2931 ( .A(n1941), .B(n1942), .Z(n40304) );
  NANDN U2932 ( .A(n40334), .B(n4068), .Z(n1943) );
  NANDN U2933 ( .A(n40294), .B(n42115), .Z(n1944) );
  AND U2934 ( .A(n1943), .B(n1944), .Z(n40336) );
  NANDN U2935 ( .A(n40330), .B(n42047), .Z(n1945) );
  NANDN U2936 ( .A(n40367), .B(n4067), .Z(n1946) );
  NAND U2937 ( .A(n1945), .B(n1946), .Z(n40378) );
  NANDN U2938 ( .A(n40408), .B(n4068), .Z(n1947) );
  NANDN U2939 ( .A(n40368), .B(n42115), .Z(n1948) );
  AND U2940 ( .A(n1947), .B(n1948), .Z(n40410) );
  NANDN U2941 ( .A(n40404), .B(n42047), .Z(n1949) );
  NANDN U2942 ( .A(n40441), .B(n4067), .Z(n1950) );
  NAND U2943 ( .A(n1949), .B(n1950), .Z(n40452) );
  NANDN U2944 ( .A(n40482), .B(n4068), .Z(n1951) );
  NANDN U2945 ( .A(n40445), .B(n42115), .Z(n1952) );
  AND U2946 ( .A(n1951), .B(n1952), .Z(n40484) );
  NANDN U2947 ( .A(n40478), .B(n42047), .Z(n1953) );
  NANDN U2948 ( .A(n40515), .B(n4067), .Z(n1954) );
  NAND U2949 ( .A(n1953), .B(n1954), .Z(n40526) );
  NANDN U2950 ( .A(n40556), .B(n4068), .Z(n1955) );
  NANDN U2951 ( .A(n40519), .B(n42115), .Z(n1956) );
  AND U2952 ( .A(n1955), .B(n1956), .Z(n40558) );
  NANDN U2953 ( .A(n40552), .B(n42047), .Z(n1957) );
  NANDN U2954 ( .A(n40589), .B(n4067), .Z(n1958) );
  NAND U2955 ( .A(n1957), .B(n1958), .Z(n40600) );
  NANDN U2956 ( .A(n40630), .B(n4068), .Z(n1959) );
  NANDN U2957 ( .A(n40593), .B(n42115), .Z(n1960) );
  AND U2958 ( .A(n1959), .B(n1960), .Z(n40632) );
  NANDN U2959 ( .A(n40626), .B(n42047), .Z(n1961) );
  NANDN U2960 ( .A(n40663), .B(n4067), .Z(n1962) );
  NAND U2961 ( .A(n1961), .B(n1962), .Z(n40674) );
  NANDN U2962 ( .A(n40704), .B(n4068), .Z(n1963) );
  NANDN U2963 ( .A(n40664), .B(n42115), .Z(n1964) );
  AND U2964 ( .A(n1963), .B(n1964), .Z(n40706) );
  NANDN U2965 ( .A(n40700), .B(n42047), .Z(n1965) );
  NANDN U2966 ( .A(n40737), .B(n4067), .Z(n1966) );
  NAND U2967 ( .A(n1965), .B(n1966), .Z(n40748) );
  NANDN U2968 ( .A(n40775), .B(n4068), .Z(n1967) );
  NANDN U2969 ( .A(n40738), .B(n42115), .Z(n1968) );
  AND U2970 ( .A(n1967), .B(n1968), .Z(n40780) );
  NANDN U2971 ( .A(n40774), .B(n42047), .Z(n1969) );
  NANDN U2972 ( .A(n40811), .B(n4067), .Z(n1970) );
  NAND U2973 ( .A(n1969), .B(n1970), .Z(n40822) );
  NANDN U2974 ( .A(n40849), .B(n4068), .Z(n1971) );
  NANDN U2975 ( .A(n40815), .B(n42115), .Z(n1972) );
  AND U2976 ( .A(n1971), .B(n1972), .Z(n40854) );
  NANDN U2977 ( .A(n40848), .B(n42047), .Z(n1973) );
  NANDN U2978 ( .A(n40885), .B(n4067), .Z(n1974) );
  NAND U2979 ( .A(n1973), .B(n1974), .Z(n40896) );
  NANDN U2980 ( .A(n40926), .B(n4068), .Z(n1975) );
  NANDN U2981 ( .A(n40886), .B(n42115), .Z(n1976) );
  AND U2982 ( .A(n1975), .B(n1976), .Z(n40928) );
  NANDN U2983 ( .A(n40922), .B(n42047), .Z(n1977) );
  NANDN U2984 ( .A(n40959), .B(n4067), .Z(n1978) );
  NAND U2985 ( .A(n1977), .B(n1978), .Z(n40970) );
  NANDN U2986 ( .A(n41000), .B(n4068), .Z(n1979) );
  NANDN U2987 ( .A(n40960), .B(n42115), .Z(n1980) );
  AND U2988 ( .A(n1979), .B(n1980), .Z(n41002) );
  NANDN U2989 ( .A(n40996), .B(n42047), .Z(n1981) );
  NANDN U2990 ( .A(n41033), .B(n4067), .Z(n1982) );
  NAND U2991 ( .A(n1981), .B(n1982), .Z(n41044) );
  NANDN U2992 ( .A(n41071), .B(n4068), .Z(n1983) );
  NANDN U2993 ( .A(n41034), .B(n42115), .Z(n1984) );
  AND U2994 ( .A(n1983), .B(n1984), .Z(n41076) );
  NANDN U2995 ( .A(n41070), .B(n42047), .Z(n1985) );
  NANDN U2996 ( .A(n41107), .B(n4067), .Z(n1986) );
  NAND U2997 ( .A(n1985), .B(n1986), .Z(n41118) );
  NANDN U2998 ( .A(n41148), .B(n4068), .Z(n1987) );
  NANDN U2999 ( .A(n41108), .B(n42115), .Z(n1988) );
  AND U3000 ( .A(n1987), .B(n1988), .Z(n41150) );
  NANDN U3001 ( .A(n41144), .B(n42047), .Z(n1989) );
  NANDN U3002 ( .A(n41181), .B(n4067), .Z(n1990) );
  NAND U3003 ( .A(n1989), .B(n1990), .Z(n41192) );
  NANDN U3004 ( .A(n41219), .B(n4068), .Z(n1991) );
  NANDN U3005 ( .A(n41185), .B(n42115), .Z(n1992) );
  AND U3006 ( .A(n1991), .B(n1992), .Z(n41224) );
  NANDN U3007 ( .A(n41218), .B(n42047), .Z(n1993) );
  NANDN U3008 ( .A(n41255), .B(n4067), .Z(n1994) );
  NAND U3009 ( .A(n1993), .B(n1994), .Z(n41266) );
  NANDN U3010 ( .A(n41293), .B(n4068), .Z(n1995) );
  NANDN U3011 ( .A(n41259), .B(n42115), .Z(n1996) );
  AND U3012 ( .A(n1995), .B(n1996), .Z(n41298) );
  NANDN U3013 ( .A(n41292), .B(n42047), .Z(n1997) );
  NANDN U3014 ( .A(n41329), .B(n4067), .Z(n1998) );
  NAND U3015 ( .A(n1997), .B(n1998), .Z(n41340) );
  NANDN U3016 ( .A(n41367), .B(n4068), .Z(n1999) );
  NANDN U3017 ( .A(n41333), .B(n42115), .Z(n2000) );
  AND U3018 ( .A(n1999), .B(n2000), .Z(n41372) );
  NANDN U3019 ( .A(n41366), .B(n42047), .Z(n2001) );
  NANDN U3020 ( .A(n41403), .B(n4067), .Z(n2002) );
  NAND U3021 ( .A(n2001), .B(n2002), .Z(n41414) );
  NANDN U3022 ( .A(n41444), .B(n4068), .Z(n2003) );
  NANDN U3023 ( .A(n41407), .B(n42115), .Z(n2004) );
  AND U3024 ( .A(n2003), .B(n2004), .Z(n41446) );
  NANDN U3025 ( .A(n41440), .B(n42047), .Z(n2005) );
  NANDN U3026 ( .A(n41477), .B(n4067), .Z(n2006) );
  NAND U3027 ( .A(n2005), .B(n2006), .Z(n41488) );
  NANDN U3028 ( .A(n41518), .B(n4068), .Z(n2007) );
  NANDN U3029 ( .A(n41481), .B(n42115), .Z(n2008) );
  AND U3030 ( .A(n2007), .B(n2008), .Z(n41520) );
  NANDN U3031 ( .A(n41514), .B(n42047), .Z(n2009) );
  NANDN U3032 ( .A(n41551), .B(n4067), .Z(n2010) );
  NAND U3033 ( .A(n2009), .B(n2010), .Z(n41562) );
  NANDN U3034 ( .A(n41592), .B(n4068), .Z(n2011) );
  NANDN U3035 ( .A(n41555), .B(n42115), .Z(n2012) );
  AND U3036 ( .A(n2011), .B(n2012), .Z(n41594) );
  NANDN U3037 ( .A(n41588), .B(n42047), .Z(n2013) );
  NANDN U3038 ( .A(n41625), .B(n4067), .Z(n2014) );
  NAND U3039 ( .A(n2013), .B(n2014), .Z(n41636) );
  NANDN U3040 ( .A(n41666), .B(n4068), .Z(n2015) );
  NANDN U3041 ( .A(n41626), .B(n42115), .Z(n2016) );
  AND U3042 ( .A(n2015), .B(n2016), .Z(n41668) );
  NANDN U3043 ( .A(n41662), .B(n42047), .Z(n2017) );
  NANDN U3044 ( .A(n41699), .B(n4067), .Z(n2018) );
  NAND U3045 ( .A(n2017), .B(n2018), .Z(n41710) );
  NANDN U3046 ( .A(n41737), .B(n4068), .Z(n2019) );
  NANDN U3047 ( .A(n41700), .B(n42115), .Z(n2020) );
  AND U3048 ( .A(n2019), .B(n2020), .Z(n41742) );
  NANDN U3049 ( .A(n41736), .B(n42047), .Z(n2021) );
  NANDN U3050 ( .A(n41773), .B(n4067), .Z(n2022) );
  NAND U3051 ( .A(n2021), .B(n2022), .Z(n41784) );
  NANDN U3052 ( .A(n41811), .B(n4068), .Z(n2023) );
  NANDN U3053 ( .A(n41777), .B(n42115), .Z(n2024) );
  AND U3054 ( .A(n2023), .B(n2024), .Z(n41816) );
  NANDN U3055 ( .A(n41810), .B(n42047), .Z(n2025) );
  NANDN U3056 ( .A(n41847), .B(n4067), .Z(n2026) );
  NAND U3057 ( .A(n2025), .B(n2026), .Z(n41858) );
  OR U3058 ( .A(n4064), .B(n4330), .Z(n2027) );
  NANDN U3059 ( .A(n4303), .B(n42047), .Z(n2028) );
  AND U3060 ( .A(n2027), .B(n2028), .Z(n4336) );
  XOR U3061 ( .A(n41929), .B(n41928), .Z(n41930) );
  XOR U3062 ( .A(n41963), .B(n41962), .Z(n41964) );
  XOR U3063 ( .A(n42016), .B(n42015), .Z(n42017) );
  XNOR U3064 ( .A(n42058), .B(n42057), .Z(n42042) );
  XOR U3065 ( .A(n41919), .B(n41918), .Z(n41910) );
  XOR U3066 ( .A(n42022), .B(n42021), .Z(n42023) );
  XOR U3067 ( .A(n42103), .B(n42102), .Z(n42104) );
  NANDN U3068 ( .A(n4268), .B(n4267), .Z(n2029) );
  NANDN U3069 ( .A(n4265), .B(n4266), .Z(n2030) );
  AND U3070 ( .A(n2029), .B(n2030), .Z(n4297) );
  XOR U3071 ( .A(n41957), .B(n41956), .Z(n41958) );
  XOR U3072 ( .A(n42136), .B(n42135), .Z(n42137) );
  XOR U3073 ( .A(b[7]), .B(a[1023]), .Z(n42160) );
  XOR U3074 ( .A(n42177), .B(n42178), .Z(n42180) );
  NANDN U3075 ( .A(n4403), .B(n4068), .Z(n2031) );
  NANDN U3076 ( .A(n4367), .B(n42115), .Z(n2032) );
  AND U3077 ( .A(n2031), .B(n2032), .Z(n4392) );
  NANDN U3078 ( .A(n4485), .B(n4068), .Z(n2033) );
  NANDN U3079 ( .A(n4437), .B(n42115), .Z(n2034) );
  AND U3080 ( .A(n2033), .B(n2034), .Z(n4487) );
  NANDN U3081 ( .A(n4481), .B(n42047), .Z(n2035) );
  NANDN U3082 ( .A(n4513), .B(n4067), .Z(n2036) );
  NAND U3083 ( .A(n2035), .B(n2036), .Z(n4524) );
  NANDN U3084 ( .A(n4554), .B(n4068), .Z(n2037) );
  NANDN U3085 ( .A(n4514), .B(n42115), .Z(n2038) );
  AND U3086 ( .A(n2037), .B(n2038), .Z(n4556) );
  NANDN U3087 ( .A(n4550), .B(n42047), .Z(n2039) );
  NANDN U3088 ( .A(n4587), .B(n4067), .Z(n2040) );
  NAND U3089 ( .A(n2039), .B(n2040), .Z(n4598) );
  NANDN U3090 ( .A(n4628), .B(n4068), .Z(n2041) );
  NANDN U3091 ( .A(n4588), .B(n42115), .Z(n2042) );
  AND U3092 ( .A(n2041), .B(n2042), .Z(n4630) );
  NANDN U3093 ( .A(n4624), .B(n42047), .Z(n2043) );
  NANDN U3094 ( .A(n4661), .B(n4067), .Z(n2044) );
  NAND U3095 ( .A(n2043), .B(n2044), .Z(n4672) );
  NANDN U3096 ( .A(n4702), .B(n4068), .Z(n2045) );
  NANDN U3097 ( .A(n4665), .B(n42115), .Z(n2046) );
  AND U3098 ( .A(n2045), .B(n2046), .Z(n4704) );
  NANDN U3099 ( .A(n4698), .B(n42047), .Z(n2047) );
  NANDN U3100 ( .A(n4735), .B(n4067), .Z(n2048) );
  NAND U3101 ( .A(n2047), .B(n2048), .Z(n4746) );
  NANDN U3102 ( .A(n4776), .B(n4068), .Z(n2049) );
  NANDN U3103 ( .A(n4736), .B(n42115), .Z(n2050) );
  AND U3104 ( .A(n2049), .B(n2050), .Z(n4778) );
  NANDN U3105 ( .A(n4772), .B(n42047), .Z(n2051) );
  NANDN U3106 ( .A(n4809), .B(n4067), .Z(n2052) );
  NAND U3107 ( .A(n2051), .B(n2052), .Z(n4820) );
  NANDN U3108 ( .A(n4847), .B(n4068), .Z(n2053) );
  NANDN U3109 ( .A(n4813), .B(n42115), .Z(n2054) );
  AND U3110 ( .A(n2053), .B(n2054), .Z(n4852) );
  NANDN U3111 ( .A(n4846), .B(n42047), .Z(n2055) );
  NANDN U3112 ( .A(n4883), .B(n4067), .Z(n2056) );
  NAND U3113 ( .A(n2055), .B(n2056), .Z(n4894) );
  NANDN U3114 ( .A(n4924), .B(n4068), .Z(n2057) );
  NANDN U3115 ( .A(n4884), .B(n42115), .Z(n2058) );
  AND U3116 ( .A(n2057), .B(n2058), .Z(n4926) );
  NANDN U3117 ( .A(n4920), .B(n42047), .Z(n2059) );
  NANDN U3118 ( .A(n4957), .B(n4067), .Z(n2060) );
  NAND U3119 ( .A(n2059), .B(n2060), .Z(n4968) );
  NANDN U3120 ( .A(n4998), .B(n4068), .Z(n2061) );
  NANDN U3121 ( .A(n4958), .B(n42115), .Z(n2062) );
  AND U3122 ( .A(n2061), .B(n2062), .Z(n5000) );
  NANDN U3123 ( .A(n4994), .B(n42047), .Z(n2063) );
  NANDN U3124 ( .A(n5031), .B(n4067), .Z(n2064) );
  NAND U3125 ( .A(n2063), .B(n2064), .Z(n5042) );
  NANDN U3126 ( .A(n5069), .B(n4068), .Z(n2065) );
  NANDN U3127 ( .A(n5035), .B(n42115), .Z(n2066) );
  AND U3128 ( .A(n2065), .B(n2066), .Z(n5074) );
  NANDN U3129 ( .A(n5068), .B(n42047), .Z(n2067) );
  NANDN U3130 ( .A(n5105), .B(n4067), .Z(n2068) );
  NAND U3131 ( .A(n2067), .B(n2068), .Z(n5116) );
  NANDN U3132 ( .A(n5146), .B(n4068), .Z(n2069) );
  NANDN U3133 ( .A(n5106), .B(n42115), .Z(n2070) );
  AND U3134 ( .A(n2069), .B(n2070), .Z(n5148) );
  NANDN U3135 ( .A(n5142), .B(n42047), .Z(n2071) );
  NANDN U3136 ( .A(n5179), .B(n4067), .Z(n2072) );
  NAND U3137 ( .A(n2071), .B(n2072), .Z(n5190) );
  NANDN U3138 ( .A(n5220), .B(n4068), .Z(n2073) );
  NANDN U3139 ( .A(n5183), .B(n42115), .Z(n2074) );
  AND U3140 ( .A(n2073), .B(n2074), .Z(n5222) );
  NANDN U3141 ( .A(n5216), .B(n42047), .Z(n2075) );
  NANDN U3142 ( .A(n5253), .B(n4067), .Z(n2076) );
  NAND U3143 ( .A(n2075), .B(n2076), .Z(n5264) );
  NANDN U3144 ( .A(n5294), .B(n4068), .Z(n2077) );
  NANDN U3145 ( .A(n5254), .B(n42115), .Z(n2078) );
  AND U3146 ( .A(n2077), .B(n2078), .Z(n5296) );
  NANDN U3147 ( .A(n5290), .B(n42047), .Z(n2079) );
  NANDN U3148 ( .A(n5327), .B(n4067), .Z(n2080) );
  NAND U3149 ( .A(n2079), .B(n2080), .Z(n5338) );
  NANDN U3150 ( .A(n5365), .B(n4068), .Z(n2081) );
  NANDN U3151 ( .A(n5331), .B(n42115), .Z(n2082) );
  AND U3152 ( .A(n2081), .B(n2082), .Z(n5370) );
  NANDN U3153 ( .A(n5364), .B(n42047), .Z(n2083) );
  NANDN U3154 ( .A(n5401), .B(n4067), .Z(n2084) );
  NAND U3155 ( .A(n2083), .B(n2084), .Z(n5412) );
  NANDN U3156 ( .A(n5442), .B(n4068), .Z(n2085) );
  NANDN U3157 ( .A(n5405), .B(n42115), .Z(n2086) );
  AND U3158 ( .A(n2085), .B(n2086), .Z(n5444) );
  NANDN U3159 ( .A(n5438), .B(n42047), .Z(n2087) );
  NANDN U3160 ( .A(n5475), .B(n4067), .Z(n2088) );
  NAND U3161 ( .A(n2087), .B(n2088), .Z(n5486) );
  NANDN U3162 ( .A(n5516), .B(n4068), .Z(n2089) );
  NANDN U3163 ( .A(n5476), .B(n42115), .Z(n2090) );
  AND U3164 ( .A(n2089), .B(n2090), .Z(n5518) );
  NANDN U3165 ( .A(n5512), .B(n42047), .Z(n2091) );
  NANDN U3166 ( .A(n5549), .B(n4067), .Z(n2092) );
  NAND U3167 ( .A(n2091), .B(n2092), .Z(n5560) );
  NANDN U3168 ( .A(n5590), .B(n4068), .Z(n2093) );
  NANDN U3169 ( .A(n5553), .B(n42115), .Z(n2094) );
  AND U3170 ( .A(n2093), .B(n2094), .Z(n5592) );
  NANDN U3171 ( .A(n5586), .B(n42047), .Z(n2095) );
  NANDN U3172 ( .A(n5623), .B(n4067), .Z(n2096) );
  NAND U3173 ( .A(n2095), .B(n2096), .Z(n5634) );
  NANDN U3174 ( .A(n5661), .B(n4068), .Z(n2097) );
  NANDN U3175 ( .A(n5627), .B(n42115), .Z(n2098) );
  AND U3176 ( .A(n2097), .B(n2098), .Z(n5666) );
  NANDN U3177 ( .A(n5660), .B(n42047), .Z(n2099) );
  NANDN U3178 ( .A(n5697), .B(n4067), .Z(n2100) );
  NAND U3179 ( .A(n2099), .B(n2100), .Z(n5708) );
  NANDN U3180 ( .A(n5735), .B(n4068), .Z(n2101) );
  NANDN U3181 ( .A(n5701), .B(n42115), .Z(n2102) );
  AND U3182 ( .A(n2101), .B(n2102), .Z(n5740) );
  NANDN U3183 ( .A(n5734), .B(n42047), .Z(n2103) );
  NANDN U3184 ( .A(n5771), .B(n4067), .Z(n2104) );
  NAND U3185 ( .A(n2103), .B(n2104), .Z(n5782) );
  NANDN U3186 ( .A(n5812), .B(n4068), .Z(n2105) );
  NANDN U3187 ( .A(n5775), .B(n42115), .Z(n2106) );
  AND U3188 ( .A(n2105), .B(n2106), .Z(n5814) );
  NANDN U3189 ( .A(n5808), .B(n42047), .Z(n2107) );
  NANDN U3190 ( .A(n5845), .B(n4067), .Z(n2108) );
  NAND U3191 ( .A(n2107), .B(n2108), .Z(n5856) );
  NANDN U3192 ( .A(n5886), .B(n4068), .Z(n2109) );
  NANDN U3193 ( .A(n5849), .B(n42115), .Z(n2110) );
  AND U3194 ( .A(n2109), .B(n2110), .Z(n5888) );
  NANDN U3195 ( .A(n5882), .B(n42047), .Z(n2111) );
  NANDN U3196 ( .A(n5919), .B(n4067), .Z(n2112) );
  NAND U3197 ( .A(n2111), .B(n2112), .Z(n5930) );
  NANDN U3198 ( .A(n5957), .B(n4068), .Z(n2113) );
  NANDN U3199 ( .A(n5923), .B(n42115), .Z(n2114) );
  AND U3200 ( .A(n2113), .B(n2114), .Z(n5962) );
  NANDN U3201 ( .A(n5956), .B(n42047), .Z(n2115) );
  NANDN U3202 ( .A(n5993), .B(n4067), .Z(n2116) );
  NAND U3203 ( .A(n2115), .B(n2116), .Z(n6004) );
  NANDN U3204 ( .A(n6034), .B(n4068), .Z(n2117) );
  NANDN U3205 ( .A(n5997), .B(n42115), .Z(n2118) );
  AND U3206 ( .A(n2117), .B(n2118), .Z(n6036) );
  NANDN U3207 ( .A(n6030), .B(n42047), .Z(n2119) );
  NANDN U3208 ( .A(n6067), .B(n4067), .Z(n2120) );
  NAND U3209 ( .A(n2119), .B(n2120), .Z(n6078) );
  NANDN U3210 ( .A(n6108), .B(n4068), .Z(n2121) );
  NANDN U3211 ( .A(n6071), .B(n42115), .Z(n2122) );
  AND U3212 ( .A(n2121), .B(n2122), .Z(n6110) );
  NANDN U3213 ( .A(n6104), .B(n42047), .Z(n2123) );
  NANDN U3214 ( .A(n6141), .B(n4067), .Z(n2124) );
  NAND U3215 ( .A(n2123), .B(n2124), .Z(n6152) );
  NANDN U3216 ( .A(n6182), .B(n4068), .Z(n2125) );
  NANDN U3217 ( .A(n6142), .B(n42115), .Z(n2126) );
  AND U3218 ( .A(n2125), .B(n2126), .Z(n6184) );
  NANDN U3219 ( .A(n6178), .B(n42047), .Z(n2127) );
  NANDN U3220 ( .A(n6215), .B(n4067), .Z(n2128) );
  NAND U3221 ( .A(n2127), .B(n2128), .Z(n6226) );
  NANDN U3222 ( .A(n6256), .B(n4068), .Z(n2129) );
  NANDN U3223 ( .A(n6216), .B(n42115), .Z(n2130) );
  AND U3224 ( .A(n2129), .B(n2130), .Z(n6258) );
  NANDN U3225 ( .A(n6252), .B(n42047), .Z(n2131) );
  NANDN U3226 ( .A(n6289), .B(n4067), .Z(n2132) );
  NAND U3227 ( .A(n2131), .B(n2132), .Z(n6300) );
  NANDN U3228 ( .A(n6330), .B(n4068), .Z(n2133) );
  NANDN U3229 ( .A(n6293), .B(n42115), .Z(n2134) );
  AND U3230 ( .A(n2133), .B(n2134), .Z(n6332) );
  NANDN U3231 ( .A(n6326), .B(n42047), .Z(n2135) );
  NANDN U3232 ( .A(n6363), .B(n4067), .Z(n2136) );
  NAND U3233 ( .A(n2135), .B(n2136), .Z(n6374) );
  NANDN U3234 ( .A(n6404), .B(n4068), .Z(n2137) );
  NANDN U3235 ( .A(n6367), .B(n42115), .Z(n2138) );
  AND U3236 ( .A(n2137), .B(n2138), .Z(n6406) );
  NANDN U3237 ( .A(n6400), .B(n42047), .Z(n2139) );
  NANDN U3238 ( .A(n6437), .B(n4067), .Z(n2140) );
  NAND U3239 ( .A(n2139), .B(n2140), .Z(n6448) );
  NANDN U3240 ( .A(n6478), .B(n4068), .Z(n2141) );
  NANDN U3241 ( .A(n6438), .B(n42115), .Z(n2142) );
  AND U3242 ( .A(n2141), .B(n2142), .Z(n6480) );
  NANDN U3243 ( .A(n6474), .B(n42047), .Z(n2143) );
  NANDN U3244 ( .A(n6511), .B(n4067), .Z(n2144) );
  NAND U3245 ( .A(n2143), .B(n2144), .Z(n6522) );
  NANDN U3246 ( .A(n6552), .B(n4068), .Z(n2145) );
  NANDN U3247 ( .A(n6515), .B(n42115), .Z(n2146) );
  AND U3248 ( .A(n2145), .B(n2146), .Z(n6554) );
  NANDN U3249 ( .A(n6548), .B(n42047), .Z(n2147) );
  NANDN U3250 ( .A(n6585), .B(n4067), .Z(n2148) );
  NAND U3251 ( .A(n2147), .B(n2148), .Z(n6596) );
  NANDN U3252 ( .A(n6626), .B(n4068), .Z(n2149) );
  NANDN U3253 ( .A(n6589), .B(n42115), .Z(n2150) );
  AND U3254 ( .A(n2149), .B(n2150), .Z(n6628) );
  NANDN U3255 ( .A(n6622), .B(n42047), .Z(n2151) );
  NANDN U3256 ( .A(n6659), .B(n4067), .Z(n2152) );
  NAND U3257 ( .A(n2151), .B(n2152), .Z(n6670) );
  NANDN U3258 ( .A(n6700), .B(n4068), .Z(n2153) );
  NANDN U3259 ( .A(n6663), .B(n42115), .Z(n2154) );
  AND U3260 ( .A(n2153), .B(n2154), .Z(n6702) );
  NANDN U3261 ( .A(n6696), .B(n42047), .Z(n2155) );
  NANDN U3262 ( .A(n6733), .B(n4067), .Z(n2156) );
  NAND U3263 ( .A(n2155), .B(n2156), .Z(n6744) );
  NANDN U3264 ( .A(n6774), .B(n4068), .Z(n2157) );
  NANDN U3265 ( .A(n6734), .B(n42115), .Z(n2158) );
  AND U3266 ( .A(n2157), .B(n2158), .Z(n6776) );
  NANDN U3267 ( .A(n6770), .B(n42047), .Z(n2159) );
  NANDN U3268 ( .A(n6807), .B(n4067), .Z(n2160) );
  NAND U3269 ( .A(n2159), .B(n2160), .Z(n6818) );
  NANDN U3270 ( .A(n6845), .B(n4068), .Z(n2161) );
  NANDN U3271 ( .A(n6811), .B(n42115), .Z(n2162) );
  AND U3272 ( .A(n2161), .B(n2162), .Z(n6850) );
  NANDN U3273 ( .A(n6844), .B(n42047), .Z(n2163) );
  NANDN U3274 ( .A(n6881), .B(n4067), .Z(n2164) );
  NAND U3275 ( .A(n2163), .B(n2164), .Z(n6892) );
  NANDN U3276 ( .A(n6924), .B(n4068), .Z(n2165) );
  NANDN U3277 ( .A(n6885), .B(n42115), .Z(n2166) );
  AND U3278 ( .A(n2165), .B(n2166), .Z(n6929) );
  NANDN U3279 ( .A(n6923), .B(n42047), .Z(n2167) );
  NANDN U3280 ( .A(n6955), .B(n4067), .Z(n2168) );
  NAND U3281 ( .A(n2167), .B(n2168), .Z(n6966) );
  NANDN U3282 ( .A(n6996), .B(n4068), .Z(n2169) );
  NANDN U3283 ( .A(n6959), .B(n42115), .Z(n2170) );
  AND U3284 ( .A(n2169), .B(n2170), .Z(n6998) );
  NANDN U3285 ( .A(n6992), .B(n42047), .Z(n2171) );
  NANDN U3286 ( .A(n7034), .B(n4067), .Z(n2172) );
  NAND U3287 ( .A(n2171), .B(n2172), .Z(n7045) );
  NANDN U3288 ( .A(n7067), .B(n4068), .Z(n2173) );
  NANDN U3289 ( .A(n7035), .B(n42115), .Z(n2174) );
  AND U3290 ( .A(n2173), .B(n2174), .Z(n7072) );
  NANDN U3291 ( .A(n7066), .B(n42047), .Z(n2175) );
  NANDN U3292 ( .A(n7103), .B(n4067), .Z(n2176) );
  NAND U3293 ( .A(n2175), .B(n2176), .Z(n7114) );
  NANDN U3294 ( .A(n7144), .B(n4068), .Z(n2177) );
  NANDN U3295 ( .A(n7104), .B(n42115), .Z(n2178) );
  AND U3296 ( .A(n2177), .B(n2178), .Z(n7146) );
  NANDN U3297 ( .A(n7140), .B(n42047), .Z(n2179) );
  NANDN U3298 ( .A(n7177), .B(n4067), .Z(n2180) );
  NAND U3299 ( .A(n2179), .B(n2180), .Z(n7188) );
  NANDN U3300 ( .A(n7218), .B(n4068), .Z(n2181) );
  NANDN U3301 ( .A(n7178), .B(n42115), .Z(n2182) );
  AND U3302 ( .A(n2181), .B(n2182), .Z(n7220) );
  NANDN U3303 ( .A(n7214), .B(n42047), .Z(n2183) );
  NANDN U3304 ( .A(n7251), .B(n4067), .Z(n2184) );
  NAND U3305 ( .A(n2183), .B(n2184), .Z(n7262) );
  NANDN U3306 ( .A(n7292), .B(n4068), .Z(n2185) );
  NANDN U3307 ( .A(n7255), .B(n42115), .Z(n2186) );
  AND U3308 ( .A(n2185), .B(n2186), .Z(n7294) );
  NANDN U3309 ( .A(n7288), .B(n42047), .Z(n2187) );
  NANDN U3310 ( .A(n7325), .B(n4067), .Z(n2188) );
  NAND U3311 ( .A(n2187), .B(n2188), .Z(n7336) );
  NANDN U3312 ( .A(n7363), .B(n4068), .Z(n2189) );
  NANDN U3313 ( .A(n7329), .B(n42115), .Z(n2190) );
  AND U3314 ( .A(n2189), .B(n2190), .Z(n7368) );
  NANDN U3315 ( .A(n7362), .B(n42047), .Z(n2191) );
  NANDN U3316 ( .A(n7399), .B(n4067), .Z(n2192) );
  NAND U3317 ( .A(n2191), .B(n2192), .Z(n7410) );
  NANDN U3318 ( .A(n7440), .B(n4068), .Z(n2193) );
  NANDN U3319 ( .A(n7403), .B(n42115), .Z(n2194) );
  AND U3320 ( .A(n2193), .B(n2194), .Z(n7442) );
  NANDN U3321 ( .A(n7436), .B(n42047), .Z(n2195) );
  NANDN U3322 ( .A(n7473), .B(n4067), .Z(n2196) );
  NAND U3323 ( .A(n2195), .B(n2196), .Z(n7484) );
  NANDN U3324 ( .A(n7514), .B(n4068), .Z(n2197) );
  NANDN U3325 ( .A(n7477), .B(n42115), .Z(n2198) );
  AND U3326 ( .A(n2197), .B(n2198), .Z(n7516) );
  NANDN U3327 ( .A(n7510), .B(n42047), .Z(n2199) );
  NANDN U3328 ( .A(n7547), .B(n4067), .Z(n2200) );
  NAND U3329 ( .A(n2199), .B(n2200), .Z(n7558) );
  NANDN U3330 ( .A(n7588), .B(n4068), .Z(n2201) );
  NANDN U3331 ( .A(n7551), .B(n42115), .Z(n2202) );
  AND U3332 ( .A(n2201), .B(n2202), .Z(n7590) );
  NANDN U3333 ( .A(n7584), .B(n42047), .Z(n2203) );
  NANDN U3334 ( .A(n7621), .B(n4067), .Z(n2204) );
  NAND U3335 ( .A(n2203), .B(n2204), .Z(n7632) );
  NANDN U3336 ( .A(n7662), .B(n4068), .Z(n2205) );
  NANDN U3337 ( .A(n7625), .B(n42115), .Z(n2206) );
  AND U3338 ( .A(n2205), .B(n2206), .Z(n7664) );
  NANDN U3339 ( .A(n7658), .B(n42047), .Z(n2207) );
  NANDN U3340 ( .A(n7695), .B(n4067), .Z(n2208) );
  NAND U3341 ( .A(n2207), .B(n2208), .Z(n7706) );
  NANDN U3342 ( .A(n7736), .B(n4068), .Z(n2209) );
  NANDN U3343 ( .A(n7699), .B(n42115), .Z(n2210) );
  AND U3344 ( .A(n2209), .B(n2210), .Z(n7738) );
  NANDN U3345 ( .A(n7732), .B(n42047), .Z(n2211) );
  NANDN U3346 ( .A(n7769), .B(n4067), .Z(n2212) );
  NAND U3347 ( .A(n2211), .B(n2212), .Z(n7780) );
  NANDN U3348 ( .A(n7810), .B(n4068), .Z(n2213) );
  NANDN U3349 ( .A(n7773), .B(n42115), .Z(n2214) );
  AND U3350 ( .A(n2213), .B(n2214), .Z(n7812) );
  NANDN U3351 ( .A(n7806), .B(n42047), .Z(n2215) );
  NANDN U3352 ( .A(n7843), .B(n4067), .Z(n2216) );
  NAND U3353 ( .A(n2215), .B(n2216), .Z(n7854) );
  NANDN U3354 ( .A(n7881), .B(n4068), .Z(n2217) );
  NANDN U3355 ( .A(n7847), .B(n42115), .Z(n2218) );
  AND U3356 ( .A(n2217), .B(n2218), .Z(n7886) );
  NANDN U3357 ( .A(n7880), .B(n42047), .Z(n2219) );
  NANDN U3358 ( .A(n7917), .B(n4067), .Z(n2220) );
  NAND U3359 ( .A(n2219), .B(n2220), .Z(n7928) );
  NANDN U3360 ( .A(n7958), .B(n4068), .Z(n2221) );
  NANDN U3361 ( .A(n7921), .B(n42115), .Z(n2222) );
  AND U3362 ( .A(n2221), .B(n2222), .Z(n7960) );
  NANDN U3363 ( .A(n7954), .B(n42047), .Z(n2223) );
  NANDN U3364 ( .A(n7991), .B(n4067), .Z(n2224) );
  NAND U3365 ( .A(n2223), .B(n2224), .Z(n8002) );
  NANDN U3366 ( .A(n8032), .B(n4068), .Z(n2225) );
  NANDN U3367 ( .A(n7995), .B(n42115), .Z(n2226) );
  AND U3368 ( .A(n2225), .B(n2226), .Z(n8034) );
  NANDN U3369 ( .A(n8028), .B(n42047), .Z(n2227) );
  NANDN U3370 ( .A(n8065), .B(n4067), .Z(n2228) );
  NAND U3371 ( .A(n2227), .B(n2228), .Z(n8076) );
  NANDN U3372 ( .A(n8103), .B(n4068), .Z(n2229) );
  NANDN U3373 ( .A(n8069), .B(n42115), .Z(n2230) );
  AND U3374 ( .A(n2229), .B(n2230), .Z(n8108) );
  NANDN U3375 ( .A(n8102), .B(n42047), .Z(n2231) );
  NANDN U3376 ( .A(n8139), .B(n4067), .Z(n2232) );
  NAND U3377 ( .A(n2231), .B(n2232), .Z(n8150) );
  NANDN U3378 ( .A(n8177), .B(n4068), .Z(n2233) );
  NANDN U3379 ( .A(n8140), .B(n42115), .Z(n2234) );
  AND U3380 ( .A(n2233), .B(n2234), .Z(n8182) );
  NANDN U3381 ( .A(n8176), .B(n42047), .Z(n2235) );
  NANDN U3382 ( .A(n8213), .B(n4067), .Z(n2236) );
  NAND U3383 ( .A(n2235), .B(n2236), .Z(n8224) );
  NANDN U3384 ( .A(n8251), .B(n4068), .Z(n2237) );
  NANDN U3385 ( .A(n8217), .B(n42115), .Z(n2238) );
  AND U3386 ( .A(n2237), .B(n2238), .Z(n8256) );
  NANDN U3387 ( .A(n8250), .B(n42047), .Z(n2239) );
  NANDN U3388 ( .A(n8287), .B(n4067), .Z(n2240) );
  NAND U3389 ( .A(n2239), .B(n2240), .Z(n8298) );
  NANDN U3390 ( .A(n8328), .B(n4068), .Z(n2241) );
  NANDN U3391 ( .A(n8291), .B(n42115), .Z(n2242) );
  AND U3392 ( .A(n2241), .B(n2242), .Z(n8330) );
  NANDN U3393 ( .A(n8324), .B(n42047), .Z(n2243) );
  NANDN U3394 ( .A(n8361), .B(n4067), .Z(n2244) );
  NAND U3395 ( .A(n2243), .B(n2244), .Z(n8372) );
  NANDN U3396 ( .A(n8402), .B(n4068), .Z(n2245) );
  NANDN U3397 ( .A(n8365), .B(n42115), .Z(n2246) );
  AND U3398 ( .A(n2245), .B(n2246), .Z(n8404) );
  NANDN U3399 ( .A(n8398), .B(n42047), .Z(n2247) );
  NANDN U3400 ( .A(n8435), .B(n4067), .Z(n2248) );
  NAND U3401 ( .A(n2247), .B(n2248), .Z(n8446) );
  NANDN U3402 ( .A(n8476), .B(n4068), .Z(n2249) );
  NANDN U3403 ( .A(n8439), .B(n42115), .Z(n2250) );
  AND U3404 ( .A(n2249), .B(n2250), .Z(n8478) );
  NANDN U3405 ( .A(n8472), .B(n42047), .Z(n2251) );
  NANDN U3406 ( .A(n8509), .B(n4067), .Z(n2252) );
  NAND U3407 ( .A(n2251), .B(n2252), .Z(n8520) );
  NANDN U3408 ( .A(n8547), .B(n4068), .Z(n2253) );
  NANDN U3409 ( .A(n8513), .B(n42115), .Z(n2254) );
  AND U3410 ( .A(n2253), .B(n2254), .Z(n8552) );
  NANDN U3411 ( .A(n8546), .B(n42047), .Z(n2255) );
  NANDN U3412 ( .A(n8583), .B(n4067), .Z(n2256) );
  NAND U3413 ( .A(n2255), .B(n2256), .Z(n8594) );
  NANDN U3414 ( .A(n8624), .B(n4068), .Z(n2257) );
  NANDN U3415 ( .A(n8587), .B(n42115), .Z(n2258) );
  AND U3416 ( .A(n2257), .B(n2258), .Z(n8626) );
  NANDN U3417 ( .A(n8620), .B(n42047), .Z(n2259) );
  NANDN U3418 ( .A(n8657), .B(n4067), .Z(n2260) );
  NAND U3419 ( .A(n2259), .B(n2260), .Z(n8668) );
  NANDN U3420 ( .A(n8695), .B(n4068), .Z(n2261) );
  NANDN U3421 ( .A(n8661), .B(n42115), .Z(n2262) );
  AND U3422 ( .A(n2261), .B(n2262), .Z(n8700) );
  NANDN U3423 ( .A(n8694), .B(n42047), .Z(n2263) );
  NANDN U3424 ( .A(n8731), .B(n4067), .Z(n2264) );
  NAND U3425 ( .A(n2263), .B(n2264), .Z(n8742) );
  NANDN U3426 ( .A(n8772), .B(n4068), .Z(n2265) );
  NANDN U3427 ( .A(n8732), .B(n42115), .Z(n2266) );
  AND U3428 ( .A(n2265), .B(n2266), .Z(n8774) );
  NANDN U3429 ( .A(n8768), .B(n42047), .Z(n2267) );
  NANDN U3430 ( .A(n8805), .B(n4067), .Z(n2268) );
  NAND U3431 ( .A(n2267), .B(n2268), .Z(n8816) );
  NANDN U3432 ( .A(n8843), .B(n4068), .Z(n2269) );
  NANDN U3433 ( .A(n8806), .B(n42115), .Z(n2270) );
  AND U3434 ( .A(n2269), .B(n2270), .Z(n8848) );
  NANDN U3435 ( .A(n8842), .B(n42047), .Z(n2271) );
  NANDN U3436 ( .A(n8879), .B(n4067), .Z(n2272) );
  NAND U3437 ( .A(n2271), .B(n2272), .Z(n8890) );
  NANDN U3438 ( .A(n8920), .B(n4068), .Z(n2273) );
  NANDN U3439 ( .A(n8883), .B(n42115), .Z(n2274) );
  AND U3440 ( .A(n2273), .B(n2274), .Z(n8922) );
  NANDN U3441 ( .A(n8916), .B(n42047), .Z(n2275) );
  NANDN U3442 ( .A(n8953), .B(n4067), .Z(n2276) );
  NAND U3443 ( .A(n2275), .B(n2276), .Z(n8964) );
  NANDN U3444 ( .A(n8994), .B(n4068), .Z(n2277) );
  NANDN U3445 ( .A(n8957), .B(n42115), .Z(n2278) );
  AND U3446 ( .A(n2277), .B(n2278), .Z(n8996) );
  NANDN U3447 ( .A(n8990), .B(n42047), .Z(n2279) );
  NANDN U3448 ( .A(n9032), .B(n4067), .Z(n2280) );
  NAND U3449 ( .A(n2279), .B(n2280), .Z(n9043) );
  NANDN U3450 ( .A(n9068), .B(n4068), .Z(n2281) );
  NANDN U3451 ( .A(n9033), .B(n42115), .Z(n2282) );
  AND U3452 ( .A(n2281), .B(n2282), .Z(n9070) );
  NANDN U3453 ( .A(n9064), .B(n42047), .Z(n2283) );
  NANDN U3454 ( .A(n9101), .B(n4067), .Z(n2284) );
  NAND U3455 ( .A(n2283), .B(n2284), .Z(n9112) );
  NANDN U3456 ( .A(n9142), .B(n4068), .Z(n2285) );
  NANDN U3457 ( .A(n9105), .B(n42115), .Z(n2286) );
  AND U3458 ( .A(n2285), .B(n2286), .Z(n9144) );
  NANDN U3459 ( .A(n9138), .B(n42047), .Z(n2287) );
  NANDN U3460 ( .A(n9175), .B(n4067), .Z(n2288) );
  NAND U3461 ( .A(n2287), .B(n2288), .Z(n9186) );
  NANDN U3462 ( .A(n9216), .B(n4068), .Z(n2289) );
  NANDN U3463 ( .A(n9179), .B(n42115), .Z(n2290) );
  AND U3464 ( .A(n2289), .B(n2290), .Z(n9218) );
  NANDN U3465 ( .A(n9212), .B(n42047), .Z(n2291) );
  NANDN U3466 ( .A(n9249), .B(n4067), .Z(n2292) );
  NAND U3467 ( .A(n2291), .B(n2292), .Z(n9260) );
  NANDN U3468 ( .A(n9290), .B(n4068), .Z(n2293) );
  NANDN U3469 ( .A(n9253), .B(n42115), .Z(n2294) );
  AND U3470 ( .A(n2293), .B(n2294), .Z(n9292) );
  NANDN U3471 ( .A(n9286), .B(n42047), .Z(n2295) );
  NANDN U3472 ( .A(n9323), .B(n4067), .Z(n2296) );
  NAND U3473 ( .A(n2295), .B(n2296), .Z(n9334) );
  NANDN U3474 ( .A(n9364), .B(n4068), .Z(n2297) );
  NANDN U3475 ( .A(n9327), .B(n42115), .Z(n2298) );
  AND U3476 ( .A(n2297), .B(n2298), .Z(n9366) );
  NANDN U3477 ( .A(n9360), .B(n42047), .Z(n2299) );
  NANDN U3478 ( .A(n9397), .B(n4067), .Z(n2300) );
  NAND U3479 ( .A(n2299), .B(n2300), .Z(n9408) );
  NANDN U3480 ( .A(n9435), .B(n4068), .Z(n2301) );
  NANDN U3481 ( .A(n9398), .B(n42115), .Z(n2302) );
  AND U3482 ( .A(n2301), .B(n2302), .Z(n9440) );
  NANDN U3483 ( .A(n9434), .B(n42047), .Z(n2303) );
  NANDN U3484 ( .A(n9471), .B(n4067), .Z(n2304) );
  NAND U3485 ( .A(n2303), .B(n2304), .Z(n9482) );
  NANDN U3486 ( .A(n9509), .B(n4068), .Z(n2305) );
  NANDN U3487 ( .A(n9475), .B(n42115), .Z(n2306) );
  AND U3488 ( .A(n2305), .B(n2306), .Z(n9514) );
  NANDN U3489 ( .A(n9508), .B(n42047), .Z(n2307) );
  NANDN U3490 ( .A(n9545), .B(n4067), .Z(n2308) );
  NAND U3491 ( .A(n2307), .B(n2308), .Z(n9556) );
  NANDN U3492 ( .A(n9586), .B(n4068), .Z(n2309) );
  NANDN U3493 ( .A(n9546), .B(n42115), .Z(n2310) );
  AND U3494 ( .A(n2309), .B(n2310), .Z(n9588) );
  NANDN U3495 ( .A(n9582), .B(n42047), .Z(n2311) );
  NANDN U3496 ( .A(n9619), .B(n4067), .Z(n2312) );
  NAND U3497 ( .A(n2311), .B(n2312), .Z(n9630) );
  NANDN U3498 ( .A(n9657), .B(n4068), .Z(n2313) );
  NANDN U3499 ( .A(n9623), .B(n42115), .Z(n2314) );
  AND U3500 ( .A(n2313), .B(n2314), .Z(n9662) );
  NANDN U3501 ( .A(n9656), .B(n42047), .Z(n2315) );
  NANDN U3502 ( .A(n9698), .B(n4067), .Z(n2316) );
  NAND U3503 ( .A(n2315), .B(n2316), .Z(n9709) );
  NANDN U3504 ( .A(n9734), .B(n4068), .Z(n2317) );
  NANDN U3505 ( .A(n9702), .B(n42115), .Z(n2318) );
  AND U3506 ( .A(n2317), .B(n2318), .Z(n9736) );
  NANDN U3507 ( .A(n9730), .B(n42047), .Z(n2319) );
  NANDN U3508 ( .A(n9767), .B(n4067), .Z(n2320) );
  NAND U3509 ( .A(n2319), .B(n2320), .Z(n9778) );
  NANDN U3510 ( .A(n9808), .B(n4068), .Z(n2321) );
  NANDN U3511 ( .A(n9771), .B(n42115), .Z(n2322) );
  AND U3512 ( .A(n2321), .B(n2322), .Z(n9810) );
  NANDN U3513 ( .A(n9804), .B(n42047), .Z(n2323) );
  NANDN U3514 ( .A(n9841), .B(n4067), .Z(n2324) );
  NAND U3515 ( .A(n2323), .B(n2324), .Z(n9852) );
  NANDN U3516 ( .A(n9882), .B(n4068), .Z(n2325) );
  NANDN U3517 ( .A(n9842), .B(n42115), .Z(n2326) );
  AND U3518 ( .A(n2325), .B(n2326), .Z(n9884) );
  NANDN U3519 ( .A(n9878), .B(n42047), .Z(n2327) );
  NANDN U3520 ( .A(n9915), .B(n4067), .Z(n2328) );
  NAND U3521 ( .A(n2327), .B(n2328), .Z(n9926) );
  NANDN U3522 ( .A(n9956), .B(n4068), .Z(n2329) );
  NANDN U3523 ( .A(n9919), .B(n42115), .Z(n2330) );
  AND U3524 ( .A(n2329), .B(n2330), .Z(n9958) );
  NANDN U3525 ( .A(n9952), .B(n42047), .Z(n2331) );
  NANDN U3526 ( .A(n9989), .B(n4067), .Z(n2332) );
  NAND U3527 ( .A(n2331), .B(n2332), .Z(n10000) );
  NANDN U3528 ( .A(n10030), .B(n4068), .Z(n2333) );
  NANDN U3529 ( .A(n9993), .B(n42115), .Z(n2334) );
  AND U3530 ( .A(n2333), .B(n2334), .Z(n10032) );
  NANDN U3531 ( .A(n10026), .B(n42047), .Z(n2335) );
  NANDN U3532 ( .A(n10063), .B(n4067), .Z(n2336) );
  NAND U3533 ( .A(n2335), .B(n2336), .Z(n10074) );
  NANDN U3534 ( .A(n10104), .B(n4068), .Z(n2337) );
  NANDN U3535 ( .A(n10067), .B(n42115), .Z(n2338) );
  AND U3536 ( .A(n2337), .B(n2338), .Z(n10106) );
  NANDN U3537 ( .A(n10100), .B(n42047), .Z(n2339) );
  NANDN U3538 ( .A(n10137), .B(n4067), .Z(n2340) );
  NAND U3539 ( .A(n2339), .B(n2340), .Z(n10148) );
  NANDN U3540 ( .A(n10175), .B(n4068), .Z(n2341) );
  NANDN U3541 ( .A(n10138), .B(n42115), .Z(n2342) );
  AND U3542 ( .A(n2341), .B(n2342), .Z(n10180) );
  NANDN U3543 ( .A(n10174), .B(n42047), .Z(n2343) );
  NANDN U3544 ( .A(n10211), .B(n4067), .Z(n2344) );
  NAND U3545 ( .A(n2343), .B(n2344), .Z(n10222) );
  NANDN U3546 ( .A(n10252), .B(n4068), .Z(n2345) );
  NANDN U3547 ( .A(n10215), .B(n42115), .Z(n2346) );
  AND U3548 ( .A(n2345), .B(n2346), .Z(n10254) );
  NANDN U3549 ( .A(n10248), .B(n42047), .Z(n2347) );
  NANDN U3550 ( .A(n10285), .B(n4067), .Z(n2348) );
  NAND U3551 ( .A(n2347), .B(n2348), .Z(n10296) );
  NANDN U3552 ( .A(n10326), .B(n4068), .Z(n2349) );
  NANDN U3553 ( .A(n10289), .B(n42115), .Z(n2350) );
  AND U3554 ( .A(n2349), .B(n2350), .Z(n10328) );
  NANDN U3555 ( .A(n10322), .B(n42047), .Z(n2351) );
  NANDN U3556 ( .A(n10359), .B(n4067), .Z(n2352) );
  NAND U3557 ( .A(n2351), .B(n2352), .Z(n10370) );
  NANDN U3558 ( .A(n10400), .B(n4068), .Z(n2353) );
  NANDN U3559 ( .A(n10363), .B(n42115), .Z(n2354) );
  AND U3560 ( .A(n2353), .B(n2354), .Z(n10402) );
  NANDN U3561 ( .A(n10396), .B(n42047), .Z(n2355) );
  NANDN U3562 ( .A(n10433), .B(n4067), .Z(n2356) );
  NAND U3563 ( .A(n2355), .B(n2356), .Z(n10444) );
  NANDN U3564 ( .A(n10474), .B(n4068), .Z(n2357) );
  NANDN U3565 ( .A(n10437), .B(n42115), .Z(n2358) );
  AND U3566 ( .A(n2357), .B(n2358), .Z(n10476) );
  NANDN U3567 ( .A(n10470), .B(n42047), .Z(n2359) );
  NANDN U3568 ( .A(n10507), .B(n4067), .Z(n2360) );
  NAND U3569 ( .A(n2359), .B(n2360), .Z(n10518) );
  NANDN U3570 ( .A(n10548), .B(n4068), .Z(n2361) );
  NANDN U3571 ( .A(n10511), .B(n42115), .Z(n2362) );
  AND U3572 ( .A(n2361), .B(n2362), .Z(n10550) );
  NANDN U3573 ( .A(n10544), .B(n42047), .Z(n2363) );
  NANDN U3574 ( .A(n10581), .B(n4067), .Z(n2364) );
  NAND U3575 ( .A(n2363), .B(n2364), .Z(n10592) );
  NANDN U3576 ( .A(n10619), .B(n4068), .Z(n2365) );
  NANDN U3577 ( .A(n10585), .B(n42115), .Z(n2366) );
  AND U3578 ( .A(n2365), .B(n2366), .Z(n10624) );
  NANDN U3579 ( .A(n10618), .B(n42047), .Z(n2367) );
  NANDN U3580 ( .A(n10655), .B(n4067), .Z(n2368) );
  NAND U3581 ( .A(n2367), .B(n2368), .Z(n10666) );
  NANDN U3582 ( .A(n10696), .B(n4068), .Z(n2369) );
  NANDN U3583 ( .A(n10656), .B(n42115), .Z(n2370) );
  AND U3584 ( .A(n2369), .B(n2370), .Z(n10698) );
  NANDN U3585 ( .A(n10692), .B(n42047), .Z(n2371) );
  NANDN U3586 ( .A(n10729), .B(n4067), .Z(n2372) );
  NAND U3587 ( .A(n2371), .B(n2372), .Z(n10740) );
  NANDN U3588 ( .A(n10770), .B(n4068), .Z(n2373) );
  NANDN U3589 ( .A(n10730), .B(n42115), .Z(n2374) );
  AND U3590 ( .A(n2373), .B(n2374), .Z(n10772) );
  NANDN U3591 ( .A(n10766), .B(n42047), .Z(n2375) );
  NANDN U3592 ( .A(n10803), .B(n4067), .Z(n2376) );
  NAND U3593 ( .A(n2375), .B(n2376), .Z(n10814) );
  NANDN U3594 ( .A(n10844), .B(n4068), .Z(n2377) );
  NANDN U3595 ( .A(n10807), .B(n42115), .Z(n2378) );
  AND U3596 ( .A(n2377), .B(n2378), .Z(n10846) );
  NANDN U3597 ( .A(n10840), .B(n42047), .Z(n2379) );
  NANDN U3598 ( .A(n10877), .B(n4067), .Z(n2380) );
  NAND U3599 ( .A(n2379), .B(n2380), .Z(n10888) );
  NANDN U3600 ( .A(n10918), .B(n4068), .Z(n2381) );
  NANDN U3601 ( .A(n10881), .B(n42115), .Z(n2382) );
  AND U3602 ( .A(n2381), .B(n2382), .Z(n10920) );
  NANDN U3603 ( .A(n10914), .B(n42047), .Z(n2383) );
  NANDN U3604 ( .A(n10951), .B(n4067), .Z(n2384) );
  NAND U3605 ( .A(n2383), .B(n2384), .Z(n10962) );
  NANDN U3606 ( .A(n10992), .B(n4068), .Z(n2385) );
  NANDN U3607 ( .A(n10955), .B(n42115), .Z(n2386) );
  AND U3608 ( .A(n2385), .B(n2386), .Z(n10994) );
  NANDN U3609 ( .A(n10988), .B(n42047), .Z(n2387) );
  NANDN U3610 ( .A(n11025), .B(n4067), .Z(n2388) );
  NAND U3611 ( .A(n2387), .B(n2388), .Z(n11036) );
  NANDN U3612 ( .A(n11066), .B(n4068), .Z(n2389) );
  NANDN U3613 ( .A(n11026), .B(n42115), .Z(n2390) );
  AND U3614 ( .A(n2389), .B(n2390), .Z(n11068) );
  NANDN U3615 ( .A(n11062), .B(n42047), .Z(n2391) );
  NANDN U3616 ( .A(n11099), .B(n4067), .Z(n2392) );
  NAND U3617 ( .A(n2391), .B(n2392), .Z(n11110) );
  NANDN U3618 ( .A(n11137), .B(n4068), .Z(n2393) );
  NANDN U3619 ( .A(n11100), .B(n42115), .Z(n2394) );
  AND U3620 ( .A(n2393), .B(n2394), .Z(n11142) );
  NANDN U3621 ( .A(n11136), .B(n42047), .Z(n2395) );
  NANDN U3622 ( .A(n11173), .B(n4067), .Z(n2396) );
  NAND U3623 ( .A(n2395), .B(n2396), .Z(n11184) );
  NANDN U3624 ( .A(n11214), .B(n4068), .Z(n2397) );
  NANDN U3625 ( .A(n11177), .B(n42115), .Z(n2398) );
  AND U3626 ( .A(n2397), .B(n2398), .Z(n11216) );
  NANDN U3627 ( .A(n11210), .B(n42047), .Z(n2399) );
  NANDN U3628 ( .A(n11247), .B(n4067), .Z(n2400) );
  NAND U3629 ( .A(n2399), .B(n2400), .Z(n11258) );
  NANDN U3630 ( .A(n11285), .B(n4068), .Z(n2401) );
  NANDN U3631 ( .A(n11251), .B(n42115), .Z(n2402) );
  AND U3632 ( .A(n2401), .B(n2402), .Z(n11290) );
  NANDN U3633 ( .A(n11284), .B(n42047), .Z(n2403) );
  NANDN U3634 ( .A(n11321), .B(n4067), .Z(n2404) );
  NAND U3635 ( .A(n2403), .B(n2404), .Z(n11332) );
  NANDN U3636 ( .A(n11362), .B(n4068), .Z(n2405) );
  NANDN U3637 ( .A(n11322), .B(n42115), .Z(n2406) );
  AND U3638 ( .A(n2405), .B(n2406), .Z(n11364) );
  NANDN U3639 ( .A(n11358), .B(n42047), .Z(n2407) );
  NANDN U3640 ( .A(n11395), .B(n4067), .Z(n2408) );
  NAND U3641 ( .A(n2407), .B(n2408), .Z(n11406) );
  NANDN U3642 ( .A(n11433), .B(n4068), .Z(n2409) );
  NANDN U3643 ( .A(n11396), .B(n42115), .Z(n2410) );
  AND U3644 ( .A(n2409), .B(n2410), .Z(n11438) );
  NANDN U3645 ( .A(n11432), .B(n42047), .Z(n2411) );
  NANDN U3646 ( .A(n11469), .B(n4067), .Z(n2412) );
  NAND U3647 ( .A(n2411), .B(n2412), .Z(n11480) );
  NANDN U3648 ( .A(n11510), .B(n4068), .Z(n2413) );
  NANDN U3649 ( .A(n11473), .B(n42115), .Z(n2414) );
  AND U3650 ( .A(n2413), .B(n2414), .Z(n11512) );
  NANDN U3651 ( .A(n11506), .B(n42047), .Z(n2415) );
  NANDN U3652 ( .A(n11543), .B(n4067), .Z(n2416) );
  NAND U3653 ( .A(n2415), .B(n2416), .Z(n11554) );
  NANDN U3654 ( .A(n11581), .B(n4068), .Z(n2417) );
  NANDN U3655 ( .A(n11547), .B(n42115), .Z(n2418) );
  AND U3656 ( .A(n2417), .B(n2418), .Z(n11586) );
  NANDN U3657 ( .A(n11580), .B(n42047), .Z(n2419) );
  NANDN U3658 ( .A(n11617), .B(n4067), .Z(n2420) );
  NAND U3659 ( .A(n2419), .B(n2420), .Z(n11628) );
  NANDN U3660 ( .A(n11655), .B(n4068), .Z(n2421) );
  NANDN U3661 ( .A(n11621), .B(n42115), .Z(n2422) );
  AND U3662 ( .A(n2421), .B(n2422), .Z(n11660) );
  NANDN U3663 ( .A(n11654), .B(n42047), .Z(n2423) );
  NANDN U3664 ( .A(n11691), .B(n4067), .Z(n2424) );
  NAND U3665 ( .A(n2423), .B(n2424), .Z(n11702) );
  NANDN U3666 ( .A(n11732), .B(n4068), .Z(n2425) );
  NANDN U3667 ( .A(n11695), .B(n42115), .Z(n2426) );
  AND U3668 ( .A(n2425), .B(n2426), .Z(n11734) );
  NANDN U3669 ( .A(n11728), .B(n42047), .Z(n2427) );
  NANDN U3670 ( .A(n11765), .B(n4067), .Z(n2428) );
  NAND U3671 ( .A(n2427), .B(n2428), .Z(n11776) );
  NANDN U3672 ( .A(n11803), .B(n4068), .Z(n2429) );
  NANDN U3673 ( .A(n11769), .B(n42115), .Z(n2430) );
  AND U3674 ( .A(n2429), .B(n2430), .Z(n11808) );
  NANDN U3675 ( .A(n11802), .B(n42047), .Z(n2431) );
  NANDN U3676 ( .A(n11839), .B(n4067), .Z(n2432) );
  NAND U3677 ( .A(n2431), .B(n2432), .Z(n11850) );
  NANDN U3678 ( .A(n11880), .B(n4068), .Z(n2433) );
  NANDN U3679 ( .A(n11843), .B(n42115), .Z(n2434) );
  AND U3680 ( .A(n2433), .B(n2434), .Z(n11882) );
  NANDN U3681 ( .A(n11876), .B(n42047), .Z(n2435) );
  NANDN U3682 ( .A(n11913), .B(n4067), .Z(n2436) );
  NAND U3683 ( .A(n2435), .B(n2436), .Z(n11924) );
  NANDN U3684 ( .A(n11954), .B(n4068), .Z(n2437) );
  NANDN U3685 ( .A(n11917), .B(n42115), .Z(n2438) );
  AND U3686 ( .A(n2437), .B(n2438), .Z(n11956) );
  NANDN U3687 ( .A(n11950), .B(n42047), .Z(n2439) );
  NANDN U3688 ( .A(n11987), .B(n4067), .Z(n2440) );
  NAND U3689 ( .A(n2439), .B(n2440), .Z(n11998) );
  NANDN U3690 ( .A(n12025), .B(n4068), .Z(n2441) );
  NANDN U3691 ( .A(n11991), .B(n42115), .Z(n2442) );
  AND U3692 ( .A(n2441), .B(n2442), .Z(n12030) );
  NANDN U3693 ( .A(n12024), .B(n42047), .Z(n2443) );
  NANDN U3694 ( .A(n12061), .B(n4067), .Z(n2444) );
  NAND U3695 ( .A(n2443), .B(n2444), .Z(n12072) );
  NANDN U3696 ( .A(n12099), .B(n4068), .Z(n2445) );
  NANDN U3697 ( .A(n12065), .B(n42115), .Z(n2446) );
  AND U3698 ( .A(n2445), .B(n2446), .Z(n12104) );
  NANDN U3699 ( .A(n12098), .B(n42047), .Z(n2447) );
  NANDN U3700 ( .A(n12135), .B(n4067), .Z(n2448) );
  NAND U3701 ( .A(n2447), .B(n2448), .Z(n12146) );
  NANDN U3702 ( .A(n12176), .B(n4068), .Z(n2449) );
  NANDN U3703 ( .A(n12139), .B(n42115), .Z(n2450) );
  AND U3704 ( .A(n2449), .B(n2450), .Z(n12178) );
  NANDN U3705 ( .A(n12172), .B(n42047), .Z(n2451) );
  NANDN U3706 ( .A(n12209), .B(n4067), .Z(n2452) );
  NAND U3707 ( .A(n2451), .B(n2452), .Z(n12220) );
  NANDN U3708 ( .A(n12250), .B(n4068), .Z(n2453) );
  NANDN U3709 ( .A(n12213), .B(n42115), .Z(n2454) );
  AND U3710 ( .A(n2453), .B(n2454), .Z(n12252) );
  NANDN U3711 ( .A(n12246), .B(n42047), .Z(n2455) );
  NANDN U3712 ( .A(n12283), .B(n4067), .Z(n2456) );
  NAND U3713 ( .A(n2455), .B(n2456), .Z(n12294) );
  NANDN U3714 ( .A(n12324), .B(n4068), .Z(n2457) );
  NANDN U3715 ( .A(n12284), .B(n42115), .Z(n2458) );
  AND U3716 ( .A(n2457), .B(n2458), .Z(n12326) );
  NANDN U3717 ( .A(n12320), .B(n42047), .Z(n2459) );
  NANDN U3718 ( .A(n12357), .B(n4067), .Z(n2460) );
  NAND U3719 ( .A(n2459), .B(n2460), .Z(n12368) );
  NANDN U3720 ( .A(n12395), .B(n4068), .Z(n2461) );
  NANDN U3721 ( .A(n12361), .B(n42115), .Z(n2462) );
  AND U3722 ( .A(n2461), .B(n2462), .Z(n12400) );
  NANDN U3723 ( .A(n12394), .B(n42047), .Z(n2463) );
  NANDN U3724 ( .A(n12431), .B(n4067), .Z(n2464) );
  NAND U3725 ( .A(n2463), .B(n2464), .Z(n12442) );
  NANDN U3726 ( .A(n12472), .B(n4068), .Z(n2465) );
  NANDN U3727 ( .A(n12435), .B(n42115), .Z(n2466) );
  AND U3728 ( .A(n2465), .B(n2466), .Z(n12474) );
  NANDN U3729 ( .A(n12468), .B(n42047), .Z(n2467) );
  NANDN U3730 ( .A(n12505), .B(n4067), .Z(n2468) );
  NAND U3731 ( .A(n2467), .B(n2468), .Z(n12516) );
  NANDN U3732 ( .A(n12546), .B(n4068), .Z(n2469) );
  NANDN U3733 ( .A(n12506), .B(n42115), .Z(n2470) );
  AND U3734 ( .A(n2469), .B(n2470), .Z(n12548) );
  NANDN U3735 ( .A(n12542), .B(n42047), .Z(n2471) );
  NANDN U3736 ( .A(n12579), .B(n4067), .Z(n2472) );
  NAND U3737 ( .A(n2471), .B(n2472), .Z(n12590) );
  NANDN U3738 ( .A(n12620), .B(n4068), .Z(n2473) );
  NANDN U3739 ( .A(n12580), .B(n42115), .Z(n2474) );
  AND U3740 ( .A(n2473), .B(n2474), .Z(n12622) );
  NANDN U3741 ( .A(n12616), .B(n42047), .Z(n2475) );
  NANDN U3742 ( .A(n12653), .B(n4067), .Z(n2476) );
  NAND U3743 ( .A(n2475), .B(n2476), .Z(n12664) );
  NANDN U3744 ( .A(n12694), .B(n4068), .Z(n2477) );
  NANDN U3745 ( .A(n12657), .B(n42115), .Z(n2478) );
  AND U3746 ( .A(n2477), .B(n2478), .Z(n12696) );
  NANDN U3747 ( .A(n12690), .B(n42047), .Z(n2479) );
  NANDN U3748 ( .A(n12727), .B(n4067), .Z(n2480) );
  NAND U3749 ( .A(n2479), .B(n2480), .Z(n12738) );
  NANDN U3750 ( .A(n12768), .B(n4068), .Z(n2481) );
  NANDN U3751 ( .A(n12731), .B(n42115), .Z(n2482) );
  AND U3752 ( .A(n2481), .B(n2482), .Z(n12770) );
  NANDN U3753 ( .A(n12764), .B(n42047), .Z(n2483) );
  NANDN U3754 ( .A(n12801), .B(n4067), .Z(n2484) );
  NAND U3755 ( .A(n2483), .B(n2484), .Z(n12812) );
  NANDN U3756 ( .A(n12842), .B(n4068), .Z(n2485) );
  NANDN U3757 ( .A(n12805), .B(n42115), .Z(n2486) );
  AND U3758 ( .A(n2485), .B(n2486), .Z(n12844) );
  NANDN U3759 ( .A(n12838), .B(n42047), .Z(n2487) );
  NANDN U3760 ( .A(n12875), .B(n4067), .Z(n2488) );
  NAND U3761 ( .A(n2487), .B(n2488), .Z(n12886) );
  NANDN U3762 ( .A(n12916), .B(n4068), .Z(n2489) );
  NANDN U3763 ( .A(n12879), .B(n42115), .Z(n2490) );
  AND U3764 ( .A(n2489), .B(n2490), .Z(n12918) );
  NANDN U3765 ( .A(n12912), .B(n42047), .Z(n2491) );
  NANDN U3766 ( .A(n12949), .B(n4067), .Z(n2492) );
  NAND U3767 ( .A(n2491), .B(n2492), .Z(n12960) );
  NANDN U3768 ( .A(n12990), .B(n4068), .Z(n2493) );
  NANDN U3769 ( .A(n12950), .B(n42115), .Z(n2494) );
  AND U3770 ( .A(n2493), .B(n2494), .Z(n12992) );
  NANDN U3771 ( .A(n12986), .B(n42047), .Z(n2495) );
  NANDN U3772 ( .A(n13023), .B(n4067), .Z(n2496) );
  NAND U3773 ( .A(n2495), .B(n2496), .Z(n13034) );
  NANDN U3774 ( .A(n13064), .B(n4068), .Z(n2497) );
  NANDN U3775 ( .A(n13024), .B(n42115), .Z(n2498) );
  AND U3776 ( .A(n2497), .B(n2498), .Z(n13066) );
  NANDN U3777 ( .A(n13060), .B(n42047), .Z(n2499) );
  NANDN U3778 ( .A(n13097), .B(n4067), .Z(n2500) );
  NAND U3779 ( .A(n2499), .B(n2500), .Z(n13108) );
  NANDN U3780 ( .A(n13138), .B(n4068), .Z(n2501) );
  NANDN U3781 ( .A(n13101), .B(n42115), .Z(n2502) );
  AND U3782 ( .A(n2501), .B(n2502), .Z(n13140) );
  NANDN U3783 ( .A(n13134), .B(n42047), .Z(n2503) );
  NANDN U3784 ( .A(n13171), .B(n4067), .Z(n2504) );
  NAND U3785 ( .A(n2503), .B(n2504), .Z(n13182) );
  NANDN U3786 ( .A(n13212), .B(n4068), .Z(n2505) );
  NANDN U3787 ( .A(n13175), .B(n42115), .Z(n2506) );
  AND U3788 ( .A(n2505), .B(n2506), .Z(n13214) );
  NANDN U3789 ( .A(n13208), .B(n42047), .Z(n2507) );
  NANDN U3790 ( .A(n13245), .B(n4067), .Z(n2508) );
  NAND U3791 ( .A(n2507), .B(n2508), .Z(n13256) );
  NANDN U3792 ( .A(n13286), .B(n4068), .Z(n2509) );
  NANDN U3793 ( .A(n13249), .B(n42115), .Z(n2510) );
  AND U3794 ( .A(n2509), .B(n2510), .Z(n13288) );
  NANDN U3795 ( .A(n13282), .B(n42047), .Z(n2511) );
  NANDN U3796 ( .A(n13319), .B(n4067), .Z(n2512) );
  NAND U3797 ( .A(n2511), .B(n2512), .Z(n13330) );
  NANDN U3798 ( .A(n13360), .B(n4068), .Z(n2513) );
  NANDN U3799 ( .A(n13320), .B(n42115), .Z(n2514) );
  AND U3800 ( .A(n2513), .B(n2514), .Z(n13362) );
  NANDN U3801 ( .A(n13356), .B(n42047), .Z(n2515) );
  NANDN U3802 ( .A(n13393), .B(n4067), .Z(n2516) );
  NAND U3803 ( .A(n2515), .B(n2516), .Z(n13404) );
  NANDN U3804 ( .A(n13431), .B(n4068), .Z(n2517) );
  NANDN U3805 ( .A(n13397), .B(n42115), .Z(n2518) );
  AND U3806 ( .A(n2517), .B(n2518), .Z(n13436) );
  NANDN U3807 ( .A(n13430), .B(n42047), .Z(n2519) );
  NANDN U3808 ( .A(n13467), .B(n4067), .Z(n2520) );
  NAND U3809 ( .A(n2519), .B(n2520), .Z(n13478) );
  NANDN U3810 ( .A(n13505), .B(n4068), .Z(n2521) );
  NANDN U3811 ( .A(n13471), .B(n42115), .Z(n2522) );
  AND U3812 ( .A(n2521), .B(n2522), .Z(n13510) );
  NANDN U3813 ( .A(n13504), .B(n42047), .Z(n2523) );
  NANDN U3814 ( .A(n13541), .B(n4067), .Z(n2524) );
  NAND U3815 ( .A(n2523), .B(n2524), .Z(n13552) );
  NANDN U3816 ( .A(n13582), .B(n4068), .Z(n2525) );
  NANDN U3817 ( .A(n13545), .B(n42115), .Z(n2526) );
  AND U3818 ( .A(n2525), .B(n2526), .Z(n13584) );
  NANDN U3819 ( .A(n13578), .B(n42047), .Z(n2527) );
  NANDN U3820 ( .A(n13615), .B(n4067), .Z(n2528) );
  NAND U3821 ( .A(n2527), .B(n2528), .Z(n13626) );
  NANDN U3822 ( .A(n13656), .B(n4068), .Z(n2529) );
  NANDN U3823 ( .A(n13619), .B(n42115), .Z(n2530) );
  AND U3824 ( .A(n2529), .B(n2530), .Z(n13658) );
  NANDN U3825 ( .A(n13652), .B(n42047), .Z(n2531) );
  NANDN U3826 ( .A(n13689), .B(n4067), .Z(n2532) );
  NAND U3827 ( .A(n2531), .B(n2532), .Z(n13700) );
  NANDN U3828 ( .A(n13727), .B(n4068), .Z(n2533) );
  NANDN U3829 ( .A(n13693), .B(n42115), .Z(n2534) );
  AND U3830 ( .A(n2533), .B(n2534), .Z(n13732) );
  NANDN U3831 ( .A(n13726), .B(n42047), .Z(n2535) );
  NANDN U3832 ( .A(n13763), .B(n4067), .Z(n2536) );
  NAND U3833 ( .A(n2535), .B(n2536), .Z(n13774) );
  NANDN U3834 ( .A(n13804), .B(n4068), .Z(n2537) );
  NANDN U3835 ( .A(n13767), .B(n42115), .Z(n2538) );
  AND U3836 ( .A(n2537), .B(n2538), .Z(n13806) );
  NANDN U3837 ( .A(n13800), .B(n42047), .Z(n2539) );
  NANDN U3838 ( .A(n13837), .B(n4067), .Z(n2540) );
  NAND U3839 ( .A(n2539), .B(n2540), .Z(n13848) );
  NANDN U3840 ( .A(n13878), .B(n4068), .Z(n2541) );
  NANDN U3841 ( .A(n13841), .B(n42115), .Z(n2542) );
  AND U3842 ( .A(n2541), .B(n2542), .Z(n13880) );
  NANDN U3843 ( .A(n13874), .B(n42047), .Z(n2543) );
  NANDN U3844 ( .A(n13911), .B(n4067), .Z(n2544) );
  NAND U3845 ( .A(n2543), .B(n2544), .Z(n13922) );
  NANDN U3846 ( .A(n13952), .B(n4068), .Z(n2545) );
  NANDN U3847 ( .A(n13915), .B(n42115), .Z(n2546) );
  AND U3848 ( .A(n2545), .B(n2546), .Z(n13954) );
  NANDN U3849 ( .A(n13948), .B(n42047), .Z(n2547) );
  NANDN U3850 ( .A(n13985), .B(n4067), .Z(n2548) );
  NAND U3851 ( .A(n2547), .B(n2548), .Z(n13996) );
  NANDN U3852 ( .A(n14026), .B(n4068), .Z(n2549) );
  NANDN U3853 ( .A(n13986), .B(n42115), .Z(n2550) );
  AND U3854 ( .A(n2549), .B(n2550), .Z(n14028) );
  NANDN U3855 ( .A(n14022), .B(n42047), .Z(n2551) );
  NANDN U3856 ( .A(n14059), .B(n4067), .Z(n2552) );
  NAND U3857 ( .A(n2551), .B(n2552), .Z(n14070) );
  NANDN U3858 ( .A(n14105), .B(n4068), .Z(n2553) );
  NANDN U3859 ( .A(n14063), .B(n42115), .Z(n2554) );
  AND U3860 ( .A(n2553), .B(n2554), .Z(n14107) );
  NANDN U3861 ( .A(n14101), .B(n42047), .Z(n2555) );
  NANDN U3862 ( .A(n14138), .B(n4067), .Z(n2556) );
  NAND U3863 ( .A(n2555), .B(n2556), .Z(n14149) );
  NANDN U3864 ( .A(n14174), .B(n4068), .Z(n2557) );
  NANDN U3865 ( .A(n14139), .B(n42115), .Z(n2558) );
  AND U3866 ( .A(n2557), .B(n2558), .Z(n14176) );
  NANDN U3867 ( .A(n14170), .B(n42047), .Z(n2559) );
  NANDN U3868 ( .A(n14207), .B(n4067), .Z(n2560) );
  NAND U3869 ( .A(n2559), .B(n2560), .Z(n14218) );
  NANDN U3870 ( .A(n14253), .B(n4068), .Z(n2561) );
  NANDN U3871 ( .A(n14211), .B(n42115), .Z(n2562) );
  AND U3872 ( .A(n2561), .B(n2562), .Z(n14255) );
  NANDN U3873 ( .A(n14249), .B(n42047), .Z(n2563) );
  NANDN U3874 ( .A(n14281), .B(n4067), .Z(n2564) );
  NAND U3875 ( .A(n2563), .B(n2564), .Z(n14292) );
  NANDN U3876 ( .A(n14319), .B(n4068), .Z(n2565) );
  NANDN U3877 ( .A(n14285), .B(n42115), .Z(n2566) );
  AND U3878 ( .A(n2565), .B(n2566), .Z(n14324) );
  NANDN U3879 ( .A(n14318), .B(n42047), .Z(n2567) );
  NANDN U3880 ( .A(n14355), .B(n4067), .Z(n2568) );
  NAND U3881 ( .A(n2567), .B(n2568), .Z(n14366) );
  NANDN U3882 ( .A(n14396), .B(n4068), .Z(n2569) );
  NANDN U3883 ( .A(n14359), .B(n42115), .Z(n2570) );
  AND U3884 ( .A(n2569), .B(n2570), .Z(n14398) );
  NANDN U3885 ( .A(n14392), .B(n42047), .Z(n2571) );
  NANDN U3886 ( .A(n14429), .B(n4067), .Z(n2572) );
  NAND U3887 ( .A(n2571), .B(n2572), .Z(n14440) );
  NANDN U3888 ( .A(n14470), .B(n4068), .Z(n2573) );
  NANDN U3889 ( .A(n14433), .B(n42115), .Z(n2574) );
  AND U3890 ( .A(n2573), .B(n2574), .Z(n14472) );
  NANDN U3891 ( .A(n14466), .B(n42047), .Z(n2575) );
  NANDN U3892 ( .A(n14503), .B(n4067), .Z(n2576) );
  NAND U3893 ( .A(n2575), .B(n2576), .Z(n14514) );
  NANDN U3894 ( .A(n14541), .B(n4068), .Z(n2577) );
  NANDN U3895 ( .A(n14504), .B(n42115), .Z(n2578) );
  AND U3896 ( .A(n2577), .B(n2578), .Z(n14546) );
  NANDN U3897 ( .A(n14540), .B(n42047), .Z(n2579) );
  NANDN U3898 ( .A(n14577), .B(n4067), .Z(n2580) );
  NAND U3899 ( .A(n2579), .B(n2580), .Z(n14588) );
  NANDN U3900 ( .A(n14618), .B(n4068), .Z(n2581) );
  NANDN U3901 ( .A(n14581), .B(n42115), .Z(n2582) );
  AND U3902 ( .A(n2581), .B(n2582), .Z(n14620) );
  NANDN U3903 ( .A(n14614), .B(n42047), .Z(n2583) );
  NANDN U3904 ( .A(n14651), .B(n4067), .Z(n2584) );
  NAND U3905 ( .A(n2583), .B(n2584), .Z(n14662) );
  NANDN U3906 ( .A(n14692), .B(n4068), .Z(n2585) );
  NANDN U3907 ( .A(n14655), .B(n42115), .Z(n2586) );
  AND U3908 ( .A(n2585), .B(n2586), .Z(n14694) );
  NANDN U3909 ( .A(n14688), .B(n42047), .Z(n2587) );
  NANDN U3910 ( .A(n14725), .B(n4067), .Z(n2588) );
  NAND U3911 ( .A(n2587), .B(n2588), .Z(n14736) );
  NANDN U3912 ( .A(n14766), .B(n4068), .Z(n2589) );
  NANDN U3913 ( .A(n14729), .B(n42115), .Z(n2590) );
  AND U3914 ( .A(n2589), .B(n2590), .Z(n14768) );
  NANDN U3915 ( .A(n14762), .B(n42047), .Z(n2591) );
  NANDN U3916 ( .A(n14799), .B(n4067), .Z(n2592) );
  NAND U3917 ( .A(n2591), .B(n2592), .Z(n14810) );
  NANDN U3918 ( .A(n14837), .B(n4068), .Z(n2593) );
  NANDN U3919 ( .A(n14800), .B(n42115), .Z(n2594) );
  AND U3920 ( .A(n2593), .B(n2594), .Z(n14842) );
  NANDN U3921 ( .A(n14836), .B(n42047), .Z(n2595) );
  NANDN U3922 ( .A(n14873), .B(n4067), .Z(n2596) );
  NAND U3923 ( .A(n2595), .B(n2596), .Z(n14884) );
  NANDN U3924 ( .A(n14914), .B(n4068), .Z(n2597) );
  NANDN U3925 ( .A(n14877), .B(n42115), .Z(n2598) );
  AND U3926 ( .A(n2597), .B(n2598), .Z(n14916) );
  NANDN U3927 ( .A(n14910), .B(n42047), .Z(n2599) );
  NANDN U3928 ( .A(n14947), .B(n4067), .Z(n2600) );
  NAND U3929 ( .A(n2599), .B(n2600), .Z(n14958) );
  NANDN U3930 ( .A(n14985), .B(n4068), .Z(n2601) );
  NANDN U3931 ( .A(n14951), .B(n42115), .Z(n2602) );
  AND U3932 ( .A(n2601), .B(n2602), .Z(n14990) );
  NANDN U3933 ( .A(n14984), .B(n42047), .Z(n2603) );
  NANDN U3934 ( .A(n15021), .B(n4067), .Z(n2604) );
  NAND U3935 ( .A(n2603), .B(n2604), .Z(n15032) );
  NANDN U3936 ( .A(n15062), .B(n4068), .Z(n2605) );
  NANDN U3937 ( .A(n15025), .B(n42115), .Z(n2606) );
  AND U3938 ( .A(n2605), .B(n2606), .Z(n15064) );
  NANDN U3939 ( .A(n15058), .B(n42047), .Z(n2607) );
  NANDN U3940 ( .A(n15095), .B(n4067), .Z(n2608) );
  NAND U3941 ( .A(n2607), .B(n2608), .Z(n15106) );
  NANDN U3942 ( .A(n15136), .B(n4068), .Z(n2609) );
  NANDN U3943 ( .A(n15099), .B(n42115), .Z(n2610) );
  AND U3944 ( .A(n2609), .B(n2610), .Z(n15138) );
  NANDN U3945 ( .A(n15132), .B(n42047), .Z(n2611) );
  NANDN U3946 ( .A(n15169), .B(n4067), .Z(n2612) );
  NAND U3947 ( .A(n2611), .B(n2612), .Z(n15180) );
  NANDN U3948 ( .A(n15210), .B(n4068), .Z(n2613) );
  NANDN U3949 ( .A(n15170), .B(n42115), .Z(n2614) );
  AND U3950 ( .A(n2613), .B(n2614), .Z(n15212) );
  NANDN U3951 ( .A(n15206), .B(n42047), .Z(n2615) );
  NANDN U3952 ( .A(n15243), .B(n4067), .Z(n2616) );
  NAND U3953 ( .A(n2615), .B(n2616), .Z(n15254) );
  NANDN U3954 ( .A(n15284), .B(n4068), .Z(n2617) );
  NANDN U3955 ( .A(n15244), .B(n42115), .Z(n2618) );
  AND U3956 ( .A(n2617), .B(n2618), .Z(n15286) );
  NANDN U3957 ( .A(n15280), .B(n42047), .Z(n2619) );
  NANDN U3958 ( .A(n15317), .B(n4067), .Z(n2620) );
  NAND U3959 ( .A(n2619), .B(n2620), .Z(n15328) );
  NANDN U3960 ( .A(n15355), .B(n4068), .Z(n2621) );
  NANDN U3961 ( .A(n15318), .B(n42115), .Z(n2622) );
  AND U3962 ( .A(n2621), .B(n2622), .Z(n15360) );
  NANDN U3963 ( .A(n15354), .B(n42047), .Z(n2623) );
  NANDN U3964 ( .A(n15391), .B(n4067), .Z(n2624) );
  NAND U3965 ( .A(n2623), .B(n2624), .Z(n15402) );
  NANDN U3966 ( .A(n15429), .B(n4068), .Z(n2625) );
  NANDN U3967 ( .A(n15395), .B(n42115), .Z(n2626) );
  AND U3968 ( .A(n2625), .B(n2626), .Z(n15434) );
  NANDN U3969 ( .A(n15428), .B(n42047), .Z(n2627) );
  NANDN U3970 ( .A(n15465), .B(n4067), .Z(n2628) );
  NAND U3971 ( .A(n2627), .B(n2628), .Z(n15476) );
  NANDN U3972 ( .A(n15503), .B(n4068), .Z(n2629) );
  NANDN U3973 ( .A(n15469), .B(n42115), .Z(n2630) );
  AND U3974 ( .A(n2629), .B(n2630), .Z(n15508) );
  NANDN U3975 ( .A(n15502), .B(n42047), .Z(n2631) );
  NANDN U3976 ( .A(n15539), .B(n4067), .Z(n2632) );
  NAND U3977 ( .A(n2631), .B(n2632), .Z(n15550) );
  NANDN U3978 ( .A(n15580), .B(n4068), .Z(n2633) );
  NANDN U3979 ( .A(n15543), .B(n42115), .Z(n2634) );
  AND U3980 ( .A(n2633), .B(n2634), .Z(n15582) );
  NANDN U3981 ( .A(n15576), .B(n42047), .Z(n2635) );
  NANDN U3982 ( .A(n15613), .B(n4067), .Z(n2636) );
  NAND U3983 ( .A(n2635), .B(n2636), .Z(n15624) );
  NANDN U3984 ( .A(n15651), .B(n4068), .Z(n2637) );
  NANDN U3985 ( .A(n15617), .B(n42115), .Z(n2638) );
  AND U3986 ( .A(n2637), .B(n2638), .Z(n15656) );
  NANDN U3987 ( .A(n15650), .B(n42047), .Z(n2639) );
  NANDN U3988 ( .A(n15687), .B(n4067), .Z(n2640) );
  NAND U3989 ( .A(n2639), .B(n2640), .Z(n15698) );
  NANDN U3990 ( .A(n15728), .B(n4068), .Z(n2641) );
  NANDN U3991 ( .A(n15691), .B(n42115), .Z(n2642) );
  AND U3992 ( .A(n2641), .B(n2642), .Z(n15730) );
  NANDN U3993 ( .A(n15724), .B(n42047), .Z(n2643) );
  NANDN U3994 ( .A(n15761), .B(n4067), .Z(n2644) );
  NAND U3995 ( .A(n2643), .B(n2644), .Z(n15772) );
  NANDN U3996 ( .A(n15802), .B(n4068), .Z(n2645) );
  NANDN U3997 ( .A(n15762), .B(n42115), .Z(n2646) );
  AND U3998 ( .A(n2645), .B(n2646), .Z(n15804) );
  NANDN U3999 ( .A(n15798), .B(n42047), .Z(n2647) );
  NANDN U4000 ( .A(n15835), .B(n4067), .Z(n2648) );
  NAND U4001 ( .A(n2647), .B(n2648), .Z(n15846) );
  NANDN U4002 ( .A(n15876), .B(n4068), .Z(n2649) );
  NANDN U4003 ( .A(n15836), .B(n42115), .Z(n2650) );
  AND U4004 ( .A(n2649), .B(n2650), .Z(n15878) );
  NANDN U4005 ( .A(n15872), .B(n42047), .Z(n2651) );
  NANDN U4006 ( .A(n15909), .B(n4067), .Z(n2652) );
  NAND U4007 ( .A(n2651), .B(n2652), .Z(n15920) );
  NANDN U4008 ( .A(n15950), .B(n4068), .Z(n2653) );
  NANDN U4009 ( .A(n15913), .B(n42115), .Z(n2654) );
  AND U4010 ( .A(n2653), .B(n2654), .Z(n15952) );
  NANDN U4011 ( .A(n15946), .B(n42047), .Z(n2655) );
  NANDN U4012 ( .A(n15983), .B(n4067), .Z(n2656) );
  NAND U4013 ( .A(n2655), .B(n2656), .Z(n15994) );
  NANDN U4014 ( .A(n16024), .B(n4068), .Z(n2657) );
  NANDN U4015 ( .A(n15984), .B(n42115), .Z(n2658) );
  AND U4016 ( .A(n2657), .B(n2658), .Z(n16026) );
  NANDN U4017 ( .A(n16020), .B(n42047), .Z(n2659) );
  NANDN U4018 ( .A(n16057), .B(n4067), .Z(n2660) );
  NAND U4019 ( .A(n2659), .B(n2660), .Z(n16068) );
  NANDN U4020 ( .A(n16098), .B(n4068), .Z(n2661) );
  NANDN U4021 ( .A(n16058), .B(n42115), .Z(n2662) );
  AND U4022 ( .A(n2661), .B(n2662), .Z(n16100) );
  NANDN U4023 ( .A(n16094), .B(n42047), .Z(n2663) );
  NANDN U4024 ( .A(n16131), .B(n4067), .Z(n2664) );
  NAND U4025 ( .A(n2663), .B(n2664), .Z(n16142) );
  NANDN U4026 ( .A(n16172), .B(n4068), .Z(n2665) );
  NANDN U4027 ( .A(n16135), .B(n42115), .Z(n2666) );
  AND U4028 ( .A(n2665), .B(n2666), .Z(n16174) );
  NANDN U4029 ( .A(n16168), .B(n42047), .Z(n2667) );
  NANDN U4030 ( .A(n16205), .B(n4067), .Z(n2668) );
  NAND U4031 ( .A(n2667), .B(n2668), .Z(n16216) );
  NANDN U4032 ( .A(n16243), .B(n4068), .Z(n2669) );
  NANDN U4033 ( .A(n16209), .B(n42115), .Z(n2670) );
  AND U4034 ( .A(n2669), .B(n2670), .Z(n16248) );
  NANDN U4035 ( .A(n16242), .B(n42047), .Z(n2671) );
  NANDN U4036 ( .A(n16279), .B(n4067), .Z(n2672) );
  NAND U4037 ( .A(n2671), .B(n2672), .Z(n16290) );
  NANDN U4038 ( .A(n16320), .B(n4068), .Z(n2673) );
  NANDN U4039 ( .A(n16283), .B(n42115), .Z(n2674) );
  AND U4040 ( .A(n2673), .B(n2674), .Z(n16322) );
  NANDN U4041 ( .A(n16316), .B(n42047), .Z(n2675) );
  NANDN U4042 ( .A(n16353), .B(n4067), .Z(n2676) );
  NAND U4043 ( .A(n2675), .B(n2676), .Z(n16364) );
  NANDN U4044 ( .A(n16391), .B(n4068), .Z(n2677) );
  NANDN U4045 ( .A(n16357), .B(n42115), .Z(n2678) );
  AND U4046 ( .A(n2677), .B(n2678), .Z(n16396) );
  NANDN U4047 ( .A(n16390), .B(n42047), .Z(n2679) );
  NANDN U4048 ( .A(n16427), .B(n4067), .Z(n2680) );
  NAND U4049 ( .A(n2679), .B(n2680), .Z(n16438) );
  NANDN U4050 ( .A(n16465), .B(n4068), .Z(n2681) );
  NANDN U4051 ( .A(n16431), .B(n42115), .Z(n2682) );
  AND U4052 ( .A(n2681), .B(n2682), .Z(n16470) );
  NANDN U4053 ( .A(n16464), .B(n42047), .Z(n2683) );
  NANDN U4054 ( .A(n16501), .B(n4067), .Z(n2684) );
  NAND U4055 ( .A(n2683), .B(n2684), .Z(n16512) );
  NANDN U4056 ( .A(n16539), .B(n4068), .Z(n2685) );
  NANDN U4057 ( .A(n16505), .B(n42115), .Z(n2686) );
  AND U4058 ( .A(n2685), .B(n2686), .Z(n16544) );
  NANDN U4059 ( .A(n16538), .B(n42047), .Z(n2687) );
  NANDN U4060 ( .A(n16575), .B(n4067), .Z(n2688) );
  NAND U4061 ( .A(n2687), .B(n2688), .Z(n16586) );
  NANDN U4062 ( .A(n16616), .B(n4068), .Z(n2689) );
  NANDN U4063 ( .A(n16579), .B(n42115), .Z(n2690) );
  AND U4064 ( .A(n2689), .B(n2690), .Z(n16618) );
  NANDN U4065 ( .A(n16612), .B(n42047), .Z(n2691) );
  NANDN U4066 ( .A(n16649), .B(n4067), .Z(n2692) );
  NAND U4067 ( .A(n2691), .B(n2692), .Z(n16660) );
  NANDN U4068 ( .A(n16690), .B(n4068), .Z(n2693) );
  NANDN U4069 ( .A(n16653), .B(n42115), .Z(n2694) );
  AND U4070 ( .A(n2693), .B(n2694), .Z(n16692) );
  NANDN U4071 ( .A(n16686), .B(n42047), .Z(n2695) );
  NANDN U4072 ( .A(n16723), .B(n4067), .Z(n2696) );
  NAND U4073 ( .A(n2695), .B(n2696), .Z(n16734) );
  NANDN U4074 ( .A(n16764), .B(n4068), .Z(n2697) );
  NANDN U4075 ( .A(n16727), .B(n42115), .Z(n2698) );
  AND U4076 ( .A(n2697), .B(n2698), .Z(n16766) );
  NANDN U4077 ( .A(n16760), .B(n42047), .Z(n2699) );
  NANDN U4078 ( .A(n16797), .B(n4067), .Z(n2700) );
  NAND U4079 ( .A(n2699), .B(n2700), .Z(n16808) );
  NANDN U4080 ( .A(n16838), .B(n4068), .Z(n2701) );
  NANDN U4081 ( .A(n16801), .B(n42115), .Z(n2702) );
  AND U4082 ( .A(n2701), .B(n2702), .Z(n16840) );
  NANDN U4083 ( .A(n16834), .B(n42047), .Z(n2703) );
  NANDN U4084 ( .A(n16871), .B(n4067), .Z(n2704) );
  NAND U4085 ( .A(n2703), .B(n2704), .Z(n16882) );
  NANDN U4086 ( .A(n16912), .B(n4068), .Z(n2705) );
  NANDN U4087 ( .A(n16872), .B(n42115), .Z(n2706) );
  AND U4088 ( .A(n2705), .B(n2706), .Z(n16914) );
  NANDN U4089 ( .A(n16908), .B(n42047), .Z(n2707) );
  NANDN U4090 ( .A(n16945), .B(n4067), .Z(n2708) );
  NAND U4091 ( .A(n2707), .B(n2708), .Z(n16956) );
  NANDN U4092 ( .A(n16986), .B(n4068), .Z(n2709) );
  NANDN U4093 ( .A(n16949), .B(n42115), .Z(n2710) );
  AND U4094 ( .A(n2709), .B(n2710), .Z(n16988) );
  NANDN U4095 ( .A(n16982), .B(n42047), .Z(n2711) );
  NANDN U4096 ( .A(n17019), .B(n4067), .Z(n2712) );
  NAND U4097 ( .A(n2711), .B(n2712), .Z(n17030) );
  NANDN U4098 ( .A(n17060), .B(n4068), .Z(n2713) );
  NANDN U4099 ( .A(n17023), .B(n42115), .Z(n2714) );
  AND U4100 ( .A(n2713), .B(n2714), .Z(n17062) );
  NANDN U4101 ( .A(n17056), .B(n42047), .Z(n2715) );
  NANDN U4102 ( .A(n17093), .B(n4067), .Z(n2716) );
  NAND U4103 ( .A(n2715), .B(n2716), .Z(n17104) );
  NANDN U4104 ( .A(n17134), .B(n4068), .Z(n2717) );
  NANDN U4105 ( .A(n17094), .B(n42115), .Z(n2718) );
  AND U4106 ( .A(n2717), .B(n2718), .Z(n17136) );
  NANDN U4107 ( .A(n17130), .B(n42047), .Z(n2719) );
  NANDN U4108 ( .A(n17167), .B(n4067), .Z(n2720) );
  NAND U4109 ( .A(n2719), .B(n2720), .Z(n17178) );
  NANDN U4110 ( .A(n17208), .B(n4068), .Z(n2721) );
  NANDN U4111 ( .A(n17168), .B(n42115), .Z(n2722) );
  AND U4112 ( .A(n2721), .B(n2722), .Z(n17210) );
  NANDN U4113 ( .A(n17204), .B(n42047), .Z(n2723) );
  NANDN U4114 ( .A(n17241), .B(n4067), .Z(n2724) );
  NAND U4115 ( .A(n2723), .B(n2724), .Z(n17252) );
  NANDN U4116 ( .A(n17282), .B(n4068), .Z(n2725) );
  NANDN U4117 ( .A(n17242), .B(n42115), .Z(n2726) );
  AND U4118 ( .A(n2725), .B(n2726), .Z(n17284) );
  NANDN U4119 ( .A(n17278), .B(n42047), .Z(n2727) );
  NANDN U4120 ( .A(n17315), .B(n4067), .Z(n2728) );
  NAND U4121 ( .A(n2727), .B(n2728), .Z(n17326) );
  NANDN U4122 ( .A(n17356), .B(n4068), .Z(n2729) );
  NANDN U4123 ( .A(n17319), .B(n42115), .Z(n2730) );
  AND U4124 ( .A(n2729), .B(n2730), .Z(n17358) );
  NANDN U4125 ( .A(n17352), .B(n42047), .Z(n2731) );
  NANDN U4126 ( .A(n17389), .B(n4067), .Z(n2732) );
  NAND U4127 ( .A(n2731), .B(n2732), .Z(n17400) );
  NANDN U4128 ( .A(n17430), .B(n4068), .Z(n2733) );
  NANDN U4129 ( .A(n17390), .B(n42115), .Z(n2734) );
  AND U4130 ( .A(n2733), .B(n2734), .Z(n17432) );
  NANDN U4131 ( .A(n17426), .B(n42047), .Z(n2735) );
  NANDN U4132 ( .A(n17463), .B(n4067), .Z(n2736) );
  NAND U4133 ( .A(n2735), .B(n2736), .Z(n17474) );
  NANDN U4134 ( .A(n17504), .B(n4068), .Z(n2737) );
  NANDN U4135 ( .A(n17467), .B(n42115), .Z(n2738) );
  AND U4136 ( .A(n2737), .B(n2738), .Z(n17506) );
  NANDN U4137 ( .A(n17500), .B(n42047), .Z(n2739) );
  NANDN U4138 ( .A(n17537), .B(n4067), .Z(n2740) );
  NAND U4139 ( .A(n2739), .B(n2740), .Z(n17548) );
  NANDN U4140 ( .A(n17578), .B(n4068), .Z(n2741) );
  NANDN U4141 ( .A(n17541), .B(n42115), .Z(n2742) );
  AND U4142 ( .A(n2741), .B(n2742), .Z(n17580) );
  NANDN U4143 ( .A(n17574), .B(n42047), .Z(n2743) );
  NANDN U4144 ( .A(n17611), .B(n4067), .Z(n2744) );
  NAND U4145 ( .A(n2743), .B(n2744), .Z(n17622) );
  NANDN U4146 ( .A(n17649), .B(n4068), .Z(n2745) );
  NANDN U4147 ( .A(n17615), .B(n42115), .Z(n2746) );
  AND U4148 ( .A(n2745), .B(n2746), .Z(n17654) );
  NANDN U4149 ( .A(n17648), .B(n42047), .Z(n2747) );
  NANDN U4150 ( .A(n17685), .B(n4067), .Z(n2748) );
  NAND U4151 ( .A(n2747), .B(n2748), .Z(n17696) );
  NANDN U4152 ( .A(n17726), .B(n4068), .Z(n2749) );
  NANDN U4153 ( .A(n17689), .B(n42115), .Z(n2750) );
  AND U4154 ( .A(n2749), .B(n2750), .Z(n17728) );
  NANDN U4155 ( .A(n17722), .B(n42047), .Z(n2751) );
  NANDN U4156 ( .A(n17759), .B(n4067), .Z(n2752) );
  NAND U4157 ( .A(n2751), .B(n2752), .Z(n17770) );
  NANDN U4158 ( .A(n17797), .B(n4068), .Z(n2753) );
  NANDN U4159 ( .A(n17763), .B(n42115), .Z(n2754) );
  AND U4160 ( .A(n2753), .B(n2754), .Z(n17802) );
  NANDN U4161 ( .A(n17796), .B(n42047), .Z(n2755) );
  NANDN U4162 ( .A(n17833), .B(n4067), .Z(n2756) );
  NAND U4163 ( .A(n2755), .B(n2756), .Z(n17844) );
  NANDN U4164 ( .A(n17874), .B(n4068), .Z(n2757) );
  NANDN U4165 ( .A(n17837), .B(n42115), .Z(n2758) );
  AND U4166 ( .A(n2757), .B(n2758), .Z(n17876) );
  NANDN U4167 ( .A(n17870), .B(n42047), .Z(n2759) );
  NANDN U4168 ( .A(n17907), .B(n4067), .Z(n2760) );
  NAND U4169 ( .A(n2759), .B(n2760), .Z(n17918) );
  NANDN U4170 ( .A(n17948), .B(n4068), .Z(n2761) );
  NANDN U4171 ( .A(n17911), .B(n42115), .Z(n2762) );
  AND U4172 ( .A(n2761), .B(n2762), .Z(n17950) );
  NANDN U4173 ( .A(n17944), .B(n42047), .Z(n2763) );
  NANDN U4174 ( .A(n17981), .B(n4067), .Z(n2764) );
  NAND U4175 ( .A(n2763), .B(n2764), .Z(n17992) );
  NANDN U4176 ( .A(n18022), .B(n4068), .Z(n2765) );
  NANDN U4177 ( .A(n17985), .B(n42115), .Z(n2766) );
  AND U4178 ( .A(n2765), .B(n2766), .Z(n18024) );
  NANDN U4179 ( .A(n18018), .B(n42047), .Z(n2767) );
  NANDN U4180 ( .A(n18055), .B(n4067), .Z(n2768) );
  NAND U4181 ( .A(n2767), .B(n2768), .Z(n18066) );
  NANDN U4182 ( .A(n18096), .B(n4068), .Z(n2769) );
  NANDN U4183 ( .A(n18059), .B(n42115), .Z(n2770) );
  AND U4184 ( .A(n2769), .B(n2770), .Z(n18098) );
  NANDN U4185 ( .A(n18092), .B(n42047), .Z(n2771) );
  NANDN U4186 ( .A(n18129), .B(n4067), .Z(n2772) );
  NAND U4187 ( .A(n2771), .B(n2772), .Z(n18140) );
  NANDN U4188 ( .A(n18167), .B(n4068), .Z(n2773) );
  NANDN U4189 ( .A(n18133), .B(n42115), .Z(n2774) );
  AND U4190 ( .A(n2773), .B(n2774), .Z(n18172) );
  NANDN U4191 ( .A(n18166), .B(n42047), .Z(n2775) );
  NANDN U4192 ( .A(n18203), .B(n4067), .Z(n2776) );
  NAND U4193 ( .A(n2775), .B(n2776), .Z(n18214) );
  NANDN U4194 ( .A(n18244), .B(n4068), .Z(n2777) );
  NANDN U4195 ( .A(n18207), .B(n42115), .Z(n2778) );
  AND U4196 ( .A(n2777), .B(n2778), .Z(n18246) );
  NANDN U4197 ( .A(n18240), .B(n42047), .Z(n2779) );
  NANDN U4198 ( .A(n18277), .B(n4067), .Z(n2780) );
  NAND U4199 ( .A(n2779), .B(n2780), .Z(n18288) );
  NANDN U4200 ( .A(n18318), .B(n4068), .Z(n2781) );
  NANDN U4201 ( .A(n18281), .B(n42115), .Z(n2782) );
  AND U4202 ( .A(n2781), .B(n2782), .Z(n18320) );
  NANDN U4203 ( .A(n18314), .B(n42047), .Z(n2783) );
  NANDN U4204 ( .A(n18351), .B(n4067), .Z(n2784) );
  NAND U4205 ( .A(n2783), .B(n2784), .Z(n18362) );
  NANDN U4206 ( .A(n18392), .B(n4068), .Z(n2785) );
  NANDN U4207 ( .A(n18355), .B(n42115), .Z(n2786) );
  AND U4208 ( .A(n2785), .B(n2786), .Z(n18394) );
  NANDN U4209 ( .A(n18388), .B(n42047), .Z(n2787) );
  NANDN U4210 ( .A(n18425), .B(n4067), .Z(n2788) );
  NAND U4211 ( .A(n2787), .B(n2788), .Z(n18436) );
  NANDN U4212 ( .A(n18463), .B(n4068), .Z(n2789) );
  NANDN U4213 ( .A(n18429), .B(n42115), .Z(n2790) );
  AND U4214 ( .A(n2789), .B(n2790), .Z(n18468) );
  NANDN U4215 ( .A(n18462), .B(n42047), .Z(n2791) );
  NANDN U4216 ( .A(n18499), .B(n4067), .Z(n2792) );
  NAND U4217 ( .A(n2791), .B(n2792), .Z(n18510) );
  NANDN U4218 ( .A(n18540), .B(n4068), .Z(n2793) );
  NANDN U4219 ( .A(n18503), .B(n42115), .Z(n2794) );
  AND U4220 ( .A(n2793), .B(n2794), .Z(n18542) );
  NANDN U4221 ( .A(n18536), .B(n42047), .Z(n2795) );
  NANDN U4222 ( .A(n18573), .B(n4067), .Z(n2796) );
  NAND U4223 ( .A(n2795), .B(n2796), .Z(n18584) );
  NANDN U4224 ( .A(n18611), .B(n4068), .Z(n2797) );
  NANDN U4225 ( .A(n18577), .B(n42115), .Z(n2798) );
  AND U4226 ( .A(n2797), .B(n2798), .Z(n18616) );
  NANDN U4227 ( .A(n18610), .B(n42047), .Z(n2799) );
  NANDN U4228 ( .A(n18647), .B(n4067), .Z(n2800) );
  NAND U4229 ( .A(n2799), .B(n2800), .Z(n18658) );
  NANDN U4230 ( .A(n18688), .B(n4068), .Z(n2801) );
  NANDN U4231 ( .A(n18648), .B(n42115), .Z(n2802) );
  AND U4232 ( .A(n2801), .B(n2802), .Z(n18690) );
  NANDN U4233 ( .A(n18684), .B(n42047), .Z(n2803) );
  NANDN U4234 ( .A(n18721), .B(n4067), .Z(n2804) );
  NAND U4235 ( .A(n2803), .B(n2804), .Z(n18732) );
  NANDN U4236 ( .A(n18759), .B(n4068), .Z(n2805) );
  NANDN U4237 ( .A(n18725), .B(n42115), .Z(n2806) );
  AND U4238 ( .A(n2805), .B(n2806), .Z(n18764) );
  NANDN U4239 ( .A(n18758), .B(n42047), .Z(n2807) );
  NANDN U4240 ( .A(n18795), .B(n4067), .Z(n2808) );
  NAND U4241 ( .A(n2807), .B(n2808), .Z(n18806) );
  NANDN U4242 ( .A(n18833), .B(n4068), .Z(n2809) );
  NANDN U4243 ( .A(n18796), .B(n42115), .Z(n2810) );
  AND U4244 ( .A(n2809), .B(n2810), .Z(n18838) );
  NANDN U4245 ( .A(n18832), .B(n42047), .Z(n2811) );
  NANDN U4246 ( .A(n18869), .B(n4067), .Z(n2812) );
  NAND U4247 ( .A(n2811), .B(n2812), .Z(n18880) );
  NANDN U4248 ( .A(n18907), .B(n4068), .Z(n2813) );
  NANDN U4249 ( .A(n18873), .B(n42115), .Z(n2814) );
  AND U4250 ( .A(n2813), .B(n2814), .Z(n18912) );
  NANDN U4251 ( .A(n18906), .B(n42047), .Z(n2815) );
  NANDN U4252 ( .A(n18943), .B(n4067), .Z(n2816) );
  NAND U4253 ( .A(n2815), .B(n2816), .Z(n18954) );
  NANDN U4254 ( .A(n18984), .B(n4068), .Z(n2817) );
  NANDN U4255 ( .A(n18944), .B(n42115), .Z(n2818) );
  AND U4256 ( .A(n2817), .B(n2818), .Z(n18986) );
  NANDN U4257 ( .A(n18980), .B(n42047), .Z(n2819) );
  NANDN U4258 ( .A(n19017), .B(n4067), .Z(n2820) );
  NAND U4259 ( .A(n2819), .B(n2820), .Z(n19028) );
  NANDN U4260 ( .A(n19058), .B(n4068), .Z(n2821) );
  NANDN U4261 ( .A(n19018), .B(n42115), .Z(n2822) );
  AND U4262 ( .A(n2821), .B(n2822), .Z(n19060) );
  NANDN U4263 ( .A(n19054), .B(n42047), .Z(n2823) );
  NANDN U4264 ( .A(n19091), .B(n4067), .Z(n2824) );
  NAND U4265 ( .A(n2823), .B(n2824), .Z(n19102) );
  NANDN U4266 ( .A(n19132), .B(n4068), .Z(n2825) );
  NANDN U4267 ( .A(n19092), .B(n42115), .Z(n2826) );
  AND U4268 ( .A(n2825), .B(n2826), .Z(n19134) );
  NANDN U4269 ( .A(n19128), .B(n42047), .Z(n2827) );
  NANDN U4270 ( .A(n19165), .B(n4067), .Z(n2828) );
  NAND U4271 ( .A(n2827), .B(n2828), .Z(n19176) );
  NANDN U4272 ( .A(n19206), .B(n4068), .Z(n2829) );
  NANDN U4273 ( .A(n19166), .B(n42115), .Z(n2830) );
  AND U4274 ( .A(n2829), .B(n2830), .Z(n19208) );
  NANDN U4275 ( .A(n19202), .B(n42047), .Z(n2831) );
  NANDN U4276 ( .A(n19239), .B(n4067), .Z(n2832) );
  NAND U4277 ( .A(n2831), .B(n2832), .Z(n19250) );
  NANDN U4278 ( .A(n19280), .B(n4068), .Z(n2833) );
  NANDN U4279 ( .A(n19243), .B(n42115), .Z(n2834) );
  AND U4280 ( .A(n2833), .B(n2834), .Z(n19282) );
  NANDN U4281 ( .A(n19276), .B(n42047), .Z(n2835) );
  NANDN U4282 ( .A(n19313), .B(n4067), .Z(n2836) );
  NAND U4283 ( .A(n2835), .B(n2836), .Z(n19324) );
  NANDN U4284 ( .A(n19354), .B(n4068), .Z(n2837) );
  NANDN U4285 ( .A(n19317), .B(n42115), .Z(n2838) );
  AND U4286 ( .A(n2837), .B(n2838), .Z(n19356) );
  NANDN U4287 ( .A(n19350), .B(n42047), .Z(n2839) );
  NANDN U4288 ( .A(n19387), .B(n4067), .Z(n2840) );
  NAND U4289 ( .A(n2839), .B(n2840), .Z(n19398) );
  NANDN U4290 ( .A(n19425), .B(n4068), .Z(n2841) );
  NANDN U4291 ( .A(n19391), .B(n42115), .Z(n2842) );
  AND U4292 ( .A(n2841), .B(n2842), .Z(n19430) );
  NANDN U4293 ( .A(n19424), .B(n42047), .Z(n2843) );
  NANDN U4294 ( .A(n19461), .B(n4067), .Z(n2844) );
  NAND U4295 ( .A(n2843), .B(n2844), .Z(n19472) );
  NANDN U4296 ( .A(n19502), .B(n4068), .Z(n2845) );
  NANDN U4297 ( .A(n19465), .B(n42115), .Z(n2846) );
  AND U4298 ( .A(n2845), .B(n2846), .Z(n19504) );
  NANDN U4299 ( .A(n19498), .B(n42047), .Z(n2847) );
  NANDN U4300 ( .A(n19535), .B(n4067), .Z(n2848) );
  NAND U4301 ( .A(n2847), .B(n2848), .Z(n19546) );
  NANDN U4302 ( .A(n19576), .B(n4068), .Z(n2849) );
  NANDN U4303 ( .A(n19539), .B(n42115), .Z(n2850) );
  AND U4304 ( .A(n2849), .B(n2850), .Z(n19578) );
  NANDN U4305 ( .A(n19572), .B(n42047), .Z(n2851) );
  NANDN U4306 ( .A(n19609), .B(n4067), .Z(n2852) );
  NAND U4307 ( .A(n2851), .B(n2852), .Z(n19620) );
  NANDN U4308 ( .A(n19650), .B(n4068), .Z(n2853) );
  NANDN U4309 ( .A(n19613), .B(n42115), .Z(n2854) );
  AND U4310 ( .A(n2853), .B(n2854), .Z(n19652) );
  NANDN U4311 ( .A(n19646), .B(n42047), .Z(n2855) );
  NANDN U4312 ( .A(n19683), .B(n4067), .Z(n2856) );
  NAND U4313 ( .A(n2855), .B(n2856), .Z(n19694) );
  NANDN U4314 ( .A(n19721), .B(n4068), .Z(n2857) );
  NANDN U4315 ( .A(n19687), .B(n42115), .Z(n2858) );
  AND U4316 ( .A(n2857), .B(n2858), .Z(n19726) );
  NANDN U4317 ( .A(n19720), .B(n42047), .Z(n2859) );
  NANDN U4318 ( .A(n19757), .B(n4067), .Z(n2860) );
  NAND U4319 ( .A(n2859), .B(n2860), .Z(n19768) );
  NANDN U4320 ( .A(n19798), .B(n4068), .Z(n2861) );
  NANDN U4321 ( .A(n19761), .B(n42115), .Z(n2862) );
  AND U4322 ( .A(n2861), .B(n2862), .Z(n19800) );
  NANDN U4323 ( .A(n19794), .B(n42047), .Z(n2863) );
  NANDN U4324 ( .A(n19831), .B(n4067), .Z(n2864) );
  NAND U4325 ( .A(n2863), .B(n2864), .Z(n19842) );
  NANDN U4326 ( .A(n19872), .B(n4068), .Z(n2865) );
  NANDN U4327 ( .A(n19832), .B(n42115), .Z(n2866) );
  AND U4328 ( .A(n2865), .B(n2866), .Z(n19874) );
  NANDN U4329 ( .A(n19868), .B(n42047), .Z(n2867) );
  NANDN U4330 ( .A(n19905), .B(n4067), .Z(n2868) );
  NAND U4331 ( .A(n2867), .B(n2868), .Z(n19916) );
  NANDN U4332 ( .A(n19946), .B(n4068), .Z(n2869) );
  NANDN U4333 ( .A(n19909), .B(n42115), .Z(n2870) );
  AND U4334 ( .A(n2869), .B(n2870), .Z(n19948) );
  NANDN U4335 ( .A(n19942), .B(n42047), .Z(n2871) );
  NANDN U4336 ( .A(n19979), .B(n4067), .Z(n2872) );
  NAND U4337 ( .A(n2871), .B(n2872), .Z(n19990) );
  NANDN U4338 ( .A(n20020), .B(n4068), .Z(n2873) );
  NANDN U4339 ( .A(n19980), .B(n42115), .Z(n2874) );
  AND U4340 ( .A(n2873), .B(n2874), .Z(n20022) );
  NANDN U4341 ( .A(n20016), .B(n42047), .Z(n2875) );
  NANDN U4342 ( .A(n20053), .B(n4067), .Z(n2876) );
  NAND U4343 ( .A(n2875), .B(n2876), .Z(n20064) );
  NANDN U4344 ( .A(n20094), .B(n4068), .Z(n2877) );
  NANDN U4345 ( .A(n20057), .B(n42115), .Z(n2878) );
  AND U4346 ( .A(n2877), .B(n2878), .Z(n20096) );
  NANDN U4347 ( .A(n20090), .B(n42047), .Z(n2879) );
  NANDN U4348 ( .A(n20127), .B(n4067), .Z(n2880) );
  NAND U4349 ( .A(n2879), .B(n2880), .Z(n20138) );
  NANDN U4350 ( .A(n20165), .B(n4068), .Z(n2881) );
  NANDN U4351 ( .A(n20131), .B(n42115), .Z(n2882) );
  AND U4352 ( .A(n2881), .B(n2882), .Z(n20170) );
  NANDN U4353 ( .A(n20164), .B(n42047), .Z(n2883) );
  NANDN U4354 ( .A(n20201), .B(n4067), .Z(n2884) );
  NAND U4355 ( .A(n2883), .B(n2884), .Z(n20212) );
  NANDN U4356 ( .A(n20242), .B(n4068), .Z(n2885) );
  NANDN U4357 ( .A(n20205), .B(n42115), .Z(n2886) );
  AND U4358 ( .A(n2885), .B(n2886), .Z(n20244) );
  NANDN U4359 ( .A(n20238), .B(n42047), .Z(n2887) );
  NANDN U4360 ( .A(n20275), .B(n4067), .Z(n2888) );
  NAND U4361 ( .A(n2887), .B(n2888), .Z(n20286) );
  NANDN U4362 ( .A(n20316), .B(n4068), .Z(n2889) );
  NANDN U4363 ( .A(n20279), .B(n42115), .Z(n2890) );
  AND U4364 ( .A(n2889), .B(n2890), .Z(n20318) );
  NANDN U4365 ( .A(n20312), .B(n42047), .Z(n2891) );
  NANDN U4366 ( .A(n20349), .B(n4067), .Z(n2892) );
  NAND U4367 ( .A(n2891), .B(n2892), .Z(n20360) );
  NANDN U4368 ( .A(n20390), .B(n4068), .Z(n2893) );
  NANDN U4369 ( .A(n20353), .B(n42115), .Z(n2894) );
  AND U4370 ( .A(n2893), .B(n2894), .Z(n20392) );
  NANDN U4371 ( .A(n20386), .B(n42047), .Z(n2895) );
  NANDN U4372 ( .A(n20423), .B(n4067), .Z(n2896) );
  NAND U4373 ( .A(n2895), .B(n2896), .Z(n20434) );
  NANDN U4374 ( .A(n20464), .B(n4068), .Z(n2897) );
  NANDN U4375 ( .A(n20424), .B(n42115), .Z(n2898) );
  AND U4376 ( .A(n2897), .B(n2898), .Z(n20466) );
  NANDN U4377 ( .A(n20460), .B(n42047), .Z(n2899) );
  NANDN U4378 ( .A(n20497), .B(n4067), .Z(n2900) );
  NAND U4379 ( .A(n2899), .B(n2900), .Z(n20508) );
  NANDN U4380 ( .A(n20538), .B(n4068), .Z(n2901) );
  NANDN U4381 ( .A(n20501), .B(n42115), .Z(n2902) );
  AND U4382 ( .A(n2901), .B(n2902), .Z(n20540) );
  NANDN U4383 ( .A(n20534), .B(n42047), .Z(n2903) );
  NANDN U4384 ( .A(n20571), .B(n4067), .Z(n2904) );
  NAND U4385 ( .A(n2903), .B(n2904), .Z(n20582) );
  NANDN U4386 ( .A(n20612), .B(n4068), .Z(n2905) );
  NANDN U4387 ( .A(n20572), .B(n42115), .Z(n2906) );
  AND U4388 ( .A(n2905), .B(n2906), .Z(n20614) );
  NANDN U4389 ( .A(n20608), .B(n42047), .Z(n2907) );
  NANDN U4390 ( .A(n20645), .B(n4067), .Z(n2908) );
  NAND U4391 ( .A(n2907), .B(n2908), .Z(n20656) );
  NANDN U4392 ( .A(n20686), .B(n4068), .Z(n2909) );
  NANDN U4393 ( .A(n20649), .B(n42115), .Z(n2910) );
  AND U4394 ( .A(n2909), .B(n2910), .Z(n20688) );
  NANDN U4395 ( .A(n20682), .B(n42047), .Z(n2911) );
  NANDN U4396 ( .A(n20719), .B(n4067), .Z(n2912) );
  NAND U4397 ( .A(n2911), .B(n2912), .Z(n20730) );
  NANDN U4398 ( .A(n20760), .B(n4068), .Z(n2913) );
  NANDN U4399 ( .A(n20723), .B(n42115), .Z(n2914) );
  AND U4400 ( .A(n2913), .B(n2914), .Z(n20762) );
  NANDN U4401 ( .A(n20756), .B(n42047), .Z(n2915) );
  NANDN U4402 ( .A(n20793), .B(n4067), .Z(n2916) );
  NAND U4403 ( .A(n2915), .B(n2916), .Z(n20804) );
  NANDN U4404 ( .A(n20834), .B(n4068), .Z(n2917) );
  NANDN U4405 ( .A(n20797), .B(n42115), .Z(n2918) );
  AND U4406 ( .A(n2917), .B(n2918), .Z(n20836) );
  NANDN U4407 ( .A(n20830), .B(n42047), .Z(n2919) );
  NANDN U4408 ( .A(n20867), .B(n4067), .Z(n2920) );
  NAND U4409 ( .A(n2919), .B(n2920), .Z(n20878) );
  NANDN U4410 ( .A(n20908), .B(n4068), .Z(n2921) );
  NANDN U4411 ( .A(n20871), .B(n42115), .Z(n2922) );
  AND U4412 ( .A(n2921), .B(n2922), .Z(n20910) );
  NANDN U4413 ( .A(n20904), .B(n42047), .Z(n2923) );
  NANDN U4414 ( .A(n20941), .B(n4067), .Z(n2924) );
  NAND U4415 ( .A(n2923), .B(n2924), .Z(n20952) );
  NANDN U4416 ( .A(n20982), .B(n4068), .Z(n2925) );
  NANDN U4417 ( .A(n20945), .B(n42115), .Z(n2926) );
  AND U4418 ( .A(n2925), .B(n2926), .Z(n20984) );
  NANDN U4419 ( .A(n20978), .B(n42047), .Z(n2927) );
  NANDN U4420 ( .A(n21015), .B(n4067), .Z(n2928) );
  NAND U4421 ( .A(n2927), .B(n2928), .Z(n21026) );
  NANDN U4422 ( .A(n21053), .B(n4068), .Z(n2929) );
  NANDN U4423 ( .A(n21019), .B(n42115), .Z(n2930) );
  AND U4424 ( .A(n2929), .B(n2930), .Z(n21058) );
  NANDN U4425 ( .A(n21052), .B(n42047), .Z(n2931) );
  NANDN U4426 ( .A(n21089), .B(n4067), .Z(n2932) );
  NAND U4427 ( .A(n2931), .B(n2932), .Z(n21100) );
  NANDN U4428 ( .A(n21130), .B(n4068), .Z(n2933) );
  NANDN U4429 ( .A(n21093), .B(n42115), .Z(n2934) );
  AND U4430 ( .A(n2933), .B(n2934), .Z(n21132) );
  NANDN U4431 ( .A(n21126), .B(n42047), .Z(n2935) );
  NANDN U4432 ( .A(n21163), .B(n4067), .Z(n2936) );
  NAND U4433 ( .A(n2935), .B(n2936), .Z(n21174) );
  NANDN U4434 ( .A(n21201), .B(n4068), .Z(n2937) );
  NANDN U4435 ( .A(n21167), .B(n42115), .Z(n2938) );
  AND U4436 ( .A(n2937), .B(n2938), .Z(n21206) );
  NANDN U4437 ( .A(n21200), .B(n42047), .Z(n2939) );
  NANDN U4438 ( .A(n21237), .B(n4067), .Z(n2940) );
  NAND U4439 ( .A(n2939), .B(n2940), .Z(n21248) );
  NANDN U4440 ( .A(n21278), .B(n4068), .Z(n2941) );
  NANDN U4441 ( .A(n21238), .B(n42115), .Z(n2942) );
  AND U4442 ( .A(n2941), .B(n2942), .Z(n21280) );
  NANDN U4443 ( .A(n21274), .B(n42047), .Z(n2943) );
  NANDN U4444 ( .A(n21311), .B(n4067), .Z(n2944) );
  NAND U4445 ( .A(n2943), .B(n2944), .Z(n21322) );
  NANDN U4446 ( .A(n21352), .B(n4068), .Z(n2945) );
  NANDN U4447 ( .A(n21312), .B(n42115), .Z(n2946) );
  AND U4448 ( .A(n2945), .B(n2946), .Z(n21354) );
  NANDN U4449 ( .A(n21348), .B(n42047), .Z(n2947) );
  NANDN U4450 ( .A(n21385), .B(n4067), .Z(n2948) );
  NAND U4451 ( .A(n2947), .B(n2948), .Z(n21396) );
  NANDN U4452 ( .A(n21423), .B(n4068), .Z(n2949) );
  NANDN U4453 ( .A(n21389), .B(n42115), .Z(n2950) );
  AND U4454 ( .A(n2949), .B(n2950), .Z(n21428) );
  NANDN U4455 ( .A(n21422), .B(n42047), .Z(n2951) );
  NANDN U4456 ( .A(n21459), .B(n4067), .Z(n2952) );
  NAND U4457 ( .A(n2951), .B(n2952), .Z(n21470) );
  NANDN U4458 ( .A(n21500), .B(n4068), .Z(n2953) );
  NANDN U4459 ( .A(n21463), .B(n42115), .Z(n2954) );
  AND U4460 ( .A(n2953), .B(n2954), .Z(n21502) );
  NANDN U4461 ( .A(n21496), .B(n42047), .Z(n2955) );
  NANDN U4462 ( .A(n21533), .B(n4067), .Z(n2956) );
  NAND U4463 ( .A(n2955), .B(n2956), .Z(n21544) );
  NANDN U4464 ( .A(n21571), .B(n4068), .Z(n2957) );
  NANDN U4465 ( .A(n21537), .B(n42115), .Z(n2958) );
  AND U4466 ( .A(n2957), .B(n2958), .Z(n21576) );
  NANDN U4467 ( .A(n21570), .B(n42047), .Z(n2959) );
  NANDN U4468 ( .A(n21607), .B(n4067), .Z(n2960) );
  NAND U4469 ( .A(n2959), .B(n2960), .Z(n21618) );
  NANDN U4470 ( .A(n21645), .B(n4068), .Z(n2961) );
  NANDN U4471 ( .A(n21611), .B(n42115), .Z(n2962) );
  AND U4472 ( .A(n2961), .B(n2962), .Z(n21650) );
  NANDN U4473 ( .A(n21644), .B(n42047), .Z(n2963) );
  NANDN U4474 ( .A(n21681), .B(n4067), .Z(n2964) );
  NAND U4475 ( .A(n2963), .B(n2964), .Z(n21692) );
  NANDN U4476 ( .A(n21722), .B(n4068), .Z(n2965) );
  NANDN U4477 ( .A(n21685), .B(n42115), .Z(n2966) );
  AND U4478 ( .A(n2965), .B(n2966), .Z(n21724) );
  NANDN U4479 ( .A(n21718), .B(n42047), .Z(n2967) );
  NANDN U4480 ( .A(n21755), .B(n4067), .Z(n2968) );
  NAND U4481 ( .A(n2967), .B(n2968), .Z(n21766) );
  NANDN U4482 ( .A(n21793), .B(n4068), .Z(n2969) );
  NANDN U4483 ( .A(n21759), .B(n42115), .Z(n2970) );
  AND U4484 ( .A(n2969), .B(n2970), .Z(n21798) );
  NANDN U4485 ( .A(n21792), .B(n42047), .Z(n2971) );
  NANDN U4486 ( .A(n21829), .B(n4067), .Z(n2972) );
  NAND U4487 ( .A(n2971), .B(n2972), .Z(n21840) );
  NANDN U4488 ( .A(n21870), .B(n4068), .Z(n2973) );
  NANDN U4489 ( .A(n21833), .B(n42115), .Z(n2974) );
  AND U4490 ( .A(n2973), .B(n2974), .Z(n21872) );
  NANDN U4491 ( .A(n21866), .B(n42047), .Z(n2975) );
  NANDN U4492 ( .A(n21903), .B(n4067), .Z(n2976) );
  NAND U4493 ( .A(n2975), .B(n2976), .Z(n21914) );
  NANDN U4494 ( .A(n21941), .B(n4068), .Z(n2977) );
  NANDN U4495 ( .A(n21907), .B(n42115), .Z(n2978) );
  AND U4496 ( .A(n2977), .B(n2978), .Z(n21946) );
  NANDN U4497 ( .A(n21940), .B(n42047), .Z(n2979) );
  NANDN U4498 ( .A(n21977), .B(n4067), .Z(n2980) );
  NAND U4499 ( .A(n2979), .B(n2980), .Z(n21988) );
  NANDN U4500 ( .A(n22018), .B(n4068), .Z(n2981) );
  NANDN U4501 ( .A(n21981), .B(n42115), .Z(n2982) );
  AND U4502 ( .A(n2981), .B(n2982), .Z(n22020) );
  NANDN U4503 ( .A(n22014), .B(n42047), .Z(n2983) );
  NANDN U4504 ( .A(n22051), .B(n4067), .Z(n2984) );
  NAND U4505 ( .A(n2983), .B(n2984), .Z(n22062) );
  NANDN U4506 ( .A(n22092), .B(n4068), .Z(n2985) );
  NANDN U4507 ( .A(n22052), .B(n42115), .Z(n2986) );
  AND U4508 ( .A(n2985), .B(n2986), .Z(n22094) );
  NANDN U4509 ( .A(n22088), .B(n42047), .Z(n2987) );
  NANDN U4510 ( .A(n22125), .B(n4067), .Z(n2988) );
  NAND U4511 ( .A(n2987), .B(n2988), .Z(n22136) );
  NANDN U4512 ( .A(n22166), .B(n4068), .Z(n2989) );
  NANDN U4513 ( .A(n22126), .B(n42115), .Z(n2990) );
  AND U4514 ( .A(n2989), .B(n2990), .Z(n22168) );
  NANDN U4515 ( .A(n22162), .B(n42047), .Z(n2991) );
  NANDN U4516 ( .A(n22199), .B(n4067), .Z(n2992) );
  NAND U4517 ( .A(n2991), .B(n2992), .Z(n22210) );
  NANDN U4518 ( .A(n22237), .B(n4068), .Z(n2993) );
  NANDN U4519 ( .A(n22203), .B(n42115), .Z(n2994) );
  AND U4520 ( .A(n2993), .B(n2994), .Z(n22242) );
  NANDN U4521 ( .A(n22236), .B(n42047), .Z(n2995) );
  NANDN U4522 ( .A(n22273), .B(n4067), .Z(n2996) );
  NAND U4523 ( .A(n2995), .B(n2996), .Z(n22284) );
  NANDN U4524 ( .A(n22314), .B(n4068), .Z(n2997) );
  NANDN U4525 ( .A(n22277), .B(n42115), .Z(n2998) );
  AND U4526 ( .A(n2997), .B(n2998), .Z(n22316) );
  NANDN U4527 ( .A(n22310), .B(n42047), .Z(n2999) );
  NANDN U4528 ( .A(n22347), .B(n4067), .Z(n3000) );
  NAND U4529 ( .A(n2999), .B(n3000), .Z(n22358) );
  NANDN U4530 ( .A(n22388), .B(n4068), .Z(n3001) );
  NANDN U4531 ( .A(n22351), .B(n42115), .Z(n3002) );
  AND U4532 ( .A(n3001), .B(n3002), .Z(n22390) );
  NANDN U4533 ( .A(n22384), .B(n42047), .Z(n3003) );
  NANDN U4534 ( .A(n22421), .B(n4067), .Z(n3004) );
  NAND U4535 ( .A(n3003), .B(n3004), .Z(n22432) );
  NANDN U4536 ( .A(n22462), .B(n4068), .Z(n3005) );
  NANDN U4537 ( .A(n22425), .B(n42115), .Z(n3006) );
  AND U4538 ( .A(n3005), .B(n3006), .Z(n22464) );
  NANDN U4539 ( .A(n22458), .B(n42047), .Z(n3007) );
  NANDN U4540 ( .A(n22495), .B(n4067), .Z(n3008) );
  NAND U4541 ( .A(n3007), .B(n3008), .Z(n22506) );
  NANDN U4542 ( .A(n22536), .B(n4068), .Z(n3009) );
  NANDN U4543 ( .A(n22496), .B(n42115), .Z(n3010) );
  AND U4544 ( .A(n3009), .B(n3010), .Z(n22538) );
  NANDN U4545 ( .A(n22532), .B(n42047), .Z(n3011) );
  NANDN U4546 ( .A(n22569), .B(n4067), .Z(n3012) );
  NAND U4547 ( .A(n3011), .B(n3012), .Z(n22580) );
  NANDN U4548 ( .A(n22610), .B(n4068), .Z(n3013) );
  NANDN U4549 ( .A(n22573), .B(n42115), .Z(n3014) );
  AND U4550 ( .A(n3013), .B(n3014), .Z(n22612) );
  NANDN U4551 ( .A(n22606), .B(n42047), .Z(n3015) );
  NANDN U4552 ( .A(n22643), .B(n4067), .Z(n3016) );
  NAND U4553 ( .A(n3015), .B(n3016), .Z(n22654) );
  NANDN U4554 ( .A(n22684), .B(n4068), .Z(n3017) );
  NANDN U4555 ( .A(n22647), .B(n42115), .Z(n3018) );
  AND U4556 ( .A(n3017), .B(n3018), .Z(n22686) );
  NANDN U4557 ( .A(n22680), .B(n42047), .Z(n3019) );
  NANDN U4558 ( .A(n22717), .B(n4067), .Z(n3020) );
  NAND U4559 ( .A(n3019), .B(n3020), .Z(n22728) );
  NANDN U4560 ( .A(n22763), .B(n4068), .Z(n3021) );
  NANDN U4561 ( .A(n22718), .B(n42115), .Z(n3022) );
  AND U4562 ( .A(n3021), .B(n3022), .Z(n22765) );
  NANDN U4563 ( .A(n22759), .B(n42047), .Z(n3023) );
  NANDN U4564 ( .A(n22791), .B(n4067), .Z(n3024) );
  NAND U4565 ( .A(n3023), .B(n3024), .Z(n22802) );
  NANDN U4566 ( .A(n22829), .B(n4068), .Z(n3025) );
  NANDN U4567 ( .A(n22792), .B(n42115), .Z(n3026) );
  AND U4568 ( .A(n3025), .B(n3026), .Z(n22834) );
  NANDN U4569 ( .A(n22828), .B(n42047), .Z(n3027) );
  NANDN U4570 ( .A(n22865), .B(n4067), .Z(n3028) );
  NAND U4571 ( .A(n3027), .B(n3028), .Z(n22876) );
  NANDN U4572 ( .A(n22903), .B(n4068), .Z(n3029) );
  NANDN U4573 ( .A(n22869), .B(n42115), .Z(n3030) );
  AND U4574 ( .A(n3029), .B(n3030), .Z(n22908) );
  NANDN U4575 ( .A(n22902), .B(n42047), .Z(n3031) );
  NANDN U4576 ( .A(n22939), .B(n4067), .Z(n3032) );
  NAND U4577 ( .A(n3031), .B(n3032), .Z(n22950) );
  NANDN U4578 ( .A(n22980), .B(n4068), .Z(n3033) );
  NANDN U4579 ( .A(n22943), .B(n42115), .Z(n3034) );
  AND U4580 ( .A(n3033), .B(n3034), .Z(n22982) );
  NANDN U4581 ( .A(n22976), .B(n42047), .Z(n3035) );
  NANDN U4582 ( .A(n23013), .B(n4067), .Z(n3036) );
  NAND U4583 ( .A(n3035), .B(n3036), .Z(n23024) );
  NANDN U4584 ( .A(n23054), .B(n4068), .Z(n3037) );
  NANDN U4585 ( .A(n23017), .B(n42115), .Z(n3038) );
  AND U4586 ( .A(n3037), .B(n3038), .Z(n23056) );
  NANDN U4587 ( .A(n23050), .B(n42047), .Z(n3039) );
  NANDN U4588 ( .A(n23087), .B(n4067), .Z(n3040) );
  NAND U4589 ( .A(n3039), .B(n3040), .Z(n23098) );
  NANDN U4590 ( .A(n23128), .B(n4068), .Z(n3041) );
  NANDN U4591 ( .A(n23088), .B(n42115), .Z(n3042) );
  AND U4592 ( .A(n3041), .B(n3042), .Z(n23130) );
  NANDN U4593 ( .A(n23124), .B(n42047), .Z(n3043) );
  NANDN U4594 ( .A(n23161), .B(n4067), .Z(n3044) );
  NAND U4595 ( .A(n3043), .B(n3044), .Z(n23172) );
  NANDN U4596 ( .A(n23199), .B(n4068), .Z(n3045) );
  NANDN U4597 ( .A(n23165), .B(n42115), .Z(n3046) );
  AND U4598 ( .A(n3045), .B(n3046), .Z(n23204) );
  NANDN U4599 ( .A(n23198), .B(n42047), .Z(n3047) );
  NANDN U4600 ( .A(n23235), .B(n4067), .Z(n3048) );
  NAND U4601 ( .A(n3047), .B(n3048), .Z(n23246) );
  NANDN U4602 ( .A(n23273), .B(n4068), .Z(n3049) );
  NANDN U4603 ( .A(n23239), .B(n42115), .Z(n3050) );
  AND U4604 ( .A(n3049), .B(n3050), .Z(n23278) );
  NANDN U4605 ( .A(n23272), .B(n42047), .Z(n3051) );
  NANDN U4606 ( .A(n23309), .B(n4067), .Z(n3052) );
  NAND U4607 ( .A(n3051), .B(n3052), .Z(n23320) );
  NANDN U4608 ( .A(n23350), .B(n4068), .Z(n3053) );
  NANDN U4609 ( .A(n23313), .B(n42115), .Z(n3054) );
  AND U4610 ( .A(n3053), .B(n3054), .Z(n23352) );
  NANDN U4611 ( .A(n23346), .B(n42047), .Z(n3055) );
  NANDN U4612 ( .A(n23383), .B(n4067), .Z(n3056) );
  NAND U4613 ( .A(n3055), .B(n3056), .Z(n23394) );
  NANDN U4614 ( .A(n23421), .B(n4068), .Z(n3057) );
  NANDN U4615 ( .A(n23384), .B(n42115), .Z(n3058) );
  AND U4616 ( .A(n3057), .B(n3058), .Z(n23426) );
  NANDN U4617 ( .A(n23420), .B(n42047), .Z(n3059) );
  NANDN U4618 ( .A(n23457), .B(n4067), .Z(n3060) );
  NAND U4619 ( .A(n3059), .B(n3060), .Z(n23468) );
  NANDN U4620 ( .A(n23498), .B(n4068), .Z(n3061) );
  NANDN U4621 ( .A(n23458), .B(n42115), .Z(n3062) );
  AND U4622 ( .A(n3061), .B(n3062), .Z(n23500) );
  NANDN U4623 ( .A(n23494), .B(n42047), .Z(n3063) );
  NANDN U4624 ( .A(n23531), .B(n4067), .Z(n3064) );
  NAND U4625 ( .A(n3063), .B(n3064), .Z(n23542) );
  NANDN U4626 ( .A(n23572), .B(n4068), .Z(n3065) );
  NANDN U4627 ( .A(n23535), .B(n42115), .Z(n3066) );
  AND U4628 ( .A(n3065), .B(n3066), .Z(n23574) );
  NANDN U4629 ( .A(n23568), .B(n42047), .Z(n3067) );
  NANDN U4630 ( .A(n23605), .B(n4067), .Z(n3068) );
  NAND U4631 ( .A(n3067), .B(n3068), .Z(n23616) );
  NANDN U4632 ( .A(n23646), .B(n4068), .Z(n3069) );
  NANDN U4633 ( .A(n23606), .B(n42115), .Z(n3070) );
  AND U4634 ( .A(n3069), .B(n3070), .Z(n23648) );
  NANDN U4635 ( .A(n23642), .B(n42047), .Z(n3071) );
  NANDN U4636 ( .A(n23679), .B(n4067), .Z(n3072) );
  NAND U4637 ( .A(n3071), .B(n3072), .Z(n23690) );
  NANDN U4638 ( .A(n23717), .B(n4068), .Z(n3073) );
  NANDN U4639 ( .A(n23683), .B(n42115), .Z(n3074) );
  AND U4640 ( .A(n3073), .B(n3074), .Z(n23722) );
  NANDN U4641 ( .A(n23716), .B(n42047), .Z(n3075) );
  NANDN U4642 ( .A(n23753), .B(n4067), .Z(n3076) );
  NAND U4643 ( .A(n3075), .B(n3076), .Z(n23764) );
  NANDN U4644 ( .A(n23794), .B(n4068), .Z(n3077) );
  NANDN U4645 ( .A(n23757), .B(n42115), .Z(n3078) );
  AND U4646 ( .A(n3077), .B(n3078), .Z(n23796) );
  NANDN U4647 ( .A(n23790), .B(n42047), .Z(n3079) );
  NANDN U4648 ( .A(n23827), .B(n4067), .Z(n3080) );
  NAND U4649 ( .A(n3079), .B(n3080), .Z(n23838) );
  NANDN U4650 ( .A(n23868), .B(n4068), .Z(n3081) );
  NANDN U4651 ( .A(n23828), .B(n42115), .Z(n3082) );
  AND U4652 ( .A(n3081), .B(n3082), .Z(n23870) );
  NANDN U4653 ( .A(n23864), .B(n42047), .Z(n3083) );
  NANDN U4654 ( .A(n23901), .B(n4067), .Z(n3084) );
  NAND U4655 ( .A(n3083), .B(n3084), .Z(n23912) );
  NANDN U4656 ( .A(n23939), .B(n4068), .Z(n3085) );
  NANDN U4657 ( .A(n23905), .B(n42115), .Z(n3086) );
  AND U4658 ( .A(n3085), .B(n3086), .Z(n23944) );
  NANDN U4659 ( .A(n23938), .B(n42047), .Z(n3087) );
  NANDN U4660 ( .A(n23975), .B(n4067), .Z(n3088) );
  NAND U4661 ( .A(n3087), .B(n3088), .Z(n23986) );
  NANDN U4662 ( .A(n24016), .B(n4068), .Z(n3089) );
  NANDN U4663 ( .A(n23979), .B(n42115), .Z(n3090) );
  AND U4664 ( .A(n3089), .B(n3090), .Z(n24018) );
  NANDN U4665 ( .A(n24012), .B(n42047), .Z(n3091) );
  NANDN U4666 ( .A(n24049), .B(n4067), .Z(n3092) );
  NAND U4667 ( .A(n3091), .B(n3092), .Z(n24060) );
  NANDN U4668 ( .A(n24087), .B(n4068), .Z(n3093) );
  NANDN U4669 ( .A(n24053), .B(n42115), .Z(n3094) );
  AND U4670 ( .A(n3093), .B(n3094), .Z(n24092) );
  NANDN U4671 ( .A(n24086), .B(n42047), .Z(n3095) );
  NANDN U4672 ( .A(n24123), .B(n4067), .Z(n3096) );
  NAND U4673 ( .A(n3095), .B(n3096), .Z(n24134) );
  NANDN U4674 ( .A(n24164), .B(n4068), .Z(n3097) );
  NANDN U4675 ( .A(n24124), .B(n42115), .Z(n3098) );
  AND U4676 ( .A(n3097), .B(n3098), .Z(n24166) );
  NANDN U4677 ( .A(n24160), .B(n42047), .Z(n3099) );
  NANDN U4678 ( .A(n24197), .B(n4067), .Z(n3100) );
  NAND U4679 ( .A(n3099), .B(n3100), .Z(n24208) );
  NANDN U4680 ( .A(n24238), .B(n4068), .Z(n3101) );
  NANDN U4681 ( .A(n24201), .B(n42115), .Z(n3102) );
  AND U4682 ( .A(n3101), .B(n3102), .Z(n24240) );
  NANDN U4683 ( .A(n24234), .B(n42047), .Z(n3103) );
  NANDN U4684 ( .A(n24271), .B(n4067), .Z(n3104) );
  NAND U4685 ( .A(n3103), .B(n3104), .Z(n24282) );
  NANDN U4686 ( .A(n24312), .B(n4068), .Z(n3105) );
  NANDN U4687 ( .A(n24275), .B(n42115), .Z(n3106) );
  AND U4688 ( .A(n3105), .B(n3106), .Z(n24314) );
  NANDN U4689 ( .A(n24308), .B(n42047), .Z(n3107) );
  NANDN U4690 ( .A(n24345), .B(n4067), .Z(n3108) );
  NAND U4691 ( .A(n3107), .B(n3108), .Z(n24356) );
  NANDN U4692 ( .A(n24386), .B(n4068), .Z(n3109) );
  NANDN U4693 ( .A(n24349), .B(n42115), .Z(n3110) );
  AND U4694 ( .A(n3109), .B(n3110), .Z(n24388) );
  NANDN U4695 ( .A(n24382), .B(n42047), .Z(n3111) );
  NANDN U4696 ( .A(n24419), .B(n4067), .Z(n3112) );
  NAND U4697 ( .A(n3111), .B(n3112), .Z(n24430) );
  NANDN U4698 ( .A(n24460), .B(n4068), .Z(n3113) );
  NANDN U4699 ( .A(n24423), .B(n42115), .Z(n3114) );
  AND U4700 ( .A(n3113), .B(n3114), .Z(n24462) );
  NANDN U4701 ( .A(n24456), .B(n42047), .Z(n3115) );
  NANDN U4702 ( .A(n24493), .B(n4067), .Z(n3116) );
  NAND U4703 ( .A(n3115), .B(n3116), .Z(n24504) );
  NANDN U4704 ( .A(n24531), .B(n4068), .Z(n3117) );
  NANDN U4705 ( .A(n24497), .B(n42115), .Z(n3118) );
  AND U4706 ( .A(n3117), .B(n3118), .Z(n24536) );
  NANDN U4707 ( .A(n24530), .B(n42047), .Z(n3119) );
  NANDN U4708 ( .A(n24567), .B(n4067), .Z(n3120) );
  NAND U4709 ( .A(n3119), .B(n3120), .Z(n24578) );
  NANDN U4710 ( .A(n24605), .B(n4068), .Z(n3121) );
  NANDN U4711 ( .A(n24571), .B(n42115), .Z(n3122) );
  AND U4712 ( .A(n3121), .B(n3122), .Z(n24610) );
  NANDN U4713 ( .A(n24604), .B(n42047), .Z(n3123) );
  NANDN U4714 ( .A(n24641), .B(n4067), .Z(n3124) );
  NAND U4715 ( .A(n3123), .B(n3124), .Z(n24652) );
  NANDN U4716 ( .A(n24682), .B(n4068), .Z(n3125) );
  NANDN U4717 ( .A(n24645), .B(n42115), .Z(n3126) );
  AND U4718 ( .A(n3125), .B(n3126), .Z(n24684) );
  NANDN U4719 ( .A(n24678), .B(n42047), .Z(n3127) );
  NANDN U4720 ( .A(n24715), .B(n4067), .Z(n3128) );
  NAND U4721 ( .A(n3127), .B(n3128), .Z(n24726) );
  NANDN U4722 ( .A(n24756), .B(n4068), .Z(n3129) );
  NANDN U4723 ( .A(n24716), .B(n42115), .Z(n3130) );
  AND U4724 ( .A(n3129), .B(n3130), .Z(n24758) );
  NANDN U4725 ( .A(n24752), .B(n42047), .Z(n3131) );
  NANDN U4726 ( .A(n24789), .B(n4067), .Z(n3132) );
  NAND U4727 ( .A(n3131), .B(n3132), .Z(n24800) );
  NANDN U4728 ( .A(n24830), .B(n4068), .Z(n3133) );
  NANDN U4729 ( .A(n24790), .B(n42115), .Z(n3134) );
  AND U4730 ( .A(n3133), .B(n3134), .Z(n24832) );
  NANDN U4731 ( .A(n24826), .B(n42047), .Z(n3135) );
  NANDN U4732 ( .A(n24863), .B(n4067), .Z(n3136) );
  NAND U4733 ( .A(n3135), .B(n3136), .Z(n24874) );
  NANDN U4734 ( .A(n24901), .B(n4068), .Z(n3137) );
  NANDN U4735 ( .A(n24867), .B(n42115), .Z(n3138) );
  AND U4736 ( .A(n3137), .B(n3138), .Z(n24906) );
  NANDN U4737 ( .A(n24900), .B(n42047), .Z(n3139) );
  NANDN U4738 ( .A(n24937), .B(n4067), .Z(n3140) );
  NAND U4739 ( .A(n3139), .B(n3140), .Z(n24948) );
  NANDN U4740 ( .A(n24978), .B(n4068), .Z(n3141) );
  NANDN U4741 ( .A(n24941), .B(n42115), .Z(n3142) );
  AND U4742 ( .A(n3141), .B(n3142), .Z(n24980) );
  NANDN U4743 ( .A(n24974), .B(n42047), .Z(n3143) );
  NANDN U4744 ( .A(n25011), .B(n4067), .Z(n3144) );
  NAND U4745 ( .A(n3143), .B(n3144), .Z(n25022) );
  NANDN U4746 ( .A(n25052), .B(n4068), .Z(n3145) );
  NANDN U4747 ( .A(n25015), .B(n42115), .Z(n3146) );
  AND U4748 ( .A(n3145), .B(n3146), .Z(n25054) );
  NANDN U4749 ( .A(n25048), .B(n42047), .Z(n3147) );
  NANDN U4750 ( .A(n25085), .B(n4067), .Z(n3148) );
  NAND U4751 ( .A(n3147), .B(n3148), .Z(n25096) );
  NANDN U4752 ( .A(n25126), .B(n4068), .Z(n3149) );
  NANDN U4753 ( .A(n25089), .B(n42115), .Z(n3150) );
  AND U4754 ( .A(n3149), .B(n3150), .Z(n25128) );
  NANDN U4755 ( .A(n25122), .B(n42047), .Z(n3151) );
  NANDN U4756 ( .A(n25159), .B(n4067), .Z(n3152) );
  NAND U4757 ( .A(n3151), .B(n3152), .Z(n25170) );
  NANDN U4758 ( .A(n25200), .B(n4068), .Z(n3153) );
  NANDN U4759 ( .A(n25163), .B(n42115), .Z(n3154) );
  AND U4760 ( .A(n3153), .B(n3154), .Z(n25202) );
  NANDN U4761 ( .A(n25196), .B(n42047), .Z(n3155) );
  NANDN U4762 ( .A(n25233), .B(n4067), .Z(n3156) );
  NAND U4763 ( .A(n3155), .B(n3156), .Z(n25244) );
  NANDN U4764 ( .A(n25271), .B(n4068), .Z(n3157) );
  NANDN U4765 ( .A(n25234), .B(n42115), .Z(n3158) );
  AND U4766 ( .A(n3157), .B(n3158), .Z(n25276) );
  NANDN U4767 ( .A(n25270), .B(n42047), .Z(n3159) );
  NANDN U4768 ( .A(n25307), .B(n4067), .Z(n3160) );
  NAND U4769 ( .A(n3159), .B(n3160), .Z(n25318) );
  NANDN U4770 ( .A(n25348), .B(n4068), .Z(n3161) );
  NANDN U4771 ( .A(n25311), .B(n42115), .Z(n3162) );
  AND U4772 ( .A(n3161), .B(n3162), .Z(n25350) );
  NANDN U4773 ( .A(n25344), .B(n42047), .Z(n3163) );
  NANDN U4774 ( .A(n25381), .B(n4067), .Z(n3164) );
  NAND U4775 ( .A(n3163), .B(n3164), .Z(n25392) );
  NANDN U4776 ( .A(n25422), .B(n4068), .Z(n3165) );
  NANDN U4777 ( .A(n25382), .B(n42115), .Z(n3166) );
  AND U4778 ( .A(n3165), .B(n3166), .Z(n25424) );
  NANDN U4779 ( .A(n25418), .B(n42047), .Z(n3167) );
  NANDN U4780 ( .A(n25455), .B(n4067), .Z(n3168) );
  NAND U4781 ( .A(n3167), .B(n3168), .Z(n25466) );
  NANDN U4782 ( .A(n25493), .B(n4068), .Z(n3169) );
  NANDN U4783 ( .A(n25459), .B(n42115), .Z(n3170) );
  AND U4784 ( .A(n3169), .B(n3170), .Z(n25498) );
  NANDN U4785 ( .A(n25492), .B(n42047), .Z(n3171) );
  NANDN U4786 ( .A(n25529), .B(n4067), .Z(n3172) );
  NAND U4787 ( .A(n3171), .B(n3172), .Z(n25540) );
  NANDN U4788 ( .A(n25567), .B(n4068), .Z(n3173) );
  NANDN U4789 ( .A(n25530), .B(n42115), .Z(n3174) );
  AND U4790 ( .A(n3173), .B(n3174), .Z(n25572) );
  NANDN U4791 ( .A(n25566), .B(n42047), .Z(n3175) );
  NANDN U4792 ( .A(n25603), .B(n4067), .Z(n3176) );
  NAND U4793 ( .A(n3175), .B(n3176), .Z(n25614) );
  NANDN U4794 ( .A(n25644), .B(n4068), .Z(n3177) );
  NANDN U4795 ( .A(n25604), .B(n42115), .Z(n3178) );
  AND U4796 ( .A(n3177), .B(n3178), .Z(n25646) );
  NANDN U4797 ( .A(n25640), .B(n42047), .Z(n3179) );
  NANDN U4798 ( .A(n25677), .B(n4067), .Z(n3180) );
  NAND U4799 ( .A(n3179), .B(n3180), .Z(n25688) );
  NANDN U4800 ( .A(n25718), .B(n4068), .Z(n3181) );
  NANDN U4801 ( .A(n25681), .B(n42115), .Z(n3182) );
  AND U4802 ( .A(n3181), .B(n3182), .Z(n25720) );
  NANDN U4803 ( .A(n25714), .B(n42047), .Z(n3183) );
  NANDN U4804 ( .A(n25751), .B(n4067), .Z(n3184) );
  NAND U4805 ( .A(n3183), .B(n3184), .Z(n25762) );
  NANDN U4806 ( .A(n25789), .B(n4068), .Z(n3185) );
  NANDN U4807 ( .A(n25755), .B(n42115), .Z(n3186) );
  AND U4808 ( .A(n3185), .B(n3186), .Z(n25794) );
  NANDN U4809 ( .A(n25788), .B(n42047), .Z(n3187) );
  NANDN U4810 ( .A(n25825), .B(n4067), .Z(n3188) );
  NAND U4811 ( .A(n3187), .B(n3188), .Z(n25836) );
  NANDN U4812 ( .A(n25866), .B(n4068), .Z(n3189) );
  NANDN U4813 ( .A(n25829), .B(n42115), .Z(n3190) );
  AND U4814 ( .A(n3189), .B(n3190), .Z(n25868) );
  NANDN U4815 ( .A(n25862), .B(n42047), .Z(n3191) );
  NANDN U4816 ( .A(n25899), .B(n4067), .Z(n3192) );
  NAND U4817 ( .A(n3191), .B(n3192), .Z(n25910) );
  NANDN U4818 ( .A(n25940), .B(n4068), .Z(n3193) );
  NANDN U4819 ( .A(n25900), .B(n42115), .Z(n3194) );
  AND U4820 ( .A(n3193), .B(n3194), .Z(n25942) );
  NANDN U4821 ( .A(n25936), .B(n42047), .Z(n3195) );
  NANDN U4822 ( .A(n25973), .B(n4067), .Z(n3196) );
  NAND U4823 ( .A(n3195), .B(n3196), .Z(n25984) );
  NANDN U4824 ( .A(n26014), .B(n4068), .Z(n3197) );
  NANDN U4825 ( .A(n25974), .B(n42115), .Z(n3198) );
  AND U4826 ( .A(n3197), .B(n3198), .Z(n26016) );
  NANDN U4827 ( .A(n26010), .B(n42047), .Z(n3199) );
  NANDN U4828 ( .A(n26047), .B(n4067), .Z(n3200) );
  NAND U4829 ( .A(n3199), .B(n3200), .Z(n26058) );
  NANDN U4830 ( .A(n26088), .B(n4068), .Z(n3201) );
  NANDN U4831 ( .A(n26051), .B(n42115), .Z(n3202) );
  AND U4832 ( .A(n3201), .B(n3202), .Z(n26090) );
  NANDN U4833 ( .A(n26084), .B(n42047), .Z(n3203) );
  NANDN U4834 ( .A(n26121), .B(n4067), .Z(n3204) );
  NAND U4835 ( .A(n3203), .B(n3204), .Z(n26132) );
  NANDN U4836 ( .A(n26159), .B(n4068), .Z(n3205) );
  NANDN U4837 ( .A(n26125), .B(n42115), .Z(n3206) );
  AND U4838 ( .A(n3205), .B(n3206), .Z(n26164) );
  NANDN U4839 ( .A(n26158), .B(n42047), .Z(n3207) );
  NANDN U4840 ( .A(n26195), .B(n4067), .Z(n3208) );
  NAND U4841 ( .A(n3207), .B(n3208), .Z(n26206) );
  NANDN U4842 ( .A(n26233), .B(n4068), .Z(n3209) );
  NANDN U4843 ( .A(n26199), .B(n42115), .Z(n3210) );
  AND U4844 ( .A(n3209), .B(n3210), .Z(n26238) );
  NANDN U4845 ( .A(n26232), .B(n42047), .Z(n3211) );
  NANDN U4846 ( .A(n26269), .B(n4067), .Z(n3212) );
  NAND U4847 ( .A(n3211), .B(n3212), .Z(n26280) );
  NANDN U4848 ( .A(n26310), .B(n4068), .Z(n3213) );
  NANDN U4849 ( .A(n26273), .B(n42115), .Z(n3214) );
  AND U4850 ( .A(n3213), .B(n3214), .Z(n26312) );
  NANDN U4851 ( .A(n26306), .B(n42047), .Z(n3215) );
  NANDN U4852 ( .A(n26343), .B(n4067), .Z(n3216) );
  NAND U4853 ( .A(n3215), .B(n3216), .Z(n26354) );
  NANDN U4854 ( .A(n26381), .B(n4068), .Z(n3217) );
  NANDN U4855 ( .A(n26347), .B(n42115), .Z(n3218) );
  AND U4856 ( .A(n3217), .B(n3218), .Z(n26386) );
  NANDN U4857 ( .A(n26380), .B(n42047), .Z(n3219) );
  NANDN U4858 ( .A(n26417), .B(n4067), .Z(n3220) );
  NAND U4859 ( .A(n3219), .B(n3220), .Z(n26428) );
  NANDN U4860 ( .A(n26455), .B(n4068), .Z(n3221) );
  NANDN U4861 ( .A(n26421), .B(n42115), .Z(n3222) );
  AND U4862 ( .A(n3221), .B(n3222), .Z(n26460) );
  NANDN U4863 ( .A(n26454), .B(n42047), .Z(n3223) );
  NANDN U4864 ( .A(n26491), .B(n4067), .Z(n3224) );
  NAND U4865 ( .A(n3223), .B(n3224), .Z(n26502) );
  NANDN U4866 ( .A(n26532), .B(n4068), .Z(n3225) );
  NANDN U4867 ( .A(n26495), .B(n42115), .Z(n3226) );
  AND U4868 ( .A(n3225), .B(n3226), .Z(n26534) );
  NANDN U4869 ( .A(n26528), .B(n42047), .Z(n3227) );
  NANDN U4870 ( .A(n26565), .B(n4067), .Z(n3228) );
  NAND U4871 ( .A(n3227), .B(n3228), .Z(n26576) );
  NANDN U4872 ( .A(n26603), .B(n4068), .Z(n3229) );
  NANDN U4873 ( .A(n26569), .B(n42115), .Z(n3230) );
  AND U4874 ( .A(n3229), .B(n3230), .Z(n26608) );
  NANDN U4875 ( .A(n26602), .B(n42047), .Z(n3231) );
  NANDN U4876 ( .A(n26639), .B(n4067), .Z(n3232) );
  NAND U4877 ( .A(n3231), .B(n3232), .Z(n26650) );
  NANDN U4878 ( .A(n26680), .B(n4068), .Z(n3233) );
  NANDN U4879 ( .A(n26640), .B(n42115), .Z(n3234) );
  AND U4880 ( .A(n3233), .B(n3234), .Z(n26682) );
  NANDN U4881 ( .A(n26676), .B(n42047), .Z(n3235) );
  NANDN U4882 ( .A(n26713), .B(n4067), .Z(n3236) );
  NAND U4883 ( .A(n3235), .B(n3236), .Z(n26724) );
  NANDN U4884 ( .A(n26751), .B(n4068), .Z(n3237) );
  NANDN U4885 ( .A(n26717), .B(n42115), .Z(n3238) );
  AND U4886 ( .A(n3237), .B(n3238), .Z(n26756) );
  NANDN U4887 ( .A(n26750), .B(n42047), .Z(n3239) );
  NANDN U4888 ( .A(n26787), .B(n4067), .Z(n3240) );
  NAND U4889 ( .A(n3239), .B(n3240), .Z(n26798) );
  NANDN U4890 ( .A(n26828), .B(n4068), .Z(n3241) );
  NANDN U4891 ( .A(n26788), .B(n42115), .Z(n3242) );
  AND U4892 ( .A(n3241), .B(n3242), .Z(n26830) );
  NANDN U4893 ( .A(n26824), .B(n42047), .Z(n3243) );
  NANDN U4894 ( .A(n26861), .B(n4067), .Z(n3244) );
  NAND U4895 ( .A(n3243), .B(n3244), .Z(n26872) );
  NANDN U4896 ( .A(n26902), .B(n4068), .Z(n3245) );
  NANDN U4897 ( .A(n26865), .B(n42115), .Z(n3246) );
  AND U4898 ( .A(n3245), .B(n3246), .Z(n26904) );
  NANDN U4899 ( .A(n26898), .B(n42047), .Z(n3247) );
  NANDN U4900 ( .A(n26935), .B(n4067), .Z(n3248) );
  NAND U4901 ( .A(n3247), .B(n3248), .Z(n26946) );
  NANDN U4902 ( .A(n26976), .B(n4068), .Z(n3249) );
  NANDN U4903 ( .A(n26939), .B(n42115), .Z(n3250) );
  AND U4904 ( .A(n3249), .B(n3250), .Z(n26978) );
  NANDN U4905 ( .A(n26972), .B(n42047), .Z(n3251) );
  NANDN U4906 ( .A(n27009), .B(n4067), .Z(n3252) );
  NAND U4907 ( .A(n3251), .B(n3252), .Z(n27020) );
  NANDN U4908 ( .A(n27050), .B(n4068), .Z(n3253) );
  NANDN U4909 ( .A(n27010), .B(n42115), .Z(n3254) );
  AND U4910 ( .A(n3253), .B(n3254), .Z(n27052) );
  NANDN U4911 ( .A(n27046), .B(n42047), .Z(n3255) );
  NANDN U4912 ( .A(n27083), .B(n4067), .Z(n3256) );
  NAND U4913 ( .A(n3255), .B(n3256), .Z(n27094) );
  NANDN U4914 ( .A(n27124), .B(n4068), .Z(n3257) );
  NANDN U4915 ( .A(n27084), .B(n42115), .Z(n3258) );
  AND U4916 ( .A(n3257), .B(n3258), .Z(n27126) );
  NANDN U4917 ( .A(n27120), .B(n42047), .Z(n3259) );
  NANDN U4918 ( .A(n27157), .B(n4067), .Z(n3260) );
  NAND U4919 ( .A(n3259), .B(n3260), .Z(n27168) );
  NANDN U4920 ( .A(n27198), .B(n4068), .Z(n3261) );
  NANDN U4921 ( .A(n27158), .B(n42115), .Z(n3262) );
  AND U4922 ( .A(n3261), .B(n3262), .Z(n27200) );
  NANDN U4923 ( .A(n27194), .B(n42047), .Z(n3263) );
  NANDN U4924 ( .A(n27231), .B(n4067), .Z(n3264) );
  NAND U4925 ( .A(n3263), .B(n3264), .Z(n27242) );
  NANDN U4926 ( .A(n27272), .B(n4068), .Z(n3265) );
  NANDN U4927 ( .A(n27235), .B(n42115), .Z(n3266) );
  AND U4928 ( .A(n3265), .B(n3266), .Z(n27274) );
  NANDN U4929 ( .A(n27268), .B(n42047), .Z(n3267) );
  NANDN U4930 ( .A(n27305), .B(n4067), .Z(n3268) );
  NAND U4931 ( .A(n3267), .B(n3268), .Z(n27316) );
  NANDN U4932 ( .A(n27346), .B(n4068), .Z(n3269) );
  NANDN U4933 ( .A(n27306), .B(n42115), .Z(n3270) );
  AND U4934 ( .A(n3269), .B(n3270), .Z(n27348) );
  NANDN U4935 ( .A(n27342), .B(n42047), .Z(n3271) );
  NANDN U4936 ( .A(n27379), .B(n4067), .Z(n3272) );
  NAND U4937 ( .A(n3271), .B(n3272), .Z(n27390) );
  NANDN U4938 ( .A(n27420), .B(n4068), .Z(n3273) );
  NANDN U4939 ( .A(n27383), .B(n42115), .Z(n3274) );
  AND U4940 ( .A(n3273), .B(n3274), .Z(n27422) );
  NANDN U4941 ( .A(n27416), .B(n42047), .Z(n3275) );
  NANDN U4942 ( .A(n27453), .B(n4067), .Z(n3276) );
  NAND U4943 ( .A(n3275), .B(n3276), .Z(n27464) );
  NANDN U4944 ( .A(n27494), .B(n4068), .Z(n3277) );
  NANDN U4945 ( .A(n27457), .B(n42115), .Z(n3278) );
  AND U4946 ( .A(n3277), .B(n3278), .Z(n27496) );
  NANDN U4947 ( .A(n27490), .B(n42047), .Z(n3279) );
  NANDN U4948 ( .A(n27527), .B(n4067), .Z(n3280) );
  NAND U4949 ( .A(n3279), .B(n3280), .Z(n27538) );
  NANDN U4950 ( .A(n27568), .B(n4068), .Z(n3281) );
  NANDN U4951 ( .A(n27531), .B(n42115), .Z(n3282) );
  AND U4952 ( .A(n3281), .B(n3282), .Z(n27570) );
  NANDN U4953 ( .A(n27564), .B(n42047), .Z(n3283) );
  NANDN U4954 ( .A(n27601), .B(n4067), .Z(n3284) );
  NAND U4955 ( .A(n3283), .B(n3284), .Z(n27612) );
  NANDN U4956 ( .A(n27642), .B(n4068), .Z(n3285) );
  NANDN U4957 ( .A(n27605), .B(n42115), .Z(n3286) );
  AND U4958 ( .A(n3285), .B(n3286), .Z(n27644) );
  NANDN U4959 ( .A(n27638), .B(n42047), .Z(n3287) );
  NANDN U4960 ( .A(n27675), .B(n4067), .Z(n3288) );
  NAND U4961 ( .A(n3287), .B(n3288), .Z(n27686) );
  NANDN U4962 ( .A(n27716), .B(n4068), .Z(n3289) );
  NANDN U4963 ( .A(n27676), .B(n42115), .Z(n3290) );
  AND U4964 ( .A(n3289), .B(n3290), .Z(n27718) );
  NANDN U4965 ( .A(n27712), .B(n42047), .Z(n3291) );
  NANDN U4966 ( .A(n27749), .B(n4067), .Z(n3292) );
  NAND U4967 ( .A(n3291), .B(n3292), .Z(n27760) );
  NANDN U4968 ( .A(n27790), .B(n4068), .Z(n3293) );
  NANDN U4969 ( .A(n27750), .B(n42115), .Z(n3294) );
  AND U4970 ( .A(n3293), .B(n3294), .Z(n27792) );
  NANDN U4971 ( .A(n27786), .B(n42047), .Z(n3295) );
  NANDN U4972 ( .A(n27823), .B(n4067), .Z(n3296) );
  NAND U4973 ( .A(n3295), .B(n3296), .Z(n27834) );
  NANDN U4974 ( .A(n27864), .B(n4068), .Z(n3297) );
  NANDN U4975 ( .A(n27827), .B(n42115), .Z(n3298) );
  AND U4976 ( .A(n3297), .B(n3298), .Z(n27866) );
  NANDN U4977 ( .A(n27860), .B(n42047), .Z(n3299) );
  NANDN U4978 ( .A(n27897), .B(n4067), .Z(n3300) );
  NAND U4979 ( .A(n3299), .B(n3300), .Z(n27908) );
  NANDN U4980 ( .A(n27935), .B(n4068), .Z(n3301) );
  NANDN U4981 ( .A(n27898), .B(n42115), .Z(n3302) );
  AND U4982 ( .A(n3301), .B(n3302), .Z(n27940) );
  NANDN U4983 ( .A(n27934), .B(n42047), .Z(n3303) );
  NANDN U4984 ( .A(n27971), .B(n4067), .Z(n3304) );
  NAND U4985 ( .A(n3303), .B(n3304), .Z(n27982) );
  NANDN U4986 ( .A(n28012), .B(n4068), .Z(n3305) );
  NANDN U4987 ( .A(n27972), .B(n42115), .Z(n3306) );
  AND U4988 ( .A(n3305), .B(n3306), .Z(n28014) );
  NANDN U4989 ( .A(n28008), .B(n42047), .Z(n3307) );
  NANDN U4990 ( .A(n28045), .B(n4067), .Z(n3308) );
  NAND U4991 ( .A(n3307), .B(n3308), .Z(n28056) );
  NANDN U4992 ( .A(n28086), .B(n4068), .Z(n3309) );
  NANDN U4993 ( .A(n28046), .B(n42115), .Z(n3310) );
  AND U4994 ( .A(n3309), .B(n3310), .Z(n28088) );
  NANDN U4995 ( .A(n28082), .B(n42047), .Z(n3311) );
  NANDN U4996 ( .A(n28119), .B(n4067), .Z(n3312) );
  NAND U4997 ( .A(n3311), .B(n3312), .Z(n28130) );
  NANDN U4998 ( .A(n28160), .B(n4068), .Z(n3313) );
  NANDN U4999 ( .A(n28123), .B(n42115), .Z(n3314) );
  AND U5000 ( .A(n3313), .B(n3314), .Z(n28162) );
  NANDN U5001 ( .A(n28156), .B(n42047), .Z(n3315) );
  NANDN U5002 ( .A(n28193), .B(n4067), .Z(n3316) );
  NAND U5003 ( .A(n3315), .B(n3316), .Z(n28204) );
  NANDN U5004 ( .A(n28234), .B(n4068), .Z(n3317) );
  NANDN U5005 ( .A(n28197), .B(n42115), .Z(n3318) );
  AND U5006 ( .A(n3317), .B(n3318), .Z(n28236) );
  NANDN U5007 ( .A(n28230), .B(n42047), .Z(n3319) );
  NANDN U5008 ( .A(n28267), .B(n4067), .Z(n3320) );
  NAND U5009 ( .A(n3319), .B(n3320), .Z(n28278) );
  NANDN U5010 ( .A(n28308), .B(n4068), .Z(n3321) );
  NANDN U5011 ( .A(n28271), .B(n42115), .Z(n3322) );
  AND U5012 ( .A(n3321), .B(n3322), .Z(n28310) );
  NANDN U5013 ( .A(n28304), .B(n42047), .Z(n3323) );
  NANDN U5014 ( .A(n28341), .B(n4067), .Z(n3324) );
  NAND U5015 ( .A(n3323), .B(n3324), .Z(n28352) );
  NANDN U5016 ( .A(n28382), .B(n4068), .Z(n3325) );
  NANDN U5017 ( .A(n28345), .B(n42115), .Z(n3326) );
  AND U5018 ( .A(n3325), .B(n3326), .Z(n28384) );
  NANDN U5019 ( .A(n28378), .B(n42047), .Z(n3327) );
  NANDN U5020 ( .A(n28415), .B(n4067), .Z(n3328) );
  NAND U5021 ( .A(n3327), .B(n3328), .Z(n28426) );
  NANDN U5022 ( .A(n28453), .B(n4068), .Z(n3329) );
  NANDN U5023 ( .A(n28416), .B(n42115), .Z(n3330) );
  AND U5024 ( .A(n3329), .B(n3330), .Z(n28458) );
  NANDN U5025 ( .A(n28452), .B(n42047), .Z(n3331) );
  NANDN U5026 ( .A(n28489), .B(n4067), .Z(n3332) );
  NAND U5027 ( .A(n3331), .B(n3332), .Z(n28500) );
  NANDN U5028 ( .A(n28530), .B(n4068), .Z(n3333) );
  NANDN U5029 ( .A(n28493), .B(n42115), .Z(n3334) );
  AND U5030 ( .A(n3333), .B(n3334), .Z(n28532) );
  NANDN U5031 ( .A(n28526), .B(n42047), .Z(n3335) );
  NANDN U5032 ( .A(n28563), .B(n4067), .Z(n3336) );
  NAND U5033 ( .A(n3335), .B(n3336), .Z(n28574) );
  NANDN U5034 ( .A(n28604), .B(n4068), .Z(n3337) );
  NANDN U5035 ( .A(n28564), .B(n42115), .Z(n3338) );
  AND U5036 ( .A(n3337), .B(n3338), .Z(n28606) );
  NANDN U5037 ( .A(n28600), .B(n42047), .Z(n3339) );
  NANDN U5038 ( .A(n28637), .B(n4067), .Z(n3340) );
  NAND U5039 ( .A(n3339), .B(n3340), .Z(n28648) );
  NANDN U5040 ( .A(n28678), .B(n4068), .Z(n3341) );
  NANDN U5041 ( .A(n28641), .B(n42115), .Z(n3342) );
  AND U5042 ( .A(n3341), .B(n3342), .Z(n28680) );
  NANDN U5043 ( .A(n28674), .B(n42047), .Z(n3343) );
  NANDN U5044 ( .A(n28711), .B(n4067), .Z(n3344) );
  NAND U5045 ( .A(n3343), .B(n3344), .Z(n28722) );
  NANDN U5046 ( .A(n28752), .B(n4068), .Z(n3345) );
  NANDN U5047 ( .A(n28715), .B(n42115), .Z(n3346) );
  AND U5048 ( .A(n3345), .B(n3346), .Z(n28754) );
  NANDN U5049 ( .A(n28748), .B(n42047), .Z(n3347) );
  NANDN U5050 ( .A(n28785), .B(n4067), .Z(n3348) );
  NAND U5051 ( .A(n3347), .B(n3348), .Z(n28796) );
  NANDN U5052 ( .A(n28823), .B(n4068), .Z(n3349) );
  NANDN U5053 ( .A(n28789), .B(n42115), .Z(n3350) );
  AND U5054 ( .A(n3349), .B(n3350), .Z(n28828) );
  NANDN U5055 ( .A(n28822), .B(n42047), .Z(n3351) );
  NANDN U5056 ( .A(n28859), .B(n4067), .Z(n3352) );
  NAND U5057 ( .A(n3351), .B(n3352), .Z(n28870) );
  NANDN U5058 ( .A(n28900), .B(n4068), .Z(n3353) );
  NANDN U5059 ( .A(n28860), .B(n42115), .Z(n3354) );
  AND U5060 ( .A(n3353), .B(n3354), .Z(n28902) );
  NANDN U5061 ( .A(n28896), .B(n42047), .Z(n3355) );
  NANDN U5062 ( .A(n28933), .B(n4067), .Z(n3356) );
  NAND U5063 ( .A(n3355), .B(n3356), .Z(n28944) );
  NANDN U5064 ( .A(n28974), .B(n4068), .Z(n3357) );
  NANDN U5065 ( .A(n28934), .B(n42115), .Z(n3358) );
  AND U5066 ( .A(n3357), .B(n3358), .Z(n28976) );
  NANDN U5067 ( .A(n28970), .B(n42047), .Z(n3359) );
  NANDN U5068 ( .A(n29007), .B(n4067), .Z(n3360) );
  NAND U5069 ( .A(n3359), .B(n3360), .Z(n29018) );
  NANDN U5070 ( .A(n29045), .B(n4068), .Z(n3361) );
  NANDN U5071 ( .A(n29011), .B(n42115), .Z(n3362) );
  AND U5072 ( .A(n3361), .B(n3362), .Z(n29050) );
  NANDN U5073 ( .A(n29044), .B(n42047), .Z(n3363) );
  NANDN U5074 ( .A(n29081), .B(n4067), .Z(n3364) );
  NAND U5075 ( .A(n3363), .B(n3364), .Z(n29092) );
  NANDN U5076 ( .A(n29122), .B(n4068), .Z(n3365) );
  NANDN U5077 ( .A(n29082), .B(n42115), .Z(n3366) );
  AND U5078 ( .A(n3365), .B(n3366), .Z(n29124) );
  NANDN U5079 ( .A(n29118), .B(n42047), .Z(n3367) );
  NANDN U5080 ( .A(n29155), .B(n4067), .Z(n3368) );
  NAND U5081 ( .A(n3367), .B(n3368), .Z(n29166) );
  NANDN U5082 ( .A(n29196), .B(n4068), .Z(n3369) );
  NANDN U5083 ( .A(n29159), .B(n42115), .Z(n3370) );
  AND U5084 ( .A(n3369), .B(n3370), .Z(n29198) );
  NANDN U5085 ( .A(n29192), .B(n42047), .Z(n3371) );
  NANDN U5086 ( .A(n29229), .B(n4067), .Z(n3372) );
  NAND U5087 ( .A(n3371), .B(n3372), .Z(n29240) );
  NANDN U5088 ( .A(n29270), .B(n4068), .Z(n3373) );
  NANDN U5089 ( .A(n29230), .B(n42115), .Z(n3374) );
  AND U5090 ( .A(n3373), .B(n3374), .Z(n29272) );
  NANDN U5091 ( .A(n29266), .B(n42047), .Z(n3375) );
  NANDN U5092 ( .A(n29303), .B(n4067), .Z(n3376) );
  NAND U5093 ( .A(n3375), .B(n3376), .Z(n29314) );
  NANDN U5094 ( .A(n29344), .B(n4068), .Z(n3377) );
  NANDN U5095 ( .A(n29307), .B(n42115), .Z(n3378) );
  AND U5096 ( .A(n3377), .B(n3378), .Z(n29346) );
  NANDN U5097 ( .A(n29340), .B(n42047), .Z(n3379) );
  NANDN U5098 ( .A(n29377), .B(n4067), .Z(n3380) );
  NAND U5099 ( .A(n3379), .B(n3380), .Z(n29388) );
  NANDN U5100 ( .A(n29418), .B(n4068), .Z(n3381) );
  NANDN U5101 ( .A(n29381), .B(n42115), .Z(n3382) );
  AND U5102 ( .A(n3381), .B(n3382), .Z(n29420) );
  NANDN U5103 ( .A(n29414), .B(n42047), .Z(n3383) );
  NANDN U5104 ( .A(n29451), .B(n4067), .Z(n3384) );
  NAND U5105 ( .A(n3383), .B(n3384), .Z(n29462) );
  NANDN U5106 ( .A(n29489), .B(n4068), .Z(n3385) );
  NANDN U5107 ( .A(n29455), .B(n42115), .Z(n3386) );
  AND U5108 ( .A(n3385), .B(n3386), .Z(n29494) );
  NANDN U5109 ( .A(n29488), .B(n42047), .Z(n3387) );
  NANDN U5110 ( .A(n29525), .B(n4067), .Z(n3388) );
  NAND U5111 ( .A(n3387), .B(n3388), .Z(n29536) );
  NANDN U5112 ( .A(n29567), .B(n4068), .Z(n3389) );
  NANDN U5113 ( .A(n29526), .B(n42115), .Z(n3390) );
  AND U5114 ( .A(n3389), .B(n3390), .Z(n29569) );
  NANDN U5115 ( .A(n29562), .B(n42047), .Z(n3391) );
  NANDN U5116 ( .A(n29600), .B(n4067), .Z(n3392) );
  NAND U5117 ( .A(n3391), .B(n3392), .Z(n29611) );
  NANDN U5118 ( .A(n29641), .B(n4068), .Z(n3393) );
  NANDN U5119 ( .A(n29604), .B(n42115), .Z(n3394) );
  AND U5120 ( .A(n3393), .B(n3394), .Z(n29643) );
  NANDN U5121 ( .A(n29637), .B(n42047), .Z(n3395) );
  NANDN U5122 ( .A(n29674), .B(n4067), .Z(n3396) );
  NAND U5123 ( .A(n3395), .B(n3396), .Z(n29685) );
  NANDN U5124 ( .A(n29712), .B(n4068), .Z(n3397) );
  NANDN U5125 ( .A(n29678), .B(n42115), .Z(n3398) );
  AND U5126 ( .A(n3397), .B(n3398), .Z(n29717) );
  NANDN U5127 ( .A(n29711), .B(n42047), .Z(n3399) );
  NANDN U5128 ( .A(n29748), .B(n4067), .Z(n3400) );
  NAND U5129 ( .A(n3399), .B(n3400), .Z(n29759) );
  NANDN U5130 ( .A(n29786), .B(n4068), .Z(n3401) );
  NANDN U5131 ( .A(n29752), .B(n42115), .Z(n3402) );
  AND U5132 ( .A(n3401), .B(n3402), .Z(n29791) );
  NANDN U5133 ( .A(n29785), .B(n42047), .Z(n3403) );
  NANDN U5134 ( .A(n29822), .B(n4067), .Z(n3404) );
  NAND U5135 ( .A(n3403), .B(n3404), .Z(n29833) );
  NANDN U5136 ( .A(n29863), .B(n4068), .Z(n3405) );
  NANDN U5137 ( .A(n29826), .B(n42115), .Z(n3406) );
  AND U5138 ( .A(n3405), .B(n3406), .Z(n29865) );
  NANDN U5139 ( .A(n29859), .B(n42047), .Z(n3407) );
  NANDN U5140 ( .A(n29896), .B(n4067), .Z(n3408) );
  NAND U5141 ( .A(n3407), .B(n3408), .Z(n29907) );
  NANDN U5142 ( .A(n29934), .B(n4068), .Z(n3409) );
  NANDN U5143 ( .A(n29897), .B(n42115), .Z(n3410) );
  AND U5144 ( .A(n3409), .B(n3410), .Z(n29939) );
  NANDN U5145 ( .A(n29933), .B(n42047), .Z(n3411) );
  NANDN U5146 ( .A(n29970), .B(n4067), .Z(n3412) );
  NAND U5147 ( .A(n3411), .B(n3412), .Z(n29981) );
  NANDN U5148 ( .A(n30011), .B(n4068), .Z(n3413) );
  NANDN U5149 ( .A(n29974), .B(n42115), .Z(n3414) );
  AND U5150 ( .A(n3413), .B(n3414), .Z(n30013) );
  NANDN U5151 ( .A(n30007), .B(n42047), .Z(n3415) );
  NANDN U5152 ( .A(n30044), .B(n4067), .Z(n3416) );
  NAND U5153 ( .A(n3415), .B(n3416), .Z(n30055) );
  NANDN U5154 ( .A(n30085), .B(n4068), .Z(n3417) );
  NANDN U5155 ( .A(n30045), .B(n42115), .Z(n3418) );
  AND U5156 ( .A(n3417), .B(n3418), .Z(n30087) );
  NANDN U5157 ( .A(n30081), .B(n42047), .Z(n3419) );
  NANDN U5158 ( .A(n30118), .B(n4067), .Z(n3420) );
  NAND U5159 ( .A(n3419), .B(n3420), .Z(n30129) );
  NANDN U5160 ( .A(n30159), .B(n4068), .Z(n3421) );
  NANDN U5161 ( .A(n30122), .B(n42115), .Z(n3422) );
  AND U5162 ( .A(n3421), .B(n3422), .Z(n30161) );
  NANDN U5163 ( .A(n30155), .B(n42047), .Z(n3423) );
  NANDN U5164 ( .A(n30192), .B(n4067), .Z(n3424) );
  NAND U5165 ( .A(n3423), .B(n3424), .Z(n30203) );
  NANDN U5166 ( .A(n30230), .B(n4068), .Z(n3425) );
  NANDN U5167 ( .A(n30193), .B(n42115), .Z(n3426) );
  AND U5168 ( .A(n3425), .B(n3426), .Z(n30235) );
  NANDN U5169 ( .A(n30229), .B(n42047), .Z(n3427) );
  NANDN U5170 ( .A(n30266), .B(n4067), .Z(n3428) );
  NAND U5171 ( .A(n3427), .B(n3428), .Z(n30277) );
  NANDN U5172 ( .A(n30304), .B(n4068), .Z(n3429) );
  NANDN U5173 ( .A(n30270), .B(n42115), .Z(n3430) );
  AND U5174 ( .A(n3429), .B(n3430), .Z(n30309) );
  NANDN U5175 ( .A(n30303), .B(n42047), .Z(n3431) );
  NANDN U5176 ( .A(n30340), .B(n4067), .Z(n3432) );
  NAND U5177 ( .A(n3431), .B(n3432), .Z(n30351) );
  NANDN U5178 ( .A(n30381), .B(n4068), .Z(n3433) );
  NANDN U5179 ( .A(n30344), .B(n42115), .Z(n3434) );
  AND U5180 ( .A(n3433), .B(n3434), .Z(n30383) );
  NANDN U5181 ( .A(n30377), .B(n42047), .Z(n3435) );
  NANDN U5182 ( .A(n30414), .B(n4067), .Z(n3436) );
  NAND U5183 ( .A(n3435), .B(n3436), .Z(n30425) );
  NANDN U5184 ( .A(n30452), .B(n4068), .Z(n3437) );
  NANDN U5185 ( .A(n30418), .B(n42115), .Z(n3438) );
  AND U5186 ( .A(n3437), .B(n3438), .Z(n30457) );
  NANDN U5187 ( .A(n30451), .B(n42047), .Z(n3439) );
  NANDN U5188 ( .A(n30488), .B(n4067), .Z(n3440) );
  NAND U5189 ( .A(n3439), .B(n3440), .Z(n30499) );
  NANDN U5190 ( .A(n30529), .B(n4068), .Z(n3441) );
  NANDN U5191 ( .A(n30492), .B(n42115), .Z(n3442) );
  AND U5192 ( .A(n3441), .B(n3442), .Z(n30531) );
  NANDN U5193 ( .A(n30525), .B(n42047), .Z(n3443) );
  NANDN U5194 ( .A(n30562), .B(n4067), .Z(n3444) );
  NAND U5195 ( .A(n3443), .B(n3444), .Z(n30573) );
  NANDN U5196 ( .A(n30603), .B(n4068), .Z(n3445) );
  NANDN U5197 ( .A(n30563), .B(n42115), .Z(n3446) );
  AND U5198 ( .A(n3445), .B(n3446), .Z(n30605) );
  NANDN U5199 ( .A(n30599), .B(n42047), .Z(n3447) );
  NANDN U5200 ( .A(n30636), .B(n4067), .Z(n3448) );
  NAND U5201 ( .A(n3447), .B(n3448), .Z(n30647) );
  NANDN U5202 ( .A(n30677), .B(n4068), .Z(n3449) );
  NANDN U5203 ( .A(n30640), .B(n42115), .Z(n3450) );
  AND U5204 ( .A(n3449), .B(n3450), .Z(n30679) );
  NANDN U5205 ( .A(n30673), .B(n42047), .Z(n3451) );
  NANDN U5206 ( .A(n30710), .B(n4067), .Z(n3452) );
  NAND U5207 ( .A(n3451), .B(n3452), .Z(n30721) );
  NANDN U5208 ( .A(n30748), .B(n4068), .Z(n3453) );
  NANDN U5209 ( .A(n30711), .B(n42115), .Z(n3454) );
  AND U5210 ( .A(n3453), .B(n3454), .Z(n30753) );
  NANDN U5211 ( .A(n30747), .B(n42047), .Z(n3455) );
  NANDN U5212 ( .A(n30784), .B(n4067), .Z(n3456) );
  NAND U5213 ( .A(n3455), .B(n3456), .Z(n30795) );
  NANDN U5214 ( .A(n30822), .B(n4068), .Z(n3457) );
  NANDN U5215 ( .A(n30788), .B(n42115), .Z(n3458) );
  AND U5216 ( .A(n3457), .B(n3458), .Z(n30827) );
  NANDN U5217 ( .A(n30821), .B(n42047), .Z(n3459) );
  NANDN U5218 ( .A(n30858), .B(n4067), .Z(n3460) );
  NAND U5219 ( .A(n3459), .B(n3460), .Z(n30869) );
  NANDN U5220 ( .A(n30899), .B(n4068), .Z(n3461) );
  NANDN U5221 ( .A(n30862), .B(n42115), .Z(n3462) );
  AND U5222 ( .A(n3461), .B(n3462), .Z(n30901) );
  NANDN U5223 ( .A(n30895), .B(n42047), .Z(n3463) );
  NANDN U5224 ( .A(n30932), .B(n4067), .Z(n3464) );
  NAND U5225 ( .A(n3463), .B(n3464), .Z(n30943) );
  NANDN U5226 ( .A(n30970), .B(n4068), .Z(n3465) );
  NANDN U5227 ( .A(n30936), .B(n42115), .Z(n3466) );
  AND U5228 ( .A(n3465), .B(n3466), .Z(n30975) );
  NANDN U5229 ( .A(n30969), .B(n42047), .Z(n3467) );
  NANDN U5230 ( .A(n31006), .B(n4067), .Z(n3468) );
  NAND U5231 ( .A(n3467), .B(n3468), .Z(n31017) );
  NANDN U5232 ( .A(n31047), .B(n4068), .Z(n3469) );
  NANDN U5233 ( .A(n31010), .B(n42115), .Z(n3470) );
  AND U5234 ( .A(n3469), .B(n3470), .Z(n31049) );
  NANDN U5235 ( .A(n31043), .B(n42047), .Z(n3471) );
  NANDN U5236 ( .A(n31080), .B(n4067), .Z(n3472) );
  NAND U5237 ( .A(n3471), .B(n3472), .Z(n31091) );
  NANDN U5238 ( .A(n31121), .B(n4068), .Z(n3473) );
  NANDN U5239 ( .A(n31084), .B(n42115), .Z(n3474) );
  AND U5240 ( .A(n3473), .B(n3474), .Z(n31123) );
  NANDN U5241 ( .A(n31117), .B(n42047), .Z(n3475) );
  NANDN U5242 ( .A(n31154), .B(n4067), .Z(n3476) );
  NAND U5243 ( .A(n3475), .B(n3476), .Z(n31165) );
  NANDN U5244 ( .A(n31195), .B(n4068), .Z(n3477) );
  NANDN U5245 ( .A(n31155), .B(n42115), .Z(n3478) );
  AND U5246 ( .A(n3477), .B(n3478), .Z(n31197) );
  NANDN U5247 ( .A(n31191), .B(n42047), .Z(n3479) );
  NANDN U5248 ( .A(n31228), .B(n4067), .Z(n3480) );
  NAND U5249 ( .A(n3479), .B(n3480), .Z(n31239) );
  NANDN U5250 ( .A(n31269), .B(n4068), .Z(n3481) );
  NANDN U5251 ( .A(n31232), .B(n42115), .Z(n3482) );
  AND U5252 ( .A(n3481), .B(n3482), .Z(n31271) );
  NANDN U5253 ( .A(n31265), .B(n42047), .Z(n3483) );
  NANDN U5254 ( .A(n31302), .B(n4067), .Z(n3484) );
  NAND U5255 ( .A(n3483), .B(n3484), .Z(n31313) );
  NANDN U5256 ( .A(n31340), .B(n4068), .Z(n3485) );
  NANDN U5257 ( .A(n31306), .B(n42115), .Z(n3486) );
  AND U5258 ( .A(n3485), .B(n3486), .Z(n31345) );
  NANDN U5259 ( .A(n31339), .B(n42047), .Z(n3487) );
  NANDN U5260 ( .A(n31376), .B(n4067), .Z(n3488) );
  NAND U5261 ( .A(n3487), .B(n3488), .Z(n31387) );
  NANDN U5262 ( .A(n31417), .B(n4068), .Z(n3489) );
  NANDN U5263 ( .A(n31380), .B(n42115), .Z(n3490) );
  AND U5264 ( .A(n3489), .B(n3490), .Z(n31419) );
  NANDN U5265 ( .A(n31413), .B(n42047), .Z(n3491) );
  NANDN U5266 ( .A(n31450), .B(n4067), .Z(n3492) );
  NAND U5267 ( .A(n3491), .B(n3492), .Z(n31461) );
  NANDN U5268 ( .A(n31491), .B(n4068), .Z(n3493) );
  NANDN U5269 ( .A(n31454), .B(n42115), .Z(n3494) );
  AND U5270 ( .A(n3493), .B(n3494), .Z(n31493) );
  NANDN U5271 ( .A(n31487), .B(n42047), .Z(n3495) );
  NANDN U5272 ( .A(n31524), .B(n4067), .Z(n3496) );
  NAND U5273 ( .A(n3495), .B(n3496), .Z(n31535) );
  NANDN U5274 ( .A(n31562), .B(n4068), .Z(n3497) );
  NANDN U5275 ( .A(n31525), .B(n42115), .Z(n3498) );
  AND U5276 ( .A(n3497), .B(n3498), .Z(n31567) );
  NANDN U5277 ( .A(n31561), .B(n42047), .Z(n3499) );
  NANDN U5278 ( .A(n31598), .B(n4067), .Z(n3500) );
  NAND U5279 ( .A(n3499), .B(n3500), .Z(n31609) );
  NANDN U5280 ( .A(n31639), .B(n4068), .Z(n3501) );
  NANDN U5281 ( .A(n31602), .B(n42115), .Z(n3502) );
  AND U5282 ( .A(n3501), .B(n3502), .Z(n31641) );
  NANDN U5283 ( .A(n31635), .B(n42047), .Z(n3503) );
  NANDN U5284 ( .A(n31672), .B(n4067), .Z(n3504) );
  NAND U5285 ( .A(n3503), .B(n3504), .Z(n31683) );
  NANDN U5286 ( .A(n31713), .B(n4068), .Z(n3505) );
  NANDN U5287 ( .A(n31673), .B(n42115), .Z(n3506) );
  AND U5288 ( .A(n3505), .B(n3506), .Z(n31715) );
  NANDN U5289 ( .A(n31709), .B(n42047), .Z(n3507) );
  NANDN U5290 ( .A(n31746), .B(n4067), .Z(n3508) );
  NAND U5291 ( .A(n3507), .B(n3508), .Z(n31757) );
  NANDN U5292 ( .A(n31787), .B(n4068), .Z(n3509) );
  NANDN U5293 ( .A(n31747), .B(n42115), .Z(n3510) );
  AND U5294 ( .A(n3509), .B(n3510), .Z(n31789) );
  NANDN U5295 ( .A(n31783), .B(n42047), .Z(n3511) );
  NANDN U5296 ( .A(n31820), .B(n4067), .Z(n3512) );
  NAND U5297 ( .A(n3511), .B(n3512), .Z(n31831) );
  NANDN U5298 ( .A(n31858), .B(n4068), .Z(n3513) );
  NANDN U5299 ( .A(n31824), .B(n42115), .Z(n3514) );
  AND U5300 ( .A(n3513), .B(n3514), .Z(n31863) );
  NANDN U5301 ( .A(n31857), .B(n42047), .Z(n3515) );
  NANDN U5302 ( .A(n31894), .B(n4067), .Z(n3516) );
  NAND U5303 ( .A(n3515), .B(n3516), .Z(n31905) );
  NANDN U5304 ( .A(n31935), .B(n4068), .Z(n3517) );
  NANDN U5305 ( .A(n31898), .B(n42115), .Z(n3518) );
  AND U5306 ( .A(n3517), .B(n3518), .Z(n31937) );
  NANDN U5307 ( .A(n31931), .B(n42047), .Z(n3519) );
  NANDN U5308 ( .A(n31968), .B(n4067), .Z(n3520) );
  NAND U5309 ( .A(n3519), .B(n3520), .Z(n31979) );
  NANDN U5310 ( .A(n32006), .B(n4068), .Z(n3521) );
  NANDN U5311 ( .A(n31972), .B(n42115), .Z(n3522) );
  AND U5312 ( .A(n3521), .B(n3522), .Z(n32011) );
  NANDN U5313 ( .A(n32005), .B(n42047), .Z(n3523) );
  NANDN U5314 ( .A(n32042), .B(n4067), .Z(n3524) );
  NAND U5315 ( .A(n3523), .B(n3524), .Z(n32053) );
  NANDN U5316 ( .A(n32083), .B(n4068), .Z(n3525) );
  NANDN U5317 ( .A(n32046), .B(n42115), .Z(n3526) );
  AND U5318 ( .A(n3525), .B(n3526), .Z(n32085) );
  NANDN U5319 ( .A(n32079), .B(n42047), .Z(n3527) );
  NANDN U5320 ( .A(n32116), .B(n4067), .Z(n3528) );
  NAND U5321 ( .A(n3527), .B(n3528), .Z(n32127) );
  NANDN U5322 ( .A(n32157), .B(n4068), .Z(n3529) );
  NANDN U5323 ( .A(n32120), .B(n42115), .Z(n3530) );
  AND U5324 ( .A(n3529), .B(n3530), .Z(n32159) );
  NANDN U5325 ( .A(n32153), .B(n42047), .Z(n3531) );
  NANDN U5326 ( .A(n32190), .B(n4067), .Z(n3532) );
  NAND U5327 ( .A(n3531), .B(n3532), .Z(n32201) );
  NANDN U5328 ( .A(n32231), .B(n4068), .Z(n3533) );
  NANDN U5329 ( .A(n32194), .B(n42115), .Z(n3534) );
  AND U5330 ( .A(n3533), .B(n3534), .Z(n32233) );
  NANDN U5331 ( .A(n32227), .B(n42047), .Z(n3535) );
  NANDN U5332 ( .A(n32264), .B(n4067), .Z(n3536) );
  NAND U5333 ( .A(n3535), .B(n3536), .Z(n32275) );
  NANDN U5334 ( .A(n32302), .B(n4068), .Z(n3537) );
  NANDN U5335 ( .A(n32268), .B(n42115), .Z(n3538) );
  AND U5336 ( .A(n3537), .B(n3538), .Z(n32307) );
  NANDN U5337 ( .A(n32301), .B(n42047), .Z(n3539) );
  NANDN U5338 ( .A(n32338), .B(n4067), .Z(n3540) );
  NAND U5339 ( .A(n3539), .B(n3540), .Z(n32349) );
  NANDN U5340 ( .A(n32376), .B(n4068), .Z(n3541) );
  NANDN U5341 ( .A(n32339), .B(n42115), .Z(n3542) );
  AND U5342 ( .A(n3541), .B(n3542), .Z(n32381) );
  NANDN U5343 ( .A(n32375), .B(n42047), .Z(n3543) );
  NANDN U5344 ( .A(n32412), .B(n4067), .Z(n3544) );
  NAND U5345 ( .A(n3543), .B(n3544), .Z(n32423) );
  NANDN U5346 ( .A(n32453), .B(n4068), .Z(n3545) );
  NANDN U5347 ( .A(n32416), .B(n42115), .Z(n3546) );
  AND U5348 ( .A(n3545), .B(n3546), .Z(n32455) );
  NANDN U5349 ( .A(n32449), .B(n42047), .Z(n3547) );
  NANDN U5350 ( .A(n32486), .B(n4067), .Z(n3548) );
  NAND U5351 ( .A(n3547), .B(n3548), .Z(n32497) );
  NANDN U5352 ( .A(n32527), .B(n4068), .Z(n3549) );
  NANDN U5353 ( .A(n32490), .B(n42115), .Z(n3550) );
  AND U5354 ( .A(n3549), .B(n3550), .Z(n32529) );
  NANDN U5355 ( .A(n32523), .B(n42047), .Z(n3551) );
  NANDN U5356 ( .A(n32560), .B(n4067), .Z(n3552) );
  NAND U5357 ( .A(n3551), .B(n3552), .Z(n32571) );
  NANDN U5358 ( .A(n32598), .B(n4068), .Z(n3553) );
  NANDN U5359 ( .A(n32564), .B(n42115), .Z(n3554) );
  AND U5360 ( .A(n3553), .B(n3554), .Z(n32603) );
  NANDN U5361 ( .A(n32597), .B(n42047), .Z(n3555) );
  NANDN U5362 ( .A(n32634), .B(n4067), .Z(n3556) );
  NAND U5363 ( .A(n3555), .B(n3556), .Z(n32645) );
  NANDN U5364 ( .A(n32672), .B(n4068), .Z(n3557) );
  NANDN U5365 ( .A(n32635), .B(n42115), .Z(n3558) );
  AND U5366 ( .A(n3557), .B(n3558), .Z(n32677) );
  NANDN U5367 ( .A(n32671), .B(n42047), .Z(n3559) );
  NANDN U5368 ( .A(n32708), .B(n4067), .Z(n3560) );
  NAND U5369 ( .A(n3559), .B(n3560), .Z(n32719) );
  NANDN U5370 ( .A(n32746), .B(n4068), .Z(n3561) );
  NANDN U5371 ( .A(n32709), .B(n42115), .Z(n3562) );
  AND U5372 ( .A(n3561), .B(n3562), .Z(n32751) );
  NANDN U5373 ( .A(n32745), .B(n42047), .Z(n3563) );
  NANDN U5374 ( .A(n32782), .B(n4067), .Z(n3564) );
  NAND U5375 ( .A(n3563), .B(n3564), .Z(n32793) );
  NANDN U5376 ( .A(n32820), .B(n4068), .Z(n3565) );
  NANDN U5377 ( .A(n32783), .B(n42115), .Z(n3566) );
  AND U5378 ( .A(n3565), .B(n3566), .Z(n32825) );
  NANDN U5379 ( .A(n32819), .B(n42047), .Z(n3567) );
  NANDN U5380 ( .A(n32856), .B(n4067), .Z(n3568) );
  NAND U5381 ( .A(n3567), .B(n3568), .Z(n32867) );
  NANDN U5382 ( .A(n32897), .B(n4068), .Z(n3569) );
  NANDN U5383 ( .A(n32857), .B(n42115), .Z(n3570) );
  AND U5384 ( .A(n3569), .B(n3570), .Z(n32899) );
  NANDN U5385 ( .A(n32893), .B(n42047), .Z(n3571) );
  NANDN U5386 ( .A(n32930), .B(n4067), .Z(n3572) );
  NAND U5387 ( .A(n3571), .B(n3572), .Z(n32941) );
  NANDN U5388 ( .A(n32971), .B(n4068), .Z(n3573) );
  NANDN U5389 ( .A(n32934), .B(n42115), .Z(n3574) );
  AND U5390 ( .A(n3573), .B(n3574), .Z(n32973) );
  NANDN U5391 ( .A(n32967), .B(n42047), .Z(n3575) );
  NANDN U5392 ( .A(n33004), .B(n4067), .Z(n3576) );
  NAND U5393 ( .A(n3575), .B(n3576), .Z(n33015) );
  NANDN U5394 ( .A(n33045), .B(n4068), .Z(n3577) );
  NANDN U5395 ( .A(n33008), .B(n42115), .Z(n3578) );
  AND U5396 ( .A(n3577), .B(n3578), .Z(n33047) );
  NANDN U5397 ( .A(n33041), .B(n42047), .Z(n3579) );
  NANDN U5398 ( .A(n33078), .B(n4067), .Z(n3580) );
  NAND U5399 ( .A(n3579), .B(n3580), .Z(n33089) );
  NANDN U5400 ( .A(n33116), .B(n4068), .Z(n3581) );
  NANDN U5401 ( .A(n33082), .B(n42115), .Z(n3582) );
  AND U5402 ( .A(n3581), .B(n3582), .Z(n33121) );
  NANDN U5403 ( .A(n33115), .B(n42047), .Z(n3583) );
  NANDN U5404 ( .A(n33152), .B(n4067), .Z(n3584) );
  NAND U5405 ( .A(n3583), .B(n3584), .Z(n33163) );
  NANDN U5406 ( .A(n33190), .B(n4068), .Z(n3585) );
  NANDN U5407 ( .A(n33156), .B(n42115), .Z(n3586) );
  AND U5408 ( .A(n3585), .B(n3586), .Z(n33195) );
  NANDN U5409 ( .A(n33189), .B(n42047), .Z(n3587) );
  NANDN U5410 ( .A(n33226), .B(n4067), .Z(n3588) );
  NAND U5411 ( .A(n3587), .B(n3588), .Z(n33237) );
  NANDN U5412 ( .A(n33267), .B(n4068), .Z(n3589) );
  NANDN U5413 ( .A(n33227), .B(n42115), .Z(n3590) );
  AND U5414 ( .A(n3589), .B(n3590), .Z(n33269) );
  NANDN U5415 ( .A(n33263), .B(n42047), .Z(n3591) );
  NANDN U5416 ( .A(n33300), .B(n4067), .Z(n3592) );
  NAND U5417 ( .A(n3591), .B(n3592), .Z(n33311) );
  NANDN U5418 ( .A(n33341), .B(n4068), .Z(n3593) );
  NANDN U5419 ( .A(n33301), .B(n42115), .Z(n3594) );
  AND U5420 ( .A(n3593), .B(n3594), .Z(n33343) );
  NANDN U5421 ( .A(n33337), .B(n42047), .Z(n3595) );
  NANDN U5422 ( .A(n33374), .B(n4067), .Z(n3596) );
  NAND U5423 ( .A(n3595), .B(n3596), .Z(n33385) );
  NANDN U5424 ( .A(n33415), .B(n4068), .Z(n3597) );
  NANDN U5425 ( .A(n33378), .B(n42115), .Z(n3598) );
  AND U5426 ( .A(n3597), .B(n3598), .Z(n33417) );
  NANDN U5427 ( .A(n33411), .B(n42047), .Z(n3599) );
  NANDN U5428 ( .A(n33448), .B(n4067), .Z(n3600) );
  NAND U5429 ( .A(n3599), .B(n3600), .Z(n33459) );
  NANDN U5430 ( .A(n33489), .B(n4068), .Z(n3601) );
  NANDN U5431 ( .A(n33449), .B(n42115), .Z(n3602) );
  AND U5432 ( .A(n3601), .B(n3602), .Z(n33491) );
  NANDN U5433 ( .A(n33485), .B(n42047), .Z(n3603) );
  NANDN U5434 ( .A(n33522), .B(n4067), .Z(n3604) );
  NAND U5435 ( .A(n3603), .B(n3604), .Z(n33533) );
  NANDN U5436 ( .A(n33563), .B(n4068), .Z(n3605) );
  NANDN U5437 ( .A(n33523), .B(n42115), .Z(n3606) );
  AND U5438 ( .A(n3605), .B(n3606), .Z(n33565) );
  NANDN U5439 ( .A(n33559), .B(n42047), .Z(n3607) );
  NANDN U5440 ( .A(n33596), .B(n4067), .Z(n3608) );
  NAND U5441 ( .A(n3607), .B(n3608), .Z(n33607) );
  NANDN U5442 ( .A(n33634), .B(n4068), .Z(n3609) );
  NANDN U5443 ( .A(n33600), .B(n42115), .Z(n3610) );
  AND U5444 ( .A(n3609), .B(n3610), .Z(n33639) );
  NANDN U5445 ( .A(n33633), .B(n42047), .Z(n3611) );
  NANDN U5446 ( .A(n33670), .B(n4067), .Z(n3612) );
  NAND U5447 ( .A(n3611), .B(n3612), .Z(n33681) );
  NANDN U5448 ( .A(n33711), .B(n4068), .Z(n3613) );
  NANDN U5449 ( .A(n33674), .B(n42115), .Z(n3614) );
  AND U5450 ( .A(n3613), .B(n3614), .Z(n33713) );
  NANDN U5451 ( .A(n33707), .B(n42047), .Z(n3615) );
  NANDN U5452 ( .A(n33744), .B(n4067), .Z(n3616) );
  NAND U5453 ( .A(n3615), .B(n3616), .Z(n33755) );
  NANDN U5454 ( .A(n33782), .B(n4068), .Z(n3617) );
  NANDN U5455 ( .A(n33748), .B(n42115), .Z(n3618) );
  AND U5456 ( .A(n3617), .B(n3618), .Z(n33787) );
  NANDN U5457 ( .A(n33781), .B(n42047), .Z(n3619) );
  NANDN U5458 ( .A(n33818), .B(n4067), .Z(n3620) );
  NAND U5459 ( .A(n3619), .B(n3620), .Z(n33829) );
  NANDN U5460 ( .A(n33859), .B(n4068), .Z(n3621) );
  NANDN U5461 ( .A(n33822), .B(n42115), .Z(n3622) );
  AND U5462 ( .A(n3621), .B(n3622), .Z(n33861) );
  NANDN U5463 ( .A(n33855), .B(n42047), .Z(n3623) );
  NANDN U5464 ( .A(n33892), .B(n4067), .Z(n3624) );
  NAND U5465 ( .A(n3623), .B(n3624), .Z(n33903) );
  NANDN U5466 ( .A(n33933), .B(n4068), .Z(n3625) );
  NANDN U5467 ( .A(n33893), .B(n42115), .Z(n3626) );
  AND U5468 ( .A(n3625), .B(n3626), .Z(n33935) );
  NANDN U5469 ( .A(n33929), .B(n42047), .Z(n3627) );
  NANDN U5470 ( .A(n33966), .B(n4067), .Z(n3628) );
  NAND U5471 ( .A(n3627), .B(n3628), .Z(n33977) );
  NANDN U5472 ( .A(n34007), .B(n4068), .Z(n3629) );
  NANDN U5473 ( .A(n33967), .B(n42115), .Z(n3630) );
  AND U5474 ( .A(n3629), .B(n3630), .Z(n34009) );
  NANDN U5475 ( .A(n34003), .B(n42047), .Z(n3631) );
  NANDN U5476 ( .A(n34040), .B(n4067), .Z(n3632) );
  NAND U5477 ( .A(n3631), .B(n3632), .Z(n34051) );
  NANDN U5478 ( .A(n34078), .B(n4068), .Z(n3633) );
  NANDN U5479 ( .A(n34044), .B(n42115), .Z(n3634) );
  AND U5480 ( .A(n3633), .B(n3634), .Z(n34083) );
  NANDN U5481 ( .A(n34077), .B(n42047), .Z(n3635) );
  NANDN U5482 ( .A(n34114), .B(n4067), .Z(n3636) );
  NAND U5483 ( .A(n3635), .B(n3636), .Z(n34125) );
  NANDN U5484 ( .A(n34155), .B(n4068), .Z(n3637) );
  NANDN U5485 ( .A(n34115), .B(n42115), .Z(n3638) );
  AND U5486 ( .A(n3637), .B(n3638), .Z(n34157) );
  NANDN U5487 ( .A(n34151), .B(n42047), .Z(n3639) );
  NANDN U5488 ( .A(n34188), .B(n4067), .Z(n3640) );
  NAND U5489 ( .A(n3639), .B(n3640), .Z(n34199) );
  NANDN U5490 ( .A(n34229), .B(n4068), .Z(n3641) );
  NANDN U5491 ( .A(n34189), .B(n42115), .Z(n3642) );
  AND U5492 ( .A(n3641), .B(n3642), .Z(n34231) );
  NANDN U5493 ( .A(n34225), .B(n42047), .Z(n3643) );
  NANDN U5494 ( .A(n34262), .B(n4067), .Z(n3644) );
  NAND U5495 ( .A(n3643), .B(n3644), .Z(n34273) );
  NANDN U5496 ( .A(n34300), .B(n4068), .Z(n3645) );
  NANDN U5497 ( .A(n34266), .B(n42115), .Z(n3646) );
  AND U5498 ( .A(n3645), .B(n3646), .Z(n34305) );
  NANDN U5499 ( .A(n34299), .B(n42047), .Z(n3647) );
  NANDN U5500 ( .A(n34336), .B(n4067), .Z(n3648) );
  NAND U5501 ( .A(n3647), .B(n3648), .Z(n34347) );
  NANDN U5502 ( .A(n34374), .B(n4068), .Z(n3649) );
  NANDN U5503 ( .A(n34340), .B(n42115), .Z(n3650) );
  AND U5504 ( .A(n3649), .B(n3650), .Z(n34379) );
  NANDN U5505 ( .A(n34373), .B(n42047), .Z(n3651) );
  NANDN U5506 ( .A(n34410), .B(n4067), .Z(n3652) );
  NAND U5507 ( .A(n3651), .B(n3652), .Z(n34421) );
  NANDN U5508 ( .A(n34448), .B(n4068), .Z(n3653) );
  NANDN U5509 ( .A(n34411), .B(n42115), .Z(n3654) );
  AND U5510 ( .A(n3653), .B(n3654), .Z(n34453) );
  NANDN U5511 ( .A(n34447), .B(n42047), .Z(n3655) );
  NANDN U5512 ( .A(n34484), .B(n4067), .Z(n3656) );
  NAND U5513 ( .A(n3655), .B(n3656), .Z(n34495) );
  NANDN U5514 ( .A(n34525), .B(n4068), .Z(n3657) );
  NANDN U5515 ( .A(n34485), .B(n42115), .Z(n3658) );
  AND U5516 ( .A(n3657), .B(n3658), .Z(n34527) );
  NANDN U5517 ( .A(n34521), .B(n42047), .Z(n3659) );
  NANDN U5518 ( .A(n34558), .B(n4067), .Z(n3660) );
  NAND U5519 ( .A(n3659), .B(n3660), .Z(n34569) );
  NANDN U5520 ( .A(n34596), .B(n4068), .Z(n3661) );
  NANDN U5521 ( .A(n34562), .B(n42115), .Z(n3662) );
  AND U5522 ( .A(n3661), .B(n3662), .Z(n34601) );
  NANDN U5523 ( .A(n34595), .B(n42047), .Z(n3663) );
  NANDN U5524 ( .A(n34632), .B(n4067), .Z(n3664) );
  NAND U5525 ( .A(n3663), .B(n3664), .Z(n34643) );
  NANDN U5526 ( .A(n34670), .B(n4068), .Z(n3665) );
  NANDN U5527 ( .A(n34636), .B(n42115), .Z(n3666) );
  AND U5528 ( .A(n3665), .B(n3666), .Z(n34675) );
  NANDN U5529 ( .A(n34669), .B(n42047), .Z(n3667) );
  NANDN U5530 ( .A(n34706), .B(n4067), .Z(n3668) );
  NAND U5531 ( .A(n3667), .B(n3668), .Z(n34717) );
  NANDN U5532 ( .A(n34744), .B(n4068), .Z(n3669) );
  NANDN U5533 ( .A(n34707), .B(n42115), .Z(n3670) );
  AND U5534 ( .A(n3669), .B(n3670), .Z(n34749) );
  NANDN U5535 ( .A(n34743), .B(n42047), .Z(n3671) );
  NANDN U5536 ( .A(n34780), .B(n4067), .Z(n3672) );
  NAND U5537 ( .A(n3671), .B(n3672), .Z(n34791) );
  NANDN U5538 ( .A(n34818), .B(n4068), .Z(n3673) );
  NANDN U5539 ( .A(n34781), .B(n42115), .Z(n3674) );
  AND U5540 ( .A(n3673), .B(n3674), .Z(n34823) );
  NANDN U5541 ( .A(n34817), .B(n42047), .Z(n3675) );
  NANDN U5542 ( .A(n34854), .B(n4067), .Z(n3676) );
  NAND U5543 ( .A(n3675), .B(n3676), .Z(n34865) );
  NANDN U5544 ( .A(n34892), .B(n4068), .Z(n3677) );
  NANDN U5545 ( .A(n34855), .B(n42115), .Z(n3678) );
  AND U5546 ( .A(n3677), .B(n3678), .Z(n34897) );
  NANDN U5547 ( .A(n34891), .B(n42047), .Z(n3679) );
  NANDN U5548 ( .A(n34928), .B(n4067), .Z(n3680) );
  NAND U5549 ( .A(n3679), .B(n3680), .Z(n34939) );
  NANDN U5550 ( .A(n34969), .B(n4068), .Z(n3681) );
  NANDN U5551 ( .A(n34929), .B(n42115), .Z(n3682) );
  AND U5552 ( .A(n3681), .B(n3682), .Z(n34971) );
  NANDN U5553 ( .A(n34965), .B(n42047), .Z(n3683) );
  NANDN U5554 ( .A(n35002), .B(n4067), .Z(n3684) );
  NAND U5555 ( .A(n3683), .B(n3684), .Z(n35013) );
  NANDN U5556 ( .A(n35043), .B(n4068), .Z(n3685) );
  NANDN U5557 ( .A(n35006), .B(n42115), .Z(n3686) );
  AND U5558 ( .A(n3685), .B(n3686), .Z(n35045) );
  NANDN U5559 ( .A(n35039), .B(n42047), .Z(n3687) );
  NANDN U5560 ( .A(n35076), .B(n4067), .Z(n3688) );
  NAND U5561 ( .A(n3687), .B(n3688), .Z(n35087) );
  NANDN U5562 ( .A(n35114), .B(n4068), .Z(n3689) );
  NANDN U5563 ( .A(n35077), .B(n42115), .Z(n3690) );
  AND U5564 ( .A(n3689), .B(n3690), .Z(n35119) );
  NANDN U5565 ( .A(n35113), .B(n42047), .Z(n3691) );
  NANDN U5566 ( .A(n35150), .B(n4067), .Z(n3692) );
  NAND U5567 ( .A(n3691), .B(n3692), .Z(n35161) );
  NANDN U5568 ( .A(n35191), .B(n4068), .Z(n3693) );
  NANDN U5569 ( .A(n35154), .B(n42115), .Z(n3694) );
  AND U5570 ( .A(n3693), .B(n3694), .Z(n35193) );
  NANDN U5571 ( .A(n35187), .B(n42047), .Z(n3695) );
  NANDN U5572 ( .A(n35224), .B(n4067), .Z(n3696) );
  NAND U5573 ( .A(n3695), .B(n3696), .Z(n35235) );
  NANDN U5574 ( .A(n35265), .B(n4068), .Z(n3697) );
  NANDN U5575 ( .A(n35228), .B(n42115), .Z(n3698) );
  AND U5576 ( .A(n3697), .B(n3698), .Z(n35267) );
  NANDN U5577 ( .A(n35261), .B(n42047), .Z(n3699) );
  NANDN U5578 ( .A(n35298), .B(n4067), .Z(n3700) );
  NAND U5579 ( .A(n3699), .B(n3700), .Z(n35309) );
  NANDN U5580 ( .A(n35336), .B(n4068), .Z(n3701) );
  NANDN U5581 ( .A(n35299), .B(n42115), .Z(n3702) );
  AND U5582 ( .A(n3701), .B(n3702), .Z(n35341) );
  NANDN U5583 ( .A(n35335), .B(n42047), .Z(n3703) );
  NANDN U5584 ( .A(n35372), .B(n4067), .Z(n3704) );
  NAND U5585 ( .A(n3703), .B(n3704), .Z(n35383) );
  NANDN U5586 ( .A(n35410), .B(n4068), .Z(n3705) );
  NANDN U5587 ( .A(n35373), .B(n42115), .Z(n3706) );
  AND U5588 ( .A(n3705), .B(n3706), .Z(n35415) );
  NANDN U5589 ( .A(n35409), .B(n42047), .Z(n3707) );
  NANDN U5590 ( .A(n35446), .B(n4067), .Z(n3708) );
  NAND U5591 ( .A(n3707), .B(n3708), .Z(n35457) );
  NANDN U5592 ( .A(n35484), .B(n4068), .Z(n3709) );
  NANDN U5593 ( .A(n35447), .B(n42115), .Z(n3710) );
  AND U5594 ( .A(n3709), .B(n3710), .Z(n35489) );
  NANDN U5595 ( .A(n35483), .B(n42047), .Z(n3711) );
  NANDN U5596 ( .A(n35520), .B(n4067), .Z(n3712) );
  NAND U5597 ( .A(n3711), .B(n3712), .Z(n35531) );
  NANDN U5598 ( .A(n35558), .B(n4068), .Z(n3713) );
  NANDN U5599 ( .A(n35521), .B(n42115), .Z(n3714) );
  AND U5600 ( .A(n3713), .B(n3714), .Z(n35563) );
  NANDN U5601 ( .A(n35557), .B(n42047), .Z(n3715) );
  NANDN U5602 ( .A(n35594), .B(n4067), .Z(n3716) );
  NAND U5603 ( .A(n3715), .B(n3716), .Z(n35605) );
  NANDN U5604 ( .A(n35635), .B(n4068), .Z(n3717) );
  NANDN U5605 ( .A(n35598), .B(n42115), .Z(n3718) );
  AND U5606 ( .A(n3717), .B(n3718), .Z(n35637) );
  NANDN U5607 ( .A(n35631), .B(n42047), .Z(n3719) );
  NANDN U5608 ( .A(n35668), .B(n4067), .Z(n3720) );
  NAND U5609 ( .A(n3719), .B(n3720), .Z(n35679) );
  NANDN U5610 ( .A(n35706), .B(n4068), .Z(n3721) );
  NANDN U5611 ( .A(n35669), .B(n42115), .Z(n3722) );
  AND U5612 ( .A(n3721), .B(n3722), .Z(n35711) );
  NANDN U5613 ( .A(n35705), .B(n42047), .Z(n3723) );
  NANDN U5614 ( .A(n35742), .B(n4067), .Z(n3724) );
  NAND U5615 ( .A(n3723), .B(n3724), .Z(n35753) );
  NANDN U5616 ( .A(n35780), .B(n4068), .Z(n3725) );
  NANDN U5617 ( .A(n35743), .B(n42115), .Z(n3726) );
  AND U5618 ( .A(n3725), .B(n3726), .Z(n35785) );
  NANDN U5619 ( .A(n35779), .B(n42047), .Z(n3727) );
  NANDN U5620 ( .A(n35816), .B(n4067), .Z(n3728) );
  NAND U5621 ( .A(n3727), .B(n3728), .Z(n35827) );
  NANDN U5622 ( .A(n35857), .B(n4068), .Z(n3729) );
  NANDN U5623 ( .A(n35820), .B(n42115), .Z(n3730) );
  AND U5624 ( .A(n3729), .B(n3730), .Z(n35859) );
  NANDN U5625 ( .A(n35853), .B(n42047), .Z(n3731) );
  NANDN U5626 ( .A(n35890), .B(n4067), .Z(n3732) );
  NAND U5627 ( .A(n3731), .B(n3732), .Z(n35901) );
  NANDN U5628 ( .A(n35928), .B(n4068), .Z(n3733) );
  NANDN U5629 ( .A(n35894), .B(n42115), .Z(n3734) );
  AND U5630 ( .A(n3733), .B(n3734), .Z(n35933) );
  NANDN U5631 ( .A(n35927), .B(n42047), .Z(n3735) );
  NANDN U5632 ( .A(n35964), .B(n4067), .Z(n3736) );
  NAND U5633 ( .A(n3735), .B(n3736), .Z(n35975) );
  NANDN U5634 ( .A(n36002), .B(n4068), .Z(n3737) );
  NANDN U5635 ( .A(n35968), .B(n42115), .Z(n3738) );
  AND U5636 ( .A(n3737), .B(n3738), .Z(n36007) );
  NANDN U5637 ( .A(n36001), .B(n42047), .Z(n3739) );
  NANDN U5638 ( .A(n36038), .B(n4067), .Z(n3740) );
  NAND U5639 ( .A(n3739), .B(n3740), .Z(n36049) );
  NANDN U5640 ( .A(n36079), .B(n4068), .Z(n3741) );
  NANDN U5641 ( .A(n36042), .B(n42115), .Z(n3742) );
  AND U5642 ( .A(n3741), .B(n3742), .Z(n36081) );
  NANDN U5643 ( .A(n36075), .B(n42047), .Z(n3743) );
  NANDN U5644 ( .A(n36112), .B(n4067), .Z(n3744) );
  NAND U5645 ( .A(n3743), .B(n3744), .Z(n36123) );
  NANDN U5646 ( .A(n36153), .B(n4068), .Z(n3745) );
  NANDN U5647 ( .A(n36113), .B(n42115), .Z(n3746) );
  AND U5648 ( .A(n3745), .B(n3746), .Z(n36155) );
  NANDN U5649 ( .A(n36149), .B(n42047), .Z(n3747) );
  NANDN U5650 ( .A(n36186), .B(n4067), .Z(n3748) );
  NAND U5651 ( .A(n3747), .B(n3748), .Z(n36197) );
  NANDN U5652 ( .A(n36224), .B(n4068), .Z(n3749) );
  NANDN U5653 ( .A(n36190), .B(n42115), .Z(n3750) );
  AND U5654 ( .A(n3749), .B(n3750), .Z(n36229) );
  NANDN U5655 ( .A(n36223), .B(n42047), .Z(n3751) );
  NANDN U5656 ( .A(n36260), .B(n4067), .Z(n3752) );
  NAND U5657 ( .A(n3751), .B(n3752), .Z(n36271) );
  NANDN U5658 ( .A(n36306), .B(n4068), .Z(n3753) );
  NANDN U5659 ( .A(n36261), .B(n42115), .Z(n3754) );
  AND U5660 ( .A(n3753), .B(n3754), .Z(n36308) );
  NANDN U5661 ( .A(n36302), .B(n42047), .Z(n3755) );
  NANDN U5662 ( .A(n36334), .B(n4067), .Z(n3756) );
  NAND U5663 ( .A(n3755), .B(n3756), .Z(n36345) );
  NANDN U5664 ( .A(n36372), .B(n4068), .Z(n3757) );
  NANDN U5665 ( .A(n36335), .B(n42115), .Z(n3758) );
  AND U5666 ( .A(n3757), .B(n3758), .Z(n36377) );
  NANDN U5667 ( .A(n36371), .B(n42047), .Z(n3759) );
  NANDN U5668 ( .A(n36408), .B(n4067), .Z(n3760) );
  NAND U5669 ( .A(n3759), .B(n3760), .Z(n36419) );
  NANDN U5670 ( .A(n36449), .B(n4068), .Z(n3761) );
  NANDN U5671 ( .A(n36412), .B(n42115), .Z(n3762) );
  AND U5672 ( .A(n3761), .B(n3762), .Z(n36451) );
  NANDN U5673 ( .A(n36445), .B(n42047), .Z(n3763) );
  NANDN U5674 ( .A(n36482), .B(n4067), .Z(n3764) );
  NAND U5675 ( .A(n3763), .B(n3764), .Z(n36493) );
  NANDN U5676 ( .A(n36523), .B(n4068), .Z(n3765) );
  NANDN U5677 ( .A(n36486), .B(n42115), .Z(n3766) );
  AND U5678 ( .A(n3765), .B(n3766), .Z(n36525) );
  NANDN U5679 ( .A(n36519), .B(n42047), .Z(n3767) );
  NANDN U5680 ( .A(n36556), .B(n4067), .Z(n3768) );
  NAND U5681 ( .A(n3767), .B(n3768), .Z(n36567) );
  NANDN U5682 ( .A(n36597), .B(n4068), .Z(n3769) );
  NANDN U5683 ( .A(n36560), .B(n42115), .Z(n3770) );
  AND U5684 ( .A(n3769), .B(n3770), .Z(n36599) );
  NANDN U5685 ( .A(n36593), .B(n42047), .Z(n3771) );
  NANDN U5686 ( .A(n36630), .B(n4067), .Z(n3772) );
  NAND U5687 ( .A(n3771), .B(n3772), .Z(n36641) );
  NANDN U5688 ( .A(n36671), .B(n4068), .Z(n3773) );
  NANDN U5689 ( .A(n36631), .B(n42115), .Z(n3774) );
  AND U5690 ( .A(n3773), .B(n3774), .Z(n36673) );
  NANDN U5691 ( .A(n36667), .B(n42047), .Z(n3775) );
  NANDN U5692 ( .A(n36704), .B(n4067), .Z(n3776) );
  NAND U5693 ( .A(n3775), .B(n3776), .Z(n36715) );
  NANDN U5694 ( .A(n36742), .B(n4068), .Z(n3777) );
  NANDN U5695 ( .A(n36708), .B(n42115), .Z(n3778) );
  AND U5696 ( .A(n3777), .B(n3778), .Z(n36747) );
  NANDN U5697 ( .A(n36741), .B(n42047), .Z(n3779) );
  NANDN U5698 ( .A(n36778), .B(n4067), .Z(n3780) );
  NAND U5699 ( .A(n3779), .B(n3780), .Z(n36789) );
  NANDN U5700 ( .A(n36816), .B(n4068), .Z(n3781) );
  NANDN U5701 ( .A(n36782), .B(n42115), .Z(n3782) );
  AND U5702 ( .A(n3781), .B(n3782), .Z(n36821) );
  NANDN U5703 ( .A(n36815), .B(n42047), .Z(n3783) );
  NANDN U5704 ( .A(n36852), .B(n4067), .Z(n3784) );
  NAND U5705 ( .A(n3783), .B(n3784), .Z(n36863) );
  NANDN U5706 ( .A(n36893), .B(n4068), .Z(n3785) );
  NANDN U5707 ( .A(n36856), .B(n42115), .Z(n3786) );
  AND U5708 ( .A(n3785), .B(n3786), .Z(n36895) );
  NANDN U5709 ( .A(n36889), .B(n42047), .Z(n3787) );
  NANDN U5710 ( .A(n36926), .B(n4067), .Z(n3788) );
  NAND U5711 ( .A(n3787), .B(n3788), .Z(n36937) );
  NANDN U5712 ( .A(n36967), .B(n4068), .Z(n3789) );
  NANDN U5713 ( .A(n36927), .B(n42115), .Z(n3790) );
  AND U5714 ( .A(n3789), .B(n3790), .Z(n36969) );
  NANDN U5715 ( .A(n36963), .B(n42047), .Z(n3791) );
  NANDN U5716 ( .A(n37000), .B(n4067), .Z(n3792) );
  NAND U5717 ( .A(n3791), .B(n3792), .Z(n37011) );
  NANDN U5718 ( .A(n37041), .B(n4068), .Z(n3793) );
  NANDN U5719 ( .A(n37001), .B(n42115), .Z(n3794) );
  AND U5720 ( .A(n3793), .B(n3794), .Z(n37043) );
  NANDN U5721 ( .A(n37037), .B(n42047), .Z(n3795) );
  NANDN U5722 ( .A(n37074), .B(n4067), .Z(n3796) );
  NAND U5723 ( .A(n3795), .B(n3796), .Z(n37085) );
  NANDN U5724 ( .A(n37112), .B(n4068), .Z(n3797) );
  NANDN U5725 ( .A(n37078), .B(n42115), .Z(n3798) );
  AND U5726 ( .A(n3797), .B(n3798), .Z(n37117) );
  NANDN U5727 ( .A(n37111), .B(n42047), .Z(n3799) );
  NANDN U5728 ( .A(n37148), .B(n4067), .Z(n3800) );
  NAND U5729 ( .A(n3799), .B(n3800), .Z(n37159) );
  NANDN U5730 ( .A(n37189), .B(n4068), .Z(n3801) );
  NANDN U5731 ( .A(n37152), .B(n42115), .Z(n3802) );
  AND U5732 ( .A(n3801), .B(n3802), .Z(n37191) );
  NANDN U5733 ( .A(n37185), .B(n42047), .Z(n3803) );
  NANDN U5734 ( .A(n37222), .B(n4067), .Z(n3804) );
  NAND U5735 ( .A(n3803), .B(n3804), .Z(n37233) );
  NANDN U5736 ( .A(n37263), .B(n4068), .Z(n3805) );
  NANDN U5737 ( .A(n37226), .B(n42115), .Z(n3806) );
  AND U5738 ( .A(n3805), .B(n3806), .Z(n37265) );
  NANDN U5739 ( .A(n37259), .B(n42047), .Z(n3807) );
  NANDN U5740 ( .A(n37296), .B(n4067), .Z(n3808) );
  NAND U5741 ( .A(n3807), .B(n3808), .Z(n37307) );
  NANDN U5742 ( .A(n37334), .B(n4068), .Z(n3809) );
  NANDN U5743 ( .A(n37297), .B(n42115), .Z(n3810) );
  AND U5744 ( .A(n3809), .B(n3810), .Z(n37339) );
  NANDN U5745 ( .A(n37333), .B(n42047), .Z(n3811) );
  NANDN U5746 ( .A(n37370), .B(n4067), .Z(n3812) );
  NAND U5747 ( .A(n3811), .B(n3812), .Z(n37381) );
  NANDN U5748 ( .A(n37411), .B(n4068), .Z(n3813) );
  NANDN U5749 ( .A(n37371), .B(n42115), .Z(n3814) );
  AND U5750 ( .A(n3813), .B(n3814), .Z(n37413) );
  NANDN U5751 ( .A(n37407), .B(n42047), .Z(n3815) );
  NANDN U5752 ( .A(n37444), .B(n4067), .Z(n3816) );
  NAND U5753 ( .A(n3815), .B(n3816), .Z(n37455) );
  NANDN U5754 ( .A(n37482), .B(n4068), .Z(n3817) );
  NANDN U5755 ( .A(n37445), .B(n42115), .Z(n3818) );
  AND U5756 ( .A(n3817), .B(n3818), .Z(n37487) );
  NANDN U5757 ( .A(n37481), .B(n42047), .Z(n3819) );
  NANDN U5758 ( .A(n37518), .B(n4067), .Z(n3820) );
  NAND U5759 ( .A(n3819), .B(n3820), .Z(n37529) );
  NANDN U5760 ( .A(n37559), .B(n4068), .Z(n3821) );
  NANDN U5761 ( .A(n37519), .B(n42115), .Z(n3822) );
  AND U5762 ( .A(n3821), .B(n3822), .Z(n37561) );
  NANDN U5763 ( .A(n37555), .B(n42047), .Z(n3823) );
  NANDN U5764 ( .A(n37592), .B(n4067), .Z(n3824) );
  NAND U5765 ( .A(n3823), .B(n3824), .Z(n37603) );
  NANDN U5766 ( .A(n37630), .B(n4068), .Z(n3825) );
  NANDN U5767 ( .A(n37596), .B(n42115), .Z(n3826) );
  AND U5768 ( .A(n3825), .B(n3826), .Z(n37635) );
  NANDN U5769 ( .A(n37629), .B(n42047), .Z(n3827) );
  NANDN U5770 ( .A(n37666), .B(n4067), .Z(n3828) );
  NAND U5771 ( .A(n3827), .B(n3828), .Z(n37677) );
  NANDN U5772 ( .A(n37707), .B(n4068), .Z(n3829) );
  NANDN U5773 ( .A(n37670), .B(n42115), .Z(n3830) );
  AND U5774 ( .A(n3829), .B(n3830), .Z(n37709) );
  NANDN U5775 ( .A(n37703), .B(n42047), .Z(n3831) );
  NANDN U5776 ( .A(n37740), .B(n4067), .Z(n3832) );
  NAND U5777 ( .A(n3831), .B(n3832), .Z(n37751) );
  NANDN U5778 ( .A(n37778), .B(n4068), .Z(n3833) );
  NANDN U5779 ( .A(n37744), .B(n42115), .Z(n3834) );
  AND U5780 ( .A(n3833), .B(n3834), .Z(n37783) );
  NANDN U5781 ( .A(n37777), .B(n42047), .Z(n3835) );
  NANDN U5782 ( .A(n37814), .B(n4067), .Z(n3836) );
  NAND U5783 ( .A(n3835), .B(n3836), .Z(n37825) );
  NANDN U5784 ( .A(n37855), .B(n4068), .Z(n3837) );
  NANDN U5785 ( .A(n37818), .B(n42115), .Z(n3838) );
  AND U5786 ( .A(n3837), .B(n3838), .Z(n37857) );
  NANDN U5787 ( .A(n37851), .B(n42047), .Z(n3839) );
  NANDN U5788 ( .A(n37888), .B(n4067), .Z(n3840) );
  NAND U5789 ( .A(n3839), .B(n3840), .Z(n37899) );
  NANDN U5790 ( .A(n37929), .B(n4068), .Z(n3841) );
  NANDN U5791 ( .A(n37889), .B(n42115), .Z(n3842) );
  AND U5792 ( .A(n3841), .B(n3842), .Z(n37931) );
  NANDN U5793 ( .A(n37925), .B(n42047), .Z(n3843) );
  NANDN U5794 ( .A(n37962), .B(n4067), .Z(n3844) );
  NAND U5795 ( .A(n3843), .B(n3844), .Z(n37973) );
  NANDN U5796 ( .A(n38003), .B(n4068), .Z(n3845) );
  NANDN U5797 ( .A(n37963), .B(n42115), .Z(n3846) );
  AND U5798 ( .A(n3845), .B(n3846), .Z(n38005) );
  NANDN U5799 ( .A(n37999), .B(n42047), .Z(n3847) );
  NANDN U5800 ( .A(n38036), .B(n4067), .Z(n3848) );
  NAND U5801 ( .A(n3847), .B(n3848), .Z(n38047) );
  NANDN U5802 ( .A(n38077), .B(n4068), .Z(n3849) );
  NANDN U5803 ( .A(n38040), .B(n42115), .Z(n3850) );
  AND U5804 ( .A(n3849), .B(n3850), .Z(n38079) );
  NANDN U5805 ( .A(n38073), .B(n42047), .Z(n3851) );
  NANDN U5806 ( .A(n38110), .B(n4067), .Z(n3852) );
  NAND U5807 ( .A(n3851), .B(n3852), .Z(n38121) );
  NANDN U5808 ( .A(n38151), .B(n4068), .Z(n3853) );
  NANDN U5809 ( .A(n38114), .B(n42115), .Z(n3854) );
  AND U5810 ( .A(n3853), .B(n3854), .Z(n38153) );
  NANDN U5811 ( .A(n38147), .B(n42047), .Z(n3855) );
  NANDN U5812 ( .A(n38184), .B(n4067), .Z(n3856) );
  NAND U5813 ( .A(n3855), .B(n3856), .Z(n38195) );
  NANDN U5814 ( .A(n38225), .B(n4068), .Z(n3857) );
  NANDN U5815 ( .A(n38188), .B(n42115), .Z(n3858) );
  AND U5816 ( .A(n3857), .B(n3858), .Z(n38227) );
  NANDN U5817 ( .A(n38221), .B(n42047), .Z(n3859) );
  NANDN U5818 ( .A(n38258), .B(n4067), .Z(n3860) );
  NAND U5819 ( .A(n3859), .B(n3860), .Z(n38269) );
  NANDN U5820 ( .A(n38296), .B(n4068), .Z(n3861) );
  NANDN U5821 ( .A(n38262), .B(n42115), .Z(n3862) );
  AND U5822 ( .A(n3861), .B(n3862), .Z(n38301) );
  NANDN U5823 ( .A(n38295), .B(n42047), .Z(n3863) );
  NANDN U5824 ( .A(n38332), .B(n4067), .Z(n3864) );
  NAND U5825 ( .A(n3863), .B(n3864), .Z(n38343) );
  NANDN U5826 ( .A(n38373), .B(n4068), .Z(n3865) );
  NANDN U5827 ( .A(n38333), .B(n42115), .Z(n3866) );
  AND U5828 ( .A(n3865), .B(n3866), .Z(n38375) );
  NANDN U5829 ( .A(n38369), .B(n42047), .Z(n3867) );
  NANDN U5830 ( .A(n38406), .B(n4067), .Z(n3868) );
  NAND U5831 ( .A(n3867), .B(n3868), .Z(n38417) );
  NANDN U5832 ( .A(n38447), .B(n4068), .Z(n3869) );
  NANDN U5833 ( .A(n38407), .B(n42115), .Z(n3870) );
  AND U5834 ( .A(n3869), .B(n3870), .Z(n38449) );
  NANDN U5835 ( .A(n38443), .B(n42047), .Z(n3871) );
  NANDN U5836 ( .A(n38480), .B(n4067), .Z(n3872) );
  NAND U5837 ( .A(n3871), .B(n3872), .Z(n38491) );
  NANDN U5838 ( .A(n38518), .B(n4068), .Z(n3873) );
  NANDN U5839 ( .A(n38481), .B(n42115), .Z(n3874) );
  AND U5840 ( .A(n3873), .B(n3874), .Z(n38523) );
  NANDN U5841 ( .A(n38517), .B(n42047), .Z(n3875) );
  NANDN U5842 ( .A(n38554), .B(n4067), .Z(n3876) );
  NAND U5843 ( .A(n3875), .B(n3876), .Z(n38565) );
  NANDN U5844 ( .A(n38595), .B(n4068), .Z(n3877) );
  NANDN U5845 ( .A(n38558), .B(n42115), .Z(n3878) );
  AND U5846 ( .A(n3877), .B(n3878), .Z(n38597) );
  NANDN U5847 ( .A(n38591), .B(n42047), .Z(n3879) );
  NANDN U5848 ( .A(n38628), .B(n4067), .Z(n3880) );
  NAND U5849 ( .A(n3879), .B(n3880), .Z(n38639) );
  NANDN U5850 ( .A(n38669), .B(n4068), .Z(n3881) );
  NANDN U5851 ( .A(n38629), .B(n42115), .Z(n3882) );
  AND U5852 ( .A(n3881), .B(n3882), .Z(n38671) );
  NANDN U5853 ( .A(n38665), .B(n42047), .Z(n3883) );
  NANDN U5854 ( .A(n38702), .B(n4067), .Z(n3884) );
  NAND U5855 ( .A(n3883), .B(n3884), .Z(n38713) );
  NANDN U5856 ( .A(n38743), .B(n4068), .Z(n3885) );
  NANDN U5857 ( .A(n38706), .B(n42115), .Z(n3886) );
  AND U5858 ( .A(n3885), .B(n3886), .Z(n38745) );
  NANDN U5859 ( .A(n38739), .B(n42047), .Z(n3887) );
  NANDN U5860 ( .A(n38776), .B(n4067), .Z(n3888) );
  NAND U5861 ( .A(n3887), .B(n3888), .Z(n38787) );
  NANDN U5862 ( .A(n38817), .B(n4068), .Z(n3889) );
  NANDN U5863 ( .A(n38780), .B(n42115), .Z(n3890) );
  AND U5864 ( .A(n3889), .B(n3890), .Z(n38819) );
  NANDN U5865 ( .A(n38813), .B(n42047), .Z(n3891) );
  NANDN U5866 ( .A(n38850), .B(n4067), .Z(n3892) );
  NAND U5867 ( .A(n3891), .B(n3892), .Z(n38861) );
  NANDN U5868 ( .A(n38891), .B(n4068), .Z(n3893) );
  NANDN U5869 ( .A(n38854), .B(n42115), .Z(n3894) );
  AND U5870 ( .A(n3893), .B(n3894), .Z(n38893) );
  NANDN U5871 ( .A(n38887), .B(n42047), .Z(n3895) );
  NANDN U5872 ( .A(n38924), .B(n4067), .Z(n3896) );
  NAND U5873 ( .A(n3895), .B(n3896), .Z(n38935) );
  NANDN U5874 ( .A(n38962), .B(n4068), .Z(n3897) );
  NANDN U5875 ( .A(n38928), .B(n42115), .Z(n3898) );
  AND U5876 ( .A(n3897), .B(n3898), .Z(n38967) );
  NANDN U5877 ( .A(n38961), .B(n42047), .Z(n3899) );
  NANDN U5878 ( .A(n38998), .B(n4067), .Z(n3900) );
  NAND U5879 ( .A(n3899), .B(n3900), .Z(n39009) );
  NANDN U5880 ( .A(n39039), .B(n4068), .Z(n3901) );
  NANDN U5881 ( .A(n39002), .B(n42115), .Z(n3902) );
  AND U5882 ( .A(n3901), .B(n3902), .Z(n39041) );
  NANDN U5883 ( .A(n39035), .B(n42047), .Z(n3903) );
  NANDN U5884 ( .A(n39072), .B(n4067), .Z(n3904) );
  NAND U5885 ( .A(n3903), .B(n3904), .Z(n39083) );
  NANDN U5886 ( .A(n39110), .B(n4068), .Z(n3905) );
  NANDN U5887 ( .A(n39076), .B(n42115), .Z(n3906) );
  AND U5888 ( .A(n3905), .B(n3906), .Z(n39115) );
  NANDN U5889 ( .A(n39109), .B(n42047), .Z(n3907) );
  NANDN U5890 ( .A(n39146), .B(n4067), .Z(n3908) );
  NAND U5891 ( .A(n3907), .B(n3908), .Z(n39157) );
  NANDN U5892 ( .A(n39184), .B(n4068), .Z(n3909) );
  NANDN U5893 ( .A(n39147), .B(n42115), .Z(n3910) );
  AND U5894 ( .A(n3909), .B(n3910), .Z(n39189) );
  NANDN U5895 ( .A(n39183), .B(n42047), .Z(n3911) );
  NANDN U5896 ( .A(n39220), .B(n4067), .Z(n3912) );
  NAND U5897 ( .A(n3911), .B(n3912), .Z(n39231) );
  NANDN U5898 ( .A(n39258), .B(n4068), .Z(n3913) );
  NANDN U5899 ( .A(n39224), .B(n42115), .Z(n3914) );
  AND U5900 ( .A(n3913), .B(n3914), .Z(n39263) );
  NANDN U5901 ( .A(n39257), .B(n42047), .Z(n3915) );
  NANDN U5902 ( .A(n39294), .B(n4067), .Z(n3916) );
  NAND U5903 ( .A(n3915), .B(n3916), .Z(n39305) );
  NANDN U5904 ( .A(n39332), .B(n4068), .Z(n3917) );
  NANDN U5905 ( .A(n39298), .B(n42115), .Z(n3918) );
  AND U5906 ( .A(n3917), .B(n3918), .Z(n39337) );
  NANDN U5907 ( .A(n39331), .B(n42047), .Z(n3919) );
  NANDN U5908 ( .A(n39368), .B(n4067), .Z(n3920) );
  NAND U5909 ( .A(n3919), .B(n3920), .Z(n39379) );
  NANDN U5910 ( .A(n39409), .B(n4068), .Z(n3921) );
  NANDN U5911 ( .A(n39372), .B(n42115), .Z(n3922) );
  AND U5912 ( .A(n3921), .B(n3922), .Z(n39411) );
  NANDN U5913 ( .A(n39405), .B(n42047), .Z(n3923) );
  NANDN U5914 ( .A(n39442), .B(n4067), .Z(n3924) );
  NAND U5915 ( .A(n3923), .B(n3924), .Z(n39453) );
  NANDN U5916 ( .A(n39483), .B(n4068), .Z(n3925) );
  NANDN U5917 ( .A(n39446), .B(n42115), .Z(n3926) );
  AND U5918 ( .A(n3925), .B(n3926), .Z(n39485) );
  NANDN U5919 ( .A(n39479), .B(n42047), .Z(n3927) );
  NANDN U5920 ( .A(n39516), .B(n4067), .Z(n3928) );
  NAND U5921 ( .A(n3927), .B(n3928), .Z(n39527) );
  NANDN U5922 ( .A(n39557), .B(n4068), .Z(n3929) );
  NANDN U5923 ( .A(n39520), .B(n42115), .Z(n3930) );
  AND U5924 ( .A(n3929), .B(n3930), .Z(n39559) );
  NANDN U5925 ( .A(n39553), .B(n42047), .Z(n3931) );
  NANDN U5926 ( .A(n39590), .B(n4067), .Z(n3932) );
  NAND U5927 ( .A(n3931), .B(n3932), .Z(n39601) );
  NANDN U5928 ( .A(n39631), .B(n4068), .Z(n3933) );
  NANDN U5929 ( .A(n39594), .B(n42115), .Z(n3934) );
  AND U5930 ( .A(n3933), .B(n3934), .Z(n39633) );
  NANDN U5931 ( .A(n39627), .B(n42047), .Z(n3935) );
  NANDN U5932 ( .A(n39664), .B(n4067), .Z(n3936) );
  NAND U5933 ( .A(n3935), .B(n3936), .Z(n39675) );
  NANDN U5934 ( .A(n39705), .B(n4068), .Z(n3937) );
  NANDN U5935 ( .A(n39665), .B(n42115), .Z(n3938) );
  AND U5936 ( .A(n3937), .B(n3938), .Z(n39707) );
  NANDN U5937 ( .A(n39701), .B(n42047), .Z(n3939) );
  NANDN U5938 ( .A(n39738), .B(n4067), .Z(n3940) );
  NAND U5939 ( .A(n3939), .B(n3940), .Z(n39749) );
  NANDN U5940 ( .A(n39779), .B(n4068), .Z(n3941) );
  NANDN U5941 ( .A(n39742), .B(n42115), .Z(n3942) );
  AND U5942 ( .A(n3941), .B(n3942), .Z(n39781) );
  NANDN U5943 ( .A(n39775), .B(n42047), .Z(n3943) );
  NANDN U5944 ( .A(n39812), .B(n4067), .Z(n3944) );
  NAND U5945 ( .A(n3943), .B(n3944), .Z(n39823) );
  NANDN U5946 ( .A(n39853), .B(n4068), .Z(n3945) );
  NANDN U5947 ( .A(n39813), .B(n42115), .Z(n3946) );
  AND U5948 ( .A(n3945), .B(n3946), .Z(n39855) );
  NANDN U5949 ( .A(n39849), .B(n42047), .Z(n3947) );
  NANDN U5950 ( .A(n39886), .B(n4067), .Z(n3948) );
  NAND U5951 ( .A(n3947), .B(n3948), .Z(n39897) );
  NANDN U5952 ( .A(n39924), .B(n4068), .Z(n3949) );
  NANDN U5953 ( .A(n39890), .B(n42115), .Z(n3950) );
  AND U5954 ( .A(n3949), .B(n3950), .Z(n39929) );
  NANDN U5955 ( .A(n39923), .B(n42047), .Z(n3951) );
  NANDN U5956 ( .A(n39960), .B(n4067), .Z(n3952) );
  NAND U5957 ( .A(n3951), .B(n3952), .Z(n39971) );
  NANDN U5958 ( .A(n39998), .B(n4068), .Z(n3953) );
  NANDN U5959 ( .A(n39964), .B(n42115), .Z(n3954) );
  AND U5960 ( .A(n3953), .B(n3954), .Z(n40003) );
  NANDN U5961 ( .A(n39997), .B(n42047), .Z(n3955) );
  NANDN U5962 ( .A(n40034), .B(n4067), .Z(n3956) );
  NAND U5963 ( .A(n3955), .B(n3956), .Z(n40045) );
  NANDN U5964 ( .A(n40072), .B(n4068), .Z(n3957) );
  NANDN U5965 ( .A(n40035), .B(n42115), .Z(n3958) );
  AND U5966 ( .A(n3957), .B(n3958), .Z(n40077) );
  NANDN U5967 ( .A(n40071), .B(n42047), .Z(n3959) );
  NANDN U5968 ( .A(n40108), .B(n4067), .Z(n3960) );
  NAND U5969 ( .A(n3959), .B(n3960), .Z(n40119) );
  NANDN U5970 ( .A(n40149), .B(n4068), .Z(n3961) );
  NANDN U5971 ( .A(n40112), .B(n42115), .Z(n3962) );
  AND U5972 ( .A(n3961), .B(n3962), .Z(n40151) );
  NANDN U5973 ( .A(n40145), .B(n42047), .Z(n3963) );
  NANDN U5974 ( .A(n40182), .B(n4067), .Z(n3964) );
  NAND U5975 ( .A(n3963), .B(n3964), .Z(n40193) );
  NANDN U5976 ( .A(n40223), .B(n4068), .Z(n3965) );
  NANDN U5977 ( .A(n40186), .B(n42115), .Z(n3966) );
  AND U5978 ( .A(n3965), .B(n3966), .Z(n40225) );
  NANDN U5979 ( .A(n40219), .B(n42047), .Z(n3967) );
  NANDN U5980 ( .A(n40256), .B(n4067), .Z(n3968) );
  NAND U5981 ( .A(n3967), .B(n3968), .Z(n40267) );
  NANDN U5982 ( .A(n40294), .B(n4068), .Z(n3969) );
  NANDN U5983 ( .A(n40260), .B(n42115), .Z(n3970) );
  AND U5984 ( .A(n3969), .B(n3970), .Z(n40299) );
  NANDN U5985 ( .A(n40293), .B(n42047), .Z(n3971) );
  NANDN U5986 ( .A(n40330), .B(n4067), .Z(n3972) );
  NAND U5987 ( .A(n3971), .B(n3972), .Z(n40341) );
  NANDN U5988 ( .A(n40368), .B(n4068), .Z(n3973) );
  NANDN U5989 ( .A(n40334), .B(n42115), .Z(n3974) );
  AND U5990 ( .A(n3973), .B(n3974), .Z(n40373) );
  NANDN U5991 ( .A(n40367), .B(n42047), .Z(n3975) );
  NANDN U5992 ( .A(n40404), .B(n4067), .Z(n3976) );
  NAND U5993 ( .A(n3975), .B(n3976), .Z(n40415) );
  NANDN U5994 ( .A(n40445), .B(n4068), .Z(n3977) );
  NANDN U5995 ( .A(n40408), .B(n42115), .Z(n3978) );
  AND U5996 ( .A(n3977), .B(n3978), .Z(n40447) );
  NANDN U5997 ( .A(n40441), .B(n42047), .Z(n3979) );
  NANDN U5998 ( .A(n40478), .B(n4067), .Z(n3980) );
  NAND U5999 ( .A(n3979), .B(n3980), .Z(n40489) );
  NANDN U6000 ( .A(n40519), .B(n4068), .Z(n3981) );
  NANDN U6001 ( .A(n40482), .B(n42115), .Z(n3982) );
  AND U6002 ( .A(n3981), .B(n3982), .Z(n40521) );
  NANDN U6003 ( .A(n40515), .B(n42047), .Z(n3983) );
  NANDN U6004 ( .A(n40552), .B(n4067), .Z(n3984) );
  NAND U6005 ( .A(n3983), .B(n3984), .Z(n40563) );
  NANDN U6006 ( .A(n40593), .B(n4068), .Z(n3985) );
  NANDN U6007 ( .A(n40556), .B(n42115), .Z(n3986) );
  AND U6008 ( .A(n3985), .B(n3986), .Z(n40595) );
  NANDN U6009 ( .A(n40589), .B(n42047), .Z(n3987) );
  NANDN U6010 ( .A(n40626), .B(n4067), .Z(n3988) );
  NAND U6011 ( .A(n3987), .B(n3988), .Z(n40637) );
  NANDN U6012 ( .A(n40664), .B(n4068), .Z(n3989) );
  NANDN U6013 ( .A(n40630), .B(n42115), .Z(n3990) );
  AND U6014 ( .A(n3989), .B(n3990), .Z(n40669) );
  NANDN U6015 ( .A(n40663), .B(n42047), .Z(n3991) );
  NANDN U6016 ( .A(n40700), .B(n4067), .Z(n3992) );
  NAND U6017 ( .A(n3991), .B(n3992), .Z(n40711) );
  NANDN U6018 ( .A(n40738), .B(n4068), .Z(n3993) );
  NANDN U6019 ( .A(n40704), .B(n42115), .Z(n3994) );
  AND U6020 ( .A(n3993), .B(n3994), .Z(n40743) );
  NANDN U6021 ( .A(n40737), .B(n42047), .Z(n3995) );
  NANDN U6022 ( .A(n40774), .B(n4067), .Z(n3996) );
  NAND U6023 ( .A(n3995), .B(n3996), .Z(n40785) );
  NANDN U6024 ( .A(n40815), .B(n4068), .Z(n3997) );
  NANDN U6025 ( .A(n40775), .B(n42115), .Z(n3998) );
  AND U6026 ( .A(n3997), .B(n3998), .Z(n40817) );
  NANDN U6027 ( .A(n40811), .B(n42047), .Z(n3999) );
  NANDN U6028 ( .A(n40848), .B(n4067), .Z(n4000) );
  NAND U6029 ( .A(n3999), .B(n4000), .Z(n40859) );
  NANDN U6030 ( .A(n40886), .B(n4068), .Z(n4001) );
  NANDN U6031 ( .A(n40849), .B(n42115), .Z(n4002) );
  AND U6032 ( .A(n4001), .B(n4002), .Z(n40891) );
  NANDN U6033 ( .A(n40885), .B(n42047), .Z(n4003) );
  NANDN U6034 ( .A(n40922), .B(n4067), .Z(n4004) );
  NAND U6035 ( .A(n4003), .B(n4004), .Z(n40933) );
  NANDN U6036 ( .A(n40960), .B(n4068), .Z(n4005) );
  NANDN U6037 ( .A(n40926), .B(n42115), .Z(n4006) );
  AND U6038 ( .A(n4005), .B(n4006), .Z(n40965) );
  NANDN U6039 ( .A(n40959), .B(n42047), .Z(n4007) );
  NANDN U6040 ( .A(n40996), .B(n4067), .Z(n4008) );
  NAND U6041 ( .A(n4007), .B(n4008), .Z(n41007) );
  NANDN U6042 ( .A(n41034), .B(n4068), .Z(n4009) );
  NANDN U6043 ( .A(n41000), .B(n42115), .Z(n4010) );
  AND U6044 ( .A(n4009), .B(n4010), .Z(n41039) );
  NANDN U6045 ( .A(n41033), .B(n42047), .Z(n4011) );
  NANDN U6046 ( .A(n41070), .B(n4067), .Z(n4012) );
  NAND U6047 ( .A(n4011), .B(n4012), .Z(n41081) );
  NANDN U6048 ( .A(n41108), .B(n4068), .Z(n4013) );
  NANDN U6049 ( .A(n41071), .B(n42115), .Z(n4014) );
  AND U6050 ( .A(n4013), .B(n4014), .Z(n41113) );
  NANDN U6051 ( .A(n41107), .B(n42047), .Z(n4015) );
  NANDN U6052 ( .A(n41144), .B(n4067), .Z(n4016) );
  NAND U6053 ( .A(n4015), .B(n4016), .Z(n41155) );
  NANDN U6054 ( .A(n41185), .B(n4068), .Z(n4017) );
  NANDN U6055 ( .A(n41148), .B(n42115), .Z(n4018) );
  AND U6056 ( .A(n4017), .B(n4018), .Z(n41187) );
  NANDN U6057 ( .A(n41181), .B(n42047), .Z(n4019) );
  NANDN U6058 ( .A(n41218), .B(n4067), .Z(n4020) );
  NAND U6059 ( .A(n4019), .B(n4020), .Z(n41229) );
  NANDN U6060 ( .A(n41259), .B(n4068), .Z(n4021) );
  NANDN U6061 ( .A(n41219), .B(n42115), .Z(n4022) );
  AND U6062 ( .A(n4021), .B(n4022), .Z(n41261) );
  NANDN U6063 ( .A(n41255), .B(n42047), .Z(n4023) );
  NANDN U6064 ( .A(n41292), .B(n4067), .Z(n4024) );
  NAND U6065 ( .A(n4023), .B(n4024), .Z(n41303) );
  NANDN U6066 ( .A(n41333), .B(n4068), .Z(n4025) );
  NANDN U6067 ( .A(n41293), .B(n42115), .Z(n4026) );
  AND U6068 ( .A(n4025), .B(n4026), .Z(n41335) );
  NANDN U6069 ( .A(n41329), .B(n42047), .Z(n4027) );
  NANDN U6070 ( .A(n41366), .B(n4067), .Z(n4028) );
  NAND U6071 ( .A(n4027), .B(n4028), .Z(n41377) );
  NANDN U6072 ( .A(n41407), .B(n4068), .Z(n4029) );
  NANDN U6073 ( .A(n41367), .B(n42115), .Z(n4030) );
  AND U6074 ( .A(n4029), .B(n4030), .Z(n41409) );
  NANDN U6075 ( .A(n41403), .B(n42047), .Z(n4031) );
  NANDN U6076 ( .A(n41440), .B(n4067), .Z(n4032) );
  NAND U6077 ( .A(n4031), .B(n4032), .Z(n41451) );
  NANDN U6078 ( .A(n41481), .B(n4068), .Z(n4033) );
  NANDN U6079 ( .A(n41444), .B(n42115), .Z(n4034) );
  AND U6080 ( .A(n4033), .B(n4034), .Z(n41483) );
  NANDN U6081 ( .A(n41477), .B(n42047), .Z(n4035) );
  NANDN U6082 ( .A(n41514), .B(n4067), .Z(n4036) );
  NAND U6083 ( .A(n4035), .B(n4036), .Z(n41525) );
  NANDN U6084 ( .A(n41555), .B(n4068), .Z(n4037) );
  NANDN U6085 ( .A(n41518), .B(n42115), .Z(n4038) );
  AND U6086 ( .A(n4037), .B(n4038), .Z(n41557) );
  NANDN U6087 ( .A(n41551), .B(n42047), .Z(n4039) );
  NANDN U6088 ( .A(n41588), .B(n4067), .Z(n4040) );
  NAND U6089 ( .A(n4039), .B(n4040), .Z(n41599) );
  NANDN U6090 ( .A(n41626), .B(n4068), .Z(n4041) );
  NANDN U6091 ( .A(n41592), .B(n42115), .Z(n4042) );
  AND U6092 ( .A(n4041), .B(n4042), .Z(n41631) );
  NANDN U6093 ( .A(n41625), .B(n42047), .Z(n4043) );
  NANDN U6094 ( .A(n41662), .B(n4067), .Z(n4044) );
  NAND U6095 ( .A(n4043), .B(n4044), .Z(n41673) );
  NANDN U6096 ( .A(n41700), .B(n4068), .Z(n4045) );
  NANDN U6097 ( .A(n41666), .B(n42115), .Z(n4046) );
  AND U6098 ( .A(n4045), .B(n4046), .Z(n41705) );
  NANDN U6099 ( .A(n41699), .B(n42047), .Z(n4047) );
  NANDN U6100 ( .A(n41736), .B(n4067), .Z(n4048) );
  NAND U6101 ( .A(n4047), .B(n4048), .Z(n41747) );
  NANDN U6102 ( .A(n41777), .B(n4068), .Z(n4049) );
  NANDN U6103 ( .A(n41737), .B(n42115), .Z(n4050) );
  AND U6104 ( .A(n4049), .B(n4050), .Z(n41779) );
  NANDN U6105 ( .A(n41773), .B(n42047), .Z(n4051) );
  NANDN U6106 ( .A(n41810), .B(n4067), .Z(n4052) );
  NAND U6107 ( .A(n4051), .B(n4052), .Z(n41821) );
  NANDN U6108 ( .A(n41848), .B(n4068), .Z(n4053) );
  NANDN U6109 ( .A(n41811), .B(n42115), .Z(n4054) );
  AND U6110 ( .A(n4053), .B(n4054), .Z(n41853) );
  NANDN U6111 ( .A(n41847), .B(n42047), .Z(n4055) );
  NANDN U6112 ( .A(n4064), .B(n41884), .Z(n4056) );
  NAND U6113 ( .A(n4055), .B(n4056), .Z(n41899) );
  XOR U6114 ( .A(n42089), .B(n42088), .Z(n42090) );
  NANDN U6115 ( .A(n4303), .B(n4067), .Z(n4057) );
  NANDN U6116 ( .A(n4269), .B(n42047), .Z(n4058) );
  AND U6117 ( .A(n4057), .B(n4058), .Z(n4308) );
  NAND U6118 ( .A(n4300), .B(n42115), .Z(n4059) );
  NANDN U6119 ( .A(n4065), .B(n4319), .Z(n4060) );
  AND U6120 ( .A(n4059), .B(n4060), .Z(n4340) );
  XOR U6121 ( .A(n41917), .B(n41916), .Z(n41918) );
  XOR U6122 ( .A(n41965), .B(n41964), .Z(n41985) );
  XNOR U6123 ( .A(n42024), .B(n42023), .Z(n41993) );
  XNOR U6124 ( .A(n42038), .B(n42037), .Z(n42029) );
  XOR U6125 ( .A(n42072), .B(n42071), .Z(n42063) );
  XOR U6126 ( .A(n4256), .B(n4254), .Z(n4061) );
  NANDN U6127 ( .A(n4255), .B(n4061), .Z(n4062) );
  NAND U6128 ( .A(n4256), .B(n4254), .Z(n4063) );
  AND U6129 ( .A(n4062), .B(n4063), .Z(n4268) );
  XOR U6130 ( .A(n41959), .B(n41958), .Z(n41951) );
  XOR U6131 ( .A(n42097), .B(n42096), .Z(n42098) );
  XOR U6132 ( .A(n42130), .B(n42129), .Z(n42131) );
  XOR U6133 ( .A(n42170), .B(n42169), .Z(n42172) );
  XNOR U6134 ( .A(n42190), .B(n42191), .Z(n42179) );
  XNOR U6135 ( .A(b[1]), .B(b[2]), .Z(n4064) );
  XNOR U6136 ( .A(b[3]), .B(b[4]), .Z(n4065) );
  IV U6137 ( .A(n42047), .Z(n4066) );
  IV U6138 ( .A(n4064), .Z(n4067) );
  IV U6139 ( .A(n4065), .Z(n4068) );
  IV U6140 ( .A(n42143), .Z(n4069) );
  IV U6141 ( .A(n42144), .Z(n4070) );
  IV U6142 ( .A(b[1]), .Z(n4071) );
  IV U6143 ( .A(b[7]), .Z(n4072) );
  IV U6144 ( .A(b[7]), .Z(n4073) );
  IV U6145 ( .A(b[7]), .Z(n4074) );
  IV U6146 ( .A(b[7]), .Z(n4075) );
  IV U6147 ( .A(b[7]), .Z(n4076) );
  IV U6148 ( .A(b[7]), .Z(n4077) );
  IV U6149 ( .A(b[7]), .Z(n4078) );
  IV U6150 ( .A(b[7]), .Z(n4079) );
  IV U6151 ( .A(b[7]), .Z(n4080) );
  IV U6152 ( .A(b[7]), .Z(n4081) );
  IV U6153 ( .A(b[7]), .Z(n4082) );
  IV U6154 ( .A(b[7]), .Z(n4083) );
  IV U6155 ( .A(b[7]), .Z(n4084) );
  IV U6156 ( .A(b[7]), .Z(n4085) );
  IV U6157 ( .A(b[7]), .Z(n4086) );
  IV U6158 ( .A(b[7]), .Z(n4087) );
  IV U6159 ( .A(b[7]), .Z(n4088) );
  IV U6160 ( .A(b[7]), .Z(n4089) );
  IV U6161 ( .A(b[7]), .Z(n4090) );
  IV U6162 ( .A(b[7]), .Z(n4091) );
  IV U6163 ( .A(b[7]), .Z(n4092) );
  IV U6164 ( .A(b[7]), .Z(n4093) );
  IV U6165 ( .A(b[7]), .Z(n4094) );
  IV U6166 ( .A(b[7]), .Z(n4095) );
  IV U6167 ( .A(b[7]), .Z(n4096) );
  IV U6168 ( .A(b[7]), .Z(n4097) );
  IV U6169 ( .A(b[7]), .Z(n4098) );
  IV U6170 ( .A(b[7]), .Z(n4099) );
  IV U6171 ( .A(b[7]), .Z(n4100) );
  IV U6172 ( .A(b[7]), .Z(n4101) );
  IV U6173 ( .A(b[7]), .Z(n4102) );
  IV U6174 ( .A(b[7]), .Z(n4103) );
  IV U6175 ( .A(b[7]), .Z(n4104) );
  IV U6176 ( .A(b[7]), .Z(n4105) );
  IV U6177 ( .A(b[7]), .Z(n4106) );
  IV U6178 ( .A(b[7]), .Z(n4107) );
  IV U6179 ( .A(b[7]), .Z(n4108) );
  IV U6180 ( .A(b[7]), .Z(n4109) );
  IV U6181 ( .A(b[7]), .Z(n4110) );
  IV U6182 ( .A(b[7]), .Z(n4111) );
  IV U6183 ( .A(b[7]), .Z(n4112) );
  IV U6184 ( .A(b[7]), .Z(n4113) );
  IV U6185 ( .A(b[7]), .Z(n4114) );
  IV U6186 ( .A(b[7]), .Z(n4115) );
  IV U6187 ( .A(b[7]), .Z(n4116) );
  IV U6188 ( .A(b[7]), .Z(n4117) );
  IV U6189 ( .A(b[7]), .Z(n4118) );
  IV U6190 ( .A(b[7]), .Z(n4119) );
  IV U6191 ( .A(b[7]), .Z(n4120) );
  IV U6192 ( .A(b[7]), .Z(n4121) );
  IV U6193 ( .A(b[7]), .Z(n4122) );
  IV U6194 ( .A(b[7]), .Z(n4123) );
  IV U6195 ( .A(b[7]), .Z(n4124) );
  IV U6196 ( .A(b[7]), .Z(n4125) );
  IV U6197 ( .A(b[7]), .Z(n4126) );
  IV U6198 ( .A(b[7]), .Z(n4127) );
  IV U6199 ( .A(b[7]), .Z(n4128) );
  IV U6200 ( .A(b[7]), .Z(n4129) );
  IV U6201 ( .A(b[7]), .Z(n4130) );
  IV U6202 ( .A(b[7]), .Z(n4131) );
  IV U6203 ( .A(b[7]), .Z(n4132) );
  IV U6204 ( .A(b[7]), .Z(n4133) );
  IV U6205 ( .A(b[7]), .Z(n4134) );
  IV U6206 ( .A(b[7]), .Z(n4135) );
  IV U6207 ( .A(b[7]), .Z(n4136) );
  IV U6208 ( .A(b[7]), .Z(n4137) );
  IV U6209 ( .A(b[7]), .Z(n4138) );
  IV U6210 ( .A(b[7]), .Z(n4139) );
  IV U6211 ( .A(b[7]), .Z(n4140) );
  IV U6212 ( .A(b[7]), .Z(n4141) );
  IV U6213 ( .A(b[7]), .Z(n4142) );
  IV U6214 ( .A(b[7]), .Z(n4143) );
  IV U6215 ( .A(b[7]), .Z(n4144) );
  IV U6216 ( .A(b[7]), .Z(n4145) );
  IV U6217 ( .A(b[7]), .Z(n4146) );
  IV U6218 ( .A(b[7]), .Z(n4147) );
  IV U6219 ( .A(b[7]), .Z(n4148) );
  IV U6220 ( .A(b[7]), .Z(n4149) );
  IV U6221 ( .A(b[7]), .Z(n4150) );
  IV U6222 ( .A(b[7]), .Z(n4151) );
  IV U6223 ( .A(b[7]), .Z(n4152) );
  IV U6224 ( .A(b[7]), .Z(n4153) );
  IV U6225 ( .A(b[7]), .Z(n4154) );
  IV U6226 ( .A(b[7]), .Z(n4155) );
  IV U6227 ( .A(b[7]), .Z(n4156) );
  IV U6228 ( .A(b[7]), .Z(n4157) );
  IV U6229 ( .A(b[7]), .Z(n4158) );
  IV U6230 ( .A(b[7]), .Z(n4159) );
  IV U6231 ( .A(b[7]), .Z(n4160) );
  IV U6232 ( .A(b[7]), .Z(n4161) );
  IV U6233 ( .A(b[7]), .Z(n4162) );
  IV U6234 ( .A(b[7]), .Z(n4163) );
  IV U6235 ( .A(b[7]), .Z(n4164) );
  IV U6236 ( .A(b[7]), .Z(n4165) );
  IV U6237 ( .A(b[7]), .Z(n4166) );
  IV U6238 ( .A(b[7]), .Z(n4167) );
  IV U6239 ( .A(b[7]), .Z(n4168) );
  IV U6240 ( .A(b[7]), .Z(n4169) );
  IV U6241 ( .A(b[7]), .Z(n4170) );
  IV U6242 ( .A(b[7]), .Z(n4171) );
  IV U6243 ( .A(b[7]), .Z(n4172) );
  IV U6244 ( .A(b[7]), .Z(n4173) );
  IV U6245 ( .A(b[7]), .Z(n4174) );
  IV U6246 ( .A(b[7]), .Z(n4175) );
  IV U6247 ( .A(b[7]), .Z(n4176) );
  IV U6248 ( .A(b[7]), .Z(n4177) );
  IV U6249 ( .A(b[7]), .Z(n4178) );
  IV U6250 ( .A(b[7]), .Z(n4179) );
  IV U6251 ( .A(b[7]), .Z(n4180) );
  IV U6252 ( .A(b[7]), .Z(n4181) );
  IV U6253 ( .A(b[7]), .Z(n4182) );
  IV U6254 ( .A(b[7]), .Z(n4183) );
  IV U6255 ( .A(b[7]), .Z(n4184) );
  IV U6256 ( .A(b[7]), .Z(n4185) );
  IV U6257 ( .A(b[7]), .Z(n4186) );
  IV U6258 ( .A(b[7]), .Z(n4187) );
  IV U6259 ( .A(b[7]), .Z(n4188) );
  IV U6260 ( .A(b[7]), .Z(n4189) );
  IV U6261 ( .A(b[7]), .Z(n4190) );
  IV U6262 ( .A(b[7]), .Z(n4191) );
  IV U6263 ( .A(b[7]), .Z(n4192) );
  IV U6264 ( .A(b[7]), .Z(n4193) );
  IV U6265 ( .A(b[7]), .Z(n4194) );
  IV U6266 ( .A(b[7]), .Z(n4195) );
  IV U6267 ( .A(b[7]), .Z(n4196) );
  IV U6268 ( .A(b[7]), .Z(n4197) );
  IV U6269 ( .A(b[7]), .Z(n4198) );
  IV U6270 ( .A(b[7]), .Z(n4199) );
  IV U6271 ( .A(b[7]), .Z(n4200) );
  IV U6272 ( .A(b[7]), .Z(n4201) );
  IV U6273 ( .A(b[7]), .Z(n4202) );
  IV U6274 ( .A(b[7]), .Z(n4203) );
  IV U6275 ( .A(b[7]), .Z(n4204) );
  IV U6276 ( .A(b[7]), .Z(n4205) );
  IV U6277 ( .A(b[7]), .Z(n4206) );
  IV U6278 ( .A(b[7]), .Z(n4207) );
  IV U6279 ( .A(b[7]), .Z(n4208) );
  IV U6280 ( .A(b[7]), .Z(n4209) );
  IV U6281 ( .A(b[7]), .Z(n4210) );
  IV U6282 ( .A(b[7]), .Z(n4211) );
  IV U6283 ( .A(b[7]), .Z(n4212) );
  IV U6284 ( .A(b[7]), .Z(n4213) );
  IV U6285 ( .A(b[7]), .Z(n4214) );
  IV U6286 ( .A(b[7]), .Z(n4215) );
  IV U6287 ( .A(b[7]), .Z(n4216) );
  IV U6288 ( .A(b[7]), .Z(n4217) );
  AND U6289 ( .A(b[0]), .B(a[0]), .Z(n4219) );
  XOR U6290 ( .A(n4219), .B(sreg[1016]), .Z(c[1016]) );
  AND U6291 ( .A(b[0]), .B(a[1]), .Z(n4226) );
  NAND U6292 ( .A(b[1]), .B(a[0]), .Z(n4218) );
  XOR U6293 ( .A(n4226), .B(n4218), .Z(n4220) );
  XNOR U6294 ( .A(sreg[1017]), .B(n4220), .Z(n4222) );
  AND U6295 ( .A(n4219), .B(sreg[1016]), .Z(n4221) );
  XOR U6296 ( .A(n4222), .B(n4221), .Z(c[1017]) );
  NANDN U6297 ( .A(n4220), .B(sreg[1017]), .Z(n4224) );
  NAND U6298 ( .A(n4222), .B(n4221), .Z(n4223) );
  AND U6299 ( .A(n4224), .B(n4223), .Z(n4244) );
  XNOR U6300 ( .A(n4244), .B(sreg[1018]), .Z(n4246) );
  AND U6301 ( .A(b[2]), .B(a[0]), .Z(n4225) );
  XNOR U6302 ( .A(n4225), .B(n4071), .Z(n4228) );
  NANDN U6303 ( .A(a[0]), .B(n4226), .Z(n4227) );
  NAND U6304 ( .A(n4228), .B(n4227), .Z(n4233) );
  AND U6305 ( .A(a[2]), .B(b[0]), .Z(n4229) );
  XNOR U6306 ( .A(n4229), .B(n4071), .Z(n4231) );
  NANDN U6307 ( .A(b[0]), .B(a[1]), .Z(n4230) );
  NAND U6308 ( .A(n4231), .B(n4230), .Z(n4232) );
  XOR U6309 ( .A(n4233), .B(n4232), .Z(n4245) );
  XOR U6310 ( .A(n4246), .B(n4245), .Z(c[1018]) );
  NOR U6311 ( .A(n4233), .B(n4232), .Z(n4256) );
  XOR U6312 ( .A(b[2]), .B(b[3]), .Z(n4234) );
  AND U6313 ( .A(n4234), .B(n4064), .Z(n42047) );
  XOR U6314 ( .A(a[0]), .B(b[3]), .Z(n4235) );
  NAND U6315 ( .A(n42047), .B(n4235), .Z(n4237) );
  IV U6316 ( .A(b[3]), .Z(n42012) );
  XNOR U6317 ( .A(a[1]), .B(n42012), .Z(n4257) );
  AND U6318 ( .A(n4257), .B(n4067), .Z(n4236) );
  ANDN U6319 ( .B(n4237), .A(n4236), .Z(n4264) );
  AND U6320 ( .A(a[3]), .B(b[0]), .Z(n4238) );
  XNOR U6321 ( .A(n4238), .B(n4071), .Z(n4240) );
  NANDN U6322 ( .A(b[0]), .B(a[2]), .Z(n4239) );
  NAND U6323 ( .A(n4240), .B(n4239), .Z(n4263) );
  XNOR U6324 ( .A(n4264), .B(n4263), .Z(n4255) );
  NAND U6325 ( .A(n4067), .B(a[0]), .Z(n4242) );
  NAND U6326 ( .A(b[1]), .B(b[2]), .Z(n4241) );
  AND U6327 ( .A(n4241), .B(b[3]), .Z(n42124) );
  AND U6328 ( .A(n4242), .B(n42124), .Z(n4254) );
  XOR U6329 ( .A(n4255), .B(n4254), .Z(n4243) );
  XOR U6330 ( .A(n4256), .B(n4243), .Z(n4249) );
  XNOR U6331 ( .A(sreg[1019]), .B(n4249), .Z(n4251) );
  NANDN U6332 ( .A(n4244), .B(sreg[1018]), .Z(n4248) );
  NAND U6333 ( .A(n4246), .B(n4245), .Z(n4247) );
  NAND U6334 ( .A(n4248), .B(n4247), .Z(n4250) );
  XOR U6335 ( .A(n4251), .B(n4250), .Z(c[1019]) );
  NANDN U6336 ( .A(n4249), .B(sreg[1019]), .Z(n4253) );
  NAND U6337 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U6338 ( .A(n4253), .B(n4252), .Z(n4284) );
  XNOR U6339 ( .A(n4284), .B(sreg[1020]), .Z(n4286) );
  XOR U6340 ( .A(a[2]), .B(n42012), .Z(n4269) );
  NANDN U6341 ( .A(n4269), .B(n4067), .Z(n4259) );
  NAND U6342 ( .A(n42047), .B(n4257), .Z(n4258) );
  AND U6343 ( .A(n4259), .B(n4258), .Z(n4281) );
  AND U6344 ( .A(a[0]), .B(n4068), .Z(n4278) );
  AND U6345 ( .A(a[4]), .B(b[0]), .Z(n4260) );
  XNOR U6346 ( .A(n4260), .B(n4071), .Z(n4262) );
  NANDN U6347 ( .A(b[0]), .B(a[3]), .Z(n4261) );
  NAND U6348 ( .A(n4262), .B(n4261), .Z(n4279) );
  XNOR U6349 ( .A(n4278), .B(n4279), .Z(n4280) );
  XNOR U6350 ( .A(n4281), .B(n4280), .Z(n4266) );
  OR U6351 ( .A(n4264), .B(n4263), .Z(n4265) );
  XNOR U6352 ( .A(n4266), .B(n4265), .Z(n4267) );
  XNOR U6353 ( .A(n4268), .B(n4267), .Z(n4285) );
  XOR U6354 ( .A(n4286), .B(n4285), .Z(c[1020]) );
  XOR U6355 ( .A(a[3]), .B(n42012), .Z(n4303) );
  NAND U6356 ( .A(b[3]), .B(b[4]), .Z(n4270) );
  AND U6357 ( .A(n4270), .B(b[5]), .Z(n42141) );
  IV U6358 ( .A(n42141), .Z(n42154) );
  NOR U6359 ( .A(n42154), .B(n4278), .Z(n4307) );
  XNOR U6360 ( .A(n4308), .B(n4307), .Z(n4310) );
  XOR U6361 ( .A(b[5]), .B(a[1]), .Z(n4300) );
  AND U6362 ( .A(n4068), .B(n4300), .Z(n4274) );
  XOR U6363 ( .A(b[5]), .B(b[4]), .Z(n4271) );
  AND U6364 ( .A(n4271), .B(n4065), .Z(n42115) );
  XOR U6365 ( .A(a[0]), .B(b[5]), .Z(n4272) );
  NAND U6366 ( .A(n42115), .B(n4272), .Z(n4273) );
  NANDN U6367 ( .A(n4274), .B(n4273), .Z(n4302) );
  AND U6368 ( .A(a[5]), .B(b[0]), .Z(n4275) );
  XNOR U6369 ( .A(n4275), .B(n4071), .Z(n4277) );
  NANDN U6370 ( .A(b[0]), .B(a[4]), .Z(n4276) );
  NAND U6371 ( .A(n4277), .B(n4276), .Z(n4301) );
  XNOR U6372 ( .A(n4302), .B(n4301), .Z(n4309) );
  XOR U6373 ( .A(n4310), .B(n4309), .Z(n4295) );
  NANDN U6374 ( .A(n4279), .B(n4278), .Z(n4283) );
  NANDN U6375 ( .A(n4281), .B(n4280), .Z(n4282) );
  AND U6376 ( .A(n4283), .B(n4282), .Z(n4294) );
  XNOR U6377 ( .A(n4295), .B(n4294), .Z(n4296) );
  XOR U6378 ( .A(n4297), .B(n4296), .Z(n4289) );
  XNOR U6379 ( .A(n4289), .B(sreg[1021]), .Z(n4291) );
  NANDN U6380 ( .A(n4284), .B(sreg[1020]), .Z(n4288) );
  NAND U6381 ( .A(n4286), .B(n4285), .Z(n4287) );
  NAND U6382 ( .A(n4288), .B(n4287), .Z(n4290) );
  XOR U6383 ( .A(n4291), .B(n4290), .Z(c[1021]) );
  NANDN U6384 ( .A(n4289), .B(sreg[1021]), .Z(n4293) );
  NAND U6385 ( .A(n4291), .B(n4290), .Z(n4292) );
  AND U6386 ( .A(n4293), .B(n4292), .Z(n4345) );
  XNOR U6387 ( .A(n4345), .B(sreg[1022]), .Z(n4347) );
  NANDN U6388 ( .A(n4295), .B(n4294), .Z(n4299) );
  NAND U6389 ( .A(n4297), .B(n4296), .Z(n4298) );
  AND U6390 ( .A(n4299), .B(n4298), .Z(n4315) );
  XOR U6391 ( .A(a[2]), .B(b[5]), .Z(n4319) );
  ANDN U6392 ( .B(n4302), .A(n4301), .Z(n4339) );
  XNOR U6393 ( .A(n4340), .B(n4339), .Z(n4342) );
  XNOR U6394 ( .A(b[3]), .B(a[4]), .Z(n4330) );
  XOR U6395 ( .A(b[5]), .B(b[6]), .Z(n42144) );
  AND U6396 ( .A(a[0]), .B(n42144), .Z(n4333) );
  AND U6397 ( .A(a[6]), .B(b[0]), .Z(n4304) );
  XNOR U6398 ( .A(n4304), .B(n4071), .Z(n4306) );
  NANDN U6399 ( .A(b[0]), .B(a[5]), .Z(n4305) );
  NAND U6400 ( .A(n4306), .B(n4305), .Z(n4334) );
  XNOR U6401 ( .A(n4333), .B(n4334), .Z(n4335) );
  XNOR U6402 ( .A(n4336), .B(n4335), .Z(n4341) );
  XOR U6403 ( .A(n4342), .B(n4341), .Z(n4314) );
  NANDN U6404 ( .A(n4308), .B(n4307), .Z(n4312) );
  NAND U6405 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U6406 ( .A(n4312), .B(n4311), .Z(n4313) );
  XOR U6407 ( .A(n4314), .B(n4313), .Z(n4316) );
  XNOR U6408 ( .A(n4315), .B(n4316), .Z(n4346) );
  XOR U6409 ( .A(n4347), .B(n4346), .Z(c[1022]) );
  NANDN U6410 ( .A(n4314), .B(n4313), .Z(n4318) );
  OR U6411 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U6412 ( .A(n4318), .B(n4317), .Z(n4376) );
  IV U6413 ( .A(b[5]), .Z(n42085) );
  XOR U6414 ( .A(a[3]), .B(n42085), .Z(n4367) );
  NANDN U6415 ( .A(n4367), .B(n4068), .Z(n4321) );
  NAND U6416 ( .A(n4319), .B(n42115), .Z(n4320) );
  AND U6417 ( .A(n4321), .B(n4320), .Z(n4357) );
  XOR U6418 ( .A(b[6]), .B(b[7]), .Z(n4322) );
  AND U6419 ( .A(n4322), .B(n4070), .Z(n42143) );
  XOR U6420 ( .A(a[0]), .B(b[7]), .Z(n4323) );
  NAND U6421 ( .A(n42143), .B(n4323), .Z(n4325) );
  XOR U6422 ( .A(b[7]), .B(a[1]), .Z(n4358) );
  AND U6423 ( .A(n4358), .B(n42144), .Z(n4324) );
  ANDN U6424 ( .B(n4325), .A(n4324), .Z(n4356) );
  XOR U6425 ( .A(n4357), .B(n4356), .Z(n4371) );
  AND U6426 ( .A(b[6]), .B(b[5]), .Z(n42186) );
  NOR U6427 ( .A(n42186), .B(n4333), .Z(n4326) );
  AND U6428 ( .A(n4326), .B(b[7]), .Z(n4369) );
  AND U6429 ( .A(a[7]), .B(b[0]), .Z(n4327) );
  XNOR U6430 ( .A(n4327), .B(n4071), .Z(n4329) );
  NANDN U6431 ( .A(b[0]), .B(a[6]), .Z(n4328) );
  NAND U6432 ( .A(n4329), .B(n4328), .Z(n4368) );
  XNOR U6433 ( .A(n4369), .B(n4368), .Z(n4370) );
  XNOR U6434 ( .A(n4371), .B(n4370), .Z(n4350) );
  OR U6435 ( .A(n4330), .B(n4066), .Z(n4332) );
  XNOR U6436 ( .A(b[3]), .B(a[5]), .Z(n4361) );
  OR U6437 ( .A(n4361), .B(n4064), .Z(n4331) );
  NAND U6438 ( .A(n4332), .B(n4331), .Z(n4351) );
  XNOR U6439 ( .A(n4350), .B(n4351), .Z(n4352) );
  NANDN U6440 ( .A(n4334), .B(n4333), .Z(n4338) );
  NANDN U6441 ( .A(n4336), .B(n4335), .Z(n4337) );
  NAND U6442 ( .A(n4338), .B(n4337), .Z(n4353) );
  XNOR U6443 ( .A(n4352), .B(n4353), .Z(n4374) );
  NANDN U6444 ( .A(n4340), .B(n4339), .Z(n4344) );
  NAND U6445 ( .A(n4342), .B(n4341), .Z(n4343) );
  NAND U6446 ( .A(n4344), .B(n4343), .Z(n4375) );
  XOR U6447 ( .A(n4374), .B(n4375), .Z(n4377) );
  XOR U6448 ( .A(n4376), .B(n4377), .Z(n4380) );
  XNOR U6449 ( .A(n4380), .B(sreg[1023]), .Z(n4382) );
  NANDN U6450 ( .A(n4345), .B(sreg[1022]), .Z(n4349) );
  NAND U6451 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U6452 ( .A(n4349), .B(n4348), .Z(n4381) );
  XOR U6453 ( .A(n4382), .B(n4381), .Z(c[1023]) );
  NANDN U6454 ( .A(n4351), .B(n4350), .Z(n4355) );
  NANDN U6455 ( .A(n4353), .B(n4352), .Z(n4354) );
  AND U6456 ( .A(n4355), .B(n4354), .Z(n4385) );
  NOR U6457 ( .A(n4357), .B(n4356), .Z(n4409) );
  NANDN U6458 ( .A(n4069), .B(n4358), .Z(n4360) );
  XOR U6459 ( .A(a[2]), .B(b[7]), .Z(n4397) );
  NANDN U6460 ( .A(n4070), .B(n4397), .Z(n4359) );
  AND U6461 ( .A(n4360), .B(n4359), .Z(n4407) );
  OR U6462 ( .A(n4361), .B(n4066), .Z(n4363) );
  XOR U6463 ( .A(a[6]), .B(b[3]), .Z(n4400) );
  NANDN U6464 ( .A(n4064), .B(n4400), .Z(n4362) );
  NAND U6465 ( .A(n4363), .B(n4362), .Z(n4408) );
  XOR U6466 ( .A(n4407), .B(n4408), .Z(n4410) );
  XOR U6467 ( .A(n4409), .B(n4410), .Z(n4414) );
  AND U6468 ( .A(a[8]), .B(b[0]), .Z(n4364) );
  XNOR U6469 ( .A(n4364), .B(n4071), .Z(n4366) );
  NANDN U6470 ( .A(b[0]), .B(a[7]), .Z(n4365) );
  NAND U6471 ( .A(n4366), .B(n4365), .Z(n4394) );
  XOR U6472 ( .A(a[4]), .B(n42085), .Z(n4403) );
  AND U6473 ( .A(a[0]), .B(b[7]), .Z(n4391) );
  XNOR U6474 ( .A(n4392), .B(n4391), .Z(n4393) );
  XNOR U6475 ( .A(n4394), .B(n4393), .Z(n4413) );
  XNOR U6476 ( .A(n4414), .B(n4413), .Z(n4415) );
  NANDN U6477 ( .A(n4369), .B(n4368), .Z(n4373) );
  NANDN U6478 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U6479 ( .A(n4373), .B(n4372), .Z(n4416) );
  XOR U6480 ( .A(n4415), .B(n4416), .Z(n4386) );
  XNOR U6481 ( .A(n4385), .B(n4386), .Z(n4387) );
  NANDN U6482 ( .A(n4375), .B(n4374), .Z(n4379) );
  OR U6483 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U6484 ( .A(n4379), .B(n4378), .Z(n4388) );
  XNOR U6485 ( .A(n4387), .B(n4388), .Z(n4421) );
  NANDN U6486 ( .A(n4380), .B(sreg[1023]), .Z(n4384) );
  NAND U6487 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U6488 ( .A(n4384), .B(n4383), .Z(n4419) );
  XNOR U6489 ( .A(n4419), .B(sreg[1024]), .Z(n4420) );
  XOR U6490 ( .A(n4421), .B(n4420), .Z(c[1024]) );
  NANDN U6491 ( .A(n4386), .B(n4385), .Z(n4390) );
  NANDN U6492 ( .A(n4388), .B(n4387), .Z(n4389) );
  AND U6493 ( .A(n4390), .B(n4389), .Z(n4427) );
  NANDN U6494 ( .A(n4392), .B(n4391), .Z(n4396) );
  NANDN U6495 ( .A(n4394), .B(n4393), .Z(n4395) );
  AND U6496 ( .A(n4396), .B(n4395), .Z(n4451) );
  NAND U6497 ( .A(n42143), .B(n4397), .Z(n4399) );
  XNOR U6498 ( .A(a[3]), .B(n4072), .Z(n4430) );
  NAND U6499 ( .A(n42144), .B(n4430), .Z(n4398) );
  AND U6500 ( .A(n4399), .B(n4398), .Z(n4445) );
  XOR U6501 ( .A(a[7]), .B(n42012), .Z(n4433) );
  NANDN U6502 ( .A(n4433), .B(n4067), .Z(n4402) );
  NAND U6503 ( .A(n42047), .B(n4400), .Z(n4401) );
  NAND U6504 ( .A(n4402), .B(n4401), .Z(n4444) );
  XNOR U6505 ( .A(n4445), .B(n4444), .Z(n4446) );
  XOR U6506 ( .A(a[5]), .B(n42085), .Z(n4437) );
  AND U6507 ( .A(a[1]), .B(b[7]), .Z(n4438) );
  XNOR U6508 ( .A(n4439), .B(n4438), .Z(n4440) );
  AND U6509 ( .A(a[9]), .B(b[0]), .Z(n4404) );
  XNOR U6510 ( .A(n4404), .B(n4071), .Z(n4406) );
  NANDN U6511 ( .A(b[0]), .B(a[8]), .Z(n4405) );
  NAND U6512 ( .A(n4406), .B(n4405), .Z(n4441) );
  XOR U6513 ( .A(n4440), .B(n4441), .Z(n4447) );
  XNOR U6514 ( .A(n4446), .B(n4447), .Z(n4450) );
  XNOR U6515 ( .A(n4451), .B(n4450), .Z(n4453) );
  NANDN U6516 ( .A(n4408), .B(n4407), .Z(n4412) );
  OR U6517 ( .A(n4410), .B(n4409), .Z(n4411) );
  AND U6518 ( .A(n4412), .B(n4411), .Z(n4452) );
  XOR U6519 ( .A(n4453), .B(n4452), .Z(n4425) );
  NANDN U6520 ( .A(n4414), .B(n4413), .Z(n4418) );
  NANDN U6521 ( .A(n4416), .B(n4415), .Z(n4417) );
  AND U6522 ( .A(n4418), .B(n4417), .Z(n4424) );
  XNOR U6523 ( .A(n4425), .B(n4424), .Z(n4426) );
  XOR U6524 ( .A(n4427), .B(n4426), .Z(n4456) );
  XNOR U6525 ( .A(n4456), .B(sreg[1025]), .Z(n4458) );
  NANDN U6526 ( .A(n4419), .B(sreg[1024]), .Z(n4423) );
  NAND U6527 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U6528 ( .A(n4423), .B(n4422), .Z(n4457) );
  XOR U6529 ( .A(n4458), .B(n4457), .Z(c[1025]) );
  NANDN U6530 ( .A(n4425), .B(n4424), .Z(n4429) );
  NAND U6531 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U6532 ( .A(n4429), .B(n4428), .Z(n4468) );
  NAND U6533 ( .A(n42143), .B(n4430), .Z(n4432) );
  XNOR U6534 ( .A(a[4]), .B(n4072), .Z(n4478) );
  NAND U6535 ( .A(n42144), .B(n4478), .Z(n4431) );
  AND U6536 ( .A(n4432), .B(n4431), .Z(n4493) );
  XOR U6537 ( .A(a[8]), .B(n42012), .Z(n4481) );
  XNOR U6538 ( .A(n4493), .B(n4492), .Z(n4495) );
  AND U6539 ( .A(a[10]), .B(b[0]), .Z(n4434) );
  XNOR U6540 ( .A(n4434), .B(n4071), .Z(n4436) );
  NANDN U6541 ( .A(b[0]), .B(a[9]), .Z(n4435) );
  NAND U6542 ( .A(n4436), .B(n4435), .Z(n4489) );
  XOR U6543 ( .A(a[6]), .B(n42085), .Z(n4485) );
  AND U6544 ( .A(a[2]), .B(b[7]), .Z(n4486) );
  XNOR U6545 ( .A(n4487), .B(n4486), .Z(n4488) );
  XNOR U6546 ( .A(n4489), .B(n4488), .Z(n4494) );
  XOR U6547 ( .A(n4495), .B(n4494), .Z(n4473) );
  NANDN U6548 ( .A(n4439), .B(n4438), .Z(n4443) );
  NANDN U6549 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U6550 ( .A(n4443), .B(n4442), .Z(n4472) );
  XNOR U6551 ( .A(n4473), .B(n4472), .Z(n4474) );
  NANDN U6552 ( .A(n4445), .B(n4444), .Z(n4449) );
  NANDN U6553 ( .A(n4447), .B(n4446), .Z(n4448) );
  NAND U6554 ( .A(n4449), .B(n4448), .Z(n4475) );
  XNOR U6555 ( .A(n4474), .B(n4475), .Z(n4466) );
  NANDN U6556 ( .A(n4451), .B(n4450), .Z(n4455) );
  NAND U6557 ( .A(n4453), .B(n4452), .Z(n4454) );
  NAND U6558 ( .A(n4455), .B(n4454), .Z(n4467) );
  XOR U6559 ( .A(n4466), .B(n4467), .Z(n4469) );
  XOR U6560 ( .A(n4468), .B(n4469), .Z(n4461) );
  XNOR U6561 ( .A(n4461), .B(sreg[1026]), .Z(n4463) );
  NANDN U6562 ( .A(n4456), .B(sreg[1025]), .Z(n4460) );
  NAND U6563 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U6564 ( .A(n4460), .B(n4459), .Z(n4462) );
  XOR U6565 ( .A(n4463), .B(n4462), .Z(c[1026]) );
  NANDN U6566 ( .A(n4461), .B(sreg[1026]), .Z(n4465) );
  NAND U6567 ( .A(n4463), .B(n4462), .Z(n4464) );
  AND U6568 ( .A(n4465), .B(n4464), .Z(n4532) );
  NANDN U6569 ( .A(n4467), .B(n4466), .Z(n4471) );
  OR U6570 ( .A(n4469), .B(n4468), .Z(n4470) );
  AND U6571 ( .A(n4471), .B(n4470), .Z(n4501) );
  NANDN U6572 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U6573 ( .A(n4475), .B(n4474), .Z(n4476) );
  AND U6574 ( .A(n4477), .B(n4476), .Z(n4499) );
  NAND U6575 ( .A(n42143), .B(n4478), .Z(n4480) );
  XNOR U6576 ( .A(a[5]), .B(n4072), .Z(n4510) );
  NAND U6577 ( .A(n42144), .B(n4510), .Z(n4479) );
  AND U6578 ( .A(n4480), .B(n4479), .Z(n4525) );
  XOR U6579 ( .A(a[9]), .B(n42012), .Z(n4513) );
  XNOR U6580 ( .A(n4525), .B(n4524), .Z(n4527) );
  AND U6581 ( .A(a[11]), .B(b[0]), .Z(n4482) );
  XNOR U6582 ( .A(n4482), .B(n4071), .Z(n4484) );
  NANDN U6583 ( .A(b[0]), .B(a[10]), .Z(n4483) );
  NAND U6584 ( .A(n4484), .B(n4483), .Z(n4521) );
  XOR U6585 ( .A(a[7]), .B(n42085), .Z(n4514) );
  AND U6586 ( .A(a[3]), .B(b[7]), .Z(n4518) );
  XNOR U6587 ( .A(n4519), .B(n4518), .Z(n4520) );
  XNOR U6588 ( .A(n4521), .B(n4520), .Z(n4526) );
  XOR U6589 ( .A(n4527), .B(n4526), .Z(n4505) );
  NANDN U6590 ( .A(n4487), .B(n4486), .Z(n4491) );
  NANDN U6591 ( .A(n4489), .B(n4488), .Z(n4490) );
  AND U6592 ( .A(n4491), .B(n4490), .Z(n4504) );
  XNOR U6593 ( .A(n4505), .B(n4504), .Z(n4506) );
  NANDN U6594 ( .A(n4493), .B(n4492), .Z(n4497) );
  NAND U6595 ( .A(n4495), .B(n4494), .Z(n4496) );
  NAND U6596 ( .A(n4497), .B(n4496), .Z(n4507) );
  XNOR U6597 ( .A(n4506), .B(n4507), .Z(n4498) );
  XNOR U6598 ( .A(n4499), .B(n4498), .Z(n4500) );
  XNOR U6599 ( .A(n4501), .B(n4500), .Z(n4530) );
  XNOR U6600 ( .A(sreg[1027]), .B(n4530), .Z(n4531) );
  XNOR U6601 ( .A(n4532), .B(n4531), .Z(c[1027]) );
  NANDN U6602 ( .A(n4499), .B(n4498), .Z(n4503) );
  NANDN U6603 ( .A(n4501), .B(n4500), .Z(n4502) );
  AND U6604 ( .A(n4503), .B(n4502), .Z(n4538) );
  NANDN U6605 ( .A(n4505), .B(n4504), .Z(n4509) );
  NANDN U6606 ( .A(n4507), .B(n4506), .Z(n4508) );
  AND U6607 ( .A(n4509), .B(n4508), .Z(n4536) );
  NAND U6608 ( .A(n42143), .B(n4510), .Z(n4512) );
  XNOR U6609 ( .A(a[6]), .B(n4072), .Z(n4547) );
  NAND U6610 ( .A(n42144), .B(n4547), .Z(n4511) );
  AND U6611 ( .A(n4512), .B(n4511), .Z(n4562) );
  XOR U6612 ( .A(a[10]), .B(n42012), .Z(n4550) );
  XNOR U6613 ( .A(n4562), .B(n4561), .Z(n4564) );
  XOR U6614 ( .A(a[8]), .B(n42085), .Z(n4554) );
  AND U6615 ( .A(a[4]), .B(b[7]), .Z(n4555) );
  XNOR U6616 ( .A(n4556), .B(n4555), .Z(n4557) );
  AND U6617 ( .A(a[12]), .B(b[0]), .Z(n4515) );
  XNOR U6618 ( .A(n4515), .B(n4071), .Z(n4517) );
  NANDN U6619 ( .A(b[0]), .B(a[11]), .Z(n4516) );
  NAND U6620 ( .A(n4517), .B(n4516), .Z(n4558) );
  XNOR U6621 ( .A(n4557), .B(n4558), .Z(n4563) );
  XOR U6622 ( .A(n4564), .B(n4563), .Z(n4542) );
  NANDN U6623 ( .A(n4519), .B(n4518), .Z(n4523) );
  NANDN U6624 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U6625 ( .A(n4523), .B(n4522), .Z(n4541) );
  XNOR U6626 ( .A(n4542), .B(n4541), .Z(n4543) );
  NANDN U6627 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U6628 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U6629 ( .A(n4529), .B(n4528), .Z(n4544) );
  XNOR U6630 ( .A(n4543), .B(n4544), .Z(n4535) );
  XNOR U6631 ( .A(n4536), .B(n4535), .Z(n4537) );
  XNOR U6632 ( .A(n4538), .B(n4537), .Z(n4567) );
  XNOR U6633 ( .A(sreg[1028]), .B(n4567), .Z(n4569) );
  NANDN U6634 ( .A(sreg[1027]), .B(n4530), .Z(n4534) );
  NAND U6635 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U6636 ( .A(n4534), .B(n4533), .Z(n4568) );
  XNOR U6637 ( .A(n4569), .B(n4568), .Z(c[1028]) );
  NANDN U6638 ( .A(n4536), .B(n4535), .Z(n4540) );
  NANDN U6639 ( .A(n4538), .B(n4537), .Z(n4539) );
  AND U6640 ( .A(n4540), .B(n4539), .Z(n4575) );
  NANDN U6641 ( .A(n4542), .B(n4541), .Z(n4546) );
  NANDN U6642 ( .A(n4544), .B(n4543), .Z(n4545) );
  AND U6643 ( .A(n4546), .B(n4545), .Z(n4573) );
  NAND U6644 ( .A(n42143), .B(n4547), .Z(n4549) );
  XNOR U6645 ( .A(a[7]), .B(n4072), .Z(n4584) );
  NAND U6646 ( .A(n42144), .B(n4584), .Z(n4548) );
  AND U6647 ( .A(n4549), .B(n4548), .Z(n4599) );
  XOR U6648 ( .A(a[11]), .B(n42012), .Z(n4587) );
  XNOR U6649 ( .A(n4599), .B(n4598), .Z(n4601) );
  AND U6650 ( .A(a[13]), .B(b[0]), .Z(n4551) );
  XNOR U6651 ( .A(n4551), .B(n4071), .Z(n4553) );
  NANDN U6652 ( .A(b[0]), .B(a[12]), .Z(n4552) );
  NAND U6653 ( .A(n4553), .B(n4552), .Z(n4595) );
  XOR U6654 ( .A(a[9]), .B(n42085), .Z(n4588) );
  AND U6655 ( .A(a[5]), .B(b[7]), .Z(n4592) );
  XNOR U6656 ( .A(n4593), .B(n4592), .Z(n4594) );
  XNOR U6657 ( .A(n4595), .B(n4594), .Z(n4600) );
  XOR U6658 ( .A(n4601), .B(n4600), .Z(n4579) );
  NANDN U6659 ( .A(n4556), .B(n4555), .Z(n4560) );
  NANDN U6660 ( .A(n4558), .B(n4557), .Z(n4559) );
  AND U6661 ( .A(n4560), .B(n4559), .Z(n4578) );
  XNOR U6662 ( .A(n4579), .B(n4578), .Z(n4580) );
  NANDN U6663 ( .A(n4562), .B(n4561), .Z(n4566) );
  NAND U6664 ( .A(n4564), .B(n4563), .Z(n4565) );
  NAND U6665 ( .A(n4566), .B(n4565), .Z(n4581) );
  XNOR U6666 ( .A(n4580), .B(n4581), .Z(n4572) );
  XNOR U6667 ( .A(n4573), .B(n4572), .Z(n4574) );
  XNOR U6668 ( .A(n4575), .B(n4574), .Z(n4604) );
  XNOR U6669 ( .A(sreg[1029]), .B(n4604), .Z(n4606) );
  NANDN U6670 ( .A(sreg[1028]), .B(n4567), .Z(n4571) );
  NAND U6671 ( .A(n4569), .B(n4568), .Z(n4570) );
  NAND U6672 ( .A(n4571), .B(n4570), .Z(n4605) );
  XNOR U6673 ( .A(n4606), .B(n4605), .Z(c[1029]) );
  NANDN U6674 ( .A(n4573), .B(n4572), .Z(n4577) );
  NANDN U6675 ( .A(n4575), .B(n4574), .Z(n4576) );
  AND U6676 ( .A(n4577), .B(n4576), .Z(n4612) );
  NANDN U6677 ( .A(n4579), .B(n4578), .Z(n4583) );
  NANDN U6678 ( .A(n4581), .B(n4580), .Z(n4582) );
  AND U6679 ( .A(n4583), .B(n4582), .Z(n4610) );
  NAND U6680 ( .A(n42143), .B(n4584), .Z(n4586) );
  XNOR U6681 ( .A(a[8]), .B(n4073), .Z(n4621) );
  NAND U6682 ( .A(n42144), .B(n4621), .Z(n4585) );
  AND U6683 ( .A(n4586), .B(n4585), .Z(n4636) );
  XOR U6684 ( .A(a[12]), .B(n42012), .Z(n4624) );
  XNOR U6685 ( .A(n4636), .B(n4635), .Z(n4638) );
  XOR U6686 ( .A(a[10]), .B(n42085), .Z(n4628) );
  AND U6687 ( .A(a[6]), .B(b[7]), .Z(n4629) );
  XNOR U6688 ( .A(n4630), .B(n4629), .Z(n4631) );
  AND U6689 ( .A(a[14]), .B(b[0]), .Z(n4589) );
  XNOR U6690 ( .A(n4589), .B(n4071), .Z(n4591) );
  NANDN U6691 ( .A(b[0]), .B(a[13]), .Z(n4590) );
  NAND U6692 ( .A(n4591), .B(n4590), .Z(n4632) );
  XNOR U6693 ( .A(n4631), .B(n4632), .Z(n4637) );
  XOR U6694 ( .A(n4638), .B(n4637), .Z(n4616) );
  NANDN U6695 ( .A(n4593), .B(n4592), .Z(n4597) );
  NANDN U6696 ( .A(n4595), .B(n4594), .Z(n4596) );
  AND U6697 ( .A(n4597), .B(n4596), .Z(n4615) );
  XNOR U6698 ( .A(n4616), .B(n4615), .Z(n4617) );
  NANDN U6699 ( .A(n4599), .B(n4598), .Z(n4603) );
  NAND U6700 ( .A(n4601), .B(n4600), .Z(n4602) );
  NAND U6701 ( .A(n4603), .B(n4602), .Z(n4618) );
  XNOR U6702 ( .A(n4617), .B(n4618), .Z(n4609) );
  XNOR U6703 ( .A(n4610), .B(n4609), .Z(n4611) );
  XNOR U6704 ( .A(n4612), .B(n4611), .Z(n4641) );
  XNOR U6705 ( .A(sreg[1030]), .B(n4641), .Z(n4643) );
  NANDN U6706 ( .A(sreg[1029]), .B(n4604), .Z(n4608) );
  NAND U6707 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U6708 ( .A(n4608), .B(n4607), .Z(n4642) );
  XNOR U6709 ( .A(n4643), .B(n4642), .Z(c[1030]) );
  NANDN U6710 ( .A(n4610), .B(n4609), .Z(n4614) );
  NANDN U6711 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U6712 ( .A(n4614), .B(n4613), .Z(n4649) );
  NANDN U6713 ( .A(n4616), .B(n4615), .Z(n4620) );
  NANDN U6714 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U6715 ( .A(n4620), .B(n4619), .Z(n4647) );
  NAND U6716 ( .A(n42143), .B(n4621), .Z(n4623) );
  XNOR U6717 ( .A(a[9]), .B(n4073), .Z(n4658) );
  NAND U6718 ( .A(n42144), .B(n4658), .Z(n4622) );
  AND U6719 ( .A(n4623), .B(n4622), .Z(n4673) );
  XOR U6720 ( .A(a[13]), .B(n42012), .Z(n4661) );
  XNOR U6721 ( .A(n4673), .B(n4672), .Z(n4675) );
  AND U6722 ( .A(a[15]), .B(b[0]), .Z(n4625) );
  XNOR U6723 ( .A(n4625), .B(n4071), .Z(n4627) );
  NANDN U6724 ( .A(b[0]), .B(a[14]), .Z(n4626) );
  NAND U6725 ( .A(n4627), .B(n4626), .Z(n4669) );
  XOR U6726 ( .A(a[11]), .B(n42085), .Z(n4665) );
  AND U6727 ( .A(a[7]), .B(b[7]), .Z(n4666) );
  XNOR U6728 ( .A(n4667), .B(n4666), .Z(n4668) );
  XNOR U6729 ( .A(n4669), .B(n4668), .Z(n4674) );
  XOR U6730 ( .A(n4675), .B(n4674), .Z(n4653) );
  NANDN U6731 ( .A(n4630), .B(n4629), .Z(n4634) );
  NANDN U6732 ( .A(n4632), .B(n4631), .Z(n4633) );
  AND U6733 ( .A(n4634), .B(n4633), .Z(n4652) );
  XNOR U6734 ( .A(n4653), .B(n4652), .Z(n4654) );
  NANDN U6735 ( .A(n4636), .B(n4635), .Z(n4640) );
  NAND U6736 ( .A(n4638), .B(n4637), .Z(n4639) );
  NAND U6737 ( .A(n4640), .B(n4639), .Z(n4655) );
  XNOR U6738 ( .A(n4654), .B(n4655), .Z(n4646) );
  XNOR U6739 ( .A(n4647), .B(n4646), .Z(n4648) );
  XNOR U6740 ( .A(n4649), .B(n4648), .Z(n4678) );
  XNOR U6741 ( .A(sreg[1031]), .B(n4678), .Z(n4680) );
  NANDN U6742 ( .A(sreg[1030]), .B(n4641), .Z(n4645) );
  NAND U6743 ( .A(n4643), .B(n4642), .Z(n4644) );
  NAND U6744 ( .A(n4645), .B(n4644), .Z(n4679) );
  XNOR U6745 ( .A(n4680), .B(n4679), .Z(c[1031]) );
  NANDN U6746 ( .A(n4647), .B(n4646), .Z(n4651) );
  NANDN U6747 ( .A(n4649), .B(n4648), .Z(n4650) );
  AND U6748 ( .A(n4651), .B(n4650), .Z(n4686) );
  NANDN U6749 ( .A(n4653), .B(n4652), .Z(n4657) );
  NANDN U6750 ( .A(n4655), .B(n4654), .Z(n4656) );
  AND U6751 ( .A(n4657), .B(n4656), .Z(n4684) );
  NAND U6752 ( .A(n42143), .B(n4658), .Z(n4660) );
  XNOR U6753 ( .A(a[10]), .B(n4073), .Z(n4695) );
  NAND U6754 ( .A(n42144), .B(n4695), .Z(n4659) );
  AND U6755 ( .A(n4660), .B(n4659), .Z(n4710) );
  XOR U6756 ( .A(a[14]), .B(n42012), .Z(n4698) );
  XNOR U6757 ( .A(n4710), .B(n4709), .Z(n4712) );
  AND U6758 ( .A(a[16]), .B(b[0]), .Z(n4662) );
  XNOR U6759 ( .A(n4662), .B(n4071), .Z(n4664) );
  NANDN U6760 ( .A(b[0]), .B(a[15]), .Z(n4663) );
  NAND U6761 ( .A(n4664), .B(n4663), .Z(n4706) );
  XOR U6762 ( .A(a[12]), .B(n42085), .Z(n4702) );
  AND U6763 ( .A(a[8]), .B(b[7]), .Z(n4703) );
  XNOR U6764 ( .A(n4704), .B(n4703), .Z(n4705) );
  XNOR U6765 ( .A(n4706), .B(n4705), .Z(n4711) );
  XOR U6766 ( .A(n4712), .B(n4711), .Z(n4690) );
  NANDN U6767 ( .A(n4667), .B(n4666), .Z(n4671) );
  NANDN U6768 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U6769 ( .A(n4671), .B(n4670), .Z(n4689) );
  XNOR U6770 ( .A(n4690), .B(n4689), .Z(n4691) );
  NANDN U6771 ( .A(n4673), .B(n4672), .Z(n4677) );
  NAND U6772 ( .A(n4675), .B(n4674), .Z(n4676) );
  NAND U6773 ( .A(n4677), .B(n4676), .Z(n4692) );
  XNOR U6774 ( .A(n4691), .B(n4692), .Z(n4683) );
  XNOR U6775 ( .A(n4684), .B(n4683), .Z(n4685) );
  XNOR U6776 ( .A(n4686), .B(n4685), .Z(n4715) );
  XNOR U6777 ( .A(sreg[1032]), .B(n4715), .Z(n4717) );
  NANDN U6778 ( .A(sreg[1031]), .B(n4678), .Z(n4682) );
  NAND U6779 ( .A(n4680), .B(n4679), .Z(n4681) );
  NAND U6780 ( .A(n4682), .B(n4681), .Z(n4716) );
  XNOR U6781 ( .A(n4717), .B(n4716), .Z(c[1032]) );
  NANDN U6782 ( .A(n4684), .B(n4683), .Z(n4688) );
  NANDN U6783 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U6784 ( .A(n4688), .B(n4687), .Z(n4723) );
  NANDN U6785 ( .A(n4690), .B(n4689), .Z(n4694) );
  NANDN U6786 ( .A(n4692), .B(n4691), .Z(n4693) );
  AND U6787 ( .A(n4694), .B(n4693), .Z(n4721) );
  NAND U6788 ( .A(n42143), .B(n4695), .Z(n4697) );
  XNOR U6789 ( .A(a[11]), .B(n4073), .Z(n4732) );
  NAND U6790 ( .A(n42144), .B(n4732), .Z(n4696) );
  AND U6791 ( .A(n4697), .B(n4696), .Z(n4747) );
  XOR U6792 ( .A(a[15]), .B(n42012), .Z(n4735) );
  XNOR U6793 ( .A(n4747), .B(n4746), .Z(n4749) );
  AND U6794 ( .A(a[17]), .B(b[0]), .Z(n4699) );
  XNOR U6795 ( .A(n4699), .B(n4071), .Z(n4701) );
  NANDN U6796 ( .A(b[0]), .B(a[16]), .Z(n4700) );
  NAND U6797 ( .A(n4701), .B(n4700), .Z(n4743) );
  XOR U6798 ( .A(a[13]), .B(n42085), .Z(n4736) );
  AND U6799 ( .A(a[9]), .B(b[7]), .Z(n4740) );
  XNOR U6800 ( .A(n4741), .B(n4740), .Z(n4742) );
  XNOR U6801 ( .A(n4743), .B(n4742), .Z(n4748) );
  XOR U6802 ( .A(n4749), .B(n4748), .Z(n4727) );
  NANDN U6803 ( .A(n4704), .B(n4703), .Z(n4708) );
  NANDN U6804 ( .A(n4706), .B(n4705), .Z(n4707) );
  AND U6805 ( .A(n4708), .B(n4707), .Z(n4726) );
  XNOR U6806 ( .A(n4727), .B(n4726), .Z(n4728) );
  NANDN U6807 ( .A(n4710), .B(n4709), .Z(n4714) );
  NAND U6808 ( .A(n4712), .B(n4711), .Z(n4713) );
  NAND U6809 ( .A(n4714), .B(n4713), .Z(n4729) );
  XNOR U6810 ( .A(n4728), .B(n4729), .Z(n4720) );
  XNOR U6811 ( .A(n4721), .B(n4720), .Z(n4722) );
  XNOR U6812 ( .A(n4723), .B(n4722), .Z(n4752) );
  XNOR U6813 ( .A(sreg[1033]), .B(n4752), .Z(n4754) );
  NANDN U6814 ( .A(sreg[1032]), .B(n4715), .Z(n4719) );
  NAND U6815 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U6816 ( .A(n4719), .B(n4718), .Z(n4753) );
  XNOR U6817 ( .A(n4754), .B(n4753), .Z(c[1033]) );
  NANDN U6818 ( .A(n4721), .B(n4720), .Z(n4725) );
  NANDN U6819 ( .A(n4723), .B(n4722), .Z(n4724) );
  AND U6820 ( .A(n4725), .B(n4724), .Z(n4760) );
  NANDN U6821 ( .A(n4727), .B(n4726), .Z(n4731) );
  NANDN U6822 ( .A(n4729), .B(n4728), .Z(n4730) );
  AND U6823 ( .A(n4731), .B(n4730), .Z(n4758) );
  NAND U6824 ( .A(n42143), .B(n4732), .Z(n4734) );
  XNOR U6825 ( .A(a[12]), .B(n4073), .Z(n4769) );
  NAND U6826 ( .A(n42144), .B(n4769), .Z(n4733) );
  AND U6827 ( .A(n4734), .B(n4733), .Z(n4784) );
  XOR U6828 ( .A(a[16]), .B(n42012), .Z(n4772) );
  XNOR U6829 ( .A(n4784), .B(n4783), .Z(n4786) );
  XOR U6830 ( .A(a[14]), .B(n42085), .Z(n4776) );
  AND U6831 ( .A(a[10]), .B(b[7]), .Z(n4777) );
  XNOR U6832 ( .A(n4778), .B(n4777), .Z(n4779) );
  AND U6833 ( .A(a[18]), .B(b[0]), .Z(n4737) );
  XNOR U6834 ( .A(n4737), .B(n4071), .Z(n4739) );
  NANDN U6835 ( .A(b[0]), .B(a[17]), .Z(n4738) );
  NAND U6836 ( .A(n4739), .B(n4738), .Z(n4780) );
  XNOR U6837 ( .A(n4779), .B(n4780), .Z(n4785) );
  XOR U6838 ( .A(n4786), .B(n4785), .Z(n4764) );
  NANDN U6839 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U6840 ( .A(n4743), .B(n4742), .Z(n4744) );
  AND U6841 ( .A(n4745), .B(n4744), .Z(n4763) );
  XNOR U6842 ( .A(n4764), .B(n4763), .Z(n4765) );
  NANDN U6843 ( .A(n4747), .B(n4746), .Z(n4751) );
  NAND U6844 ( .A(n4749), .B(n4748), .Z(n4750) );
  NAND U6845 ( .A(n4751), .B(n4750), .Z(n4766) );
  XNOR U6846 ( .A(n4765), .B(n4766), .Z(n4757) );
  XNOR U6847 ( .A(n4758), .B(n4757), .Z(n4759) );
  XNOR U6848 ( .A(n4760), .B(n4759), .Z(n4789) );
  XNOR U6849 ( .A(sreg[1034]), .B(n4789), .Z(n4791) );
  NANDN U6850 ( .A(sreg[1033]), .B(n4752), .Z(n4756) );
  NAND U6851 ( .A(n4754), .B(n4753), .Z(n4755) );
  NAND U6852 ( .A(n4756), .B(n4755), .Z(n4790) );
  XNOR U6853 ( .A(n4791), .B(n4790), .Z(c[1034]) );
  NANDN U6854 ( .A(n4758), .B(n4757), .Z(n4762) );
  NANDN U6855 ( .A(n4760), .B(n4759), .Z(n4761) );
  AND U6856 ( .A(n4762), .B(n4761), .Z(n4797) );
  NANDN U6857 ( .A(n4764), .B(n4763), .Z(n4768) );
  NANDN U6858 ( .A(n4766), .B(n4765), .Z(n4767) );
  AND U6859 ( .A(n4768), .B(n4767), .Z(n4795) );
  NAND U6860 ( .A(n42143), .B(n4769), .Z(n4771) );
  XNOR U6861 ( .A(a[13]), .B(n4073), .Z(n4806) );
  NAND U6862 ( .A(n42144), .B(n4806), .Z(n4770) );
  AND U6863 ( .A(n4771), .B(n4770), .Z(n4821) );
  XOR U6864 ( .A(a[17]), .B(n42012), .Z(n4809) );
  XNOR U6865 ( .A(n4821), .B(n4820), .Z(n4823) );
  AND U6866 ( .A(a[19]), .B(b[0]), .Z(n4773) );
  XNOR U6867 ( .A(n4773), .B(n4071), .Z(n4775) );
  NANDN U6868 ( .A(b[0]), .B(a[18]), .Z(n4774) );
  NAND U6869 ( .A(n4775), .B(n4774), .Z(n4817) );
  XOR U6870 ( .A(a[15]), .B(n42085), .Z(n4813) );
  AND U6871 ( .A(a[11]), .B(b[7]), .Z(n4814) );
  XNOR U6872 ( .A(n4815), .B(n4814), .Z(n4816) );
  XNOR U6873 ( .A(n4817), .B(n4816), .Z(n4822) );
  XOR U6874 ( .A(n4823), .B(n4822), .Z(n4801) );
  NANDN U6875 ( .A(n4778), .B(n4777), .Z(n4782) );
  NANDN U6876 ( .A(n4780), .B(n4779), .Z(n4781) );
  AND U6877 ( .A(n4782), .B(n4781), .Z(n4800) );
  XNOR U6878 ( .A(n4801), .B(n4800), .Z(n4802) );
  NANDN U6879 ( .A(n4784), .B(n4783), .Z(n4788) );
  NAND U6880 ( .A(n4786), .B(n4785), .Z(n4787) );
  NAND U6881 ( .A(n4788), .B(n4787), .Z(n4803) );
  XNOR U6882 ( .A(n4802), .B(n4803), .Z(n4794) );
  XNOR U6883 ( .A(n4795), .B(n4794), .Z(n4796) );
  XNOR U6884 ( .A(n4797), .B(n4796), .Z(n4826) );
  XNOR U6885 ( .A(sreg[1035]), .B(n4826), .Z(n4828) );
  NANDN U6886 ( .A(sreg[1034]), .B(n4789), .Z(n4793) );
  NAND U6887 ( .A(n4791), .B(n4790), .Z(n4792) );
  NAND U6888 ( .A(n4793), .B(n4792), .Z(n4827) );
  XNOR U6889 ( .A(n4828), .B(n4827), .Z(c[1035]) );
  NANDN U6890 ( .A(n4795), .B(n4794), .Z(n4799) );
  NANDN U6891 ( .A(n4797), .B(n4796), .Z(n4798) );
  AND U6892 ( .A(n4799), .B(n4798), .Z(n4834) );
  NANDN U6893 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U6894 ( .A(n4803), .B(n4802), .Z(n4804) );
  AND U6895 ( .A(n4805), .B(n4804), .Z(n4832) );
  NAND U6896 ( .A(n42143), .B(n4806), .Z(n4808) );
  XNOR U6897 ( .A(a[14]), .B(n4073), .Z(n4843) );
  NAND U6898 ( .A(n42144), .B(n4843), .Z(n4807) );
  AND U6899 ( .A(n4808), .B(n4807), .Z(n4858) );
  XOR U6900 ( .A(a[18]), .B(n42012), .Z(n4846) );
  XNOR U6901 ( .A(n4858), .B(n4857), .Z(n4860) );
  AND U6902 ( .A(a[20]), .B(b[0]), .Z(n4810) );
  XNOR U6903 ( .A(n4810), .B(n4071), .Z(n4812) );
  NANDN U6904 ( .A(b[0]), .B(a[19]), .Z(n4811) );
  NAND U6905 ( .A(n4812), .B(n4811), .Z(n4854) );
  XOR U6906 ( .A(a[16]), .B(n42085), .Z(n4847) );
  AND U6907 ( .A(a[12]), .B(b[7]), .Z(n4851) );
  XNOR U6908 ( .A(n4852), .B(n4851), .Z(n4853) );
  XNOR U6909 ( .A(n4854), .B(n4853), .Z(n4859) );
  XOR U6910 ( .A(n4860), .B(n4859), .Z(n4838) );
  NANDN U6911 ( .A(n4815), .B(n4814), .Z(n4819) );
  NANDN U6912 ( .A(n4817), .B(n4816), .Z(n4818) );
  AND U6913 ( .A(n4819), .B(n4818), .Z(n4837) );
  XNOR U6914 ( .A(n4838), .B(n4837), .Z(n4839) );
  NANDN U6915 ( .A(n4821), .B(n4820), .Z(n4825) );
  NAND U6916 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U6917 ( .A(n4825), .B(n4824), .Z(n4840) );
  XNOR U6918 ( .A(n4839), .B(n4840), .Z(n4831) );
  XNOR U6919 ( .A(n4832), .B(n4831), .Z(n4833) );
  XNOR U6920 ( .A(n4834), .B(n4833), .Z(n4863) );
  XNOR U6921 ( .A(sreg[1036]), .B(n4863), .Z(n4865) );
  NANDN U6922 ( .A(sreg[1035]), .B(n4826), .Z(n4830) );
  NAND U6923 ( .A(n4828), .B(n4827), .Z(n4829) );
  NAND U6924 ( .A(n4830), .B(n4829), .Z(n4864) );
  XNOR U6925 ( .A(n4865), .B(n4864), .Z(c[1036]) );
  NANDN U6926 ( .A(n4832), .B(n4831), .Z(n4836) );
  NANDN U6927 ( .A(n4834), .B(n4833), .Z(n4835) );
  AND U6928 ( .A(n4836), .B(n4835), .Z(n4871) );
  NANDN U6929 ( .A(n4838), .B(n4837), .Z(n4842) );
  NANDN U6930 ( .A(n4840), .B(n4839), .Z(n4841) );
  AND U6931 ( .A(n4842), .B(n4841), .Z(n4869) );
  NAND U6932 ( .A(n42143), .B(n4843), .Z(n4845) );
  XNOR U6933 ( .A(a[15]), .B(n4074), .Z(n4880) );
  NAND U6934 ( .A(n42144), .B(n4880), .Z(n4844) );
  AND U6935 ( .A(n4845), .B(n4844), .Z(n4895) );
  XOR U6936 ( .A(a[19]), .B(n42012), .Z(n4883) );
  XNOR U6937 ( .A(n4895), .B(n4894), .Z(n4897) );
  XOR U6938 ( .A(a[17]), .B(n42085), .Z(n4884) );
  AND U6939 ( .A(a[13]), .B(b[7]), .Z(n4888) );
  XNOR U6940 ( .A(n4889), .B(n4888), .Z(n4890) );
  AND U6941 ( .A(a[21]), .B(b[0]), .Z(n4848) );
  XNOR U6942 ( .A(n4848), .B(n4071), .Z(n4850) );
  NANDN U6943 ( .A(b[0]), .B(a[20]), .Z(n4849) );
  NAND U6944 ( .A(n4850), .B(n4849), .Z(n4891) );
  XNOR U6945 ( .A(n4890), .B(n4891), .Z(n4896) );
  XOR U6946 ( .A(n4897), .B(n4896), .Z(n4875) );
  NANDN U6947 ( .A(n4852), .B(n4851), .Z(n4856) );
  NANDN U6948 ( .A(n4854), .B(n4853), .Z(n4855) );
  AND U6949 ( .A(n4856), .B(n4855), .Z(n4874) );
  XNOR U6950 ( .A(n4875), .B(n4874), .Z(n4876) );
  NANDN U6951 ( .A(n4858), .B(n4857), .Z(n4862) );
  NAND U6952 ( .A(n4860), .B(n4859), .Z(n4861) );
  NAND U6953 ( .A(n4862), .B(n4861), .Z(n4877) );
  XNOR U6954 ( .A(n4876), .B(n4877), .Z(n4868) );
  XNOR U6955 ( .A(n4869), .B(n4868), .Z(n4870) );
  XNOR U6956 ( .A(n4871), .B(n4870), .Z(n4900) );
  XNOR U6957 ( .A(sreg[1037]), .B(n4900), .Z(n4902) );
  NANDN U6958 ( .A(sreg[1036]), .B(n4863), .Z(n4867) );
  NAND U6959 ( .A(n4865), .B(n4864), .Z(n4866) );
  NAND U6960 ( .A(n4867), .B(n4866), .Z(n4901) );
  XNOR U6961 ( .A(n4902), .B(n4901), .Z(c[1037]) );
  NANDN U6962 ( .A(n4869), .B(n4868), .Z(n4873) );
  NANDN U6963 ( .A(n4871), .B(n4870), .Z(n4872) );
  AND U6964 ( .A(n4873), .B(n4872), .Z(n4908) );
  NANDN U6965 ( .A(n4875), .B(n4874), .Z(n4879) );
  NANDN U6966 ( .A(n4877), .B(n4876), .Z(n4878) );
  AND U6967 ( .A(n4879), .B(n4878), .Z(n4906) );
  NAND U6968 ( .A(n42143), .B(n4880), .Z(n4882) );
  XNOR U6969 ( .A(a[16]), .B(n4074), .Z(n4917) );
  NAND U6970 ( .A(n42144), .B(n4917), .Z(n4881) );
  AND U6971 ( .A(n4882), .B(n4881), .Z(n4932) );
  XOR U6972 ( .A(a[20]), .B(n42012), .Z(n4920) );
  XNOR U6973 ( .A(n4932), .B(n4931), .Z(n4934) );
  XOR U6974 ( .A(a[18]), .B(n42085), .Z(n4924) );
  AND U6975 ( .A(a[14]), .B(b[7]), .Z(n4925) );
  XNOR U6976 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U6977 ( .A(a[22]), .B(b[0]), .Z(n4885) );
  XNOR U6978 ( .A(n4885), .B(n4071), .Z(n4887) );
  NANDN U6979 ( .A(b[0]), .B(a[21]), .Z(n4886) );
  NAND U6980 ( .A(n4887), .B(n4886), .Z(n4928) );
  XNOR U6981 ( .A(n4927), .B(n4928), .Z(n4933) );
  XOR U6982 ( .A(n4934), .B(n4933), .Z(n4912) );
  NANDN U6983 ( .A(n4889), .B(n4888), .Z(n4893) );
  NANDN U6984 ( .A(n4891), .B(n4890), .Z(n4892) );
  AND U6985 ( .A(n4893), .B(n4892), .Z(n4911) );
  XNOR U6986 ( .A(n4912), .B(n4911), .Z(n4913) );
  NANDN U6987 ( .A(n4895), .B(n4894), .Z(n4899) );
  NAND U6988 ( .A(n4897), .B(n4896), .Z(n4898) );
  NAND U6989 ( .A(n4899), .B(n4898), .Z(n4914) );
  XNOR U6990 ( .A(n4913), .B(n4914), .Z(n4905) );
  XNOR U6991 ( .A(n4906), .B(n4905), .Z(n4907) );
  XNOR U6992 ( .A(n4908), .B(n4907), .Z(n4937) );
  XNOR U6993 ( .A(sreg[1038]), .B(n4937), .Z(n4939) );
  NANDN U6994 ( .A(sreg[1037]), .B(n4900), .Z(n4904) );
  NAND U6995 ( .A(n4902), .B(n4901), .Z(n4903) );
  NAND U6996 ( .A(n4904), .B(n4903), .Z(n4938) );
  XNOR U6997 ( .A(n4939), .B(n4938), .Z(c[1038]) );
  NANDN U6998 ( .A(n4906), .B(n4905), .Z(n4910) );
  NANDN U6999 ( .A(n4908), .B(n4907), .Z(n4909) );
  AND U7000 ( .A(n4910), .B(n4909), .Z(n4945) );
  NANDN U7001 ( .A(n4912), .B(n4911), .Z(n4916) );
  NANDN U7002 ( .A(n4914), .B(n4913), .Z(n4915) );
  AND U7003 ( .A(n4916), .B(n4915), .Z(n4943) );
  NAND U7004 ( .A(n42143), .B(n4917), .Z(n4919) );
  XNOR U7005 ( .A(a[17]), .B(n4074), .Z(n4954) );
  NAND U7006 ( .A(n42144), .B(n4954), .Z(n4918) );
  AND U7007 ( .A(n4919), .B(n4918), .Z(n4969) );
  XOR U7008 ( .A(a[21]), .B(n42012), .Z(n4957) );
  XNOR U7009 ( .A(n4969), .B(n4968), .Z(n4971) );
  AND U7010 ( .A(a[23]), .B(b[0]), .Z(n4921) );
  XNOR U7011 ( .A(n4921), .B(n4071), .Z(n4923) );
  NANDN U7012 ( .A(b[0]), .B(a[22]), .Z(n4922) );
  NAND U7013 ( .A(n4923), .B(n4922), .Z(n4965) );
  XOR U7014 ( .A(a[19]), .B(n42085), .Z(n4958) );
  AND U7015 ( .A(a[15]), .B(b[7]), .Z(n4962) );
  XNOR U7016 ( .A(n4963), .B(n4962), .Z(n4964) );
  XNOR U7017 ( .A(n4965), .B(n4964), .Z(n4970) );
  XOR U7018 ( .A(n4971), .B(n4970), .Z(n4949) );
  NANDN U7019 ( .A(n4926), .B(n4925), .Z(n4930) );
  NANDN U7020 ( .A(n4928), .B(n4927), .Z(n4929) );
  AND U7021 ( .A(n4930), .B(n4929), .Z(n4948) );
  XNOR U7022 ( .A(n4949), .B(n4948), .Z(n4950) );
  NANDN U7023 ( .A(n4932), .B(n4931), .Z(n4936) );
  NAND U7024 ( .A(n4934), .B(n4933), .Z(n4935) );
  NAND U7025 ( .A(n4936), .B(n4935), .Z(n4951) );
  XNOR U7026 ( .A(n4950), .B(n4951), .Z(n4942) );
  XNOR U7027 ( .A(n4943), .B(n4942), .Z(n4944) );
  XNOR U7028 ( .A(n4945), .B(n4944), .Z(n4974) );
  XNOR U7029 ( .A(sreg[1039]), .B(n4974), .Z(n4976) );
  NANDN U7030 ( .A(sreg[1038]), .B(n4937), .Z(n4941) );
  NAND U7031 ( .A(n4939), .B(n4938), .Z(n4940) );
  NAND U7032 ( .A(n4941), .B(n4940), .Z(n4975) );
  XNOR U7033 ( .A(n4976), .B(n4975), .Z(c[1039]) );
  NANDN U7034 ( .A(n4943), .B(n4942), .Z(n4947) );
  NANDN U7035 ( .A(n4945), .B(n4944), .Z(n4946) );
  AND U7036 ( .A(n4947), .B(n4946), .Z(n4982) );
  NANDN U7037 ( .A(n4949), .B(n4948), .Z(n4953) );
  NANDN U7038 ( .A(n4951), .B(n4950), .Z(n4952) );
  AND U7039 ( .A(n4953), .B(n4952), .Z(n4980) );
  NAND U7040 ( .A(n42143), .B(n4954), .Z(n4956) );
  XNOR U7041 ( .A(a[18]), .B(n4074), .Z(n4991) );
  NAND U7042 ( .A(n42144), .B(n4991), .Z(n4955) );
  AND U7043 ( .A(n4956), .B(n4955), .Z(n5006) );
  XOR U7044 ( .A(a[22]), .B(n42012), .Z(n4994) );
  XNOR U7045 ( .A(n5006), .B(n5005), .Z(n5008) );
  XOR U7046 ( .A(a[20]), .B(n42085), .Z(n4998) );
  AND U7047 ( .A(a[16]), .B(b[7]), .Z(n4999) );
  XNOR U7048 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U7049 ( .A(a[24]), .B(b[0]), .Z(n4959) );
  XNOR U7050 ( .A(n4959), .B(n4071), .Z(n4961) );
  NANDN U7051 ( .A(b[0]), .B(a[23]), .Z(n4960) );
  NAND U7052 ( .A(n4961), .B(n4960), .Z(n5002) );
  XNOR U7053 ( .A(n5001), .B(n5002), .Z(n5007) );
  XOR U7054 ( .A(n5008), .B(n5007), .Z(n4986) );
  NANDN U7055 ( .A(n4963), .B(n4962), .Z(n4967) );
  NANDN U7056 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U7057 ( .A(n4967), .B(n4966), .Z(n4985) );
  XNOR U7058 ( .A(n4986), .B(n4985), .Z(n4987) );
  NANDN U7059 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U7060 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U7061 ( .A(n4973), .B(n4972), .Z(n4988) );
  XNOR U7062 ( .A(n4987), .B(n4988), .Z(n4979) );
  XNOR U7063 ( .A(n4980), .B(n4979), .Z(n4981) );
  XNOR U7064 ( .A(n4982), .B(n4981), .Z(n5011) );
  XNOR U7065 ( .A(sreg[1040]), .B(n5011), .Z(n5013) );
  NANDN U7066 ( .A(sreg[1039]), .B(n4974), .Z(n4978) );
  NAND U7067 ( .A(n4976), .B(n4975), .Z(n4977) );
  NAND U7068 ( .A(n4978), .B(n4977), .Z(n5012) );
  XNOR U7069 ( .A(n5013), .B(n5012), .Z(c[1040]) );
  NANDN U7070 ( .A(n4980), .B(n4979), .Z(n4984) );
  NANDN U7071 ( .A(n4982), .B(n4981), .Z(n4983) );
  AND U7072 ( .A(n4984), .B(n4983), .Z(n5019) );
  NANDN U7073 ( .A(n4986), .B(n4985), .Z(n4990) );
  NANDN U7074 ( .A(n4988), .B(n4987), .Z(n4989) );
  AND U7075 ( .A(n4990), .B(n4989), .Z(n5017) );
  NAND U7076 ( .A(n42143), .B(n4991), .Z(n4993) );
  XNOR U7077 ( .A(a[19]), .B(n4074), .Z(n5028) );
  NAND U7078 ( .A(n42144), .B(n5028), .Z(n4992) );
  AND U7079 ( .A(n4993), .B(n4992), .Z(n5043) );
  XOR U7080 ( .A(a[23]), .B(n42012), .Z(n5031) );
  XNOR U7081 ( .A(n5043), .B(n5042), .Z(n5045) );
  AND U7082 ( .A(a[25]), .B(b[0]), .Z(n4995) );
  XNOR U7083 ( .A(n4995), .B(n4071), .Z(n4997) );
  NANDN U7084 ( .A(b[0]), .B(a[24]), .Z(n4996) );
  NAND U7085 ( .A(n4997), .B(n4996), .Z(n5039) );
  XOR U7086 ( .A(a[21]), .B(n42085), .Z(n5035) );
  AND U7087 ( .A(a[17]), .B(b[7]), .Z(n5036) );
  XNOR U7088 ( .A(n5037), .B(n5036), .Z(n5038) );
  XNOR U7089 ( .A(n5039), .B(n5038), .Z(n5044) );
  XOR U7090 ( .A(n5045), .B(n5044), .Z(n5023) );
  NANDN U7091 ( .A(n5000), .B(n4999), .Z(n5004) );
  NANDN U7092 ( .A(n5002), .B(n5001), .Z(n5003) );
  AND U7093 ( .A(n5004), .B(n5003), .Z(n5022) );
  XNOR U7094 ( .A(n5023), .B(n5022), .Z(n5024) );
  NANDN U7095 ( .A(n5006), .B(n5005), .Z(n5010) );
  NAND U7096 ( .A(n5008), .B(n5007), .Z(n5009) );
  NAND U7097 ( .A(n5010), .B(n5009), .Z(n5025) );
  XNOR U7098 ( .A(n5024), .B(n5025), .Z(n5016) );
  XNOR U7099 ( .A(n5017), .B(n5016), .Z(n5018) );
  XNOR U7100 ( .A(n5019), .B(n5018), .Z(n5048) );
  XNOR U7101 ( .A(sreg[1041]), .B(n5048), .Z(n5050) );
  NANDN U7102 ( .A(sreg[1040]), .B(n5011), .Z(n5015) );
  NAND U7103 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U7104 ( .A(n5015), .B(n5014), .Z(n5049) );
  XNOR U7105 ( .A(n5050), .B(n5049), .Z(c[1041]) );
  NANDN U7106 ( .A(n5017), .B(n5016), .Z(n5021) );
  NANDN U7107 ( .A(n5019), .B(n5018), .Z(n5020) );
  AND U7108 ( .A(n5021), .B(n5020), .Z(n5056) );
  NANDN U7109 ( .A(n5023), .B(n5022), .Z(n5027) );
  NANDN U7110 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U7111 ( .A(n5027), .B(n5026), .Z(n5054) );
  NAND U7112 ( .A(n42143), .B(n5028), .Z(n5030) );
  XNOR U7113 ( .A(a[20]), .B(n4074), .Z(n5065) );
  NAND U7114 ( .A(n42144), .B(n5065), .Z(n5029) );
  AND U7115 ( .A(n5030), .B(n5029), .Z(n5080) );
  XOR U7116 ( .A(a[24]), .B(n42012), .Z(n5068) );
  XNOR U7117 ( .A(n5080), .B(n5079), .Z(n5082) );
  AND U7118 ( .A(a[26]), .B(b[0]), .Z(n5032) );
  XNOR U7119 ( .A(n5032), .B(n4071), .Z(n5034) );
  NANDN U7120 ( .A(b[0]), .B(a[25]), .Z(n5033) );
  NAND U7121 ( .A(n5034), .B(n5033), .Z(n5076) );
  XOR U7122 ( .A(a[22]), .B(n42085), .Z(n5069) );
  AND U7123 ( .A(a[18]), .B(b[7]), .Z(n5073) );
  XNOR U7124 ( .A(n5074), .B(n5073), .Z(n5075) );
  XNOR U7125 ( .A(n5076), .B(n5075), .Z(n5081) );
  XOR U7126 ( .A(n5082), .B(n5081), .Z(n5060) );
  NANDN U7127 ( .A(n5037), .B(n5036), .Z(n5041) );
  NANDN U7128 ( .A(n5039), .B(n5038), .Z(n5040) );
  AND U7129 ( .A(n5041), .B(n5040), .Z(n5059) );
  XNOR U7130 ( .A(n5060), .B(n5059), .Z(n5061) );
  NANDN U7131 ( .A(n5043), .B(n5042), .Z(n5047) );
  NAND U7132 ( .A(n5045), .B(n5044), .Z(n5046) );
  NAND U7133 ( .A(n5047), .B(n5046), .Z(n5062) );
  XNOR U7134 ( .A(n5061), .B(n5062), .Z(n5053) );
  XNOR U7135 ( .A(n5054), .B(n5053), .Z(n5055) );
  XNOR U7136 ( .A(n5056), .B(n5055), .Z(n5085) );
  XNOR U7137 ( .A(sreg[1042]), .B(n5085), .Z(n5087) );
  NANDN U7138 ( .A(sreg[1041]), .B(n5048), .Z(n5052) );
  NAND U7139 ( .A(n5050), .B(n5049), .Z(n5051) );
  NAND U7140 ( .A(n5052), .B(n5051), .Z(n5086) );
  XNOR U7141 ( .A(n5087), .B(n5086), .Z(c[1042]) );
  NANDN U7142 ( .A(n5054), .B(n5053), .Z(n5058) );
  NANDN U7143 ( .A(n5056), .B(n5055), .Z(n5057) );
  AND U7144 ( .A(n5058), .B(n5057), .Z(n5093) );
  NANDN U7145 ( .A(n5060), .B(n5059), .Z(n5064) );
  NANDN U7146 ( .A(n5062), .B(n5061), .Z(n5063) );
  AND U7147 ( .A(n5064), .B(n5063), .Z(n5091) );
  NAND U7148 ( .A(n42143), .B(n5065), .Z(n5067) );
  XNOR U7149 ( .A(a[21]), .B(n4074), .Z(n5102) );
  NAND U7150 ( .A(n42144), .B(n5102), .Z(n5066) );
  AND U7151 ( .A(n5067), .B(n5066), .Z(n5117) );
  XOR U7152 ( .A(a[25]), .B(n42012), .Z(n5105) );
  XNOR U7153 ( .A(n5117), .B(n5116), .Z(n5119) );
  XOR U7154 ( .A(a[23]), .B(n42085), .Z(n5106) );
  AND U7155 ( .A(a[19]), .B(b[7]), .Z(n5110) );
  XNOR U7156 ( .A(n5111), .B(n5110), .Z(n5112) );
  AND U7157 ( .A(a[27]), .B(b[0]), .Z(n5070) );
  XNOR U7158 ( .A(n5070), .B(n4071), .Z(n5072) );
  NANDN U7159 ( .A(b[0]), .B(a[26]), .Z(n5071) );
  NAND U7160 ( .A(n5072), .B(n5071), .Z(n5113) );
  XNOR U7161 ( .A(n5112), .B(n5113), .Z(n5118) );
  XOR U7162 ( .A(n5119), .B(n5118), .Z(n5097) );
  NANDN U7163 ( .A(n5074), .B(n5073), .Z(n5078) );
  NANDN U7164 ( .A(n5076), .B(n5075), .Z(n5077) );
  AND U7165 ( .A(n5078), .B(n5077), .Z(n5096) );
  XNOR U7166 ( .A(n5097), .B(n5096), .Z(n5098) );
  NANDN U7167 ( .A(n5080), .B(n5079), .Z(n5084) );
  NAND U7168 ( .A(n5082), .B(n5081), .Z(n5083) );
  NAND U7169 ( .A(n5084), .B(n5083), .Z(n5099) );
  XNOR U7170 ( .A(n5098), .B(n5099), .Z(n5090) );
  XNOR U7171 ( .A(n5091), .B(n5090), .Z(n5092) );
  XNOR U7172 ( .A(n5093), .B(n5092), .Z(n5122) );
  XNOR U7173 ( .A(sreg[1043]), .B(n5122), .Z(n5124) );
  NANDN U7174 ( .A(sreg[1042]), .B(n5085), .Z(n5089) );
  NAND U7175 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U7176 ( .A(n5089), .B(n5088), .Z(n5123) );
  XNOR U7177 ( .A(n5124), .B(n5123), .Z(c[1043]) );
  NANDN U7178 ( .A(n5091), .B(n5090), .Z(n5095) );
  NANDN U7179 ( .A(n5093), .B(n5092), .Z(n5094) );
  AND U7180 ( .A(n5095), .B(n5094), .Z(n5130) );
  NANDN U7181 ( .A(n5097), .B(n5096), .Z(n5101) );
  NANDN U7182 ( .A(n5099), .B(n5098), .Z(n5100) );
  AND U7183 ( .A(n5101), .B(n5100), .Z(n5128) );
  NAND U7184 ( .A(n42143), .B(n5102), .Z(n5104) );
  XNOR U7185 ( .A(a[22]), .B(n4075), .Z(n5139) );
  NAND U7186 ( .A(n42144), .B(n5139), .Z(n5103) );
  AND U7187 ( .A(n5104), .B(n5103), .Z(n5154) );
  XOR U7188 ( .A(a[26]), .B(n42012), .Z(n5142) );
  XNOR U7189 ( .A(n5154), .B(n5153), .Z(n5156) );
  XOR U7190 ( .A(a[24]), .B(n42085), .Z(n5146) );
  AND U7191 ( .A(a[20]), .B(b[7]), .Z(n5147) );
  XNOR U7192 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U7193 ( .A(a[28]), .B(b[0]), .Z(n5107) );
  XNOR U7194 ( .A(n5107), .B(n4071), .Z(n5109) );
  NANDN U7195 ( .A(b[0]), .B(a[27]), .Z(n5108) );
  NAND U7196 ( .A(n5109), .B(n5108), .Z(n5150) );
  XNOR U7197 ( .A(n5149), .B(n5150), .Z(n5155) );
  XOR U7198 ( .A(n5156), .B(n5155), .Z(n5134) );
  NANDN U7199 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U7200 ( .A(n5113), .B(n5112), .Z(n5114) );
  AND U7201 ( .A(n5115), .B(n5114), .Z(n5133) );
  XNOR U7202 ( .A(n5134), .B(n5133), .Z(n5135) );
  NANDN U7203 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U7204 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U7205 ( .A(n5121), .B(n5120), .Z(n5136) );
  XNOR U7206 ( .A(n5135), .B(n5136), .Z(n5127) );
  XNOR U7207 ( .A(n5128), .B(n5127), .Z(n5129) );
  XNOR U7208 ( .A(n5130), .B(n5129), .Z(n5159) );
  XNOR U7209 ( .A(sreg[1044]), .B(n5159), .Z(n5161) );
  NANDN U7210 ( .A(sreg[1043]), .B(n5122), .Z(n5126) );
  NAND U7211 ( .A(n5124), .B(n5123), .Z(n5125) );
  NAND U7212 ( .A(n5126), .B(n5125), .Z(n5160) );
  XNOR U7213 ( .A(n5161), .B(n5160), .Z(c[1044]) );
  NANDN U7214 ( .A(n5128), .B(n5127), .Z(n5132) );
  NANDN U7215 ( .A(n5130), .B(n5129), .Z(n5131) );
  AND U7216 ( .A(n5132), .B(n5131), .Z(n5167) );
  NANDN U7217 ( .A(n5134), .B(n5133), .Z(n5138) );
  NANDN U7218 ( .A(n5136), .B(n5135), .Z(n5137) );
  AND U7219 ( .A(n5138), .B(n5137), .Z(n5165) );
  NAND U7220 ( .A(n42143), .B(n5139), .Z(n5141) );
  XNOR U7221 ( .A(a[23]), .B(n4075), .Z(n5176) );
  NAND U7222 ( .A(n42144), .B(n5176), .Z(n5140) );
  AND U7223 ( .A(n5141), .B(n5140), .Z(n5191) );
  XOR U7224 ( .A(a[27]), .B(n42012), .Z(n5179) );
  XNOR U7225 ( .A(n5191), .B(n5190), .Z(n5193) );
  AND U7226 ( .A(a[29]), .B(b[0]), .Z(n5143) );
  XNOR U7227 ( .A(n5143), .B(n4071), .Z(n5145) );
  NANDN U7228 ( .A(b[0]), .B(a[28]), .Z(n5144) );
  NAND U7229 ( .A(n5145), .B(n5144), .Z(n5187) );
  XOR U7230 ( .A(a[25]), .B(n42085), .Z(n5183) );
  AND U7231 ( .A(a[21]), .B(b[7]), .Z(n5184) );
  XNOR U7232 ( .A(n5185), .B(n5184), .Z(n5186) );
  XNOR U7233 ( .A(n5187), .B(n5186), .Z(n5192) );
  XOR U7234 ( .A(n5193), .B(n5192), .Z(n5171) );
  NANDN U7235 ( .A(n5148), .B(n5147), .Z(n5152) );
  NANDN U7236 ( .A(n5150), .B(n5149), .Z(n5151) );
  AND U7237 ( .A(n5152), .B(n5151), .Z(n5170) );
  XNOR U7238 ( .A(n5171), .B(n5170), .Z(n5172) );
  NANDN U7239 ( .A(n5154), .B(n5153), .Z(n5158) );
  NAND U7240 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U7241 ( .A(n5158), .B(n5157), .Z(n5173) );
  XNOR U7242 ( .A(n5172), .B(n5173), .Z(n5164) );
  XNOR U7243 ( .A(n5165), .B(n5164), .Z(n5166) );
  XNOR U7244 ( .A(n5167), .B(n5166), .Z(n5196) );
  XNOR U7245 ( .A(sreg[1045]), .B(n5196), .Z(n5198) );
  NANDN U7246 ( .A(sreg[1044]), .B(n5159), .Z(n5163) );
  NAND U7247 ( .A(n5161), .B(n5160), .Z(n5162) );
  NAND U7248 ( .A(n5163), .B(n5162), .Z(n5197) );
  XNOR U7249 ( .A(n5198), .B(n5197), .Z(c[1045]) );
  NANDN U7250 ( .A(n5165), .B(n5164), .Z(n5169) );
  NANDN U7251 ( .A(n5167), .B(n5166), .Z(n5168) );
  AND U7252 ( .A(n5169), .B(n5168), .Z(n5204) );
  NANDN U7253 ( .A(n5171), .B(n5170), .Z(n5175) );
  NANDN U7254 ( .A(n5173), .B(n5172), .Z(n5174) );
  AND U7255 ( .A(n5175), .B(n5174), .Z(n5202) );
  NAND U7256 ( .A(n42143), .B(n5176), .Z(n5178) );
  XNOR U7257 ( .A(a[24]), .B(n4075), .Z(n5213) );
  NAND U7258 ( .A(n42144), .B(n5213), .Z(n5177) );
  AND U7259 ( .A(n5178), .B(n5177), .Z(n5228) );
  XOR U7260 ( .A(a[28]), .B(n42012), .Z(n5216) );
  XNOR U7261 ( .A(n5228), .B(n5227), .Z(n5230) );
  AND U7262 ( .A(a[30]), .B(b[0]), .Z(n5180) );
  XNOR U7263 ( .A(n5180), .B(n4071), .Z(n5182) );
  NANDN U7264 ( .A(b[0]), .B(a[29]), .Z(n5181) );
  NAND U7265 ( .A(n5182), .B(n5181), .Z(n5224) );
  XOR U7266 ( .A(a[26]), .B(n42085), .Z(n5220) );
  AND U7267 ( .A(a[22]), .B(b[7]), .Z(n5221) );
  XNOR U7268 ( .A(n5222), .B(n5221), .Z(n5223) );
  XNOR U7269 ( .A(n5224), .B(n5223), .Z(n5229) );
  XOR U7270 ( .A(n5230), .B(n5229), .Z(n5208) );
  NANDN U7271 ( .A(n5185), .B(n5184), .Z(n5189) );
  NANDN U7272 ( .A(n5187), .B(n5186), .Z(n5188) );
  AND U7273 ( .A(n5189), .B(n5188), .Z(n5207) );
  XNOR U7274 ( .A(n5208), .B(n5207), .Z(n5209) );
  NANDN U7275 ( .A(n5191), .B(n5190), .Z(n5195) );
  NAND U7276 ( .A(n5193), .B(n5192), .Z(n5194) );
  NAND U7277 ( .A(n5195), .B(n5194), .Z(n5210) );
  XNOR U7278 ( .A(n5209), .B(n5210), .Z(n5201) );
  XNOR U7279 ( .A(n5202), .B(n5201), .Z(n5203) );
  XNOR U7280 ( .A(n5204), .B(n5203), .Z(n5233) );
  XNOR U7281 ( .A(sreg[1046]), .B(n5233), .Z(n5235) );
  NANDN U7282 ( .A(sreg[1045]), .B(n5196), .Z(n5200) );
  NAND U7283 ( .A(n5198), .B(n5197), .Z(n5199) );
  NAND U7284 ( .A(n5200), .B(n5199), .Z(n5234) );
  XNOR U7285 ( .A(n5235), .B(n5234), .Z(c[1046]) );
  NANDN U7286 ( .A(n5202), .B(n5201), .Z(n5206) );
  NANDN U7287 ( .A(n5204), .B(n5203), .Z(n5205) );
  AND U7288 ( .A(n5206), .B(n5205), .Z(n5241) );
  NANDN U7289 ( .A(n5208), .B(n5207), .Z(n5212) );
  NANDN U7290 ( .A(n5210), .B(n5209), .Z(n5211) );
  AND U7291 ( .A(n5212), .B(n5211), .Z(n5239) );
  NAND U7292 ( .A(n42143), .B(n5213), .Z(n5215) );
  XNOR U7293 ( .A(a[25]), .B(n4075), .Z(n5250) );
  NAND U7294 ( .A(n42144), .B(n5250), .Z(n5214) );
  AND U7295 ( .A(n5215), .B(n5214), .Z(n5265) );
  XOR U7296 ( .A(a[29]), .B(n42012), .Z(n5253) );
  XNOR U7297 ( .A(n5265), .B(n5264), .Z(n5267) );
  AND U7298 ( .A(a[31]), .B(b[0]), .Z(n5217) );
  XNOR U7299 ( .A(n5217), .B(n4071), .Z(n5219) );
  NANDN U7300 ( .A(b[0]), .B(a[30]), .Z(n5218) );
  NAND U7301 ( .A(n5219), .B(n5218), .Z(n5261) );
  XOR U7302 ( .A(a[27]), .B(n42085), .Z(n5254) );
  AND U7303 ( .A(a[23]), .B(b[7]), .Z(n5258) );
  XNOR U7304 ( .A(n5259), .B(n5258), .Z(n5260) );
  XNOR U7305 ( .A(n5261), .B(n5260), .Z(n5266) );
  XOR U7306 ( .A(n5267), .B(n5266), .Z(n5245) );
  NANDN U7307 ( .A(n5222), .B(n5221), .Z(n5226) );
  NANDN U7308 ( .A(n5224), .B(n5223), .Z(n5225) );
  AND U7309 ( .A(n5226), .B(n5225), .Z(n5244) );
  XNOR U7310 ( .A(n5245), .B(n5244), .Z(n5246) );
  NANDN U7311 ( .A(n5228), .B(n5227), .Z(n5232) );
  NAND U7312 ( .A(n5230), .B(n5229), .Z(n5231) );
  NAND U7313 ( .A(n5232), .B(n5231), .Z(n5247) );
  XNOR U7314 ( .A(n5246), .B(n5247), .Z(n5238) );
  XNOR U7315 ( .A(n5239), .B(n5238), .Z(n5240) );
  XNOR U7316 ( .A(n5241), .B(n5240), .Z(n5270) );
  XNOR U7317 ( .A(sreg[1047]), .B(n5270), .Z(n5272) );
  NANDN U7318 ( .A(sreg[1046]), .B(n5233), .Z(n5237) );
  NAND U7319 ( .A(n5235), .B(n5234), .Z(n5236) );
  NAND U7320 ( .A(n5237), .B(n5236), .Z(n5271) );
  XNOR U7321 ( .A(n5272), .B(n5271), .Z(c[1047]) );
  NANDN U7322 ( .A(n5239), .B(n5238), .Z(n5243) );
  NANDN U7323 ( .A(n5241), .B(n5240), .Z(n5242) );
  AND U7324 ( .A(n5243), .B(n5242), .Z(n5278) );
  NANDN U7325 ( .A(n5245), .B(n5244), .Z(n5249) );
  NANDN U7326 ( .A(n5247), .B(n5246), .Z(n5248) );
  AND U7327 ( .A(n5249), .B(n5248), .Z(n5276) );
  NAND U7328 ( .A(n42143), .B(n5250), .Z(n5252) );
  XNOR U7329 ( .A(a[26]), .B(n4075), .Z(n5287) );
  NAND U7330 ( .A(n42144), .B(n5287), .Z(n5251) );
  AND U7331 ( .A(n5252), .B(n5251), .Z(n5302) );
  XOR U7332 ( .A(a[30]), .B(n42012), .Z(n5290) );
  XNOR U7333 ( .A(n5302), .B(n5301), .Z(n5304) );
  XOR U7334 ( .A(a[28]), .B(n42085), .Z(n5294) );
  AND U7335 ( .A(a[24]), .B(b[7]), .Z(n5295) );
  XNOR U7336 ( .A(n5296), .B(n5295), .Z(n5297) );
  AND U7337 ( .A(a[32]), .B(b[0]), .Z(n5255) );
  XNOR U7338 ( .A(n5255), .B(n4071), .Z(n5257) );
  NANDN U7339 ( .A(b[0]), .B(a[31]), .Z(n5256) );
  NAND U7340 ( .A(n5257), .B(n5256), .Z(n5298) );
  XNOR U7341 ( .A(n5297), .B(n5298), .Z(n5303) );
  XOR U7342 ( .A(n5304), .B(n5303), .Z(n5282) );
  NANDN U7343 ( .A(n5259), .B(n5258), .Z(n5263) );
  NANDN U7344 ( .A(n5261), .B(n5260), .Z(n5262) );
  AND U7345 ( .A(n5263), .B(n5262), .Z(n5281) );
  XNOR U7346 ( .A(n5282), .B(n5281), .Z(n5283) );
  NANDN U7347 ( .A(n5265), .B(n5264), .Z(n5269) );
  NAND U7348 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U7349 ( .A(n5269), .B(n5268), .Z(n5284) );
  XNOR U7350 ( .A(n5283), .B(n5284), .Z(n5275) );
  XNOR U7351 ( .A(n5276), .B(n5275), .Z(n5277) );
  XNOR U7352 ( .A(n5278), .B(n5277), .Z(n5307) );
  XNOR U7353 ( .A(sreg[1048]), .B(n5307), .Z(n5309) );
  NANDN U7354 ( .A(sreg[1047]), .B(n5270), .Z(n5274) );
  NAND U7355 ( .A(n5272), .B(n5271), .Z(n5273) );
  NAND U7356 ( .A(n5274), .B(n5273), .Z(n5308) );
  XNOR U7357 ( .A(n5309), .B(n5308), .Z(c[1048]) );
  NANDN U7358 ( .A(n5276), .B(n5275), .Z(n5280) );
  NANDN U7359 ( .A(n5278), .B(n5277), .Z(n5279) );
  AND U7360 ( .A(n5280), .B(n5279), .Z(n5315) );
  NANDN U7361 ( .A(n5282), .B(n5281), .Z(n5286) );
  NANDN U7362 ( .A(n5284), .B(n5283), .Z(n5285) );
  AND U7363 ( .A(n5286), .B(n5285), .Z(n5313) );
  NAND U7364 ( .A(n42143), .B(n5287), .Z(n5289) );
  XNOR U7365 ( .A(a[27]), .B(n4075), .Z(n5324) );
  NAND U7366 ( .A(n42144), .B(n5324), .Z(n5288) );
  AND U7367 ( .A(n5289), .B(n5288), .Z(n5339) );
  XOR U7368 ( .A(a[31]), .B(n42012), .Z(n5327) );
  XNOR U7369 ( .A(n5339), .B(n5338), .Z(n5341) );
  AND U7370 ( .A(a[33]), .B(b[0]), .Z(n5291) );
  XNOR U7371 ( .A(n5291), .B(n4071), .Z(n5293) );
  NANDN U7372 ( .A(b[0]), .B(a[32]), .Z(n5292) );
  NAND U7373 ( .A(n5293), .B(n5292), .Z(n5335) );
  XOR U7374 ( .A(a[29]), .B(n42085), .Z(n5331) );
  AND U7375 ( .A(a[25]), .B(b[7]), .Z(n5332) );
  XNOR U7376 ( .A(n5333), .B(n5332), .Z(n5334) );
  XNOR U7377 ( .A(n5335), .B(n5334), .Z(n5340) );
  XOR U7378 ( .A(n5341), .B(n5340), .Z(n5319) );
  NANDN U7379 ( .A(n5296), .B(n5295), .Z(n5300) );
  NANDN U7380 ( .A(n5298), .B(n5297), .Z(n5299) );
  AND U7381 ( .A(n5300), .B(n5299), .Z(n5318) );
  XNOR U7382 ( .A(n5319), .B(n5318), .Z(n5320) );
  NANDN U7383 ( .A(n5302), .B(n5301), .Z(n5306) );
  NAND U7384 ( .A(n5304), .B(n5303), .Z(n5305) );
  NAND U7385 ( .A(n5306), .B(n5305), .Z(n5321) );
  XNOR U7386 ( .A(n5320), .B(n5321), .Z(n5312) );
  XNOR U7387 ( .A(n5313), .B(n5312), .Z(n5314) );
  XNOR U7388 ( .A(n5315), .B(n5314), .Z(n5344) );
  XNOR U7389 ( .A(sreg[1049]), .B(n5344), .Z(n5346) );
  NANDN U7390 ( .A(sreg[1048]), .B(n5307), .Z(n5311) );
  NAND U7391 ( .A(n5309), .B(n5308), .Z(n5310) );
  NAND U7392 ( .A(n5311), .B(n5310), .Z(n5345) );
  XNOR U7393 ( .A(n5346), .B(n5345), .Z(c[1049]) );
  NANDN U7394 ( .A(n5313), .B(n5312), .Z(n5317) );
  NANDN U7395 ( .A(n5315), .B(n5314), .Z(n5316) );
  AND U7396 ( .A(n5317), .B(n5316), .Z(n5352) );
  NANDN U7397 ( .A(n5319), .B(n5318), .Z(n5323) );
  NANDN U7398 ( .A(n5321), .B(n5320), .Z(n5322) );
  AND U7399 ( .A(n5323), .B(n5322), .Z(n5350) );
  NAND U7400 ( .A(n42143), .B(n5324), .Z(n5326) );
  XNOR U7401 ( .A(a[28]), .B(n4075), .Z(n5361) );
  NAND U7402 ( .A(n42144), .B(n5361), .Z(n5325) );
  AND U7403 ( .A(n5326), .B(n5325), .Z(n5376) );
  XOR U7404 ( .A(a[32]), .B(n42012), .Z(n5364) );
  XNOR U7405 ( .A(n5376), .B(n5375), .Z(n5378) );
  AND U7406 ( .A(a[34]), .B(b[0]), .Z(n5328) );
  XNOR U7407 ( .A(n5328), .B(n4071), .Z(n5330) );
  NANDN U7408 ( .A(b[0]), .B(a[33]), .Z(n5329) );
  NAND U7409 ( .A(n5330), .B(n5329), .Z(n5372) );
  XOR U7410 ( .A(a[30]), .B(n42085), .Z(n5365) );
  AND U7411 ( .A(a[26]), .B(b[7]), .Z(n5369) );
  XNOR U7412 ( .A(n5370), .B(n5369), .Z(n5371) );
  XNOR U7413 ( .A(n5372), .B(n5371), .Z(n5377) );
  XOR U7414 ( .A(n5378), .B(n5377), .Z(n5356) );
  NANDN U7415 ( .A(n5333), .B(n5332), .Z(n5337) );
  NANDN U7416 ( .A(n5335), .B(n5334), .Z(n5336) );
  AND U7417 ( .A(n5337), .B(n5336), .Z(n5355) );
  XNOR U7418 ( .A(n5356), .B(n5355), .Z(n5357) );
  NANDN U7419 ( .A(n5339), .B(n5338), .Z(n5343) );
  NAND U7420 ( .A(n5341), .B(n5340), .Z(n5342) );
  NAND U7421 ( .A(n5343), .B(n5342), .Z(n5358) );
  XNOR U7422 ( .A(n5357), .B(n5358), .Z(n5349) );
  XNOR U7423 ( .A(n5350), .B(n5349), .Z(n5351) );
  XNOR U7424 ( .A(n5352), .B(n5351), .Z(n5381) );
  XNOR U7425 ( .A(sreg[1050]), .B(n5381), .Z(n5383) );
  NANDN U7426 ( .A(sreg[1049]), .B(n5344), .Z(n5348) );
  NAND U7427 ( .A(n5346), .B(n5345), .Z(n5347) );
  NAND U7428 ( .A(n5348), .B(n5347), .Z(n5382) );
  XNOR U7429 ( .A(n5383), .B(n5382), .Z(c[1050]) );
  NANDN U7430 ( .A(n5350), .B(n5349), .Z(n5354) );
  NANDN U7431 ( .A(n5352), .B(n5351), .Z(n5353) );
  AND U7432 ( .A(n5354), .B(n5353), .Z(n5389) );
  NANDN U7433 ( .A(n5356), .B(n5355), .Z(n5360) );
  NANDN U7434 ( .A(n5358), .B(n5357), .Z(n5359) );
  AND U7435 ( .A(n5360), .B(n5359), .Z(n5387) );
  NAND U7436 ( .A(n42143), .B(n5361), .Z(n5363) );
  XNOR U7437 ( .A(a[29]), .B(n4076), .Z(n5398) );
  NAND U7438 ( .A(n42144), .B(n5398), .Z(n5362) );
  AND U7439 ( .A(n5363), .B(n5362), .Z(n5413) );
  XOR U7440 ( .A(a[33]), .B(n42012), .Z(n5401) );
  XNOR U7441 ( .A(n5413), .B(n5412), .Z(n5415) );
  XOR U7442 ( .A(a[31]), .B(n42085), .Z(n5405) );
  AND U7443 ( .A(a[27]), .B(b[7]), .Z(n5406) );
  XNOR U7444 ( .A(n5407), .B(n5406), .Z(n5408) );
  AND U7445 ( .A(a[35]), .B(b[0]), .Z(n5366) );
  XNOR U7446 ( .A(n5366), .B(n4071), .Z(n5368) );
  NANDN U7447 ( .A(b[0]), .B(a[34]), .Z(n5367) );
  NAND U7448 ( .A(n5368), .B(n5367), .Z(n5409) );
  XNOR U7449 ( .A(n5408), .B(n5409), .Z(n5414) );
  XOR U7450 ( .A(n5415), .B(n5414), .Z(n5393) );
  NANDN U7451 ( .A(n5370), .B(n5369), .Z(n5374) );
  NANDN U7452 ( .A(n5372), .B(n5371), .Z(n5373) );
  AND U7453 ( .A(n5374), .B(n5373), .Z(n5392) );
  XNOR U7454 ( .A(n5393), .B(n5392), .Z(n5394) );
  NANDN U7455 ( .A(n5376), .B(n5375), .Z(n5380) );
  NAND U7456 ( .A(n5378), .B(n5377), .Z(n5379) );
  NAND U7457 ( .A(n5380), .B(n5379), .Z(n5395) );
  XNOR U7458 ( .A(n5394), .B(n5395), .Z(n5386) );
  XNOR U7459 ( .A(n5387), .B(n5386), .Z(n5388) );
  XNOR U7460 ( .A(n5389), .B(n5388), .Z(n5418) );
  XNOR U7461 ( .A(sreg[1051]), .B(n5418), .Z(n5420) );
  NANDN U7462 ( .A(sreg[1050]), .B(n5381), .Z(n5385) );
  NAND U7463 ( .A(n5383), .B(n5382), .Z(n5384) );
  NAND U7464 ( .A(n5385), .B(n5384), .Z(n5419) );
  XNOR U7465 ( .A(n5420), .B(n5419), .Z(c[1051]) );
  NANDN U7466 ( .A(n5387), .B(n5386), .Z(n5391) );
  NANDN U7467 ( .A(n5389), .B(n5388), .Z(n5390) );
  AND U7468 ( .A(n5391), .B(n5390), .Z(n5426) );
  NANDN U7469 ( .A(n5393), .B(n5392), .Z(n5397) );
  NANDN U7470 ( .A(n5395), .B(n5394), .Z(n5396) );
  AND U7471 ( .A(n5397), .B(n5396), .Z(n5424) );
  NAND U7472 ( .A(n42143), .B(n5398), .Z(n5400) );
  XNOR U7473 ( .A(a[30]), .B(n4076), .Z(n5435) );
  NAND U7474 ( .A(n42144), .B(n5435), .Z(n5399) );
  AND U7475 ( .A(n5400), .B(n5399), .Z(n5450) );
  XOR U7476 ( .A(a[34]), .B(n42012), .Z(n5438) );
  XNOR U7477 ( .A(n5450), .B(n5449), .Z(n5452) );
  AND U7478 ( .A(a[36]), .B(b[0]), .Z(n5402) );
  XNOR U7479 ( .A(n5402), .B(n4071), .Z(n5404) );
  NANDN U7480 ( .A(b[0]), .B(a[35]), .Z(n5403) );
  NAND U7481 ( .A(n5404), .B(n5403), .Z(n5446) );
  XOR U7482 ( .A(a[32]), .B(n42085), .Z(n5442) );
  AND U7483 ( .A(a[28]), .B(b[7]), .Z(n5443) );
  XNOR U7484 ( .A(n5444), .B(n5443), .Z(n5445) );
  XNOR U7485 ( .A(n5446), .B(n5445), .Z(n5451) );
  XOR U7486 ( .A(n5452), .B(n5451), .Z(n5430) );
  NANDN U7487 ( .A(n5407), .B(n5406), .Z(n5411) );
  NANDN U7488 ( .A(n5409), .B(n5408), .Z(n5410) );
  AND U7489 ( .A(n5411), .B(n5410), .Z(n5429) );
  XNOR U7490 ( .A(n5430), .B(n5429), .Z(n5431) );
  NANDN U7491 ( .A(n5413), .B(n5412), .Z(n5417) );
  NAND U7492 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U7493 ( .A(n5417), .B(n5416), .Z(n5432) );
  XNOR U7494 ( .A(n5431), .B(n5432), .Z(n5423) );
  XNOR U7495 ( .A(n5424), .B(n5423), .Z(n5425) );
  XNOR U7496 ( .A(n5426), .B(n5425), .Z(n5455) );
  XNOR U7497 ( .A(sreg[1052]), .B(n5455), .Z(n5457) );
  NANDN U7498 ( .A(sreg[1051]), .B(n5418), .Z(n5422) );
  NAND U7499 ( .A(n5420), .B(n5419), .Z(n5421) );
  NAND U7500 ( .A(n5422), .B(n5421), .Z(n5456) );
  XNOR U7501 ( .A(n5457), .B(n5456), .Z(c[1052]) );
  NANDN U7502 ( .A(n5424), .B(n5423), .Z(n5428) );
  NANDN U7503 ( .A(n5426), .B(n5425), .Z(n5427) );
  AND U7504 ( .A(n5428), .B(n5427), .Z(n5463) );
  NANDN U7505 ( .A(n5430), .B(n5429), .Z(n5434) );
  NANDN U7506 ( .A(n5432), .B(n5431), .Z(n5433) );
  AND U7507 ( .A(n5434), .B(n5433), .Z(n5461) );
  NAND U7508 ( .A(n42143), .B(n5435), .Z(n5437) );
  XNOR U7509 ( .A(a[31]), .B(n4076), .Z(n5472) );
  NAND U7510 ( .A(n42144), .B(n5472), .Z(n5436) );
  AND U7511 ( .A(n5437), .B(n5436), .Z(n5487) );
  XOR U7512 ( .A(a[35]), .B(n42012), .Z(n5475) );
  XNOR U7513 ( .A(n5487), .B(n5486), .Z(n5489) );
  AND U7514 ( .A(a[37]), .B(b[0]), .Z(n5439) );
  XNOR U7515 ( .A(n5439), .B(n4071), .Z(n5441) );
  NANDN U7516 ( .A(b[0]), .B(a[36]), .Z(n5440) );
  NAND U7517 ( .A(n5441), .B(n5440), .Z(n5483) );
  XOR U7518 ( .A(a[33]), .B(n42085), .Z(n5476) );
  AND U7519 ( .A(a[29]), .B(b[7]), .Z(n5480) );
  XNOR U7520 ( .A(n5481), .B(n5480), .Z(n5482) );
  XNOR U7521 ( .A(n5483), .B(n5482), .Z(n5488) );
  XOR U7522 ( .A(n5489), .B(n5488), .Z(n5467) );
  NANDN U7523 ( .A(n5444), .B(n5443), .Z(n5448) );
  NANDN U7524 ( .A(n5446), .B(n5445), .Z(n5447) );
  AND U7525 ( .A(n5448), .B(n5447), .Z(n5466) );
  XNOR U7526 ( .A(n5467), .B(n5466), .Z(n5468) );
  NANDN U7527 ( .A(n5450), .B(n5449), .Z(n5454) );
  NAND U7528 ( .A(n5452), .B(n5451), .Z(n5453) );
  NAND U7529 ( .A(n5454), .B(n5453), .Z(n5469) );
  XNOR U7530 ( .A(n5468), .B(n5469), .Z(n5460) );
  XNOR U7531 ( .A(n5461), .B(n5460), .Z(n5462) );
  XNOR U7532 ( .A(n5463), .B(n5462), .Z(n5492) );
  XNOR U7533 ( .A(sreg[1053]), .B(n5492), .Z(n5494) );
  NANDN U7534 ( .A(sreg[1052]), .B(n5455), .Z(n5459) );
  NAND U7535 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U7536 ( .A(n5459), .B(n5458), .Z(n5493) );
  XNOR U7537 ( .A(n5494), .B(n5493), .Z(c[1053]) );
  NANDN U7538 ( .A(n5461), .B(n5460), .Z(n5465) );
  NANDN U7539 ( .A(n5463), .B(n5462), .Z(n5464) );
  AND U7540 ( .A(n5465), .B(n5464), .Z(n5500) );
  NANDN U7541 ( .A(n5467), .B(n5466), .Z(n5471) );
  NANDN U7542 ( .A(n5469), .B(n5468), .Z(n5470) );
  AND U7543 ( .A(n5471), .B(n5470), .Z(n5498) );
  NAND U7544 ( .A(n42143), .B(n5472), .Z(n5474) );
  XNOR U7545 ( .A(a[32]), .B(n4076), .Z(n5509) );
  NAND U7546 ( .A(n42144), .B(n5509), .Z(n5473) );
  AND U7547 ( .A(n5474), .B(n5473), .Z(n5524) );
  XOR U7548 ( .A(a[36]), .B(n42012), .Z(n5512) );
  XNOR U7549 ( .A(n5524), .B(n5523), .Z(n5526) );
  XOR U7550 ( .A(a[34]), .B(n42085), .Z(n5516) );
  AND U7551 ( .A(a[30]), .B(b[7]), .Z(n5517) );
  XNOR U7552 ( .A(n5518), .B(n5517), .Z(n5519) );
  AND U7553 ( .A(a[38]), .B(b[0]), .Z(n5477) );
  XNOR U7554 ( .A(n5477), .B(n4071), .Z(n5479) );
  NANDN U7555 ( .A(b[0]), .B(a[37]), .Z(n5478) );
  NAND U7556 ( .A(n5479), .B(n5478), .Z(n5520) );
  XNOR U7557 ( .A(n5519), .B(n5520), .Z(n5525) );
  XOR U7558 ( .A(n5526), .B(n5525), .Z(n5504) );
  NANDN U7559 ( .A(n5481), .B(n5480), .Z(n5485) );
  NANDN U7560 ( .A(n5483), .B(n5482), .Z(n5484) );
  AND U7561 ( .A(n5485), .B(n5484), .Z(n5503) );
  XNOR U7562 ( .A(n5504), .B(n5503), .Z(n5505) );
  NANDN U7563 ( .A(n5487), .B(n5486), .Z(n5491) );
  NAND U7564 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U7565 ( .A(n5491), .B(n5490), .Z(n5506) );
  XNOR U7566 ( .A(n5505), .B(n5506), .Z(n5497) );
  XNOR U7567 ( .A(n5498), .B(n5497), .Z(n5499) );
  XNOR U7568 ( .A(n5500), .B(n5499), .Z(n5529) );
  XNOR U7569 ( .A(sreg[1054]), .B(n5529), .Z(n5531) );
  NANDN U7570 ( .A(sreg[1053]), .B(n5492), .Z(n5496) );
  NAND U7571 ( .A(n5494), .B(n5493), .Z(n5495) );
  NAND U7572 ( .A(n5496), .B(n5495), .Z(n5530) );
  XNOR U7573 ( .A(n5531), .B(n5530), .Z(c[1054]) );
  NANDN U7574 ( .A(n5498), .B(n5497), .Z(n5502) );
  NANDN U7575 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U7576 ( .A(n5502), .B(n5501), .Z(n5537) );
  NANDN U7577 ( .A(n5504), .B(n5503), .Z(n5508) );
  NANDN U7578 ( .A(n5506), .B(n5505), .Z(n5507) );
  AND U7579 ( .A(n5508), .B(n5507), .Z(n5535) );
  NAND U7580 ( .A(n42143), .B(n5509), .Z(n5511) );
  XNOR U7581 ( .A(a[33]), .B(n4076), .Z(n5546) );
  NAND U7582 ( .A(n42144), .B(n5546), .Z(n5510) );
  AND U7583 ( .A(n5511), .B(n5510), .Z(n5561) );
  XOR U7584 ( .A(a[37]), .B(n42012), .Z(n5549) );
  XNOR U7585 ( .A(n5561), .B(n5560), .Z(n5563) );
  AND U7586 ( .A(a[39]), .B(b[0]), .Z(n5513) );
  XNOR U7587 ( .A(n5513), .B(n4071), .Z(n5515) );
  NANDN U7588 ( .A(b[0]), .B(a[38]), .Z(n5514) );
  NAND U7589 ( .A(n5515), .B(n5514), .Z(n5557) );
  XOR U7590 ( .A(a[35]), .B(n42085), .Z(n5553) );
  AND U7591 ( .A(a[31]), .B(b[7]), .Z(n5554) );
  XNOR U7592 ( .A(n5555), .B(n5554), .Z(n5556) );
  XNOR U7593 ( .A(n5557), .B(n5556), .Z(n5562) );
  XOR U7594 ( .A(n5563), .B(n5562), .Z(n5541) );
  NANDN U7595 ( .A(n5518), .B(n5517), .Z(n5522) );
  NANDN U7596 ( .A(n5520), .B(n5519), .Z(n5521) );
  AND U7597 ( .A(n5522), .B(n5521), .Z(n5540) );
  XNOR U7598 ( .A(n5541), .B(n5540), .Z(n5542) );
  NANDN U7599 ( .A(n5524), .B(n5523), .Z(n5528) );
  NAND U7600 ( .A(n5526), .B(n5525), .Z(n5527) );
  NAND U7601 ( .A(n5528), .B(n5527), .Z(n5543) );
  XNOR U7602 ( .A(n5542), .B(n5543), .Z(n5534) );
  XNOR U7603 ( .A(n5535), .B(n5534), .Z(n5536) );
  XNOR U7604 ( .A(n5537), .B(n5536), .Z(n5566) );
  XNOR U7605 ( .A(sreg[1055]), .B(n5566), .Z(n5568) );
  NANDN U7606 ( .A(sreg[1054]), .B(n5529), .Z(n5533) );
  NAND U7607 ( .A(n5531), .B(n5530), .Z(n5532) );
  NAND U7608 ( .A(n5533), .B(n5532), .Z(n5567) );
  XNOR U7609 ( .A(n5568), .B(n5567), .Z(c[1055]) );
  NANDN U7610 ( .A(n5535), .B(n5534), .Z(n5539) );
  NANDN U7611 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U7612 ( .A(n5539), .B(n5538), .Z(n5574) );
  NANDN U7613 ( .A(n5541), .B(n5540), .Z(n5545) );
  NANDN U7614 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U7615 ( .A(n5545), .B(n5544), .Z(n5572) );
  NAND U7616 ( .A(n42143), .B(n5546), .Z(n5548) );
  XNOR U7617 ( .A(a[34]), .B(n4076), .Z(n5583) );
  NAND U7618 ( .A(n42144), .B(n5583), .Z(n5547) );
  AND U7619 ( .A(n5548), .B(n5547), .Z(n5598) );
  XOR U7620 ( .A(a[38]), .B(n42012), .Z(n5586) );
  XNOR U7621 ( .A(n5598), .B(n5597), .Z(n5600) );
  AND U7622 ( .A(a[40]), .B(b[0]), .Z(n5550) );
  XNOR U7623 ( .A(n5550), .B(n4071), .Z(n5552) );
  NANDN U7624 ( .A(b[0]), .B(a[39]), .Z(n5551) );
  NAND U7625 ( .A(n5552), .B(n5551), .Z(n5594) );
  XOR U7626 ( .A(a[36]), .B(n42085), .Z(n5590) );
  AND U7627 ( .A(a[32]), .B(b[7]), .Z(n5591) );
  XNOR U7628 ( .A(n5592), .B(n5591), .Z(n5593) );
  XNOR U7629 ( .A(n5594), .B(n5593), .Z(n5599) );
  XOR U7630 ( .A(n5600), .B(n5599), .Z(n5578) );
  NANDN U7631 ( .A(n5555), .B(n5554), .Z(n5559) );
  NANDN U7632 ( .A(n5557), .B(n5556), .Z(n5558) );
  AND U7633 ( .A(n5559), .B(n5558), .Z(n5577) );
  XNOR U7634 ( .A(n5578), .B(n5577), .Z(n5579) );
  NANDN U7635 ( .A(n5561), .B(n5560), .Z(n5565) );
  NAND U7636 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U7637 ( .A(n5565), .B(n5564), .Z(n5580) );
  XNOR U7638 ( .A(n5579), .B(n5580), .Z(n5571) );
  XNOR U7639 ( .A(n5572), .B(n5571), .Z(n5573) );
  XNOR U7640 ( .A(n5574), .B(n5573), .Z(n5603) );
  XNOR U7641 ( .A(sreg[1056]), .B(n5603), .Z(n5605) );
  NANDN U7642 ( .A(sreg[1055]), .B(n5566), .Z(n5570) );
  NAND U7643 ( .A(n5568), .B(n5567), .Z(n5569) );
  NAND U7644 ( .A(n5570), .B(n5569), .Z(n5604) );
  XNOR U7645 ( .A(n5605), .B(n5604), .Z(c[1056]) );
  NANDN U7646 ( .A(n5572), .B(n5571), .Z(n5576) );
  NANDN U7647 ( .A(n5574), .B(n5573), .Z(n5575) );
  AND U7648 ( .A(n5576), .B(n5575), .Z(n5611) );
  NANDN U7649 ( .A(n5578), .B(n5577), .Z(n5582) );
  NANDN U7650 ( .A(n5580), .B(n5579), .Z(n5581) );
  AND U7651 ( .A(n5582), .B(n5581), .Z(n5609) );
  NAND U7652 ( .A(n42143), .B(n5583), .Z(n5585) );
  XNOR U7653 ( .A(a[35]), .B(n4076), .Z(n5620) );
  NAND U7654 ( .A(n42144), .B(n5620), .Z(n5584) );
  AND U7655 ( .A(n5585), .B(n5584), .Z(n5635) );
  XOR U7656 ( .A(a[39]), .B(n42012), .Z(n5623) );
  XNOR U7657 ( .A(n5635), .B(n5634), .Z(n5637) );
  AND U7658 ( .A(a[41]), .B(b[0]), .Z(n5587) );
  XNOR U7659 ( .A(n5587), .B(n4071), .Z(n5589) );
  NANDN U7660 ( .A(b[0]), .B(a[40]), .Z(n5588) );
  NAND U7661 ( .A(n5589), .B(n5588), .Z(n5631) );
  XOR U7662 ( .A(a[37]), .B(n42085), .Z(n5627) );
  AND U7663 ( .A(a[33]), .B(b[7]), .Z(n5628) );
  XNOR U7664 ( .A(n5629), .B(n5628), .Z(n5630) );
  XNOR U7665 ( .A(n5631), .B(n5630), .Z(n5636) );
  XOR U7666 ( .A(n5637), .B(n5636), .Z(n5615) );
  NANDN U7667 ( .A(n5592), .B(n5591), .Z(n5596) );
  NANDN U7668 ( .A(n5594), .B(n5593), .Z(n5595) );
  AND U7669 ( .A(n5596), .B(n5595), .Z(n5614) );
  XNOR U7670 ( .A(n5615), .B(n5614), .Z(n5616) );
  NANDN U7671 ( .A(n5598), .B(n5597), .Z(n5602) );
  NAND U7672 ( .A(n5600), .B(n5599), .Z(n5601) );
  NAND U7673 ( .A(n5602), .B(n5601), .Z(n5617) );
  XNOR U7674 ( .A(n5616), .B(n5617), .Z(n5608) );
  XNOR U7675 ( .A(n5609), .B(n5608), .Z(n5610) );
  XNOR U7676 ( .A(n5611), .B(n5610), .Z(n5640) );
  XNOR U7677 ( .A(sreg[1057]), .B(n5640), .Z(n5642) );
  NANDN U7678 ( .A(sreg[1056]), .B(n5603), .Z(n5607) );
  NAND U7679 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U7680 ( .A(n5607), .B(n5606), .Z(n5641) );
  XNOR U7681 ( .A(n5642), .B(n5641), .Z(c[1057]) );
  NANDN U7682 ( .A(n5609), .B(n5608), .Z(n5613) );
  NANDN U7683 ( .A(n5611), .B(n5610), .Z(n5612) );
  AND U7684 ( .A(n5613), .B(n5612), .Z(n5648) );
  NANDN U7685 ( .A(n5615), .B(n5614), .Z(n5619) );
  NANDN U7686 ( .A(n5617), .B(n5616), .Z(n5618) );
  AND U7687 ( .A(n5619), .B(n5618), .Z(n5646) );
  NAND U7688 ( .A(n42143), .B(n5620), .Z(n5622) );
  XNOR U7689 ( .A(a[36]), .B(n4077), .Z(n5657) );
  NAND U7690 ( .A(n42144), .B(n5657), .Z(n5621) );
  AND U7691 ( .A(n5622), .B(n5621), .Z(n5672) );
  XOR U7692 ( .A(a[40]), .B(n42012), .Z(n5660) );
  XNOR U7693 ( .A(n5672), .B(n5671), .Z(n5674) );
  AND U7694 ( .A(a[42]), .B(b[0]), .Z(n5624) );
  XNOR U7695 ( .A(n5624), .B(n4071), .Z(n5626) );
  NANDN U7696 ( .A(b[0]), .B(a[41]), .Z(n5625) );
  NAND U7697 ( .A(n5626), .B(n5625), .Z(n5668) );
  XOR U7698 ( .A(a[38]), .B(n42085), .Z(n5661) );
  AND U7699 ( .A(a[34]), .B(b[7]), .Z(n5665) );
  XNOR U7700 ( .A(n5666), .B(n5665), .Z(n5667) );
  XNOR U7701 ( .A(n5668), .B(n5667), .Z(n5673) );
  XOR U7702 ( .A(n5674), .B(n5673), .Z(n5652) );
  NANDN U7703 ( .A(n5629), .B(n5628), .Z(n5633) );
  NANDN U7704 ( .A(n5631), .B(n5630), .Z(n5632) );
  AND U7705 ( .A(n5633), .B(n5632), .Z(n5651) );
  XNOR U7706 ( .A(n5652), .B(n5651), .Z(n5653) );
  NANDN U7707 ( .A(n5635), .B(n5634), .Z(n5639) );
  NAND U7708 ( .A(n5637), .B(n5636), .Z(n5638) );
  NAND U7709 ( .A(n5639), .B(n5638), .Z(n5654) );
  XNOR U7710 ( .A(n5653), .B(n5654), .Z(n5645) );
  XNOR U7711 ( .A(n5646), .B(n5645), .Z(n5647) );
  XNOR U7712 ( .A(n5648), .B(n5647), .Z(n5677) );
  XNOR U7713 ( .A(sreg[1058]), .B(n5677), .Z(n5679) );
  NANDN U7714 ( .A(sreg[1057]), .B(n5640), .Z(n5644) );
  NAND U7715 ( .A(n5642), .B(n5641), .Z(n5643) );
  NAND U7716 ( .A(n5644), .B(n5643), .Z(n5678) );
  XNOR U7717 ( .A(n5679), .B(n5678), .Z(c[1058]) );
  NANDN U7718 ( .A(n5646), .B(n5645), .Z(n5650) );
  NANDN U7719 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U7720 ( .A(n5650), .B(n5649), .Z(n5685) );
  NANDN U7721 ( .A(n5652), .B(n5651), .Z(n5656) );
  NANDN U7722 ( .A(n5654), .B(n5653), .Z(n5655) );
  AND U7723 ( .A(n5656), .B(n5655), .Z(n5683) );
  NAND U7724 ( .A(n42143), .B(n5657), .Z(n5659) );
  XNOR U7725 ( .A(a[37]), .B(n4077), .Z(n5694) );
  NAND U7726 ( .A(n42144), .B(n5694), .Z(n5658) );
  AND U7727 ( .A(n5659), .B(n5658), .Z(n5709) );
  XOR U7728 ( .A(a[41]), .B(n42012), .Z(n5697) );
  XNOR U7729 ( .A(n5709), .B(n5708), .Z(n5711) );
  XOR U7730 ( .A(a[39]), .B(n42085), .Z(n5701) );
  AND U7731 ( .A(a[35]), .B(b[7]), .Z(n5702) );
  XNOR U7732 ( .A(n5703), .B(n5702), .Z(n5704) );
  AND U7733 ( .A(a[43]), .B(b[0]), .Z(n5662) );
  XNOR U7734 ( .A(n5662), .B(n4071), .Z(n5664) );
  NANDN U7735 ( .A(b[0]), .B(a[42]), .Z(n5663) );
  NAND U7736 ( .A(n5664), .B(n5663), .Z(n5705) );
  XNOR U7737 ( .A(n5704), .B(n5705), .Z(n5710) );
  XOR U7738 ( .A(n5711), .B(n5710), .Z(n5689) );
  NANDN U7739 ( .A(n5666), .B(n5665), .Z(n5670) );
  NANDN U7740 ( .A(n5668), .B(n5667), .Z(n5669) );
  AND U7741 ( .A(n5670), .B(n5669), .Z(n5688) );
  XNOR U7742 ( .A(n5689), .B(n5688), .Z(n5690) );
  NANDN U7743 ( .A(n5672), .B(n5671), .Z(n5676) );
  NAND U7744 ( .A(n5674), .B(n5673), .Z(n5675) );
  NAND U7745 ( .A(n5676), .B(n5675), .Z(n5691) );
  XNOR U7746 ( .A(n5690), .B(n5691), .Z(n5682) );
  XNOR U7747 ( .A(n5683), .B(n5682), .Z(n5684) );
  XNOR U7748 ( .A(n5685), .B(n5684), .Z(n5714) );
  XNOR U7749 ( .A(sreg[1059]), .B(n5714), .Z(n5716) );
  NANDN U7750 ( .A(sreg[1058]), .B(n5677), .Z(n5681) );
  NAND U7751 ( .A(n5679), .B(n5678), .Z(n5680) );
  NAND U7752 ( .A(n5681), .B(n5680), .Z(n5715) );
  XNOR U7753 ( .A(n5716), .B(n5715), .Z(c[1059]) );
  NANDN U7754 ( .A(n5683), .B(n5682), .Z(n5687) );
  NANDN U7755 ( .A(n5685), .B(n5684), .Z(n5686) );
  AND U7756 ( .A(n5687), .B(n5686), .Z(n5722) );
  NANDN U7757 ( .A(n5689), .B(n5688), .Z(n5693) );
  NANDN U7758 ( .A(n5691), .B(n5690), .Z(n5692) );
  AND U7759 ( .A(n5693), .B(n5692), .Z(n5720) );
  NAND U7760 ( .A(n42143), .B(n5694), .Z(n5696) );
  XNOR U7761 ( .A(a[38]), .B(n4077), .Z(n5731) );
  NAND U7762 ( .A(n42144), .B(n5731), .Z(n5695) );
  AND U7763 ( .A(n5696), .B(n5695), .Z(n5746) );
  XOR U7764 ( .A(a[42]), .B(n42012), .Z(n5734) );
  XNOR U7765 ( .A(n5746), .B(n5745), .Z(n5748) );
  AND U7766 ( .A(a[44]), .B(b[0]), .Z(n5698) );
  XNOR U7767 ( .A(n5698), .B(n4071), .Z(n5700) );
  NANDN U7768 ( .A(b[0]), .B(a[43]), .Z(n5699) );
  NAND U7769 ( .A(n5700), .B(n5699), .Z(n5742) );
  XOR U7770 ( .A(a[40]), .B(n42085), .Z(n5735) );
  AND U7771 ( .A(a[36]), .B(b[7]), .Z(n5739) );
  XNOR U7772 ( .A(n5740), .B(n5739), .Z(n5741) );
  XNOR U7773 ( .A(n5742), .B(n5741), .Z(n5747) );
  XOR U7774 ( .A(n5748), .B(n5747), .Z(n5726) );
  NANDN U7775 ( .A(n5703), .B(n5702), .Z(n5707) );
  NANDN U7776 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U7777 ( .A(n5707), .B(n5706), .Z(n5725) );
  XNOR U7778 ( .A(n5726), .B(n5725), .Z(n5727) );
  NANDN U7779 ( .A(n5709), .B(n5708), .Z(n5713) );
  NAND U7780 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U7781 ( .A(n5713), .B(n5712), .Z(n5728) );
  XNOR U7782 ( .A(n5727), .B(n5728), .Z(n5719) );
  XNOR U7783 ( .A(n5720), .B(n5719), .Z(n5721) );
  XNOR U7784 ( .A(n5722), .B(n5721), .Z(n5751) );
  XNOR U7785 ( .A(sreg[1060]), .B(n5751), .Z(n5753) );
  NANDN U7786 ( .A(sreg[1059]), .B(n5714), .Z(n5718) );
  NAND U7787 ( .A(n5716), .B(n5715), .Z(n5717) );
  NAND U7788 ( .A(n5718), .B(n5717), .Z(n5752) );
  XNOR U7789 ( .A(n5753), .B(n5752), .Z(c[1060]) );
  NANDN U7790 ( .A(n5720), .B(n5719), .Z(n5724) );
  NANDN U7791 ( .A(n5722), .B(n5721), .Z(n5723) );
  AND U7792 ( .A(n5724), .B(n5723), .Z(n5759) );
  NANDN U7793 ( .A(n5726), .B(n5725), .Z(n5730) );
  NANDN U7794 ( .A(n5728), .B(n5727), .Z(n5729) );
  AND U7795 ( .A(n5730), .B(n5729), .Z(n5757) );
  NAND U7796 ( .A(n42143), .B(n5731), .Z(n5733) );
  XNOR U7797 ( .A(a[39]), .B(n4077), .Z(n5768) );
  NAND U7798 ( .A(n42144), .B(n5768), .Z(n5732) );
  AND U7799 ( .A(n5733), .B(n5732), .Z(n5783) );
  XOR U7800 ( .A(a[43]), .B(n42012), .Z(n5771) );
  XNOR U7801 ( .A(n5783), .B(n5782), .Z(n5785) );
  XOR U7802 ( .A(a[41]), .B(n42085), .Z(n5775) );
  AND U7803 ( .A(a[37]), .B(b[7]), .Z(n5776) );
  XNOR U7804 ( .A(n5777), .B(n5776), .Z(n5778) );
  AND U7805 ( .A(a[45]), .B(b[0]), .Z(n5736) );
  XNOR U7806 ( .A(n5736), .B(n4071), .Z(n5738) );
  NANDN U7807 ( .A(b[0]), .B(a[44]), .Z(n5737) );
  NAND U7808 ( .A(n5738), .B(n5737), .Z(n5779) );
  XNOR U7809 ( .A(n5778), .B(n5779), .Z(n5784) );
  XOR U7810 ( .A(n5785), .B(n5784), .Z(n5763) );
  NANDN U7811 ( .A(n5740), .B(n5739), .Z(n5744) );
  NANDN U7812 ( .A(n5742), .B(n5741), .Z(n5743) );
  AND U7813 ( .A(n5744), .B(n5743), .Z(n5762) );
  XNOR U7814 ( .A(n5763), .B(n5762), .Z(n5764) );
  NANDN U7815 ( .A(n5746), .B(n5745), .Z(n5750) );
  NAND U7816 ( .A(n5748), .B(n5747), .Z(n5749) );
  NAND U7817 ( .A(n5750), .B(n5749), .Z(n5765) );
  XNOR U7818 ( .A(n5764), .B(n5765), .Z(n5756) );
  XNOR U7819 ( .A(n5757), .B(n5756), .Z(n5758) );
  XNOR U7820 ( .A(n5759), .B(n5758), .Z(n5788) );
  XNOR U7821 ( .A(sreg[1061]), .B(n5788), .Z(n5790) );
  NANDN U7822 ( .A(sreg[1060]), .B(n5751), .Z(n5755) );
  NAND U7823 ( .A(n5753), .B(n5752), .Z(n5754) );
  NAND U7824 ( .A(n5755), .B(n5754), .Z(n5789) );
  XNOR U7825 ( .A(n5790), .B(n5789), .Z(c[1061]) );
  NANDN U7826 ( .A(n5757), .B(n5756), .Z(n5761) );
  NANDN U7827 ( .A(n5759), .B(n5758), .Z(n5760) );
  AND U7828 ( .A(n5761), .B(n5760), .Z(n5796) );
  NANDN U7829 ( .A(n5763), .B(n5762), .Z(n5767) );
  NANDN U7830 ( .A(n5765), .B(n5764), .Z(n5766) );
  AND U7831 ( .A(n5767), .B(n5766), .Z(n5794) );
  NAND U7832 ( .A(n42143), .B(n5768), .Z(n5770) );
  XNOR U7833 ( .A(a[40]), .B(n4077), .Z(n5805) );
  NAND U7834 ( .A(n42144), .B(n5805), .Z(n5769) );
  AND U7835 ( .A(n5770), .B(n5769), .Z(n5820) );
  XOR U7836 ( .A(a[44]), .B(n42012), .Z(n5808) );
  XNOR U7837 ( .A(n5820), .B(n5819), .Z(n5822) );
  AND U7838 ( .A(a[46]), .B(b[0]), .Z(n5772) );
  XNOR U7839 ( .A(n5772), .B(n4071), .Z(n5774) );
  NANDN U7840 ( .A(b[0]), .B(a[45]), .Z(n5773) );
  NAND U7841 ( .A(n5774), .B(n5773), .Z(n5816) );
  XOR U7842 ( .A(a[42]), .B(n42085), .Z(n5812) );
  AND U7843 ( .A(a[38]), .B(b[7]), .Z(n5813) );
  XNOR U7844 ( .A(n5814), .B(n5813), .Z(n5815) );
  XNOR U7845 ( .A(n5816), .B(n5815), .Z(n5821) );
  XOR U7846 ( .A(n5822), .B(n5821), .Z(n5800) );
  NANDN U7847 ( .A(n5777), .B(n5776), .Z(n5781) );
  NANDN U7848 ( .A(n5779), .B(n5778), .Z(n5780) );
  AND U7849 ( .A(n5781), .B(n5780), .Z(n5799) );
  XNOR U7850 ( .A(n5800), .B(n5799), .Z(n5801) );
  NANDN U7851 ( .A(n5783), .B(n5782), .Z(n5787) );
  NAND U7852 ( .A(n5785), .B(n5784), .Z(n5786) );
  NAND U7853 ( .A(n5787), .B(n5786), .Z(n5802) );
  XNOR U7854 ( .A(n5801), .B(n5802), .Z(n5793) );
  XNOR U7855 ( .A(n5794), .B(n5793), .Z(n5795) );
  XNOR U7856 ( .A(n5796), .B(n5795), .Z(n5825) );
  XNOR U7857 ( .A(sreg[1062]), .B(n5825), .Z(n5827) );
  NANDN U7858 ( .A(sreg[1061]), .B(n5788), .Z(n5792) );
  NAND U7859 ( .A(n5790), .B(n5789), .Z(n5791) );
  NAND U7860 ( .A(n5792), .B(n5791), .Z(n5826) );
  XNOR U7861 ( .A(n5827), .B(n5826), .Z(c[1062]) );
  NANDN U7862 ( .A(n5794), .B(n5793), .Z(n5798) );
  NANDN U7863 ( .A(n5796), .B(n5795), .Z(n5797) );
  AND U7864 ( .A(n5798), .B(n5797), .Z(n5833) );
  NANDN U7865 ( .A(n5800), .B(n5799), .Z(n5804) );
  NANDN U7866 ( .A(n5802), .B(n5801), .Z(n5803) );
  AND U7867 ( .A(n5804), .B(n5803), .Z(n5831) );
  NAND U7868 ( .A(n42143), .B(n5805), .Z(n5807) );
  XNOR U7869 ( .A(a[41]), .B(n4077), .Z(n5842) );
  NAND U7870 ( .A(n42144), .B(n5842), .Z(n5806) );
  AND U7871 ( .A(n5807), .B(n5806), .Z(n5857) );
  XOR U7872 ( .A(a[45]), .B(n42012), .Z(n5845) );
  XNOR U7873 ( .A(n5857), .B(n5856), .Z(n5859) );
  AND U7874 ( .A(a[47]), .B(b[0]), .Z(n5809) );
  XNOR U7875 ( .A(n5809), .B(n4071), .Z(n5811) );
  NANDN U7876 ( .A(b[0]), .B(a[46]), .Z(n5810) );
  NAND U7877 ( .A(n5811), .B(n5810), .Z(n5853) );
  XOR U7878 ( .A(a[43]), .B(n42085), .Z(n5849) );
  AND U7879 ( .A(a[39]), .B(b[7]), .Z(n5850) );
  XNOR U7880 ( .A(n5851), .B(n5850), .Z(n5852) );
  XNOR U7881 ( .A(n5853), .B(n5852), .Z(n5858) );
  XOR U7882 ( .A(n5859), .B(n5858), .Z(n5837) );
  NANDN U7883 ( .A(n5814), .B(n5813), .Z(n5818) );
  NANDN U7884 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U7885 ( .A(n5818), .B(n5817), .Z(n5836) );
  XNOR U7886 ( .A(n5837), .B(n5836), .Z(n5838) );
  NANDN U7887 ( .A(n5820), .B(n5819), .Z(n5824) );
  NAND U7888 ( .A(n5822), .B(n5821), .Z(n5823) );
  NAND U7889 ( .A(n5824), .B(n5823), .Z(n5839) );
  XNOR U7890 ( .A(n5838), .B(n5839), .Z(n5830) );
  XNOR U7891 ( .A(n5831), .B(n5830), .Z(n5832) );
  XNOR U7892 ( .A(n5833), .B(n5832), .Z(n5862) );
  XNOR U7893 ( .A(sreg[1063]), .B(n5862), .Z(n5864) );
  NANDN U7894 ( .A(sreg[1062]), .B(n5825), .Z(n5829) );
  NAND U7895 ( .A(n5827), .B(n5826), .Z(n5828) );
  NAND U7896 ( .A(n5829), .B(n5828), .Z(n5863) );
  XNOR U7897 ( .A(n5864), .B(n5863), .Z(c[1063]) );
  NANDN U7898 ( .A(n5831), .B(n5830), .Z(n5835) );
  NANDN U7899 ( .A(n5833), .B(n5832), .Z(n5834) );
  AND U7900 ( .A(n5835), .B(n5834), .Z(n5870) );
  NANDN U7901 ( .A(n5837), .B(n5836), .Z(n5841) );
  NANDN U7902 ( .A(n5839), .B(n5838), .Z(n5840) );
  AND U7903 ( .A(n5841), .B(n5840), .Z(n5868) );
  NAND U7904 ( .A(n42143), .B(n5842), .Z(n5844) );
  XNOR U7905 ( .A(a[42]), .B(n4077), .Z(n5879) );
  NAND U7906 ( .A(n42144), .B(n5879), .Z(n5843) );
  AND U7907 ( .A(n5844), .B(n5843), .Z(n5894) );
  XOR U7908 ( .A(a[46]), .B(n42012), .Z(n5882) );
  XNOR U7909 ( .A(n5894), .B(n5893), .Z(n5896) );
  AND U7910 ( .A(a[48]), .B(b[0]), .Z(n5846) );
  XNOR U7911 ( .A(n5846), .B(n4071), .Z(n5848) );
  NANDN U7912 ( .A(b[0]), .B(a[47]), .Z(n5847) );
  NAND U7913 ( .A(n5848), .B(n5847), .Z(n5890) );
  XOR U7914 ( .A(a[44]), .B(n42085), .Z(n5886) );
  AND U7915 ( .A(a[40]), .B(b[7]), .Z(n5887) );
  XNOR U7916 ( .A(n5888), .B(n5887), .Z(n5889) );
  XNOR U7917 ( .A(n5890), .B(n5889), .Z(n5895) );
  XOR U7918 ( .A(n5896), .B(n5895), .Z(n5874) );
  NANDN U7919 ( .A(n5851), .B(n5850), .Z(n5855) );
  NANDN U7920 ( .A(n5853), .B(n5852), .Z(n5854) );
  AND U7921 ( .A(n5855), .B(n5854), .Z(n5873) );
  XNOR U7922 ( .A(n5874), .B(n5873), .Z(n5875) );
  NANDN U7923 ( .A(n5857), .B(n5856), .Z(n5861) );
  NAND U7924 ( .A(n5859), .B(n5858), .Z(n5860) );
  NAND U7925 ( .A(n5861), .B(n5860), .Z(n5876) );
  XNOR U7926 ( .A(n5875), .B(n5876), .Z(n5867) );
  XNOR U7927 ( .A(n5868), .B(n5867), .Z(n5869) );
  XNOR U7928 ( .A(n5870), .B(n5869), .Z(n5899) );
  XNOR U7929 ( .A(sreg[1064]), .B(n5899), .Z(n5901) );
  NANDN U7930 ( .A(sreg[1063]), .B(n5862), .Z(n5866) );
  NAND U7931 ( .A(n5864), .B(n5863), .Z(n5865) );
  NAND U7932 ( .A(n5866), .B(n5865), .Z(n5900) );
  XNOR U7933 ( .A(n5901), .B(n5900), .Z(c[1064]) );
  NANDN U7934 ( .A(n5868), .B(n5867), .Z(n5872) );
  NANDN U7935 ( .A(n5870), .B(n5869), .Z(n5871) );
  AND U7936 ( .A(n5872), .B(n5871), .Z(n5907) );
  NANDN U7937 ( .A(n5874), .B(n5873), .Z(n5878) );
  NANDN U7938 ( .A(n5876), .B(n5875), .Z(n5877) );
  AND U7939 ( .A(n5878), .B(n5877), .Z(n5905) );
  NAND U7940 ( .A(n42143), .B(n5879), .Z(n5881) );
  XNOR U7941 ( .A(a[43]), .B(n4078), .Z(n5916) );
  NAND U7942 ( .A(n42144), .B(n5916), .Z(n5880) );
  AND U7943 ( .A(n5881), .B(n5880), .Z(n5931) );
  XOR U7944 ( .A(a[47]), .B(n42012), .Z(n5919) );
  XNOR U7945 ( .A(n5931), .B(n5930), .Z(n5933) );
  AND U7946 ( .A(a[49]), .B(b[0]), .Z(n5883) );
  XNOR U7947 ( .A(n5883), .B(n4071), .Z(n5885) );
  NANDN U7948 ( .A(b[0]), .B(a[48]), .Z(n5884) );
  NAND U7949 ( .A(n5885), .B(n5884), .Z(n5927) );
  XOR U7950 ( .A(a[45]), .B(n42085), .Z(n5923) );
  AND U7951 ( .A(a[41]), .B(b[7]), .Z(n5924) );
  XNOR U7952 ( .A(n5925), .B(n5924), .Z(n5926) );
  XNOR U7953 ( .A(n5927), .B(n5926), .Z(n5932) );
  XOR U7954 ( .A(n5933), .B(n5932), .Z(n5911) );
  NANDN U7955 ( .A(n5888), .B(n5887), .Z(n5892) );
  NANDN U7956 ( .A(n5890), .B(n5889), .Z(n5891) );
  AND U7957 ( .A(n5892), .B(n5891), .Z(n5910) );
  XNOR U7958 ( .A(n5911), .B(n5910), .Z(n5912) );
  NANDN U7959 ( .A(n5894), .B(n5893), .Z(n5898) );
  NAND U7960 ( .A(n5896), .B(n5895), .Z(n5897) );
  NAND U7961 ( .A(n5898), .B(n5897), .Z(n5913) );
  XNOR U7962 ( .A(n5912), .B(n5913), .Z(n5904) );
  XNOR U7963 ( .A(n5905), .B(n5904), .Z(n5906) );
  XNOR U7964 ( .A(n5907), .B(n5906), .Z(n5936) );
  XNOR U7965 ( .A(sreg[1065]), .B(n5936), .Z(n5938) );
  NANDN U7966 ( .A(sreg[1064]), .B(n5899), .Z(n5903) );
  NAND U7967 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U7968 ( .A(n5903), .B(n5902), .Z(n5937) );
  XNOR U7969 ( .A(n5938), .B(n5937), .Z(c[1065]) );
  NANDN U7970 ( .A(n5905), .B(n5904), .Z(n5909) );
  NANDN U7971 ( .A(n5907), .B(n5906), .Z(n5908) );
  AND U7972 ( .A(n5909), .B(n5908), .Z(n5944) );
  NANDN U7973 ( .A(n5911), .B(n5910), .Z(n5915) );
  NANDN U7974 ( .A(n5913), .B(n5912), .Z(n5914) );
  AND U7975 ( .A(n5915), .B(n5914), .Z(n5942) );
  NAND U7976 ( .A(n42143), .B(n5916), .Z(n5918) );
  XNOR U7977 ( .A(a[44]), .B(n4078), .Z(n5953) );
  NAND U7978 ( .A(n42144), .B(n5953), .Z(n5917) );
  AND U7979 ( .A(n5918), .B(n5917), .Z(n5968) );
  XOR U7980 ( .A(a[48]), .B(n42012), .Z(n5956) );
  XNOR U7981 ( .A(n5968), .B(n5967), .Z(n5970) );
  AND U7982 ( .A(a[50]), .B(b[0]), .Z(n5920) );
  XNOR U7983 ( .A(n5920), .B(n4071), .Z(n5922) );
  NANDN U7984 ( .A(b[0]), .B(a[49]), .Z(n5921) );
  NAND U7985 ( .A(n5922), .B(n5921), .Z(n5964) );
  XOR U7986 ( .A(a[46]), .B(n42085), .Z(n5957) );
  AND U7987 ( .A(a[42]), .B(b[7]), .Z(n5961) );
  XNOR U7988 ( .A(n5962), .B(n5961), .Z(n5963) );
  XNOR U7989 ( .A(n5964), .B(n5963), .Z(n5969) );
  XOR U7990 ( .A(n5970), .B(n5969), .Z(n5948) );
  NANDN U7991 ( .A(n5925), .B(n5924), .Z(n5929) );
  NANDN U7992 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U7993 ( .A(n5929), .B(n5928), .Z(n5947) );
  XNOR U7994 ( .A(n5948), .B(n5947), .Z(n5949) );
  NANDN U7995 ( .A(n5931), .B(n5930), .Z(n5935) );
  NAND U7996 ( .A(n5933), .B(n5932), .Z(n5934) );
  NAND U7997 ( .A(n5935), .B(n5934), .Z(n5950) );
  XNOR U7998 ( .A(n5949), .B(n5950), .Z(n5941) );
  XNOR U7999 ( .A(n5942), .B(n5941), .Z(n5943) );
  XNOR U8000 ( .A(n5944), .B(n5943), .Z(n5973) );
  XNOR U8001 ( .A(sreg[1066]), .B(n5973), .Z(n5975) );
  NANDN U8002 ( .A(sreg[1065]), .B(n5936), .Z(n5940) );
  NAND U8003 ( .A(n5938), .B(n5937), .Z(n5939) );
  NAND U8004 ( .A(n5940), .B(n5939), .Z(n5974) );
  XNOR U8005 ( .A(n5975), .B(n5974), .Z(c[1066]) );
  NANDN U8006 ( .A(n5942), .B(n5941), .Z(n5946) );
  NANDN U8007 ( .A(n5944), .B(n5943), .Z(n5945) );
  AND U8008 ( .A(n5946), .B(n5945), .Z(n5981) );
  NANDN U8009 ( .A(n5948), .B(n5947), .Z(n5952) );
  NANDN U8010 ( .A(n5950), .B(n5949), .Z(n5951) );
  AND U8011 ( .A(n5952), .B(n5951), .Z(n5979) );
  NAND U8012 ( .A(n42143), .B(n5953), .Z(n5955) );
  XNOR U8013 ( .A(a[45]), .B(n4078), .Z(n5990) );
  NAND U8014 ( .A(n42144), .B(n5990), .Z(n5954) );
  AND U8015 ( .A(n5955), .B(n5954), .Z(n6005) );
  XOR U8016 ( .A(a[49]), .B(n42012), .Z(n5993) );
  XNOR U8017 ( .A(n6005), .B(n6004), .Z(n6007) );
  XOR U8018 ( .A(a[47]), .B(n42085), .Z(n5997) );
  AND U8019 ( .A(a[43]), .B(b[7]), .Z(n5998) );
  XNOR U8020 ( .A(n5999), .B(n5998), .Z(n6000) );
  AND U8021 ( .A(a[51]), .B(b[0]), .Z(n5958) );
  XNOR U8022 ( .A(n5958), .B(n4071), .Z(n5960) );
  NANDN U8023 ( .A(b[0]), .B(a[50]), .Z(n5959) );
  NAND U8024 ( .A(n5960), .B(n5959), .Z(n6001) );
  XNOR U8025 ( .A(n6000), .B(n6001), .Z(n6006) );
  XOR U8026 ( .A(n6007), .B(n6006), .Z(n5985) );
  NANDN U8027 ( .A(n5962), .B(n5961), .Z(n5966) );
  NANDN U8028 ( .A(n5964), .B(n5963), .Z(n5965) );
  AND U8029 ( .A(n5966), .B(n5965), .Z(n5984) );
  XNOR U8030 ( .A(n5985), .B(n5984), .Z(n5986) );
  NANDN U8031 ( .A(n5968), .B(n5967), .Z(n5972) );
  NAND U8032 ( .A(n5970), .B(n5969), .Z(n5971) );
  NAND U8033 ( .A(n5972), .B(n5971), .Z(n5987) );
  XNOR U8034 ( .A(n5986), .B(n5987), .Z(n5978) );
  XNOR U8035 ( .A(n5979), .B(n5978), .Z(n5980) );
  XNOR U8036 ( .A(n5981), .B(n5980), .Z(n6010) );
  XNOR U8037 ( .A(sreg[1067]), .B(n6010), .Z(n6012) );
  NANDN U8038 ( .A(sreg[1066]), .B(n5973), .Z(n5977) );
  NAND U8039 ( .A(n5975), .B(n5974), .Z(n5976) );
  NAND U8040 ( .A(n5977), .B(n5976), .Z(n6011) );
  XNOR U8041 ( .A(n6012), .B(n6011), .Z(c[1067]) );
  NANDN U8042 ( .A(n5979), .B(n5978), .Z(n5983) );
  NANDN U8043 ( .A(n5981), .B(n5980), .Z(n5982) );
  AND U8044 ( .A(n5983), .B(n5982), .Z(n6018) );
  NANDN U8045 ( .A(n5985), .B(n5984), .Z(n5989) );
  NANDN U8046 ( .A(n5987), .B(n5986), .Z(n5988) );
  AND U8047 ( .A(n5989), .B(n5988), .Z(n6016) );
  NAND U8048 ( .A(n42143), .B(n5990), .Z(n5992) );
  XNOR U8049 ( .A(a[46]), .B(n4078), .Z(n6027) );
  NAND U8050 ( .A(n42144), .B(n6027), .Z(n5991) );
  AND U8051 ( .A(n5992), .B(n5991), .Z(n6042) );
  XOR U8052 ( .A(a[50]), .B(n42012), .Z(n6030) );
  XNOR U8053 ( .A(n6042), .B(n6041), .Z(n6044) );
  AND U8054 ( .A(a[52]), .B(b[0]), .Z(n5994) );
  XNOR U8055 ( .A(n5994), .B(n4071), .Z(n5996) );
  NANDN U8056 ( .A(b[0]), .B(a[51]), .Z(n5995) );
  NAND U8057 ( .A(n5996), .B(n5995), .Z(n6038) );
  XOR U8058 ( .A(a[48]), .B(n42085), .Z(n6034) );
  AND U8059 ( .A(a[44]), .B(b[7]), .Z(n6035) );
  XNOR U8060 ( .A(n6036), .B(n6035), .Z(n6037) );
  XNOR U8061 ( .A(n6038), .B(n6037), .Z(n6043) );
  XOR U8062 ( .A(n6044), .B(n6043), .Z(n6022) );
  NANDN U8063 ( .A(n5999), .B(n5998), .Z(n6003) );
  NANDN U8064 ( .A(n6001), .B(n6000), .Z(n6002) );
  AND U8065 ( .A(n6003), .B(n6002), .Z(n6021) );
  XNOR U8066 ( .A(n6022), .B(n6021), .Z(n6023) );
  NANDN U8067 ( .A(n6005), .B(n6004), .Z(n6009) );
  NAND U8068 ( .A(n6007), .B(n6006), .Z(n6008) );
  NAND U8069 ( .A(n6009), .B(n6008), .Z(n6024) );
  XNOR U8070 ( .A(n6023), .B(n6024), .Z(n6015) );
  XNOR U8071 ( .A(n6016), .B(n6015), .Z(n6017) );
  XNOR U8072 ( .A(n6018), .B(n6017), .Z(n6047) );
  XNOR U8073 ( .A(sreg[1068]), .B(n6047), .Z(n6049) );
  NANDN U8074 ( .A(sreg[1067]), .B(n6010), .Z(n6014) );
  NAND U8075 ( .A(n6012), .B(n6011), .Z(n6013) );
  NAND U8076 ( .A(n6014), .B(n6013), .Z(n6048) );
  XNOR U8077 ( .A(n6049), .B(n6048), .Z(c[1068]) );
  NANDN U8078 ( .A(n6016), .B(n6015), .Z(n6020) );
  NANDN U8079 ( .A(n6018), .B(n6017), .Z(n6019) );
  AND U8080 ( .A(n6020), .B(n6019), .Z(n6055) );
  NANDN U8081 ( .A(n6022), .B(n6021), .Z(n6026) );
  NANDN U8082 ( .A(n6024), .B(n6023), .Z(n6025) );
  AND U8083 ( .A(n6026), .B(n6025), .Z(n6053) );
  NAND U8084 ( .A(n42143), .B(n6027), .Z(n6029) );
  XNOR U8085 ( .A(a[47]), .B(n4078), .Z(n6064) );
  NAND U8086 ( .A(n42144), .B(n6064), .Z(n6028) );
  AND U8087 ( .A(n6029), .B(n6028), .Z(n6079) );
  XOR U8088 ( .A(a[51]), .B(n42012), .Z(n6067) );
  XNOR U8089 ( .A(n6079), .B(n6078), .Z(n6081) );
  AND U8090 ( .A(a[53]), .B(b[0]), .Z(n6031) );
  XNOR U8091 ( .A(n6031), .B(n4071), .Z(n6033) );
  NANDN U8092 ( .A(b[0]), .B(a[52]), .Z(n6032) );
  NAND U8093 ( .A(n6033), .B(n6032), .Z(n6075) );
  XOR U8094 ( .A(a[49]), .B(n42085), .Z(n6071) );
  AND U8095 ( .A(a[45]), .B(b[7]), .Z(n6072) );
  XNOR U8096 ( .A(n6073), .B(n6072), .Z(n6074) );
  XNOR U8097 ( .A(n6075), .B(n6074), .Z(n6080) );
  XOR U8098 ( .A(n6081), .B(n6080), .Z(n6059) );
  NANDN U8099 ( .A(n6036), .B(n6035), .Z(n6040) );
  NANDN U8100 ( .A(n6038), .B(n6037), .Z(n6039) );
  AND U8101 ( .A(n6040), .B(n6039), .Z(n6058) );
  XNOR U8102 ( .A(n6059), .B(n6058), .Z(n6060) );
  NANDN U8103 ( .A(n6042), .B(n6041), .Z(n6046) );
  NAND U8104 ( .A(n6044), .B(n6043), .Z(n6045) );
  NAND U8105 ( .A(n6046), .B(n6045), .Z(n6061) );
  XNOR U8106 ( .A(n6060), .B(n6061), .Z(n6052) );
  XNOR U8107 ( .A(n6053), .B(n6052), .Z(n6054) );
  XNOR U8108 ( .A(n6055), .B(n6054), .Z(n6084) );
  XNOR U8109 ( .A(sreg[1069]), .B(n6084), .Z(n6086) );
  NANDN U8110 ( .A(sreg[1068]), .B(n6047), .Z(n6051) );
  NAND U8111 ( .A(n6049), .B(n6048), .Z(n6050) );
  NAND U8112 ( .A(n6051), .B(n6050), .Z(n6085) );
  XNOR U8113 ( .A(n6086), .B(n6085), .Z(c[1069]) );
  NANDN U8114 ( .A(n6053), .B(n6052), .Z(n6057) );
  NANDN U8115 ( .A(n6055), .B(n6054), .Z(n6056) );
  AND U8116 ( .A(n6057), .B(n6056), .Z(n6092) );
  NANDN U8117 ( .A(n6059), .B(n6058), .Z(n6063) );
  NANDN U8118 ( .A(n6061), .B(n6060), .Z(n6062) );
  AND U8119 ( .A(n6063), .B(n6062), .Z(n6090) );
  NAND U8120 ( .A(n42143), .B(n6064), .Z(n6066) );
  XNOR U8121 ( .A(a[48]), .B(n4078), .Z(n6101) );
  NAND U8122 ( .A(n42144), .B(n6101), .Z(n6065) );
  AND U8123 ( .A(n6066), .B(n6065), .Z(n6116) );
  XOR U8124 ( .A(a[52]), .B(n42012), .Z(n6104) );
  XNOR U8125 ( .A(n6116), .B(n6115), .Z(n6118) );
  AND U8126 ( .A(a[54]), .B(b[0]), .Z(n6068) );
  XNOR U8127 ( .A(n6068), .B(n4071), .Z(n6070) );
  NANDN U8128 ( .A(b[0]), .B(a[53]), .Z(n6069) );
  NAND U8129 ( .A(n6070), .B(n6069), .Z(n6112) );
  XOR U8130 ( .A(a[50]), .B(n42085), .Z(n6108) );
  AND U8131 ( .A(a[46]), .B(b[7]), .Z(n6109) );
  XNOR U8132 ( .A(n6110), .B(n6109), .Z(n6111) );
  XNOR U8133 ( .A(n6112), .B(n6111), .Z(n6117) );
  XOR U8134 ( .A(n6118), .B(n6117), .Z(n6096) );
  NANDN U8135 ( .A(n6073), .B(n6072), .Z(n6077) );
  NANDN U8136 ( .A(n6075), .B(n6074), .Z(n6076) );
  AND U8137 ( .A(n6077), .B(n6076), .Z(n6095) );
  XNOR U8138 ( .A(n6096), .B(n6095), .Z(n6097) );
  NANDN U8139 ( .A(n6079), .B(n6078), .Z(n6083) );
  NAND U8140 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U8141 ( .A(n6083), .B(n6082), .Z(n6098) );
  XNOR U8142 ( .A(n6097), .B(n6098), .Z(n6089) );
  XNOR U8143 ( .A(n6090), .B(n6089), .Z(n6091) );
  XNOR U8144 ( .A(n6092), .B(n6091), .Z(n6121) );
  XNOR U8145 ( .A(sreg[1070]), .B(n6121), .Z(n6123) );
  NANDN U8146 ( .A(sreg[1069]), .B(n6084), .Z(n6088) );
  NAND U8147 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U8148 ( .A(n6088), .B(n6087), .Z(n6122) );
  XNOR U8149 ( .A(n6123), .B(n6122), .Z(c[1070]) );
  NANDN U8150 ( .A(n6090), .B(n6089), .Z(n6094) );
  NANDN U8151 ( .A(n6092), .B(n6091), .Z(n6093) );
  AND U8152 ( .A(n6094), .B(n6093), .Z(n6129) );
  NANDN U8153 ( .A(n6096), .B(n6095), .Z(n6100) );
  NANDN U8154 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U8155 ( .A(n6100), .B(n6099), .Z(n6127) );
  NAND U8156 ( .A(n42143), .B(n6101), .Z(n6103) );
  XNOR U8157 ( .A(a[49]), .B(n4078), .Z(n6138) );
  NAND U8158 ( .A(n42144), .B(n6138), .Z(n6102) );
  AND U8159 ( .A(n6103), .B(n6102), .Z(n6153) );
  XOR U8160 ( .A(a[53]), .B(n42012), .Z(n6141) );
  XNOR U8161 ( .A(n6153), .B(n6152), .Z(n6155) );
  AND U8162 ( .A(a[55]), .B(b[0]), .Z(n6105) );
  XNOR U8163 ( .A(n6105), .B(n4071), .Z(n6107) );
  NANDN U8164 ( .A(b[0]), .B(a[54]), .Z(n6106) );
  NAND U8165 ( .A(n6107), .B(n6106), .Z(n6149) );
  XOR U8166 ( .A(a[51]), .B(n42085), .Z(n6142) );
  AND U8167 ( .A(a[47]), .B(b[7]), .Z(n6146) );
  XNOR U8168 ( .A(n6147), .B(n6146), .Z(n6148) );
  XNOR U8169 ( .A(n6149), .B(n6148), .Z(n6154) );
  XOR U8170 ( .A(n6155), .B(n6154), .Z(n6133) );
  NANDN U8171 ( .A(n6110), .B(n6109), .Z(n6114) );
  NANDN U8172 ( .A(n6112), .B(n6111), .Z(n6113) );
  AND U8173 ( .A(n6114), .B(n6113), .Z(n6132) );
  XNOR U8174 ( .A(n6133), .B(n6132), .Z(n6134) );
  NANDN U8175 ( .A(n6116), .B(n6115), .Z(n6120) );
  NAND U8176 ( .A(n6118), .B(n6117), .Z(n6119) );
  NAND U8177 ( .A(n6120), .B(n6119), .Z(n6135) );
  XNOR U8178 ( .A(n6134), .B(n6135), .Z(n6126) );
  XNOR U8179 ( .A(n6127), .B(n6126), .Z(n6128) );
  XNOR U8180 ( .A(n6129), .B(n6128), .Z(n6158) );
  XNOR U8181 ( .A(sreg[1071]), .B(n6158), .Z(n6160) );
  NANDN U8182 ( .A(sreg[1070]), .B(n6121), .Z(n6125) );
  NAND U8183 ( .A(n6123), .B(n6122), .Z(n6124) );
  NAND U8184 ( .A(n6125), .B(n6124), .Z(n6159) );
  XNOR U8185 ( .A(n6160), .B(n6159), .Z(c[1071]) );
  NANDN U8186 ( .A(n6127), .B(n6126), .Z(n6131) );
  NANDN U8187 ( .A(n6129), .B(n6128), .Z(n6130) );
  AND U8188 ( .A(n6131), .B(n6130), .Z(n6166) );
  NANDN U8189 ( .A(n6133), .B(n6132), .Z(n6137) );
  NANDN U8190 ( .A(n6135), .B(n6134), .Z(n6136) );
  AND U8191 ( .A(n6137), .B(n6136), .Z(n6164) );
  NAND U8192 ( .A(n42143), .B(n6138), .Z(n6140) );
  XNOR U8193 ( .A(a[50]), .B(n4079), .Z(n6175) );
  NAND U8194 ( .A(n42144), .B(n6175), .Z(n6139) );
  AND U8195 ( .A(n6140), .B(n6139), .Z(n6190) );
  XOR U8196 ( .A(a[54]), .B(n42012), .Z(n6178) );
  XNOR U8197 ( .A(n6190), .B(n6189), .Z(n6192) );
  XOR U8198 ( .A(a[52]), .B(n42085), .Z(n6182) );
  AND U8199 ( .A(a[48]), .B(b[7]), .Z(n6183) );
  XNOR U8200 ( .A(n6184), .B(n6183), .Z(n6185) );
  AND U8201 ( .A(a[56]), .B(b[0]), .Z(n6143) );
  XNOR U8202 ( .A(n6143), .B(n4071), .Z(n6145) );
  NANDN U8203 ( .A(b[0]), .B(a[55]), .Z(n6144) );
  NAND U8204 ( .A(n6145), .B(n6144), .Z(n6186) );
  XNOR U8205 ( .A(n6185), .B(n6186), .Z(n6191) );
  XOR U8206 ( .A(n6192), .B(n6191), .Z(n6170) );
  NANDN U8207 ( .A(n6147), .B(n6146), .Z(n6151) );
  NANDN U8208 ( .A(n6149), .B(n6148), .Z(n6150) );
  AND U8209 ( .A(n6151), .B(n6150), .Z(n6169) );
  XNOR U8210 ( .A(n6170), .B(n6169), .Z(n6171) );
  NANDN U8211 ( .A(n6153), .B(n6152), .Z(n6157) );
  NAND U8212 ( .A(n6155), .B(n6154), .Z(n6156) );
  NAND U8213 ( .A(n6157), .B(n6156), .Z(n6172) );
  XNOR U8214 ( .A(n6171), .B(n6172), .Z(n6163) );
  XNOR U8215 ( .A(n6164), .B(n6163), .Z(n6165) );
  XNOR U8216 ( .A(n6166), .B(n6165), .Z(n6195) );
  XNOR U8217 ( .A(sreg[1072]), .B(n6195), .Z(n6197) );
  NANDN U8218 ( .A(sreg[1071]), .B(n6158), .Z(n6162) );
  NAND U8219 ( .A(n6160), .B(n6159), .Z(n6161) );
  NAND U8220 ( .A(n6162), .B(n6161), .Z(n6196) );
  XNOR U8221 ( .A(n6197), .B(n6196), .Z(c[1072]) );
  NANDN U8222 ( .A(n6164), .B(n6163), .Z(n6168) );
  NANDN U8223 ( .A(n6166), .B(n6165), .Z(n6167) );
  AND U8224 ( .A(n6168), .B(n6167), .Z(n6203) );
  NANDN U8225 ( .A(n6170), .B(n6169), .Z(n6174) );
  NANDN U8226 ( .A(n6172), .B(n6171), .Z(n6173) );
  AND U8227 ( .A(n6174), .B(n6173), .Z(n6201) );
  NAND U8228 ( .A(n42143), .B(n6175), .Z(n6177) );
  XNOR U8229 ( .A(a[51]), .B(n4079), .Z(n6212) );
  NAND U8230 ( .A(n42144), .B(n6212), .Z(n6176) );
  AND U8231 ( .A(n6177), .B(n6176), .Z(n6227) );
  XOR U8232 ( .A(a[55]), .B(n42012), .Z(n6215) );
  XNOR U8233 ( .A(n6227), .B(n6226), .Z(n6229) );
  AND U8234 ( .A(a[57]), .B(b[0]), .Z(n6179) );
  XNOR U8235 ( .A(n6179), .B(n4071), .Z(n6181) );
  NANDN U8236 ( .A(b[0]), .B(a[56]), .Z(n6180) );
  NAND U8237 ( .A(n6181), .B(n6180), .Z(n6223) );
  XOR U8238 ( .A(a[53]), .B(n42085), .Z(n6216) );
  AND U8239 ( .A(a[49]), .B(b[7]), .Z(n6220) );
  XNOR U8240 ( .A(n6221), .B(n6220), .Z(n6222) );
  XNOR U8241 ( .A(n6223), .B(n6222), .Z(n6228) );
  XOR U8242 ( .A(n6229), .B(n6228), .Z(n6207) );
  NANDN U8243 ( .A(n6184), .B(n6183), .Z(n6188) );
  NANDN U8244 ( .A(n6186), .B(n6185), .Z(n6187) );
  AND U8245 ( .A(n6188), .B(n6187), .Z(n6206) );
  XNOR U8246 ( .A(n6207), .B(n6206), .Z(n6208) );
  NANDN U8247 ( .A(n6190), .B(n6189), .Z(n6194) );
  NAND U8248 ( .A(n6192), .B(n6191), .Z(n6193) );
  NAND U8249 ( .A(n6194), .B(n6193), .Z(n6209) );
  XNOR U8250 ( .A(n6208), .B(n6209), .Z(n6200) );
  XNOR U8251 ( .A(n6201), .B(n6200), .Z(n6202) );
  XNOR U8252 ( .A(n6203), .B(n6202), .Z(n6232) );
  XNOR U8253 ( .A(sreg[1073]), .B(n6232), .Z(n6234) );
  NANDN U8254 ( .A(sreg[1072]), .B(n6195), .Z(n6199) );
  NAND U8255 ( .A(n6197), .B(n6196), .Z(n6198) );
  NAND U8256 ( .A(n6199), .B(n6198), .Z(n6233) );
  XNOR U8257 ( .A(n6234), .B(n6233), .Z(c[1073]) );
  NANDN U8258 ( .A(n6201), .B(n6200), .Z(n6205) );
  NANDN U8259 ( .A(n6203), .B(n6202), .Z(n6204) );
  AND U8260 ( .A(n6205), .B(n6204), .Z(n6240) );
  NANDN U8261 ( .A(n6207), .B(n6206), .Z(n6211) );
  NANDN U8262 ( .A(n6209), .B(n6208), .Z(n6210) );
  AND U8263 ( .A(n6211), .B(n6210), .Z(n6238) );
  NAND U8264 ( .A(n42143), .B(n6212), .Z(n6214) );
  XNOR U8265 ( .A(a[52]), .B(n4079), .Z(n6249) );
  NAND U8266 ( .A(n42144), .B(n6249), .Z(n6213) );
  AND U8267 ( .A(n6214), .B(n6213), .Z(n6264) );
  XOR U8268 ( .A(a[56]), .B(n42012), .Z(n6252) );
  XNOR U8269 ( .A(n6264), .B(n6263), .Z(n6266) );
  XOR U8270 ( .A(a[54]), .B(n42085), .Z(n6256) );
  AND U8271 ( .A(a[50]), .B(b[7]), .Z(n6257) );
  XNOR U8272 ( .A(n6258), .B(n6257), .Z(n6259) );
  AND U8273 ( .A(a[58]), .B(b[0]), .Z(n6217) );
  XNOR U8274 ( .A(n6217), .B(n4071), .Z(n6219) );
  NANDN U8275 ( .A(b[0]), .B(a[57]), .Z(n6218) );
  NAND U8276 ( .A(n6219), .B(n6218), .Z(n6260) );
  XNOR U8277 ( .A(n6259), .B(n6260), .Z(n6265) );
  XOR U8278 ( .A(n6266), .B(n6265), .Z(n6244) );
  NANDN U8279 ( .A(n6221), .B(n6220), .Z(n6225) );
  NANDN U8280 ( .A(n6223), .B(n6222), .Z(n6224) );
  AND U8281 ( .A(n6225), .B(n6224), .Z(n6243) );
  XNOR U8282 ( .A(n6244), .B(n6243), .Z(n6245) );
  NANDN U8283 ( .A(n6227), .B(n6226), .Z(n6231) );
  NAND U8284 ( .A(n6229), .B(n6228), .Z(n6230) );
  NAND U8285 ( .A(n6231), .B(n6230), .Z(n6246) );
  XNOR U8286 ( .A(n6245), .B(n6246), .Z(n6237) );
  XNOR U8287 ( .A(n6238), .B(n6237), .Z(n6239) );
  XNOR U8288 ( .A(n6240), .B(n6239), .Z(n6269) );
  XNOR U8289 ( .A(sreg[1074]), .B(n6269), .Z(n6271) );
  NANDN U8290 ( .A(sreg[1073]), .B(n6232), .Z(n6236) );
  NAND U8291 ( .A(n6234), .B(n6233), .Z(n6235) );
  NAND U8292 ( .A(n6236), .B(n6235), .Z(n6270) );
  XNOR U8293 ( .A(n6271), .B(n6270), .Z(c[1074]) );
  NANDN U8294 ( .A(n6238), .B(n6237), .Z(n6242) );
  NANDN U8295 ( .A(n6240), .B(n6239), .Z(n6241) );
  AND U8296 ( .A(n6242), .B(n6241), .Z(n6277) );
  NANDN U8297 ( .A(n6244), .B(n6243), .Z(n6248) );
  NANDN U8298 ( .A(n6246), .B(n6245), .Z(n6247) );
  AND U8299 ( .A(n6248), .B(n6247), .Z(n6275) );
  NAND U8300 ( .A(n42143), .B(n6249), .Z(n6251) );
  XNOR U8301 ( .A(a[53]), .B(n4079), .Z(n6286) );
  NAND U8302 ( .A(n42144), .B(n6286), .Z(n6250) );
  AND U8303 ( .A(n6251), .B(n6250), .Z(n6301) );
  XOR U8304 ( .A(a[57]), .B(n42012), .Z(n6289) );
  XNOR U8305 ( .A(n6301), .B(n6300), .Z(n6303) );
  AND U8306 ( .A(a[59]), .B(b[0]), .Z(n6253) );
  XNOR U8307 ( .A(n6253), .B(n4071), .Z(n6255) );
  NANDN U8308 ( .A(b[0]), .B(a[58]), .Z(n6254) );
  NAND U8309 ( .A(n6255), .B(n6254), .Z(n6297) );
  XOR U8310 ( .A(a[55]), .B(n42085), .Z(n6293) );
  AND U8311 ( .A(a[51]), .B(b[7]), .Z(n6294) );
  XNOR U8312 ( .A(n6295), .B(n6294), .Z(n6296) );
  XNOR U8313 ( .A(n6297), .B(n6296), .Z(n6302) );
  XOR U8314 ( .A(n6303), .B(n6302), .Z(n6281) );
  NANDN U8315 ( .A(n6258), .B(n6257), .Z(n6262) );
  NANDN U8316 ( .A(n6260), .B(n6259), .Z(n6261) );
  AND U8317 ( .A(n6262), .B(n6261), .Z(n6280) );
  XNOR U8318 ( .A(n6281), .B(n6280), .Z(n6282) );
  NANDN U8319 ( .A(n6264), .B(n6263), .Z(n6268) );
  NAND U8320 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U8321 ( .A(n6268), .B(n6267), .Z(n6283) );
  XNOR U8322 ( .A(n6282), .B(n6283), .Z(n6274) );
  XNOR U8323 ( .A(n6275), .B(n6274), .Z(n6276) );
  XNOR U8324 ( .A(n6277), .B(n6276), .Z(n6306) );
  XNOR U8325 ( .A(sreg[1075]), .B(n6306), .Z(n6308) );
  NANDN U8326 ( .A(sreg[1074]), .B(n6269), .Z(n6273) );
  NAND U8327 ( .A(n6271), .B(n6270), .Z(n6272) );
  NAND U8328 ( .A(n6273), .B(n6272), .Z(n6307) );
  XNOR U8329 ( .A(n6308), .B(n6307), .Z(c[1075]) );
  NANDN U8330 ( .A(n6275), .B(n6274), .Z(n6279) );
  NANDN U8331 ( .A(n6277), .B(n6276), .Z(n6278) );
  AND U8332 ( .A(n6279), .B(n6278), .Z(n6314) );
  NANDN U8333 ( .A(n6281), .B(n6280), .Z(n6285) );
  NANDN U8334 ( .A(n6283), .B(n6282), .Z(n6284) );
  AND U8335 ( .A(n6285), .B(n6284), .Z(n6312) );
  NAND U8336 ( .A(n42143), .B(n6286), .Z(n6288) );
  XNOR U8337 ( .A(a[54]), .B(n4079), .Z(n6323) );
  NAND U8338 ( .A(n42144), .B(n6323), .Z(n6287) );
  AND U8339 ( .A(n6288), .B(n6287), .Z(n6338) );
  XOR U8340 ( .A(a[58]), .B(n42012), .Z(n6326) );
  XNOR U8341 ( .A(n6338), .B(n6337), .Z(n6340) );
  AND U8342 ( .A(a[60]), .B(b[0]), .Z(n6290) );
  XNOR U8343 ( .A(n6290), .B(n4071), .Z(n6292) );
  NANDN U8344 ( .A(b[0]), .B(a[59]), .Z(n6291) );
  NAND U8345 ( .A(n6292), .B(n6291), .Z(n6334) );
  XOR U8346 ( .A(a[56]), .B(n42085), .Z(n6330) );
  AND U8347 ( .A(a[52]), .B(b[7]), .Z(n6331) );
  XNOR U8348 ( .A(n6332), .B(n6331), .Z(n6333) );
  XNOR U8349 ( .A(n6334), .B(n6333), .Z(n6339) );
  XOR U8350 ( .A(n6340), .B(n6339), .Z(n6318) );
  NANDN U8351 ( .A(n6295), .B(n6294), .Z(n6299) );
  NANDN U8352 ( .A(n6297), .B(n6296), .Z(n6298) );
  AND U8353 ( .A(n6299), .B(n6298), .Z(n6317) );
  XNOR U8354 ( .A(n6318), .B(n6317), .Z(n6319) );
  NANDN U8355 ( .A(n6301), .B(n6300), .Z(n6305) );
  NAND U8356 ( .A(n6303), .B(n6302), .Z(n6304) );
  NAND U8357 ( .A(n6305), .B(n6304), .Z(n6320) );
  XNOR U8358 ( .A(n6319), .B(n6320), .Z(n6311) );
  XNOR U8359 ( .A(n6312), .B(n6311), .Z(n6313) );
  XNOR U8360 ( .A(n6314), .B(n6313), .Z(n6343) );
  XNOR U8361 ( .A(sreg[1076]), .B(n6343), .Z(n6345) );
  NANDN U8362 ( .A(sreg[1075]), .B(n6306), .Z(n6310) );
  NAND U8363 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U8364 ( .A(n6310), .B(n6309), .Z(n6344) );
  XNOR U8365 ( .A(n6345), .B(n6344), .Z(c[1076]) );
  NANDN U8366 ( .A(n6312), .B(n6311), .Z(n6316) );
  NANDN U8367 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U8368 ( .A(n6316), .B(n6315), .Z(n6351) );
  NANDN U8369 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U8370 ( .A(n6320), .B(n6319), .Z(n6321) );
  AND U8371 ( .A(n6322), .B(n6321), .Z(n6349) );
  NAND U8372 ( .A(n42143), .B(n6323), .Z(n6325) );
  XNOR U8373 ( .A(a[55]), .B(n4079), .Z(n6360) );
  NAND U8374 ( .A(n42144), .B(n6360), .Z(n6324) );
  AND U8375 ( .A(n6325), .B(n6324), .Z(n6375) );
  XOR U8376 ( .A(a[59]), .B(n42012), .Z(n6363) );
  XNOR U8377 ( .A(n6375), .B(n6374), .Z(n6377) );
  AND U8378 ( .A(a[61]), .B(b[0]), .Z(n6327) );
  XNOR U8379 ( .A(n6327), .B(n4071), .Z(n6329) );
  NANDN U8380 ( .A(b[0]), .B(a[60]), .Z(n6328) );
  NAND U8381 ( .A(n6329), .B(n6328), .Z(n6371) );
  XOR U8382 ( .A(a[57]), .B(n42085), .Z(n6367) );
  AND U8383 ( .A(a[53]), .B(b[7]), .Z(n6368) );
  XNOR U8384 ( .A(n6369), .B(n6368), .Z(n6370) );
  XNOR U8385 ( .A(n6371), .B(n6370), .Z(n6376) );
  XOR U8386 ( .A(n6377), .B(n6376), .Z(n6355) );
  NANDN U8387 ( .A(n6332), .B(n6331), .Z(n6336) );
  NANDN U8388 ( .A(n6334), .B(n6333), .Z(n6335) );
  AND U8389 ( .A(n6336), .B(n6335), .Z(n6354) );
  XNOR U8390 ( .A(n6355), .B(n6354), .Z(n6356) );
  NANDN U8391 ( .A(n6338), .B(n6337), .Z(n6342) );
  NAND U8392 ( .A(n6340), .B(n6339), .Z(n6341) );
  NAND U8393 ( .A(n6342), .B(n6341), .Z(n6357) );
  XNOR U8394 ( .A(n6356), .B(n6357), .Z(n6348) );
  XNOR U8395 ( .A(n6349), .B(n6348), .Z(n6350) );
  XNOR U8396 ( .A(n6351), .B(n6350), .Z(n6380) );
  XNOR U8397 ( .A(sreg[1077]), .B(n6380), .Z(n6382) );
  NANDN U8398 ( .A(sreg[1076]), .B(n6343), .Z(n6347) );
  NAND U8399 ( .A(n6345), .B(n6344), .Z(n6346) );
  NAND U8400 ( .A(n6347), .B(n6346), .Z(n6381) );
  XNOR U8401 ( .A(n6382), .B(n6381), .Z(c[1077]) );
  NANDN U8402 ( .A(n6349), .B(n6348), .Z(n6353) );
  NANDN U8403 ( .A(n6351), .B(n6350), .Z(n6352) );
  AND U8404 ( .A(n6353), .B(n6352), .Z(n6388) );
  NANDN U8405 ( .A(n6355), .B(n6354), .Z(n6359) );
  NANDN U8406 ( .A(n6357), .B(n6356), .Z(n6358) );
  AND U8407 ( .A(n6359), .B(n6358), .Z(n6386) );
  NAND U8408 ( .A(n42143), .B(n6360), .Z(n6362) );
  XNOR U8409 ( .A(a[56]), .B(n4079), .Z(n6397) );
  NAND U8410 ( .A(n42144), .B(n6397), .Z(n6361) );
  AND U8411 ( .A(n6362), .B(n6361), .Z(n6412) );
  XOR U8412 ( .A(a[60]), .B(n42012), .Z(n6400) );
  XNOR U8413 ( .A(n6412), .B(n6411), .Z(n6414) );
  AND U8414 ( .A(b[0]), .B(a[62]), .Z(n6364) );
  XOR U8415 ( .A(b[1]), .B(n6364), .Z(n6366) );
  NANDN U8416 ( .A(b[0]), .B(a[61]), .Z(n6365) );
  AND U8417 ( .A(n6366), .B(n6365), .Z(n6407) );
  XOR U8418 ( .A(a[58]), .B(n42085), .Z(n6404) );
  AND U8419 ( .A(a[54]), .B(b[7]), .Z(n6405) );
  XOR U8420 ( .A(n6406), .B(n6405), .Z(n6408) );
  XNOR U8421 ( .A(n6407), .B(n6408), .Z(n6413) );
  XOR U8422 ( .A(n6414), .B(n6413), .Z(n6392) );
  NANDN U8423 ( .A(n6369), .B(n6368), .Z(n6373) );
  NANDN U8424 ( .A(n6371), .B(n6370), .Z(n6372) );
  AND U8425 ( .A(n6373), .B(n6372), .Z(n6391) );
  XNOR U8426 ( .A(n6392), .B(n6391), .Z(n6393) );
  NANDN U8427 ( .A(n6375), .B(n6374), .Z(n6379) );
  NAND U8428 ( .A(n6377), .B(n6376), .Z(n6378) );
  NAND U8429 ( .A(n6379), .B(n6378), .Z(n6394) );
  XNOR U8430 ( .A(n6393), .B(n6394), .Z(n6385) );
  XNOR U8431 ( .A(n6386), .B(n6385), .Z(n6387) );
  XNOR U8432 ( .A(n6388), .B(n6387), .Z(n6417) );
  XNOR U8433 ( .A(sreg[1078]), .B(n6417), .Z(n6419) );
  NANDN U8434 ( .A(sreg[1077]), .B(n6380), .Z(n6384) );
  NAND U8435 ( .A(n6382), .B(n6381), .Z(n6383) );
  NAND U8436 ( .A(n6384), .B(n6383), .Z(n6418) );
  XNOR U8437 ( .A(n6419), .B(n6418), .Z(c[1078]) );
  NANDN U8438 ( .A(n6386), .B(n6385), .Z(n6390) );
  NANDN U8439 ( .A(n6388), .B(n6387), .Z(n6389) );
  AND U8440 ( .A(n6390), .B(n6389), .Z(n6425) );
  NANDN U8441 ( .A(n6392), .B(n6391), .Z(n6396) );
  NANDN U8442 ( .A(n6394), .B(n6393), .Z(n6395) );
  AND U8443 ( .A(n6396), .B(n6395), .Z(n6423) );
  NAND U8444 ( .A(n42143), .B(n6397), .Z(n6399) );
  XNOR U8445 ( .A(a[57]), .B(n4080), .Z(n6434) );
  NAND U8446 ( .A(n42144), .B(n6434), .Z(n6398) );
  AND U8447 ( .A(n6399), .B(n6398), .Z(n6449) );
  XOR U8448 ( .A(a[61]), .B(n42012), .Z(n6437) );
  XNOR U8449 ( .A(n6449), .B(n6448), .Z(n6451) );
  AND U8450 ( .A(a[63]), .B(b[0]), .Z(n6401) );
  XNOR U8451 ( .A(n6401), .B(n4071), .Z(n6403) );
  NANDN U8452 ( .A(b[0]), .B(a[62]), .Z(n6402) );
  NAND U8453 ( .A(n6403), .B(n6402), .Z(n6445) );
  XOR U8454 ( .A(a[59]), .B(n42085), .Z(n6438) );
  AND U8455 ( .A(a[55]), .B(b[7]), .Z(n6442) );
  XNOR U8456 ( .A(n6443), .B(n6442), .Z(n6444) );
  XNOR U8457 ( .A(n6445), .B(n6444), .Z(n6450) );
  XOR U8458 ( .A(n6451), .B(n6450), .Z(n6429) );
  NANDN U8459 ( .A(n6406), .B(n6405), .Z(n6410) );
  NANDN U8460 ( .A(n6408), .B(n6407), .Z(n6409) );
  AND U8461 ( .A(n6410), .B(n6409), .Z(n6428) );
  XNOR U8462 ( .A(n6429), .B(n6428), .Z(n6430) );
  NANDN U8463 ( .A(n6412), .B(n6411), .Z(n6416) );
  NAND U8464 ( .A(n6414), .B(n6413), .Z(n6415) );
  NAND U8465 ( .A(n6416), .B(n6415), .Z(n6431) );
  XNOR U8466 ( .A(n6430), .B(n6431), .Z(n6422) );
  XNOR U8467 ( .A(n6423), .B(n6422), .Z(n6424) );
  XNOR U8468 ( .A(n6425), .B(n6424), .Z(n6454) );
  XNOR U8469 ( .A(sreg[1079]), .B(n6454), .Z(n6456) );
  NANDN U8470 ( .A(sreg[1078]), .B(n6417), .Z(n6421) );
  NAND U8471 ( .A(n6419), .B(n6418), .Z(n6420) );
  NAND U8472 ( .A(n6421), .B(n6420), .Z(n6455) );
  XNOR U8473 ( .A(n6456), .B(n6455), .Z(c[1079]) );
  NANDN U8474 ( .A(n6423), .B(n6422), .Z(n6427) );
  NANDN U8475 ( .A(n6425), .B(n6424), .Z(n6426) );
  AND U8476 ( .A(n6427), .B(n6426), .Z(n6462) );
  NANDN U8477 ( .A(n6429), .B(n6428), .Z(n6433) );
  NANDN U8478 ( .A(n6431), .B(n6430), .Z(n6432) );
  AND U8479 ( .A(n6433), .B(n6432), .Z(n6460) );
  NAND U8480 ( .A(n42143), .B(n6434), .Z(n6436) );
  XNOR U8481 ( .A(a[58]), .B(n4080), .Z(n6471) );
  NAND U8482 ( .A(n42144), .B(n6471), .Z(n6435) );
  AND U8483 ( .A(n6436), .B(n6435), .Z(n6486) );
  XOR U8484 ( .A(a[62]), .B(n42012), .Z(n6474) );
  XNOR U8485 ( .A(n6486), .B(n6485), .Z(n6488) );
  XOR U8486 ( .A(a[60]), .B(n42085), .Z(n6478) );
  AND U8487 ( .A(a[56]), .B(b[7]), .Z(n6479) );
  XNOR U8488 ( .A(n6480), .B(n6479), .Z(n6481) );
  AND U8489 ( .A(a[64]), .B(b[0]), .Z(n6439) );
  XNOR U8490 ( .A(n6439), .B(n4071), .Z(n6441) );
  NANDN U8491 ( .A(b[0]), .B(a[63]), .Z(n6440) );
  NAND U8492 ( .A(n6441), .B(n6440), .Z(n6482) );
  XNOR U8493 ( .A(n6481), .B(n6482), .Z(n6487) );
  XOR U8494 ( .A(n6488), .B(n6487), .Z(n6466) );
  NANDN U8495 ( .A(n6443), .B(n6442), .Z(n6447) );
  NANDN U8496 ( .A(n6445), .B(n6444), .Z(n6446) );
  AND U8497 ( .A(n6447), .B(n6446), .Z(n6465) );
  XNOR U8498 ( .A(n6466), .B(n6465), .Z(n6467) );
  NANDN U8499 ( .A(n6449), .B(n6448), .Z(n6453) );
  NAND U8500 ( .A(n6451), .B(n6450), .Z(n6452) );
  NAND U8501 ( .A(n6453), .B(n6452), .Z(n6468) );
  XNOR U8502 ( .A(n6467), .B(n6468), .Z(n6459) );
  XNOR U8503 ( .A(n6460), .B(n6459), .Z(n6461) );
  XNOR U8504 ( .A(n6462), .B(n6461), .Z(n6491) );
  XNOR U8505 ( .A(sreg[1080]), .B(n6491), .Z(n6493) );
  NANDN U8506 ( .A(sreg[1079]), .B(n6454), .Z(n6458) );
  NAND U8507 ( .A(n6456), .B(n6455), .Z(n6457) );
  NAND U8508 ( .A(n6458), .B(n6457), .Z(n6492) );
  XNOR U8509 ( .A(n6493), .B(n6492), .Z(c[1080]) );
  NANDN U8510 ( .A(n6460), .B(n6459), .Z(n6464) );
  NANDN U8511 ( .A(n6462), .B(n6461), .Z(n6463) );
  AND U8512 ( .A(n6464), .B(n6463), .Z(n6499) );
  NANDN U8513 ( .A(n6466), .B(n6465), .Z(n6470) );
  NANDN U8514 ( .A(n6468), .B(n6467), .Z(n6469) );
  AND U8515 ( .A(n6470), .B(n6469), .Z(n6497) );
  NAND U8516 ( .A(n42143), .B(n6471), .Z(n6473) );
  XNOR U8517 ( .A(a[59]), .B(n4080), .Z(n6508) );
  NAND U8518 ( .A(n42144), .B(n6508), .Z(n6472) );
  AND U8519 ( .A(n6473), .B(n6472), .Z(n6523) );
  XOR U8520 ( .A(a[63]), .B(n42012), .Z(n6511) );
  XNOR U8521 ( .A(n6523), .B(n6522), .Z(n6525) );
  AND U8522 ( .A(a[65]), .B(b[0]), .Z(n6475) );
  XNOR U8523 ( .A(n6475), .B(n4071), .Z(n6477) );
  NANDN U8524 ( .A(b[0]), .B(a[64]), .Z(n6476) );
  NAND U8525 ( .A(n6477), .B(n6476), .Z(n6519) );
  XOR U8526 ( .A(a[61]), .B(n42085), .Z(n6515) );
  AND U8527 ( .A(a[57]), .B(b[7]), .Z(n6516) );
  XNOR U8528 ( .A(n6517), .B(n6516), .Z(n6518) );
  XNOR U8529 ( .A(n6519), .B(n6518), .Z(n6524) );
  XOR U8530 ( .A(n6525), .B(n6524), .Z(n6503) );
  NANDN U8531 ( .A(n6480), .B(n6479), .Z(n6484) );
  NANDN U8532 ( .A(n6482), .B(n6481), .Z(n6483) );
  AND U8533 ( .A(n6484), .B(n6483), .Z(n6502) );
  XNOR U8534 ( .A(n6503), .B(n6502), .Z(n6504) );
  NANDN U8535 ( .A(n6486), .B(n6485), .Z(n6490) );
  NAND U8536 ( .A(n6488), .B(n6487), .Z(n6489) );
  NAND U8537 ( .A(n6490), .B(n6489), .Z(n6505) );
  XNOR U8538 ( .A(n6504), .B(n6505), .Z(n6496) );
  XNOR U8539 ( .A(n6497), .B(n6496), .Z(n6498) );
  XNOR U8540 ( .A(n6499), .B(n6498), .Z(n6528) );
  XNOR U8541 ( .A(sreg[1081]), .B(n6528), .Z(n6530) );
  NANDN U8542 ( .A(sreg[1080]), .B(n6491), .Z(n6495) );
  NAND U8543 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U8544 ( .A(n6495), .B(n6494), .Z(n6529) );
  XNOR U8545 ( .A(n6530), .B(n6529), .Z(c[1081]) );
  NANDN U8546 ( .A(n6497), .B(n6496), .Z(n6501) );
  NANDN U8547 ( .A(n6499), .B(n6498), .Z(n6500) );
  AND U8548 ( .A(n6501), .B(n6500), .Z(n6536) );
  NANDN U8549 ( .A(n6503), .B(n6502), .Z(n6507) );
  NANDN U8550 ( .A(n6505), .B(n6504), .Z(n6506) );
  AND U8551 ( .A(n6507), .B(n6506), .Z(n6534) );
  NAND U8552 ( .A(n42143), .B(n6508), .Z(n6510) );
  XNOR U8553 ( .A(a[60]), .B(n4080), .Z(n6545) );
  NAND U8554 ( .A(n42144), .B(n6545), .Z(n6509) );
  AND U8555 ( .A(n6510), .B(n6509), .Z(n6560) );
  XOR U8556 ( .A(a[64]), .B(n42012), .Z(n6548) );
  XNOR U8557 ( .A(n6560), .B(n6559), .Z(n6562) );
  AND U8558 ( .A(a[66]), .B(b[0]), .Z(n6512) );
  XNOR U8559 ( .A(n6512), .B(n4071), .Z(n6514) );
  NANDN U8560 ( .A(b[0]), .B(a[65]), .Z(n6513) );
  NAND U8561 ( .A(n6514), .B(n6513), .Z(n6556) );
  XOR U8562 ( .A(a[62]), .B(n42085), .Z(n6552) );
  AND U8563 ( .A(a[58]), .B(b[7]), .Z(n6553) );
  XNOR U8564 ( .A(n6554), .B(n6553), .Z(n6555) );
  XNOR U8565 ( .A(n6556), .B(n6555), .Z(n6561) );
  XOR U8566 ( .A(n6562), .B(n6561), .Z(n6540) );
  NANDN U8567 ( .A(n6517), .B(n6516), .Z(n6521) );
  NANDN U8568 ( .A(n6519), .B(n6518), .Z(n6520) );
  AND U8569 ( .A(n6521), .B(n6520), .Z(n6539) );
  XNOR U8570 ( .A(n6540), .B(n6539), .Z(n6541) );
  NANDN U8571 ( .A(n6523), .B(n6522), .Z(n6527) );
  NAND U8572 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U8573 ( .A(n6527), .B(n6526), .Z(n6542) );
  XNOR U8574 ( .A(n6541), .B(n6542), .Z(n6533) );
  XNOR U8575 ( .A(n6534), .B(n6533), .Z(n6535) );
  XNOR U8576 ( .A(n6536), .B(n6535), .Z(n6565) );
  XNOR U8577 ( .A(sreg[1082]), .B(n6565), .Z(n6567) );
  NANDN U8578 ( .A(sreg[1081]), .B(n6528), .Z(n6532) );
  NAND U8579 ( .A(n6530), .B(n6529), .Z(n6531) );
  NAND U8580 ( .A(n6532), .B(n6531), .Z(n6566) );
  XNOR U8581 ( .A(n6567), .B(n6566), .Z(c[1082]) );
  NANDN U8582 ( .A(n6534), .B(n6533), .Z(n6538) );
  NANDN U8583 ( .A(n6536), .B(n6535), .Z(n6537) );
  AND U8584 ( .A(n6538), .B(n6537), .Z(n6573) );
  NANDN U8585 ( .A(n6540), .B(n6539), .Z(n6544) );
  NANDN U8586 ( .A(n6542), .B(n6541), .Z(n6543) );
  AND U8587 ( .A(n6544), .B(n6543), .Z(n6571) );
  NAND U8588 ( .A(n42143), .B(n6545), .Z(n6547) );
  XNOR U8589 ( .A(a[61]), .B(n4080), .Z(n6582) );
  NAND U8590 ( .A(n42144), .B(n6582), .Z(n6546) );
  AND U8591 ( .A(n6547), .B(n6546), .Z(n6597) );
  XOR U8592 ( .A(a[65]), .B(n42012), .Z(n6585) );
  XNOR U8593 ( .A(n6597), .B(n6596), .Z(n6599) );
  AND U8594 ( .A(a[67]), .B(b[0]), .Z(n6549) );
  XNOR U8595 ( .A(n6549), .B(n4071), .Z(n6551) );
  NANDN U8596 ( .A(b[0]), .B(a[66]), .Z(n6550) );
  NAND U8597 ( .A(n6551), .B(n6550), .Z(n6593) );
  XOR U8598 ( .A(a[63]), .B(n42085), .Z(n6589) );
  AND U8599 ( .A(a[59]), .B(b[7]), .Z(n6590) );
  XNOR U8600 ( .A(n6591), .B(n6590), .Z(n6592) );
  XNOR U8601 ( .A(n6593), .B(n6592), .Z(n6598) );
  XOR U8602 ( .A(n6599), .B(n6598), .Z(n6577) );
  NANDN U8603 ( .A(n6554), .B(n6553), .Z(n6558) );
  NANDN U8604 ( .A(n6556), .B(n6555), .Z(n6557) );
  AND U8605 ( .A(n6558), .B(n6557), .Z(n6576) );
  XNOR U8606 ( .A(n6577), .B(n6576), .Z(n6578) );
  NANDN U8607 ( .A(n6560), .B(n6559), .Z(n6564) );
  NAND U8608 ( .A(n6562), .B(n6561), .Z(n6563) );
  NAND U8609 ( .A(n6564), .B(n6563), .Z(n6579) );
  XNOR U8610 ( .A(n6578), .B(n6579), .Z(n6570) );
  XNOR U8611 ( .A(n6571), .B(n6570), .Z(n6572) );
  XNOR U8612 ( .A(n6573), .B(n6572), .Z(n6602) );
  XNOR U8613 ( .A(sreg[1083]), .B(n6602), .Z(n6604) );
  NANDN U8614 ( .A(sreg[1082]), .B(n6565), .Z(n6569) );
  NAND U8615 ( .A(n6567), .B(n6566), .Z(n6568) );
  NAND U8616 ( .A(n6569), .B(n6568), .Z(n6603) );
  XNOR U8617 ( .A(n6604), .B(n6603), .Z(c[1083]) );
  NANDN U8618 ( .A(n6571), .B(n6570), .Z(n6575) );
  NANDN U8619 ( .A(n6573), .B(n6572), .Z(n6574) );
  AND U8620 ( .A(n6575), .B(n6574), .Z(n6610) );
  NANDN U8621 ( .A(n6577), .B(n6576), .Z(n6581) );
  NANDN U8622 ( .A(n6579), .B(n6578), .Z(n6580) );
  AND U8623 ( .A(n6581), .B(n6580), .Z(n6608) );
  NAND U8624 ( .A(n42143), .B(n6582), .Z(n6584) );
  XNOR U8625 ( .A(a[62]), .B(n4080), .Z(n6619) );
  NAND U8626 ( .A(n42144), .B(n6619), .Z(n6583) );
  AND U8627 ( .A(n6584), .B(n6583), .Z(n6634) );
  XOR U8628 ( .A(a[66]), .B(n42012), .Z(n6622) );
  XNOR U8629 ( .A(n6634), .B(n6633), .Z(n6636) );
  AND U8630 ( .A(a[68]), .B(b[0]), .Z(n6586) );
  XNOR U8631 ( .A(n6586), .B(n4071), .Z(n6588) );
  NANDN U8632 ( .A(b[0]), .B(a[67]), .Z(n6587) );
  NAND U8633 ( .A(n6588), .B(n6587), .Z(n6630) );
  XOR U8634 ( .A(a[64]), .B(n42085), .Z(n6626) );
  AND U8635 ( .A(a[60]), .B(b[7]), .Z(n6627) );
  XNOR U8636 ( .A(n6628), .B(n6627), .Z(n6629) );
  XNOR U8637 ( .A(n6630), .B(n6629), .Z(n6635) );
  XOR U8638 ( .A(n6636), .B(n6635), .Z(n6614) );
  NANDN U8639 ( .A(n6591), .B(n6590), .Z(n6595) );
  NANDN U8640 ( .A(n6593), .B(n6592), .Z(n6594) );
  AND U8641 ( .A(n6595), .B(n6594), .Z(n6613) );
  XNOR U8642 ( .A(n6614), .B(n6613), .Z(n6615) );
  NANDN U8643 ( .A(n6597), .B(n6596), .Z(n6601) );
  NAND U8644 ( .A(n6599), .B(n6598), .Z(n6600) );
  NAND U8645 ( .A(n6601), .B(n6600), .Z(n6616) );
  XNOR U8646 ( .A(n6615), .B(n6616), .Z(n6607) );
  XNOR U8647 ( .A(n6608), .B(n6607), .Z(n6609) );
  XNOR U8648 ( .A(n6610), .B(n6609), .Z(n6639) );
  XNOR U8649 ( .A(sreg[1084]), .B(n6639), .Z(n6641) );
  NANDN U8650 ( .A(sreg[1083]), .B(n6602), .Z(n6606) );
  NAND U8651 ( .A(n6604), .B(n6603), .Z(n6605) );
  NAND U8652 ( .A(n6606), .B(n6605), .Z(n6640) );
  XNOR U8653 ( .A(n6641), .B(n6640), .Z(c[1084]) );
  NANDN U8654 ( .A(n6608), .B(n6607), .Z(n6612) );
  NANDN U8655 ( .A(n6610), .B(n6609), .Z(n6611) );
  AND U8656 ( .A(n6612), .B(n6611), .Z(n6647) );
  NANDN U8657 ( .A(n6614), .B(n6613), .Z(n6618) );
  NANDN U8658 ( .A(n6616), .B(n6615), .Z(n6617) );
  AND U8659 ( .A(n6618), .B(n6617), .Z(n6645) );
  NAND U8660 ( .A(n42143), .B(n6619), .Z(n6621) );
  XNOR U8661 ( .A(a[63]), .B(n4080), .Z(n6656) );
  NAND U8662 ( .A(n42144), .B(n6656), .Z(n6620) );
  AND U8663 ( .A(n6621), .B(n6620), .Z(n6671) );
  XOR U8664 ( .A(a[67]), .B(n42012), .Z(n6659) );
  XNOR U8665 ( .A(n6671), .B(n6670), .Z(n6673) );
  AND U8666 ( .A(a[69]), .B(b[0]), .Z(n6623) );
  XNOR U8667 ( .A(n6623), .B(n4071), .Z(n6625) );
  NANDN U8668 ( .A(b[0]), .B(a[68]), .Z(n6624) );
  NAND U8669 ( .A(n6625), .B(n6624), .Z(n6667) );
  XOR U8670 ( .A(a[65]), .B(n42085), .Z(n6663) );
  AND U8671 ( .A(a[61]), .B(b[7]), .Z(n6664) );
  XNOR U8672 ( .A(n6665), .B(n6664), .Z(n6666) );
  XNOR U8673 ( .A(n6667), .B(n6666), .Z(n6672) );
  XOR U8674 ( .A(n6673), .B(n6672), .Z(n6651) );
  NANDN U8675 ( .A(n6628), .B(n6627), .Z(n6632) );
  NANDN U8676 ( .A(n6630), .B(n6629), .Z(n6631) );
  AND U8677 ( .A(n6632), .B(n6631), .Z(n6650) );
  XNOR U8678 ( .A(n6651), .B(n6650), .Z(n6652) );
  NANDN U8679 ( .A(n6634), .B(n6633), .Z(n6638) );
  NAND U8680 ( .A(n6636), .B(n6635), .Z(n6637) );
  NAND U8681 ( .A(n6638), .B(n6637), .Z(n6653) );
  XNOR U8682 ( .A(n6652), .B(n6653), .Z(n6644) );
  XNOR U8683 ( .A(n6645), .B(n6644), .Z(n6646) );
  XNOR U8684 ( .A(n6647), .B(n6646), .Z(n6676) );
  XNOR U8685 ( .A(sreg[1085]), .B(n6676), .Z(n6678) );
  NANDN U8686 ( .A(sreg[1084]), .B(n6639), .Z(n6643) );
  NAND U8687 ( .A(n6641), .B(n6640), .Z(n6642) );
  NAND U8688 ( .A(n6643), .B(n6642), .Z(n6677) );
  XNOR U8689 ( .A(n6678), .B(n6677), .Z(c[1085]) );
  NANDN U8690 ( .A(n6645), .B(n6644), .Z(n6649) );
  NANDN U8691 ( .A(n6647), .B(n6646), .Z(n6648) );
  AND U8692 ( .A(n6649), .B(n6648), .Z(n6684) );
  NANDN U8693 ( .A(n6651), .B(n6650), .Z(n6655) );
  NANDN U8694 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U8695 ( .A(n6655), .B(n6654), .Z(n6682) );
  NAND U8696 ( .A(n42143), .B(n6656), .Z(n6658) );
  XNOR U8697 ( .A(a[64]), .B(n4081), .Z(n6693) );
  NAND U8698 ( .A(n42144), .B(n6693), .Z(n6657) );
  AND U8699 ( .A(n6658), .B(n6657), .Z(n6708) );
  XOR U8700 ( .A(a[68]), .B(n42012), .Z(n6696) );
  XNOR U8701 ( .A(n6708), .B(n6707), .Z(n6710) );
  AND U8702 ( .A(a[70]), .B(b[0]), .Z(n6660) );
  XNOR U8703 ( .A(n6660), .B(n4071), .Z(n6662) );
  NANDN U8704 ( .A(b[0]), .B(a[69]), .Z(n6661) );
  NAND U8705 ( .A(n6662), .B(n6661), .Z(n6704) );
  XOR U8706 ( .A(a[66]), .B(n42085), .Z(n6700) );
  AND U8707 ( .A(a[62]), .B(b[7]), .Z(n6701) );
  XNOR U8708 ( .A(n6702), .B(n6701), .Z(n6703) );
  XNOR U8709 ( .A(n6704), .B(n6703), .Z(n6709) );
  XOR U8710 ( .A(n6710), .B(n6709), .Z(n6688) );
  NANDN U8711 ( .A(n6665), .B(n6664), .Z(n6669) );
  NANDN U8712 ( .A(n6667), .B(n6666), .Z(n6668) );
  AND U8713 ( .A(n6669), .B(n6668), .Z(n6687) );
  XNOR U8714 ( .A(n6688), .B(n6687), .Z(n6689) );
  NANDN U8715 ( .A(n6671), .B(n6670), .Z(n6675) );
  NAND U8716 ( .A(n6673), .B(n6672), .Z(n6674) );
  NAND U8717 ( .A(n6675), .B(n6674), .Z(n6690) );
  XNOR U8718 ( .A(n6689), .B(n6690), .Z(n6681) );
  XNOR U8719 ( .A(n6682), .B(n6681), .Z(n6683) );
  XNOR U8720 ( .A(n6684), .B(n6683), .Z(n6713) );
  XNOR U8721 ( .A(sreg[1086]), .B(n6713), .Z(n6715) );
  NANDN U8722 ( .A(sreg[1085]), .B(n6676), .Z(n6680) );
  NAND U8723 ( .A(n6678), .B(n6677), .Z(n6679) );
  NAND U8724 ( .A(n6680), .B(n6679), .Z(n6714) );
  XNOR U8725 ( .A(n6715), .B(n6714), .Z(c[1086]) );
  NANDN U8726 ( .A(n6682), .B(n6681), .Z(n6686) );
  NANDN U8727 ( .A(n6684), .B(n6683), .Z(n6685) );
  AND U8728 ( .A(n6686), .B(n6685), .Z(n6721) );
  NANDN U8729 ( .A(n6688), .B(n6687), .Z(n6692) );
  NANDN U8730 ( .A(n6690), .B(n6689), .Z(n6691) );
  AND U8731 ( .A(n6692), .B(n6691), .Z(n6719) );
  NAND U8732 ( .A(n42143), .B(n6693), .Z(n6695) );
  XNOR U8733 ( .A(a[65]), .B(n4081), .Z(n6730) );
  NAND U8734 ( .A(n42144), .B(n6730), .Z(n6694) );
  AND U8735 ( .A(n6695), .B(n6694), .Z(n6745) );
  XOR U8736 ( .A(a[69]), .B(n42012), .Z(n6733) );
  XNOR U8737 ( .A(n6745), .B(n6744), .Z(n6747) );
  AND U8738 ( .A(a[71]), .B(b[0]), .Z(n6697) );
  XNOR U8739 ( .A(n6697), .B(n4071), .Z(n6699) );
  NANDN U8740 ( .A(b[0]), .B(a[70]), .Z(n6698) );
  NAND U8741 ( .A(n6699), .B(n6698), .Z(n6741) );
  XOR U8742 ( .A(a[67]), .B(n42085), .Z(n6734) );
  AND U8743 ( .A(a[63]), .B(b[7]), .Z(n6738) );
  XNOR U8744 ( .A(n6739), .B(n6738), .Z(n6740) );
  XNOR U8745 ( .A(n6741), .B(n6740), .Z(n6746) );
  XOR U8746 ( .A(n6747), .B(n6746), .Z(n6725) );
  NANDN U8747 ( .A(n6702), .B(n6701), .Z(n6706) );
  NANDN U8748 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U8749 ( .A(n6706), .B(n6705), .Z(n6724) );
  XNOR U8750 ( .A(n6725), .B(n6724), .Z(n6726) );
  NANDN U8751 ( .A(n6708), .B(n6707), .Z(n6712) );
  NAND U8752 ( .A(n6710), .B(n6709), .Z(n6711) );
  NAND U8753 ( .A(n6712), .B(n6711), .Z(n6727) );
  XNOR U8754 ( .A(n6726), .B(n6727), .Z(n6718) );
  XNOR U8755 ( .A(n6719), .B(n6718), .Z(n6720) );
  XNOR U8756 ( .A(n6721), .B(n6720), .Z(n6750) );
  XNOR U8757 ( .A(sreg[1087]), .B(n6750), .Z(n6752) );
  NANDN U8758 ( .A(sreg[1086]), .B(n6713), .Z(n6717) );
  NAND U8759 ( .A(n6715), .B(n6714), .Z(n6716) );
  NAND U8760 ( .A(n6717), .B(n6716), .Z(n6751) );
  XNOR U8761 ( .A(n6752), .B(n6751), .Z(c[1087]) );
  NANDN U8762 ( .A(n6719), .B(n6718), .Z(n6723) );
  NANDN U8763 ( .A(n6721), .B(n6720), .Z(n6722) );
  AND U8764 ( .A(n6723), .B(n6722), .Z(n6758) );
  NANDN U8765 ( .A(n6725), .B(n6724), .Z(n6729) );
  NANDN U8766 ( .A(n6727), .B(n6726), .Z(n6728) );
  AND U8767 ( .A(n6729), .B(n6728), .Z(n6756) );
  NAND U8768 ( .A(n42143), .B(n6730), .Z(n6732) );
  XNOR U8769 ( .A(a[66]), .B(n4081), .Z(n6767) );
  NAND U8770 ( .A(n42144), .B(n6767), .Z(n6731) );
  AND U8771 ( .A(n6732), .B(n6731), .Z(n6782) );
  XOR U8772 ( .A(a[70]), .B(n42012), .Z(n6770) );
  XNOR U8773 ( .A(n6782), .B(n6781), .Z(n6784) );
  XOR U8774 ( .A(a[68]), .B(n42085), .Z(n6774) );
  AND U8775 ( .A(a[64]), .B(b[7]), .Z(n6775) );
  XNOR U8776 ( .A(n6776), .B(n6775), .Z(n6777) );
  AND U8777 ( .A(a[72]), .B(b[0]), .Z(n6735) );
  XNOR U8778 ( .A(n6735), .B(n4071), .Z(n6737) );
  NANDN U8779 ( .A(b[0]), .B(a[71]), .Z(n6736) );
  NAND U8780 ( .A(n6737), .B(n6736), .Z(n6778) );
  XNOR U8781 ( .A(n6777), .B(n6778), .Z(n6783) );
  XOR U8782 ( .A(n6784), .B(n6783), .Z(n6762) );
  NANDN U8783 ( .A(n6739), .B(n6738), .Z(n6743) );
  NANDN U8784 ( .A(n6741), .B(n6740), .Z(n6742) );
  AND U8785 ( .A(n6743), .B(n6742), .Z(n6761) );
  XNOR U8786 ( .A(n6762), .B(n6761), .Z(n6763) );
  NANDN U8787 ( .A(n6745), .B(n6744), .Z(n6749) );
  NAND U8788 ( .A(n6747), .B(n6746), .Z(n6748) );
  NAND U8789 ( .A(n6749), .B(n6748), .Z(n6764) );
  XNOR U8790 ( .A(n6763), .B(n6764), .Z(n6755) );
  XNOR U8791 ( .A(n6756), .B(n6755), .Z(n6757) );
  XNOR U8792 ( .A(n6758), .B(n6757), .Z(n6787) );
  XNOR U8793 ( .A(sreg[1088]), .B(n6787), .Z(n6789) );
  NANDN U8794 ( .A(sreg[1087]), .B(n6750), .Z(n6754) );
  NAND U8795 ( .A(n6752), .B(n6751), .Z(n6753) );
  NAND U8796 ( .A(n6754), .B(n6753), .Z(n6788) );
  XNOR U8797 ( .A(n6789), .B(n6788), .Z(c[1088]) );
  NANDN U8798 ( .A(n6756), .B(n6755), .Z(n6760) );
  NANDN U8799 ( .A(n6758), .B(n6757), .Z(n6759) );
  AND U8800 ( .A(n6760), .B(n6759), .Z(n6795) );
  NANDN U8801 ( .A(n6762), .B(n6761), .Z(n6766) );
  NANDN U8802 ( .A(n6764), .B(n6763), .Z(n6765) );
  AND U8803 ( .A(n6766), .B(n6765), .Z(n6793) );
  NAND U8804 ( .A(n42143), .B(n6767), .Z(n6769) );
  XNOR U8805 ( .A(a[67]), .B(n4081), .Z(n6804) );
  NAND U8806 ( .A(n42144), .B(n6804), .Z(n6768) );
  AND U8807 ( .A(n6769), .B(n6768), .Z(n6819) );
  XOR U8808 ( .A(a[71]), .B(n42012), .Z(n6807) );
  XNOR U8809 ( .A(n6819), .B(n6818), .Z(n6821) );
  AND U8810 ( .A(a[73]), .B(b[0]), .Z(n6771) );
  XNOR U8811 ( .A(n6771), .B(n4071), .Z(n6773) );
  NANDN U8812 ( .A(b[0]), .B(a[72]), .Z(n6772) );
  NAND U8813 ( .A(n6773), .B(n6772), .Z(n6815) );
  XOR U8814 ( .A(a[69]), .B(n42085), .Z(n6811) );
  AND U8815 ( .A(a[65]), .B(b[7]), .Z(n6812) );
  XNOR U8816 ( .A(n6813), .B(n6812), .Z(n6814) );
  XNOR U8817 ( .A(n6815), .B(n6814), .Z(n6820) );
  XOR U8818 ( .A(n6821), .B(n6820), .Z(n6799) );
  NANDN U8819 ( .A(n6776), .B(n6775), .Z(n6780) );
  NANDN U8820 ( .A(n6778), .B(n6777), .Z(n6779) );
  AND U8821 ( .A(n6780), .B(n6779), .Z(n6798) );
  XNOR U8822 ( .A(n6799), .B(n6798), .Z(n6800) );
  NANDN U8823 ( .A(n6782), .B(n6781), .Z(n6786) );
  NAND U8824 ( .A(n6784), .B(n6783), .Z(n6785) );
  NAND U8825 ( .A(n6786), .B(n6785), .Z(n6801) );
  XNOR U8826 ( .A(n6800), .B(n6801), .Z(n6792) );
  XNOR U8827 ( .A(n6793), .B(n6792), .Z(n6794) );
  XNOR U8828 ( .A(n6795), .B(n6794), .Z(n6824) );
  XNOR U8829 ( .A(sreg[1089]), .B(n6824), .Z(n6826) );
  NANDN U8830 ( .A(sreg[1088]), .B(n6787), .Z(n6791) );
  NAND U8831 ( .A(n6789), .B(n6788), .Z(n6790) );
  NAND U8832 ( .A(n6791), .B(n6790), .Z(n6825) );
  XNOR U8833 ( .A(n6826), .B(n6825), .Z(c[1089]) );
  NANDN U8834 ( .A(n6793), .B(n6792), .Z(n6797) );
  NANDN U8835 ( .A(n6795), .B(n6794), .Z(n6796) );
  AND U8836 ( .A(n6797), .B(n6796), .Z(n6832) );
  NANDN U8837 ( .A(n6799), .B(n6798), .Z(n6803) );
  NANDN U8838 ( .A(n6801), .B(n6800), .Z(n6802) );
  AND U8839 ( .A(n6803), .B(n6802), .Z(n6830) );
  NAND U8840 ( .A(n42143), .B(n6804), .Z(n6806) );
  XNOR U8841 ( .A(a[68]), .B(n4081), .Z(n6841) );
  NAND U8842 ( .A(n42144), .B(n6841), .Z(n6805) );
  AND U8843 ( .A(n6806), .B(n6805), .Z(n6856) );
  XOR U8844 ( .A(a[72]), .B(n42012), .Z(n6844) );
  XNOR U8845 ( .A(n6856), .B(n6855), .Z(n6858) );
  AND U8846 ( .A(a[74]), .B(b[0]), .Z(n6808) );
  XNOR U8847 ( .A(n6808), .B(n4071), .Z(n6810) );
  NANDN U8848 ( .A(b[0]), .B(a[73]), .Z(n6809) );
  NAND U8849 ( .A(n6810), .B(n6809), .Z(n6852) );
  XOR U8850 ( .A(a[70]), .B(n42085), .Z(n6845) );
  AND U8851 ( .A(a[66]), .B(b[7]), .Z(n6849) );
  XNOR U8852 ( .A(n6850), .B(n6849), .Z(n6851) );
  XNOR U8853 ( .A(n6852), .B(n6851), .Z(n6857) );
  XOR U8854 ( .A(n6858), .B(n6857), .Z(n6836) );
  NANDN U8855 ( .A(n6813), .B(n6812), .Z(n6817) );
  NANDN U8856 ( .A(n6815), .B(n6814), .Z(n6816) );
  AND U8857 ( .A(n6817), .B(n6816), .Z(n6835) );
  XNOR U8858 ( .A(n6836), .B(n6835), .Z(n6837) );
  NANDN U8859 ( .A(n6819), .B(n6818), .Z(n6823) );
  NAND U8860 ( .A(n6821), .B(n6820), .Z(n6822) );
  NAND U8861 ( .A(n6823), .B(n6822), .Z(n6838) );
  XNOR U8862 ( .A(n6837), .B(n6838), .Z(n6829) );
  XNOR U8863 ( .A(n6830), .B(n6829), .Z(n6831) );
  XNOR U8864 ( .A(n6832), .B(n6831), .Z(n6861) );
  XNOR U8865 ( .A(sreg[1090]), .B(n6861), .Z(n6863) );
  NANDN U8866 ( .A(sreg[1089]), .B(n6824), .Z(n6828) );
  NAND U8867 ( .A(n6826), .B(n6825), .Z(n6827) );
  NAND U8868 ( .A(n6828), .B(n6827), .Z(n6862) );
  XNOR U8869 ( .A(n6863), .B(n6862), .Z(c[1090]) );
  NANDN U8870 ( .A(n6830), .B(n6829), .Z(n6834) );
  NANDN U8871 ( .A(n6832), .B(n6831), .Z(n6833) );
  AND U8872 ( .A(n6834), .B(n6833), .Z(n6869) );
  NANDN U8873 ( .A(n6836), .B(n6835), .Z(n6840) );
  NANDN U8874 ( .A(n6838), .B(n6837), .Z(n6839) );
  AND U8875 ( .A(n6840), .B(n6839), .Z(n6867) );
  NAND U8876 ( .A(n42143), .B(n6841), .Z(n6843) );
  XNOR U8877 ( .A(a[69]), .B(n4081), .Z(n6878) );
  NAND U8878 ( .A(n42144), .B(n6878), .Z(n6842) );
  AND U8879 ( .A(n6843), .B(n6842), .Z(n6893) );
  XOR U8880 ( .A(a[73]), .B(n42012), .Z(n6881) );
  XNOR U8881 ( .A(n6893), .B(n6892), .Z(n6895) );
  XOR U8882 ( .A(a[71]), .B(n42085), .Z(n6885) );
  AND U8883 ( .A(a[67]), .B(b[7]), .Z(n6886) );
  XNOR U8884 ( .A(n6887), .B(n6886), .Z(n6888) );
  AND U8885 ( .A(a[75]), .B(b[0]), .Z(n6846) );
  XNOR U8886 ( .A(n6846), .B(n4071), .Z(n6848) );
  NANDN U8887 ( .A(b[0]), .B(a[74]), .Z(n6847) );
  NAND U8888 ( .A(n6848), .B(n6847), .Z(n6889) );
  XNOR U8889 ( .A(n6888), .B(n6889), .Z(n6894) );
  XOR U8890 ( .A(n6895), .B(n6894), .Z(n6873) );
  NANDN U8891 ( .A(n6850), .B(n6849), .Z(n6854) );
  NANDN U8892 ( .A(n6852), .B(n6851), .Z(n6853) );
  AND U8893 ( .A(n6854), .B(n6853), .Z(n6872) );
  XNOR U8894 ( .A(n6873), .B(n6872), .Z(n6874) );
  NANDN U8895 ( .A(n6856), .B(n6855), .Z(n6860) );
  NAND U8896 ( .A(n6858), .B(n6857), .Z(n6859) );
  NAND U8897 ( .A(n6860), .B(n6859), .Z(n6875) );
  XNOR U8898 ( .A(n6874), .B(n6875), .Z(n6866) );
  XNOR U8899 ( .A(n6867), .B(n6866), .Z(n6868) );
  XNOR U8900 ( .A(n6869), .B(n6868), .Z(n6898) );
  XNOR U8901 ( .A(sreg[1091]), .B(n6898), .Z(n6900) );
  NANDN U8902 ( .A(sreg[1090]), .B(n6861), .Z(n6865) );
  NAND U8903 ( .A(n6863), .B(n6862), .Z(n6864) );
  NAND U8904 ( .A(n6865), .B(n6864), .Z(n6899) );
  XNOR U8905 ( .A(n6900), .B(n6899), .Z(c[1091]) );
  NANDN U8906 ( .A(n6867), .B(n6866), .Z(n6871) );
  NANDN U8907 ( .A(n6869), .B(n6868), .Z(n6870) );
  AND U8908 ( .A(n6871), .B(n6870), .Z(n6910) );
  NANDN U8909 ( .A(n6873), .B(n6872), .Z(n6877) );
  NANDN U8910 ( .A(n6875), .B(n6874), .Z(n6876) );
  AND U8911 ( .A(n6877), .B(n6876), .Z(n6909) );
  NAND U8912 ( .A(n42143), .B(n6878), .Z(n6880) );
  XNOR U8913 ( .A(a[70]), .B(n4081), .Z(n6920) );
  NAND U8914 ( .A(n42144), .B(n6920), .Z(n6879) );
  AND U8915 ( .A(n6880), .B(n6879), .Z(n6935) );
  XOR U8916 ( .A(a[74]), .B(n42012), .Z(n6923) );
  XNOR U8917 ( .A(n6935), .B(n6934), .Z(n6937) );
  AND U8918 ( .A(a[76]), .B(b[0]), .Z(n6882) );
  XNOR U8919 ( .A(n6882), .B(n4071), .Z(n6884) );
  NANDN U8920 ( .A(b[0]), .B(a[75]), .Z(n6883) );
  NAND U8921 ( .A(n6884), .B(n6883), .Z(n6931) );
  XOR U8922 ( .A(a[72]), .B(n42085), .Z(n6924) );
  AND U8923 ( .A(a[68]), .B(b[7]), .Z(n6928) );
  XNOR U8924 ( .A(n6929), .B(n6928), .Z(n6930) );
  XNOR U8925 ( .A(n6931), .B(n6930), .Z(n6936) );
  XOR U8926 ( .A(n6937), .B(n6936), .Z(n6915) );
  NANDN U8927 ( .A(n6887), .B(n6886), .Z(n6891) );
  NANDN U8928 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U8929 ( .A(n6891), .B(n6890), .Z(n6914) );
  XNOR U8930 ( .A(n6915), .B(n6914), .Z(n6916) );
  NANDN U8931 ( .A(n6893), .B(n6892), .Z(n6897) );
  NAND U8932 ( .A(n6895), .B(n6894), .Z(n6896) );
  NAND U8933 ( .A(n6897), .B(n6896), .Z(n6917) );
  XNOR U8934 ( .A(n6916), .B(n6917), .Z(n6908) );
  XOR U8935 ( .A(n6909), .B(n6908), .Z(n6911) );
  XOR U8936 ( .A(n6910), .B(n6911), .Z(n6903) );
  XNOR U8937 ( .A(n6903), .B(sreg[1092]), .Z(n6905) );
  NANDN U8938 ( .A(sreg[1091]), .B(n6898), .Z(n6902) );
  NAND U8939 ( .A(n6900), .B(n6899), .Z(n6901) );
  AND U8940 ( .A(n6902), .B(n6901), .Z(n6904) );
  XOR U8941 ( .A(n6905), .B(n6904), .Z(c[1092]) );
  NANDN U8942 ( .A(n6903), .B(sreg[1092]), .Z(n6907) );
  NAND U8943 ( .A(n6905), .B(n6904), .Z(n6906) );
  AND U8944 ( .A(n6907), .B(n6906), .Z(n6974) );
  NANDN U8945 ( .A(n6909), .B(n6908), .Z(n6913) );
  OR U8946 ( .A(n6911), .B(n6910), .Z(n6912) );
  AND U8947 ( .A(n6913), .B(n6912), .Z(n6943) );
  NANDN U8948 ( .A(n6915), .B(n6914), .Z(n6919) );
  NANDN U8949 ( .A(n6917), .B(n6916), .Z(n6918) );
  AND U8950 ( .A(n6919), .B(n6918), .Z(n6941) );
  NAND U8951 ( .A(n42143), .B(n6920), .Z(n6922) );
  XNOR U8952 ( .A(a[71]), .B(n4082), .Z(n6952) );
  NAND U8953 ( .A(n42144), .B(n6952), .Z(n6921) );
  AND U8954 ( .A(n6922), .B(n6921), .Z(n6967) );
  XOR U8955 ( .A(a[75]), .B(n42012), .Z(n6955) );
  XNOR U8956 ( .A(n6967), .B(n6966), .Z(n6969) );
  XOR U8957 ( .A(a[73]), .B(n42085), .Z(n6959) );
  AND U8958 ( .A(a[69]), .B(b[7]), .Z(n6960) );
  XNOR U8959 ( .A(n6961), .B(n6960), .Z(n6962) );
  AND U8960 ( .A(a[77]), .B(b[0]), .Z(n6925) );
  XNOR U8961 ( .A(n6925), .B(n4071), .Z(n6927) );
  NANDN U8962 ( .A(b[0]), .B(a[76]), .Z(n6926) );
  NAND U8963 ( .A(n6927), .B(n6926), .Z(n6963) );
  XNOR U8964 ( .A(n6962), .B(n6963), .Z(n6968) );
  XOR U8965 ( .A(n6969), .B(n6968), .Z(n6947) );
  NANDN U8966 ( .A(n6929), .B(n6928), .Z(n6933) );
  NANDN U8967 ( .A(n6931), .B(n6930), .Z(n6932) );
  AND U8968 ( .A(n6933), .B(n6932), .Z(n6946) );
  XNOR U8969 ( .A(n6947), .B(n6946), .Z(n6948) );
  NANDN U8970 ( .A(n6935), .B(n6934), .Z(n6939) );
  NAND U8971 ( .A(n6937), .B(n6936), .Z(n6938) );
  NAND U8972 ( .A(n6939), .B(n6938), .Z(n6949) );
  XNOR U8973 ( .A(n6948), .B(n6949), .Z(n6940) );
  XNOR U8974 ( .A(n6941), .B(n6940), .Z(n6942) );
  XNOR U8975 ( .A(n6943), .B(n6942), .Z(n6972) );
  XNOR U8976 ( .A(sreg[1093]), .B(n6972), .Z(n6973) );
  XNOR U8977 ( .A(n6974), .B(n6973), .Z(c[1093]) );
  NANDN U8978 ( .A(n6941), .B(n6940), .Z(n6945) );
  NANDN U8979 ( .A(n6943), .B(n6942), .Z(n6944) );
  AND U8980 ( .A(n6945), .B(n6944), .Z(n6980) );
  NANDN U8981 ( .A(n6947), .B(n6946), .Z(n6951) );
  NANDN U8982 ( .A(n6949), .B(n6948), .Z(n6950) );
  AND U8983 ( .A(n6951), .B(n6950), .Z(n6978) );
  NAND U8984 ( .A(n42143), .B(n6952), .Z(n6954) );
  XNOR U8985 ( .A(a[72]), .B(n4082), .Z(n6989) );
  NAND U8986 ( .A(n42144), .B(n6989), .Z(n6953) );
  AND U8987 ( .A(n6954), .B(n6953), .Z(n7004) );
  XOR U8988 ( .A(a[76]), .B(n42012), .Z(n6992) );
  XNOR U8989 ( .A(n7004), .B(n7003), .Z(n7006) );
  AND U8990 ( .A(a[78]), .B(b[0]), .Z(n6956) );
  XNOR U8991 ( .A(n6956), .B(n4071), .Z(n6958) );
  NANDN U8992 ( .A(b[0]), .B(a[77]), .Z(n6957) );
  NAND U8993 ( .A(n6958), .B(n6957), .Z(n7000) );
  XOR U8994 ( .A(a[74]), .B(n42085), .Z(n6996) );
  AND U8995 ( .A(a[70]), .B(b[7]), .Z(n6997) );
  XNOR U8996 ( .A(n6998), .B(n6997), .Z(n6999) );
  XNOR U8997 ( .A(n7000), .B(n6999), .Z(n7005) );
  XOR U8998 ( .A(n7006), .B(n7005), .Z(n6984) );
  NANDN U8999 ( .A(n6961), .B(n6960), .Z(n6965) );
  NANDN U9000 ( .A(n6963), .B(n6962), .Z(n6964) );
  AND U9001 ( .A(n6965), .B(n6964), .Z(n6983) );
  XNOR U9002 ( .A(n6984), .B(n6983), .Z(n6985) );
  NANDN U9003 ( .A(n6967), .B(n6966), .Z(n6971) );
  NAND U9004 ( .A(n6969), .B(n6968), .Z(n6970) );
  NAND U9005 ( .A(n6971), .B(n6970), .Z(n6986) );
  XNOR U9006 ( .A(n6985), .B(n6986), .Z(n6977) );
  XNOR U9007 ( .A(n6978), .B(n6977), .Z(n6979) );
  XNOR U9008 ( .A(n6980), .B(n6979), .Z(n7009) );
  XNOR U9009 ( .A(sreg[1094]), .B(n7009), .Z(n7011) );
  NANDN U9010 ( .A(sreg[1093]), .B(n6972), .Z(n6976) );
  NAND U9011 ( .A(n6974), .B(n6973), .Z(n6975) );
  NAND U9012 ( .A(n6976), .B(n6975), .Z(n7010) );
  XNOR U9013 ( .A(n7011), .B(n7010), .Z(c[1094]) );
  NANDN U9014 ( .A(n6978), .B(n6977), .Z(n6982) );
  NANDN U9015 ( .A(n6980), .B(n6979), .Z(n6981) );
  AND U9016 ( .A(n6982), .B(n6981), .Z(n7021) );
  NANDN U9017 ( .A(n6984), .B(n6983), .Z(n6988) );
  NANDN U9018 ( .A(n6986), .B(n6985), .Z(n6987) );
  AND U9019 ( .A(n6988), .B(n6987), .Z(n7020) );
  NAND U9020 ( .A(n42143), .B(n6989), .Z(n6991) );
  XNOR U9021 ( .A(a[73]), .B(n4082), .Z(n7031) );
  NAND U9022 ( .A(n42144), .B(n7031), .Z(n6990) );
  AND U9023 ( .A(n6991), .B(n6990), .Z(n7046) );
  XOR U9024 ( .A(a[77]), .B(n42012), .Z(n7034) );
  XNOR U9025 ( .A(n7046), .B(n7045), .Z(n7048) );
  AND U9026 ( .A(a[79]), .B(b[0]), .Z(n6993) );
  XNOR U9027 ( .A(n6993), .B(n4071), .Z(n6995) );
  NANDN U9028 ( .A(b[0]), .B(a[78]), .Z(n6994) );
  NAND U9029 ( .A(n6995), .B(n6994), .Z(n7042) );
  XOR U9030 ( .A(a[75]), .B(n42085), .Z(n7035) );
  AND U9031 ( .A(a[71]), .B(b[7]), .Z(n7039) );
  XNOR U9032 ( .A(n7040), .B(n7039), .Z(n7041) );
  XNOR U9033 ( .A(n7042), .B(n7041), .Z(n7047) );
  XOR U9034 ( .A(n7048), .B(n7047), .Z(n7026) );
  NANDN U9035 ( .A(n6998), .B(n6997), .Z(n7002) );
  NANDN U9036 ( .A(n7000), .B(n6999), .Z(n7001) );
  AND U9037 ( .A(n7002), .B(n7001), .Z(n7025) );
  XNOR U9038 ( .A(n7026), .B(n7025), .Z(n7027) );
  NANDN U9039 ( .A(n7004), .B(n7003), .Z(n7008) );
  NAND U9040 ( .A(n7006), .B(n7005), .Z(n7007) );
  NAND U9041 ( .A(n7008), .B(n7007), .Z(n7028) );
  XNOR U9042 ( .A(n7027), .B(n7028), .Z(n7019) );
  XOR U9043 ( .A(n7020), .B(n7019), .Z(n7022) );
  XOR U9044 ( .A(n7021), .B(n7022), .Z(n7014) );
  XNOR U9045 ( .A(n7014), .B(sreg[1095]), .Z(n7016) );
  NANDN U9046 ( .A(sreg[1094]), .B(n7009), .Z(n7013) );
  NAND U9047 ( .A(n7011), .B(n7010), .Z(n7012) );
  AND U9048 ( .A(n7013), .B(n7012), .Z(n7015) );
  XOR U9049 ( .A(n7016), .B(n7015), .Z(c[1095]) );
  NANDN U9050 ( .A(n7014), .B(sreg[1095]), .Z(n7018) );
  NAND U9051 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U9052 ( .A(n7018), .B(n7017), .Z(n7085) );
  NANDN U9053 ( .A(n7020), .B(n7019), .Z(n7024) );
  OR U9054 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U9055 ( .A(n7024), .B(n7023), .Z(n7054) );
  NANDN U9056 ( .A(n7026), .B(n7025), .Z(n7030) );
  NANDN U9057 ( .A(n7028), .B(n7027), .Z(n7029) );
  AND U9058 ( .A(n7030), .B(n7029), .Z(n7052) );
  NAND U9059 ( .A(n42143), .B(n7031), .Z(n7033) );
  XNOR U9060 ( .A(a[74]), .B(n4082), .Z(n7063) );
  NAND U9061 ( .A(n42144), .B(n7063), .Z(n7032) );
  AND U9062 ( .A(n7033), .B(n7032), .Z(n7078) );
  XOR U9063 ( .A(a[78]), .B(n42012), .Z(n7066) );
  XNOR U9064 ( .A(n7078), .B(n7077), .Z(n7080) );
  XOR U9065 ( .A(a[76]), .B(n42085), .Z(n7067) );
  AND U9066 ( .A(a[72]), .B(b[7]), .Z(n7071) );
  XNOR U9067 ( .A(n7072), .B(n7071), .Z(n7073) );
  AND U9068 ( .A(a[80]), .B(b[0]), .Z(n7036) );
  XNOR U9069 ( .A(n7036), .B(n4071), .Z(n7038) );
  NANDN U9070 ( .A(b[0]), .B(a[79]), .Z(n7037) );
  NAND U9071 ( .A(n7038), .B(n7037), .Z(n7074) );
  XNOR U9072 ( .A(n7073), .B(n7074), .Z(n7079) );
  XOR U9073 ( .A(n7080), .B(n7079), .Z(n7058) );
  NANDN U9074 ( .A(n7040), .B(n7039), .Z(n7044) );
  NANDN U9075 ( .A(n7042), .B(n7041), .Z(n7043) );
  AND U9076 ( .A(n7044), .B(n7043), .Z(n7057) );
  XNOR U9077 ( .A(n7058), .B(n7057), .Z(n7059) );
  NANDN U9078 ( .A(n7046), .B(n7045), .Z(n7050) );
  NAND U9079 ( .A(n7048), .B(n7047), .Z(n7049) );
  NAND U9080 ( .A(n7050), .B(n7049), .Z(n7060) );
  XNOR U9081 ( .A(n7059), .B(n7060), .Z(n7051) );
  XNOR U9082 ( .A(n7052), .B(n7051), .Z(n7053) );
  XNOR U9083 ( .A(n7054), .B(n7053), .Z(n7083) );
  XNOR U9084 ( .A(sreg[1096]), .B(n7083), .Z(n7084) );
  XNOR U9085 ( .A(n7085), .B(n7084), .Z(c[1096]) );
  NANDN U9086 ( .A(n7052), .B(n7051), .Z(n7056) );
  NANDN U9087 ( .A(n7054), .B(n7053), .Z(n7055) );
  AND U9088 ( .A(n7056), .B(n7055), .Z(n7091) );
  NANDN U9089 ( .A(n7058), .B(n7057), .Z(n7062) );
  NANDN U9090 ( .A(n7060), .B(n7059), .Z(n7061) );
  AND U9091 ( .A(n7062), .B(n7061), .Z(n7089) );
  NAND U9092 ( .A(n42143), .B(n7063), .Z(n7065) );
  XNOR U9093 ( .A(a[75]), .B(n4082), .Z(n7100) );
  NAND U9094 ( .A(n42144), .B(n7100), .Z(n7064) );
  AND U9095 ( .A(n7065), .B(n7064), .Z(n7115) );
  XOR U9096 ( .A(a[79]), .B(n42012), .Z(n7103) );
  XNOR U9097 ( .A(n7115), .B(n7114), .Z(n7117) );
  XOR U9098 ( .A(a[77]), .B(n42085), .Z(n7104) );
  AND U9099 ( .A(a[73]), .B(b[7]), .Z(n7108) );
  XNOR U9100 ( .A(n7109), .B(n7108), .Z(n7110) );
  AND U9101 ( .A(a[81]), .B(b[0]), .Z(n7068) );
  XNOR U9102 ( .A(n7068), .B(n4071), .Z(n7070) );
  NANDN U9103 ( .A(b[0]), .B(a[80]), .Z(n7069) );
  NAND U9104 ( .A(n7070), .B(n7069), .Z(n7111) );
  XNOR U9105 ( .A(n7110), .B(n7111), .Z(n7116) );
  XOR U9106 ( .A(n7117), .B(n7116), .Z(n7095) );
  NANDN U9107 ( .A(n7072), .B(n7071), .Z(n7076) );
  NANDN U9108 ( .A(n7074), .B(n7073), .Z(n7075) );
  AND U9109 ( .A(n7076), .B(n7075), .Z(n7094) );
  XNOR U9110 ( .A(n7095), .B(n7094), .Z(n7096) );
  NANDN U9111 ( .A(n7078), .B(n7077), .Z(n7082) );
  NAND U9112 ( .A(n7080), .B(n7079), .Z(n7081) );
  NAND U9113 ( .A(n7082), .B(n7081), .Z(n7097) );
  XNOR U9114 ( .A(n7096), .B(n7097), .Z(n7088) );
  XNOR U9115 ( .A(n7089), .B(n7088), .Z(n7090) );
  XNOR U9116 ( .A(n7091), .B(n7090), .Z(n7120) );
  XNOR U9117 ( .A(sreg[1097]), .B(n7120), .Z(n7122) );
  NANDN U9118 ( .A(sreg[1096]), .B(n7083), .Z(n7087) );
  NAND U9119 ( .A(n7085), .B(n7084), .Z(n7086) );
  NAND U9120 ( .A(n7087), .B(n7086), .Z(n7121) );
  XNOR U9121 ( .A(n7122), .B(n7121), .Z(c[1097]) );
  NANDN U9122 ( .A(n7089), .B(n7088), .Z(n7093) );
  NANDN U9123 ( .A(n7091), .B(n7090), .Z(n7092) );
  AND U9124 ( .A(n7093), .B(n7092), .Z(n7128) );
  NANDN U9125 ( .A(n7095), .B(n7094), .Z(n7099) );
  NANDN U9126 ( .A(n7097), .B(n7096), .Z(n7098) );
  AND U9127 ( .A(n7099), .B(n7098), .Z(n7126) );
  NAND U9128 ( .A(n42143), .B(n7100), .Z(n7102) );
  XNOR U9129 ( .A(a[76]), .B(n4082), .Z(n7137) );
  NAND U9130 ( .A(n42144), .B(n7137), .Z(n7101) );
  AND U9131 ( .A(n7102), .B(n7101), .Z(n7152) );
  XOR U9132 ( .A(a[80]), .B(n42012), .Z(n7140) );
  XNOR U9133 ( .A(n7152), .B(n7151), .Z(n7154) );
  XOR U9134 ( .A(a[78]), .B(n42085), .Z(n7144) );
  AND U9135 ( .A(a[74]), .B(b[7]), .Z(n7145) );
  XNOR U9136 ( .A(n7146), .B(n7145), .Z(n7147) );
  AND U9137 ( .A(a[82]), .B(b[0]), .Z(n7105) );
  XNOR U9138 ( .A(n7105), .B(n4071), .Z(n7107) );
  NANDN U9139 ( .A(b[0]), .B(a[81]), .Z(n7106) );
  NAND U9140 ( .A(n7107), .B(n7106), .Z(n7148) );
  XNOR U9141 ( .A(n7147), .B(n7148), .Z(n7153) );
  XOR U9142 ( .A(n7154), .B(n7153), .Z(n7132) );
  NANDN U9143 ( .A(n7109), .B(n7108), .Z(n7113) );
  NANDN U9144 ( .A(n7111), .B(n7110), .Z(n7112) );
  AND U9145 ( .A(n7113), .B(n7112), .Z(n7131) );
  XNOR U9146 ( .A(n7132), .B(n7131), .Z(n7133) );
  NANDN U9147 ( .A(n7115), .B(n7114), .Z(n7119) );
  NAND U9148 ( .A(n7117), .B(n7116), .Z(n7118) );
  NAND U9149 ( .A(n7119), .B(n7118), .Z(n7134) );
  XNOR U9150 ( .A(n7133), .B(n7134), .Z(n7125) );
  XNOR U9151 ( .A(n7126), .B(n7125), .Z(n7127) );
  XNOR U9152 ( .A(n7128), .B(n7127), .Z(n7157) );
  XNOR U9153 ( .A(sreg[1098]), .B(n7157), .Z(n7159) );
  NANDN U9154 ( .A(sreg[1097]), .B(n7120), .Z(n7124) );
  NAND U9155 ( .A(n7122), .B(n7121), .Z(n7123) );
  NAND U9156 ( .A(n7124), .B(n7123), .Z(n7158) );
  XNOR U9157 ( .A(n7159), .B(n7158), .Z(c[1098]) );
  NANDN U9158 ( .A(n7126), .B(n7125), .Z(n7130) );
  NANDN U9159 ( .A(n7128), .B(n7127), .Z(n7129) );
  AND U9160 ( .A(n7130), .B(n7129), .Z(n7165) );
  NANDN U9161 ( .A(n7132), .B(n7131), .Z(n7136) );
  NANDN U9162 ( .A(n7134), .B(n7133), .Z(n7135) );
  AND U9163 ( .A(n7136), .B(n7135), .Z(n7163) );
  NAND U9164 ( .A(n42143), .B(n7137), .Z(n7139) );
  XNOR U9165 ( .A(a[77]), .B(n4082), .Z(n7174) );
  NAND U9166 ( .A(n42144), .B(n7174), .Z(n7138) );
  AND U9167 ( .A(n7139), .B(n7138), .Z(n7189) );
  XOR U9168 ( .A(a[81]), .B(n42012), .Z(n7177) );
  XNOR U9169 ( .A(n7189), .B(n7188), .Z(n7191) );
  AND U9170 ( .A(a[83]), .B(b[0]), .Z(n7141) );
  XNOR U9171 ( .A(n7141), .B(n4071), .Z(n7143) );
  NANDN U9172 ( .A(b[0]), .B(a[82]), .Z(n7142) );
  NAND U9173 ( .A(n7143), .B(n7142), .Z(n7185) );
  XOR U9174 ( .A(a[79]), .B(n42085), .Z(n7178) );
  AND U9175 ( .A(a[75]), .B(b[7]), .Z(n7182) );
  XNOR U9176 ( .A(n7183), .B(n7182), .Z(n7184) );
  XNOR U9177 ( .A(n7185), .B(n7184), .Z(n7190) );
  XOR U9178 ( .A(n7191), .B(n7190), .Z(n7169) );
  NANDN U9179 ( .A(n7146), .B(n7145), .Z(n7150) );
  NANDN U9180 ( .A(n7148), .B(n7147), .Z(n7149) );
  AND U9181 ( .A(n7150), .B(n7149), .Z(n7168) );
  XNOR U9182 ( .A(n7169), .B(n7168), .Z(n7170) );
  NANDN U9183 ( .A(n7152), .B(n7151), .Z(n7156) );
  NAND U9184 ( .A(n7154), .B(n7153), .Z(n7155) );
  NAND U9185 ( .A(n7156), .B(n7155), .Z(n7171) );
  XNOR U9186 ( .A(n7170), .B(n7171), .Z(n7162) );
  XNOR U9187 ( .A(n7163), .B(n7162), .Z(n7164) );
  XNOR U9188 ( .A(n7165), .B(n7164), .Z(n7194) );
  XNOR U9189 ( .A(sreg[1099]), .B(n7194), .Z(n7196) );
  NANDN U9190 ( .A(sreg[1098]), .B(n7157), .Z(n7161) );
  NAND U9191 ( .A(n7159), .B(n7158), .Z(n7160) );
  NAND U9192 ( .A(n7161), .B(n7160), .Z(n7195) );
  XNOR U9193 ( .A(n7196), .B(n7195), .Z(c[1099]) );
  NANDN U9194 ( .A(n7163), .B(n7162), .Z(n7167) );
  NANDN U9195 ( .A(n7165), .B(n7164), .Z(n7166) );
  AND U9196 ( .A(n7167), .B(n7166), .Z(n7202) );
  NANDN U9197 ( .A(n7169), .B(n7168), .Z(n7173) );
  NANDN U9198 ( .A(n7171), .B(n7170), .Z(n7172) );
  AND U9199 ( .A(n7173), .B(n7172), .Z(n7200) );
  NAND U9200 ( .A(n42143), .B(n7174), .Z(n7176) );
  XNOR U9201 ( .A(a[78]), .B(n4083), .Z(n7211) );
  NAND U9202 ( .A(n42144), .B(n7211), .Z(n7175) );
  AND U9203 ( .A(n7176), .B(n7175), .Z(n7226) );
  XOR U9204 ( .A(a[82]), .B(n42012), .Z(n7214) );
  XNOR U9205 ( .A(n7226), .B(n7225), .Z(n7228) );
  XOR U9206 ( .A(a[80]), .B(n42085), .Z(n7218) );
  AND U9207 ( .A(a[76]), .B(b[7]), .Z(n7219) );
  XNOR U9208 ( .A(n7220), .B(n7219), .Z(n7221) );
  AND U9209 ( .A(a[84]), .B(b[0]), .Z(n7179) );
  XNOR U9210 ( .A(n7179), .B(n4071), .Z(n7181) );
  NANDN U9211 ( .A(b[0]), .B(a[83]), .Z(n7180) );
  NAND U9212 ( .A(n7181), .B(n7180), .Z(n7222) );
  XNOR U9213 ( .A(n7221), .B(n7222), .Z(n7227) );
  XOR U9214 ( .A(n7228), .B(n7227), .Z(n7206) );
  NANDN U9215 ( .A(n7183), .B(n7182), .Z(n7187) );
  NANDN U9216 ( .A(n7185), .B(n7184), .Z(n7186) );
  AND U9217 ( .A(n7187), .B(n7186), .Z(n7205) );
  XNOR U9218 ( .A(n7206), .B(n7205), .Z(n7207) );
  NANDN U9219 ( .A(n7189), .B(n7188), .Z(n7193) );
  NAND U9220 ( .A(n7191), .B(n7190), .Z(n7192) );
  NAND U9221 ( .A(n7193), .B(n7192), .Z(n7208) );
  XNOR U9222 ( .A(n7207), .B(n7208), .Z(n7199) );
  XNOR U9223 ( .A(n7200), .B(n7199), .Z(n7201) );
  XNOR U9224 ( .A(n7202), .B(n7201), .Z(n7231) );
  XNOR U9225 ( .A(sreg[1100]), .B(n7231), .Z(n7233) );
  NANDN U9226 ( .A(sreg[1099]), .B(n7194), .Z(n7198) );
  NAND U9227 ( .A(n7196), .B(n7195), .Z(n7197) );
  NAND U9228 ( .A(n7198), .B(n7197), .Z(n7232) );
  XNOR U9229 ( .A(n7233), .B(n7232), .Z(c[1100]) );
  NANDN U9230 ( .A(n7200), .B(n7199), .Z(n7204) );
  NANDN U9231 ( .A(n7202), .B(n7201), .Z(n7203) );
  AND U9232 ( .A(n7204), .B(n7203), .Z(n7239) );
  NANDN U9233 ( .A(n7206), .B(n7205), .Z(n7210) );
  NANDN U9234 ( .A(n7208), .B(n7207), .Z(n7209) );
  AND U9235 ( .A(n7210), .B(n7209), .Z(n7237) );
  NAND U9236 ( .A(n42143), .B(n7211), .Z(n7213) );
  XNOR U9237 ( .A(a[79]), .B(n4083), .Z(n7248) );
  NAND U9238 ( .A(n42144), .B(n7248), .Z(n7212) );
  AND U9239 ( .A(n7213), .B(n7212), .Z(n7263) );
  XOR U9240 ( .A(a[83]), .B(n42012), .Z(n7251) );
  XNOR U9241 ( .A(n7263), .B(n7262), .Z(n7265) );
  AND U9242 ( .A(a[85]), .B(b[0]), .Z(n7215) );
  XNOR U9243 ( .A(n7215), .B(n4071), .Z(n7217) );
  NANDN U9244 ( .A(b[0]), .B(a[84]), .Z(n7216) );
  NAND U9245 ( .A(n7217), .B(n7216), .Z(n7259) );
  XOR U9246 ( .A(a[81]), .B(n42085), .Z(n7255) );
  AND U9247 ( .A(a[77]), .B(b[7]), .Z(n7256) );
  XNOR U9248 ( .A(n7257), .B(n7256), .Z(n7258) );
  XNOR U9249 ( .A(n7259), .B(n7258), .Z(n7264) );
  XOR U9250 ( .A(n7265), .B(n7264), .Z(n7243) );
  NANDN U9251 ( .A(n7220), .B(n7219), .Z(n7224) );
  NANDN U9252 ( .A(n7222), .B(n7221), .Z(n7223) );
  AND U9253 ( .A(n7224), .B(n7223), .Z(n7242) );
  XNOR U9254 ( .A(n7243), .B(n7242), .Z(n7244) );
  NANDN U9255 ( .A(n7226), .B(n7225), .Z(n7230) );
  NAND U9256 ( .A(n7228), .B(n7227), .Z(n7229) );
  NAND U9257 ( .A(n7230), .B(n7229), .Z(n7245) );
  XNOR U9258 ( .A(n7244), .B(n7245), .Z(n7236) );
  XNOR U9259 ( .A(n7237), .B(n7236), .Z(n7238) );
  XNOR U9260 ( .A(n7239), .B(n7238), .Z(n7268) );
  XNOR U9261 ( .A(sreg[1101]), .B(n7268), .Z(n7270) );
  NANDN U9262 ( .A(sreg[1100]), .B(n7231), .Z(n7235) );
  NAND U9263 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U9264 ( .A(n7235), .B(n7234), .Z(n7269) );
  XNOR U9265 ( .A(n7270), .B(n7269), .Z(c[1101]) );
  NANDN U9266 ( .A(n7237), .B(n7236), .Z(n7241) );
  NANDN U9267 ( .A(n7239), .B(n7238), .Z(n7240) );
  AND U9268 ( .A(n7241), .B(n7240), .Z(n7276) );
  NANDN U9269 ( .A(n7243), .B(n7242), .Z(n7247) );
  NANDN U9270 ( .A(n7245), .B(n7244), .Z(n7246) );
  AND U9271 ( .A(n7247), .B(n7246), .Z(n7274) );
  NAND U9272 ( .A(n42143), .B(n7248), .Z(n7250) );
  XNOR U9273 ( .A(a[80]), .B(n4083), .Z(n7285) );
  NAND U9274 ( .A(n42144), .B(n7285), .Z(n7249) );
  AND U9275 ( .A(n7250), .B(n7249), .Z(n7300) );
  XOR U9276 ( .A(a[84]), .B(n42012), .Z(n7288) );
  XNOR U9277 ( .A(n7300), .B(n7299), .Z(n7302) );
  AND U9278 ( .A(a[86]), .B(b[0]), .Z(n7252) );
  XNOR U9279 ( .A(n7252), .B(n4071), .Z(n7254) );
  NANDN U9280 ( .A(b[0]), .B(a[85]), .Z(n7253) );
  NAND U9281 ( .A(n7254), .B(n7253), .Z(n7296) );
  XOR U9282 ( .A(a[82]), .B(n42085), .Z(n7292) );
  AND U9283 ( .A(a[78]), .B(b[7]), .Z(n7293) );
  XNOR U9284 ( .A(n7294), .B(n7293), .Z(n7295) );
  XNOR U9285 ( .A(n7296), .B(n7295), .Z(n7301) );
  XOR U9286 ( .A(n7302), .B(n7301), .Z(n7280) );
  NANDN U9287 ( .A(n7257), .B(n7256), .Z(n7261) );
  NANDN U9288 ( .A(n7259), .B(n7258), .Z(n7260) );
  AND U9289 ( .A(n7261), .B(n7260), .Z(n7279) );
  XNOR U9290 ( .A(n7280), .B(n7279), .Z(n7281) );
  NANDN U9291 ( .A(n7263), .B(n7262), .Z(n7267) );
  NAND U9292 ( .A(n7265), .B(n7264), .Z(n7266) );
  NAND U9293 ( .A(n7267), .B(n7266), .Z(n7282) );
  XNOR U9294 ( .A(n7281), .B(n7282), .Z(n7273) );
  XNOR U9295 ( .A(n7274), .B(n7273), .Z(n7275) );
  XNOR U9296 ( .A(n7276), .B(n7275), .Z(n7305) );
  XNOR U9297 ( .A(sreg[1102]), .B(n7305), .Z(n7307) );
  NANDN U9298 ( .A(sreg[1101]), .B(n7268), .Z(n7272) );
  NAND U9299 ( .A(n7270), .B(n7269), .Z(n7271) );
  NAND U9300 ( .A(n7272), .B(n7271), .Z(n7306) );
  XNOR U9301 ( .A(n7307), .B(n7306), .Z(c[1102]) );
  NANDN U9302 ( .A(n7274), .B(n7273), .Z(n7278) );
  NANDN U9303 ( .A(n7276), .B(n7275), .Z(n7277) );
  AND U9304 ( .A(n7278), .B(n7277), .Z(n7313) );
  NANDN U9305 ( .A(n7280), .B(n7279), .Z(n7284) );
  NANDN U9306 ( .A(n7282), .B(n7281), .Z(n7283) );
  AND U9307 ( .A(n7284), .B(n7283), .Z(n7311) );
  NAND U9308 ( .A(n42143), .B(n7285), .Z(n7287) );
  XNOR U9309 ( .A(a[81]), .B(n4083), .Z(n7322) );
  NAND U9310 ( .A(n42144), .B(n7322), .Z(n7286) );
  AND U9311 ( .A(n7287), .B(n7286), .Z(n7337) );
  XOR U9312 ( .A(a[85]), .B(n42012), .Z(n7325) );
  XNOR U9313 ( .A(n7337), .B(n7336), .Z(n7339) );
  AND U9314 ( .A(a[87]), .B(b[0]), .Z(n7289) );
  XNOR U9315 ( .A(n7289), .B(n4071), .Z(n7291) );
  NANDN U9316 ( .A(b[0]), .B(a[86]), .Z(n7290) );
  NAND U9317 ( .A(n7291), .B(n7290), .Z(n7333) );
  XOR U9318 ( .A(a[83]), .B(n42085), .Z(n7329) );
  AND U9319 ( .A(a[79]), .B(b[7]), .Z(n7330) );
  XNOR U9320 ( .A(n7331), .B(n7330), .Z(n7332) );
  XNOR U9321 ( .A(n7333), .B(n7332), .Z(n7338) );
  XOR U9322 ( .A(n7339), .B(n7338), .Z(n7317) );
  NANDN U9323 ( .A(n7294), .B(n7293), .Z(n7298) );
  NANDN U9324 ( .A(n7296), .B(n7295), .Z(n7297) );
  AND U9325 ( .A(n7298), .B(n7297), .Z(n7316) );
  XNOR U9326 ( .A(n7317), .B(n7316), .Z(n7318) );
  NANDN U9327 ( .A(n7300), .B(n7299), .Z(n7304) );
  NAND U9328 ( .A(n7302), .B(n7301), .Z(n7303) );
  NAND U9329 ( .A(n7304), .B(n7303), .Z(n7319) );
  XNOR U9330 ( .A(n7318), .B(n7319), .Z(n7310) );
  XNOR U9331 ( .A(n7311), .B(n7310), .Z(n7312) );
  XNOR U9332 ( .A(n7313), .B(n7312), .Z(n7342) );
  XNOR U9333 ( .A(sreg[1103]), .B(n7342), .Z(n7344) );
  NANDN U9334 ( .A(sreg[1102]), .B(n7305), .Z(n7309) );
  NAND U9335 ( .A(n7307), .B(n7306), .Z(n7308) );
  NAND U9336 ( .A(n7309), .B(n7308), .Z(n7343) );
  XNOR U9337 ( .A(n7344), .B(n7343), .Z(c[1103]) );
  NANDN U9338 ( .A(n7311), .B(n7310), .Z(n7315) );
  NANDN U9339 ( .A(n7313), .B(n7312), .Z(n7314) );
  AND U9340 ( .A(n7315), .B(n7314), .Z(n7350) );
  NANDN U9341 ( .A(n7317), .B(n7316), .Z(n7321) );
  NANDN U9342 ( .A(n7319), .B(n7318), .Z(n7320) );
  AND U9343 ( .A(n7321), .B(n7320), .Z(n7348) );
  NAND U9344 ( .A(n42143), .B(n7322), .Z(n7324) );
  XNOR U9345 ( .A(a[82]), .B(n4083), .Z(n7359) );
  NAND U9346 ( .A(n42144), .B(n7359), .Z(n7323) );
  AND U9347 ( .A(n7324), .B(n7323), .Z(n7374) );
  XOR U9348 ( .A(a[86]), .B(n42012), .Z(n7362) );
  XNOR U9349 ( .A(n7374), .B(n7373), .Z(n7376) );
  AND U9350 ( .A(a[88]), .B(b[0]), .Z(n7326) );
  XNOR U9351 ( .A(n7326), .B(n4071), .Z(n7328) );
  NANDN U9352 ( .A(b[0]), .B(a[87]), .Z(n7327) );
  NAND U9353 ( .A(n7328), .B(n7327), .Z(n7370) );
  XOR U9354 ( .A(a[84]), .B(n42085), .Z(n7363) );
  AND U9355 ( .A(a[80]), .B(b[7]), .Z(n7367) );
  XNOR U9356 ( .A(n7368), .B(n7367), .Z(n7369) );
  XNOR U9357 ( .A(n7370), .B(n7369), .Z(n7375) );
  XOR U9358 ( .A(n7376), .B(n7375), .Z(n7354) );
  NANDN U9359 ( .A(n7331), .B(n7330), .Z(n7335) );
  NANDN U9360 ( .A(n7333), .B(n7332), .Z(n7334) );
  AND U9361 ( .A(n7335), .B(n7334), .Z(n7353) );
  XNOR U9362 ( .A(n7354), .B(n7353), .Z(n7355) );
  NANDN U9363 ( .A(n7337), .B(n7336), .Z(n7341) );
  NAND U9364 ( .A(n7339), .B(n7338), .Z(n7340) );
  NAND U9365 ( .A(n7341), .B(n7340), .Z(n7356) );
  XNOR U9366 ( .A(n7355), .B(n7356), .Z(n7347) );
  XNOR U9367 ( .A(n7348), .B(n7347), .Z(n7349) );
  XNOR U9368 ( .A(n7350), .B(n7349), .Z(n7379) );
  XNOR U9369 ( .A(sreg[1104]), .B(n7379), .Z(n7381) );
  NANDN U9370 ( .A(sreg[1103]), .B(n7342), .Z(n7346) );
  NAND U9371 ( .A(n7344), .B(n7343), .Z(n7345) );
  NAND U9372 ( .A(n7346), .B(n7345), .Z(n7380) );
  XNOR U9373 ( .A(n7381), .B(n7380), .Z(c[1104]) );
  NANDN U9374 ( .A(n7348), .B(n7347), .Z(n7352) );
  NANDN U9375 ( .A(n7350), .B(n7349), .Z(n7351) );
  AND U9376 ( .A(n7352), .B(n7351), .Z(n7387) );
  NANDN U9377 ( .A(n7354), .B(n7353), .Z(n7358) );
  NANDN U9378 ( .A(n7356), .B(n7355), .Z(n7357) );
  AND U9379 ( .A(n7358), .B(n7357), .Z(n7385) );
  NAND U9380 ( .A(n42143), .B(n7359), .Z(n7361) );
  XNOR U9381 ( .A(a[83]), .B(n4083), .Z(n7396) );
  NAND U9382 ( .A(n42144), .B(n7396), .Z(n7360) );
  AND U9383 ( .A(n7361), .B(n7360), .Z(n7411) );
  XOR U9384 ( .A(a[87]), .B(n42012), .Z(n7399) );
  XNOR U9385 ( .A(n7411), .B(n7410), .Z(n7413) );
  XOR U9386 ( .A(a[85]), .B(n42085), .Z(n7403) );
  AND U9387 ( .A(a[81]), .B(b[7]), .Z(n7404) );
  XNOR U9388 ( .A(n7405), .B(n7404), .Z(n7406) );
  AND U9389 ( .A(a[89]), .B(b[0]), .Z(n7364) );
  XNOR U9390 ( .A(n7364), .B(n4071), .Z(n7366) );
  NANDN U9391 ( .A(b[0]), .B(a[88]), .Z(n7365) );
  NAND U9392 ( .A(n7366), .B(n7365), .Z(n7407) );
  XNOR U9393 ( .A(n7406), .B(n7407), .Z(n7412) );
  XOR U9394 ( .A(n7413), .B(n7412), .Z(n7391) );
  NANDN U9395 ( .A(n7368), .B(n7367), .Z(n7372) );
  NANDN U9396 ( .A(n7370), .B(n7369), .Z(n7371) );
  AND U9397 ( .A(n7372), .B(n7371), .Z(n7390) );
  XNOR U9398 ( .A(n7391), .B(n7390), .Z(n7392) );
  NANDN U9399 ( .A(n7374), .B(n7373), .Z(n7378) );
  NAND U9400 ( .A(n7376), .B(n7375), .Z(n7377) );
  NAND U9401 ( .A(n7378), .B(n7377), .Z(n7393) );
  XNOR U9402 ( .A(n7392), .B(n7393), .Z(n7384) );
  XNOR U9403 ( .A(n7385), .B(n7384), .Z(n7386) );
  XNOR U9404 ( .A(n7387), .B(n7386), .Z(n7416) );
  XNOR U9405 ( .A(sreg[1105]), .B(n7416), .Z(n7418) );
  NANDN U9406 ( .A(sreg[1104]), .B(n7379), .Z(n7383) );
  NAND U9407 ( .A(n7381), .B(n7380), .Z(n7382) );
  NAND U9408 ( .A(n7383), .B(n7382), .Z(n7417) );
  XNOR U9409 ( .A(n7418), .B(n7417), .Z(c[1105]) );
  NANDN U9410 ( .A(n7385), .B(n7384), .Z(n7389) );
  NANDN U9411 ( .A(n7387), .B(n7386), .Z(n7388) );
  AND U9412 ( .A(n7389), .B(n7388), .Z(n7424) );
  NANDN U9413 ( .A(n7391), .B(n7390), .Z(n7395) );
  NANDN U9414 ( .A(n7393), .B(n7392), .Z(n7394) );
  AND U9415 ( .A(n7395), .B(n7394), .Z(n7422) );
  NAND U9416 ( .A(n42143), .B(n7396), .Z(n7398) );
  XNOR U9417 ( .A(a[84]), .B(n4083), .Z(n7433) );
  NAND U9418 ( .A(n42144), .B(n7433), .Z(n7397) );
  AND U9419 ( .A(n7398), .B(n7397), .Z(n7448) );
  XOR U9420 ( .A(a[88]), .B(n42012), .Z(n7436) );
  XNOR U9421 ( .A(n7448), .B(n7447), .Z(n7450) );
  AND U9422 ( .A(a[90]), .B(b[0]), .Z(n7400) );
  XNOR U9423 ( .A(n7400), .B(n4071), .Z(n7402) );
  NANDN U9424 ( .A(b[0]), .B(a[89]), .Z(n7401) );
  NAND U9425 ( .A(n7402), .B(n7401), .Z(n7444) );
  XOR U9426 ( .A(a[86]), .B(n42085), .Z(n7440) );
  AND U9427 ( .A(a[82]), .B(b[7]), .Z(n7441) );
  XNOR U9428 ( .A(n7442), .B(n7441), .Z(n7443) );
  XNOR U9429 ( .A(n7444), .B(n7443), .Z(n7449) );
  XOR U9430 ( .A(n7450), .B(n7449), .Z(n7428) );
  NANDN U9431 ( .A(n7405), .B(n7404), .Z(n7409) );
  NANDN U9432 ( .A(n7407), .B(n7406), .Z(n7408) );
  AND U9433 ( .A(n7409), .B(n7408), .Z(n7427) );
  XNOR U9434 ( .A(n7428), .B(n7427), .Z(n7429) );
  NANDN U9435 ( .A(n7411), .B(n7410), .Z(n7415) );
  NAND U9436 ( .A(n7413), .B(n7412), .Z(n7414) );
  NAND U9437 ( .A(n7415), .B(n7414), .Z(n7430) );
  XNOR U9438 ( .A(n7429), .B(n7430), .Z(n7421) );
  XNOR U9439 ( .A(n7422), .B(n7421), .Z(n7423) );
  XNOR U9440 ( .A(n7424), .B(n7423), .Z(n7453) );
  XNOR U9441 ( .A(sreg[1106]), .B(n7453), .Z(n7455) );
  NANDN U9442 ( .A(sreg[1105]), .B(n7416), .Z(n7420) );
  NAND U9443 ( .A(n7418), .B(n7417), .Z(n7419) );
  NAND U9444 ( .A(n7420), .B(n7419), .Z(n7454) );
  XNOR U9445 ( .A(n7455), .B(n7454), .Z(c[1106]) );
  NANDN U9446 ( .A(n7422), .B(n7421), .Z(n7426) );
  NANDN U9447 ( .A(n7424), .B(n7423), .Z(n7425) );
  AND U9448 ( .A(n7426), .B(n7425), .Z(n7461) );
  NANDN U9449 ( .A(n7428), .B(n7427), .Z(n7432) );
  NANDN U9450 ( .A(n7430), .B(n7429), .Z(n7431) );
  AND U9451 ( .A(n7432), .B(n7431), .Z(n7459) );
  NAND U9452 ( .A(n42143), .B(n7433), .Z(n7435) );
  XNOR U9453 ( .A(a[85]), .B(n4084), .Z(n7470) );
  NAND U9454 ( .A(n42144), .B(n7470), .Z(n7434) );
  AND U9455 ( .A(n7435), .B(n7434), .Z(n7485) );
  XOR U9456 ( .A(a[89]), .B(n42012), .Z(n7473) );
  XNOR U9457 ( .A(n7485), .B(n7484), .Z(n7487) );
  AND U9458 ( .A(a[91]), .B(b[0]), .Z(n7437) );
  XNOR U9459 ( .A(n7437), .B(n4071), .Z(n7439) );
  NANDN U9460 ( .A(b[0]), .B(a[90]), .Z(n7438) );
  NAND U9461 ( .A(n7439), .B(n7438), .Z(n7481) );
  XOR U9462 ( .A(a[87]), .B(n42085), .Z(n7477) );
  AND U9463 ( .A(a[83]), .B(b[7]), .Z(n7478) );
  XNOR U9464 ( .A(n7479), .B(n7478), .Z(n7480) );
  XNOR U9465 ( .A(n7481), .B(n7480), .Z(n7486) );
  XOR U9466 ( .A(n7487), .B(n7486), .Z(n7465) );
  NANDN U9467 ( .A(n7442), .B(n7441), .Z(n7446) );
  NANDN U9468 ( .A(n7444), .B(n7443), .Z(n7445) );
  AND U9469 ( .A(n7446), .B(n7445), .Z(n7464) );
  XNOR U9470 ( .A(n7465), .B(n7464), .Z(n7466) );
  NANDN U9471 ( .A(n7448), .B(n7447), .Z(n7452) );
  NAND U9472 ( .A(n7450), .B(n7449), .Z(n7451) );
  NAND U9473 ( .A(n7452), .B(n7451), .Z(n7467) );
  XNOR U9474 ( .A(n7466), .B(n7467), .Z(n7458) );
  XNOR U9475 ( .A(n7459), .B(n7458), .Z(n7460) );
  XNOR U9476 ( .A(n7461), .B(n7460), .Z(n7490) );
  XNOR U9477 ( .A(sreg[1107]), .B(n7490), .Z(n7492) );
  NANDN U9478 ( .A(sreg[1106]), .B(n7453), .Z(n7457) );
  NAND U9479 ( .A(n7455), .B(n7454), .Z(n7456) );
  NAND U9480 ( .A(n7457), .B(n7456), .Z(n7491) );
  XNOR U9481 ( .A(n7492), .B(n7491), .Z(c[1107]) );
  NANDN U9482 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U9483 ( .A(n7461), .B(n7460), .Z(n7462) );
  AND U9484 ( .A(n7463), .B(n7462), .Z(n7498) );
  NANDN U9485 ( .A(n7465), .B(n7464), .Z(n7469) );
  NANDN U9486 ( .A(n7467), .B(n7466), .Z(n7468) );
  AND U9487 ( .A(n7469), .B(n7468), .Z(n7496) );
  NAND U9488 ( .A(n42143), .B(n7470), .Z(n7472) );
  XNOR U9489 ( .A(a[86]), .B(n4084), .Z(n7507) );
  NAND U9490 ( .A(n42144), .B(n7507), .Z(n7471) );
  AND U9491 ( .A(n7472), .B(n7471), .Z(n7522) );
  XOR U9492 ( .A(a[90]), .B(n42012), .Z(n7510) );
  XNOR U9493 ( .A(n7522), .B(n7521), .Z(n7524) );
  AND U9494 ( .A(a[92]), .B(b[0]), .Z(n7474) );
  XNOR U9495 ( .A(n7474), .B(n4071), .Z(n7476) );
  NANDN U9496 ( .A(b[0]), .B(a[91]), .Z(n7475) );
  NAND U9497 ( .A(n7476), .B(n7475), .Z(n7518) );
  XOR U9498 ( .A(a[88]), .B(n42085), .Z(n7514) );
  AND U9499 ( .A(a[84]), .B(b[7]), .Z(n7515) );
  XNOR U9500 ( .A(n7516), .B(n7515), .Z(n7517) );
  XNOR U9501 ( .A(n7518), .B(n7517), .Z(n7523) );
  XOR U9502 ( .A(n7524), .B(n7523), .Z(n7502) );
  NANDN U9503 ( .A(n7479), .B(n7478), .Z(n7483) );
  NANDN U9504 ( .A(n7481), .B(n7480), .Z(n7482) );
  AND U9505 ( .A(n7483), .B(n7482), .Z(n7501) );
  XNOR U9506 ( .A(n7502), .B(n7501), .Z(n7503) );
  NANDN U9507 ( .A(n7485), .B(n7484), .Z(n7489) );
  NAND U9508 ( .A(n7487), .B(n7486), .Z(n7488) );
  NAND U9509 ( .A(n7489), .B(n7488), .Z(n7504) );
  XNOR U9510 ( .A(n7503), .B(n7504), .Z(n7495) );
  XNOR U9511 ( .A(n7496), .B(n7495), .Z(n7497) );
  XNOR U9512 ( .A(n7498), .B(n7497), .Z(n7527) );
  XNOR U9513 ( .A(sreg[1108]), .B(n7527), .Z(n7529) );
  NANDN U9514 ( .A(sreg[1107]), .B(n7490), .Z(n7494) );
  NAND U9515 ( .A(n7492), .B(n7491), .Z(n7493) );
  NAND U9516 ( .A(n7494), .B(n7493), .Z(n7528) );
  XNOR U9517 ( .A(n7529), .B(n7528), .Z(c[1108]) );
  NANDN U9518 ( .A(n7496), .B(n7495), .Z(n7500) );
  NANDN U9519 ( .A(n7498), .B(n7497), .Z(n7499) );
  AND U9520 ( .A(n7500), .B(n7499), .Z(n7535) );
  NANDN U9521 ( .A(n7502), .B(n7501), .Z(n7506) );
  NANDN U9522 ( .A(n7504), .B(n7503), .Z(n7505) );
  AND U9523 ( .A(n7506), .B(n7505), .Z(n7533) );
  NAND U9524 ( .A(n42143), .B(n7507), .Z(n7509) );
  XNOR U9525 ( .A(a[87]), .B(n4084), .Z(n7544) );
  NAND U9526 ( .A(n42144), .B(n7544), .Z(n7508) );
  AND U9527 ( .A(n7509), .B(n7508), .Z(n7559) );
  XOR U9528 ( .A(a[91]), .B(n42012), .Z(n7547) );
  XNOR U9529 ( .A(n7559), .B(n7558), .Z(n7561) );
  AND U9530 ( .A(a[93]), .B(b[0]), .Z(n7511) );
  XNOR U9531 ( .A(n7511), .B(n4071), .Z(n7513) );
  NANDN U9532 ( .A(b[0]), .B(a[92]), .Z(n7512) );
  NAND U9533 ( .A(n7513), .B(n7512), .Z(n7555) );
  XOR U9534 ( .A(a[89]), .B(n42085), .Z(n7551) );
  AND U9535 ( .A(a[85]), .B(b[7]), .Z(n7552) );
  XNOR U9536 ( .A(n7553), .B(n7552), .Z(n7554) );
  XNOR U9537 ( .A(n7555), .B(n7554), .Z(n7560) );
  XOR U9538 ( .A(n7561), .B(n7560), .Z(n7539) );
  NANDN U9539 ( .A(n7516), .B(n7515), .Z(n7520) );
  NANDN U9540 ( .A(n7518), .B(n7517), .Z(n7519) );
  AND U9541 ( .A(n7520), .B(n7519), .Z(n7538) );
  XNOR U9542 ( .A(n7539), .B(n7538), .Z(n7540) );
  NANDN U9543 ( .A(n7522), .B(n7521), .Z(n7526) );
  NAND U9544 ( .A(n7524), .B(n7523), .Z(n7525) );
  NAND U9545 ( .A(n7526), .B(n7525), .Z(n7541) );
  XNOR U9546 ( .A(n7540), .B(n7541), .Z(n7532) );
  XNOR U9547 ( .A(n7533), .B(n7532), .Z(n7534) );
  XNOR U9548 ( .A(n7535), .B(n7534), .Z(n7564) );
  XNOR U9549 ( .A(sreg[1109]), .B(n7564), .Z(n7566) );
  NANDN U9550 ( .A(sreg[1108]), .B(n7527), .Z(n7531) );
  NAND U9551 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U9552 ( .A(n7531), .B(n7530), .Z(n7565) );
  XNOR U9553 ( .A(n7566), .B(n7565), .Z(c[1109]) );
  NANDN U9554 ( .A(n7533), .B(n7532), .Z(n7537) );
  NANDN U9555 ( .A(n7535), .B(n7534), .Z(n7536) );
  AND U9556 ( .A(n7537), .B(n7536), .Z(n7572) );
  NANDN U9557 ( .A(n7539), .B(n7538), .Z(n7543) );
  NANDN U9558 ( .A(n7541), .B(n7540), .Z(n7542) );
  AND U9559 ( .A(n7543), .B(n7542), .Z(n7570) );
  NAND U9560 ( .A(n42143), .B(n7544), .Z(n7546) );
  XNOR U9561 ( .A(a[88]), .B(n4084), .Z(n7581) );
  NAND U9562 ( .A(n42144), .B(n7581), .Z(n7545) );
  AND U9563 ( .A(n7546), .B(n7545), .Z(n7596) );
  XOR U9564 ( .A(a[92]), .B(n42012), .Z(n7584) );
  XNOR U9565 ( .A(n7596), .B(n7595), .Z(n7598) );
  AND U9566 ( .A(a[94]), .B(b[0]), .Z(n7548) );
  XNOR U9567 ( .A(n7548), .B(n4071), .Z(n7550) );
  NANDN U9568 ( .A(b[0]), .B(a[93]), .Z(n7549) );
  NAND U9569 ( .A(n7550), .B(n7549), .Z(n7592) );
  XOR U9570 ( .A(a[90]), .B(n42085), .Z(n7588) );
  AND U9571 ( .A(a[86]), .B(b[7]), .Z(n7589) );
  XNOR U9572 ( .A(n7590), .B(n7589), .Z(n7591) );
  XNOR U9573 ( .A(n7592), .B(n7591), .Z(n7597) );
  XOR U9574 ( .A(n7598), .B(n7597), .Z(n7576) );
  NANDN U9575 ( .A(n7553), .B(n7552), .Z(n7557) );
  NANDN U9576 ( .A(n7555), .B(n7554), .Z(n7556) );
  AND U9577 ( .A(n7557), .B(n7556), .Z(n7575) );
  XNOR U9578 ( .A(n7576), .B(n7575), .Z(n7577) );
  NANDN U9579 ( .A(n7559), .B(n7558), .Z(n7563) );
  NAND U9580 ( .A(n7561), .B(n7560), .Z(n7562) );
  NAND U9581 ( .A(n7563), .B(n7562), .Z(n7578) );
  XNOR U9582 ( .A(n7577), .B(n7578), .Z(n7569) );
  XNOR U9583 ( .A(n7570), .B(n7569), .Z(n7571) );
  XNOR U9584 ( .A(n7572), .B(n7571), .Z(n7601) );
  XNOR U9585 ( .A(sreg[1110]), .B(n7601), .Z(n7603) );
  NANDN U9586 ( .A(sreg[1109]), .B(n7564), .Z(n7568) );
  NAND U9587 ( .A(n7566), .B(n7565), .Z(n7567) );
  NAND U9588 ( .A(n7568), .B(n7567), .Z(n7602) );
  XNOR U9589 ( .A(n7603), .B(n7602), .Z(c[1110]) );
  NANDN U9590 ( .A(n7570), .B(n7569), .Z(n7574) );
  NANDN U9591 ( .A(n7572), .B(n7571), .Z(n7573) );
  AND U9592 ( .A(n7574), .B(n7573), .Z(n7609) );
  NANDN U9593 ( .A(n7576), .B(n7575), .Z(n7580) );
  NANDN U9594 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U9595 ( .A(n7580), .B(n7579), .Z(n7607) );
  NAND U9596 ( .A(n42143), .B(n7581), .Z(n7583) );
  XNOR U9597 ( .A(a[89]), .B(n4084), .Z(n7618) );
  NAND U9598 ( .A(n42144), .B(n7618), .Z(n7582) );
  AND U9599 ( .A(n7583), .B(n7582), .Z(n7633) );
  XOR U9600 ( .A(a[93]), .B(n42012), .Z(n7621) );
  XNOR U9601 ( .A(n7633), .B(n7632), .Z(n7635) );
  AND U9602 ( .A(a[95]), .B(b[0]), .Z(n7585) );
  XNOR U9603 ( .A(n7585), .B(n4071), .Z(n7587) );
  NANDN U9604 ( .A(b[0]), .B(a[94]), .Z(n7586) );
  NAND U9605 ( .A(n7587), .B(n7586), .Z(n7629) );
  XOR U9606 ( .A(a[91]), .B(n42085), .Z(n7625) );
  AND U9607 ( .A(a[87]), .B(b[7]), .Z(n7626) );
  XNOR U9608 ( .A(n7627), .B(n7626), .Z(n7628) );
  XNOR U9609 ( .A(n7629), .B(n7628), .Z(n7634) );
  XOR U9610 ( .A(n7635), .B(n7634), .Z(n7613) );
  NANDN U9611 ( .A(n7590), .B(n7589), .Z(n7594) );
  NANDN U9612 ( .A(n7592), .B(n7591), .Z(n7593) );
  AND U9613 ( .A(n7594), .B(n7593), .Z(n7612) );
  XNOR U9614 ( .A(n7613), .B(n7612), .Z(n7614) );
  NANDN U9615 ( .A(n7596), .B(n7595), .Z(n7600) );
  NAND U9616 ( .A(n7598), .B(n7597), .Z(n7599) );
  NAND U9617 ( .A(n7600), .B(n7599), .Z(n7615) );
  XNOR U9618 ( .A(n7614), .B(n7615), .Z(n7606) );
  XNOR U9619 ( .A(n7607), .B(n7606), .Z(n7608) );
  XNOR U9620 ( .A(n7609), .B(n7608), .Z(n7638) );
  XNOR U9621 ( .A(sreg[1111]), .B(n7638), .Z(n7640) );
  NANDN U9622 ( .A(sreg[1110]), .B(n7601), .Z(n7605) );
  NAND U9623 ( .A(n7603), .B(n7602), .Z(n7604) );
  NAND U9624 ( .A(n7605), .B(n7604), .Z(n7639) );
  XNOR U9625 ( .A(n7640), .B(n7639), .Z(c[1111]) );
  NANDN U9626 ( .A(n7607), .B(n7606), .Z(n7611) );
  NANDN U9627 ( .A(n7609), .B(n7608), .Z(n7610) );
  AND U9628 ( .A(n7611), .B(n7610), .Z(n7646) );
  NANDN U9629 ( .A(n7613), .B(n7612), .Z(n7617) );
  NANDN U9630 ( .A(n7615), .B(n7614), .Z(n7616) );
  AND U9631 ( .A(n7617), .B(n7616), .Z(n7644) );
  NAND U9632 ( .A(n42143), .B(n7618), .Z(n7620) );
  XNOR U9633 ( .A(a[90]), .B(n4084), .Z(n7655) );
  NAND U9634 ( .A(n42144), .B(n7655), .Z(n7619) );
  AND U9635 ( .A(n7620), .B(n7619), .Z(n7670) );
  XOR U9636 ( .A(a[94]), .B(n42012), .Z(n7658) );
  XNOR U9637 ( .A(n7670), .B(n7669), .Z(n7672) );
  AND U9638 ( .A(a[96]), .B(b[0]), .Z(n7622) );
  XNOR U9639 ( .A(n7622), .B(n4071), .Z(n7624) );
  NANDN U9640 ( .A(b[0]), .B(a[95]), .Z(n7623) );
  NAND U9641 ( .A(n7624), .B(n7623), .Z(n7666) );
  XOR U9642 ( .A(a[92]), .B(n42085), .Z(n7662) );
  AND U9643 ( .A(a[88]), .B(b[7]), .Z(n7663) );
  XNOR U9644 ( .A(n7664), .B(n7663), .Z(n7665) );
  XNOR U9645 ( .A(n7666), .B(n7665), .Z(n7671) );
  XOR U9646 ( .A(n7672), .B(n7671), .Z(n7650) );
  NANDN U9647 ( .A(n7627), .B(n7626), .Z(n7631) );
  NANDN U9648 ( .A(n7629), .B(n7628), .Z(n7630) );
  AND U9649 ( .A(n7631), .B(n7630), .Z(n7649) );
  XNOR U9650 ( .A(n7650), .B(n7649), .Z(n7651) );
  NANDN U9651 ( .A(n7633), .B(n7632), .Z(n7637) );
  NAND U9652 ( .A(n7635), .B(n7634), .Z(n7636) );
  NAND U9653 ( .A(n7637), .B(n7636), .Z(n7652) );
  XNOR U9654 ( .A(n7651), .B(n7652), .Z(n7643) );
  XNOR U9655 ( .A(n7644), .B(n7643), .Z(n7645) );
  XNOR U9656 ( .A(n7646), .B(n7645), .Z(n7675) );
  XNOR U9657 ( .A(sreg[1112]), .B(n7675), .Z(n7677) );
  NANDN U9658 ( .A(sreg[1111]), .B(n7638), .Z(n7642) );
  NAND U9659 ( .A(n7640), .B(n7639), .Z(n7641) );
  NAND U9660 ( .A(n7642), .B(n7641), .Z(n7676) );
  XNOR U9661 ( .A(n7677), .B(n7676), .Z(c[1112]) );
  NANDN U9662 ( .A(n7644), .B(n7643), .Z(n7648) );
  NANDN U9663 ( .A(n7646), .B(n7645), .Z(n7647) );
  AND U9664 ( .A(n7648), .B(n7647), .Z(n7683) );
  NANDN U9665 ( .A(n7650), .B(n7649), .Z(n7654) );
  NANDN U9666 ( .A(n7652), .B(n7651), .Z(n7653) );
  AND U9667 ( .A(n7654), .B(n7653), .Z(n7681) );
  NAND U9668 ( .A(n42143), .B(n7655), .Z(n7657) );
  XNOR U9669 ( .A(a[91]), .B(n4084), .Z(n7692) );
  NAND U9670 ( .A(n42144), .B(n7692), .Z(n7656) );
  AND U9671 ( .A(n7657), .B(n7656), .Z(n7707) );
  XOR U9672 ( .A(a[95]), .B(n42012), .Z(n7695) );
  XNOR U9673 ( .A(n7707), .B(n7706), .Z(n7709) );
  AND U9674 ( .A(a[97]), .B(b[0]), .Z(n7659) );
  XNOR U9675 ( .A(n7659), .B(n4071), .Z(n7661) );
  NANDN U9676 ( .A(b[0]), .B(a[96]), .Z(n7660) );
  NAND U9677 ( .A(n7661), .B(n7660), .Z(n7703) );
  XOR U9678 ( .A(a[93]), .B(n42085), .Z(n7699) );
  AND U9679 ( .A(a[89]), .B(b[7]), .Z(n7700) );
  XNOR U9680 ( .A(n7701), .B(n7700), .Z(n7702) );
  XNOR U9681 ( .A(n7703), .B(n7702), .Z(n7708) );
  XOR U9682 ( .A(n7709), .B(n7708), .Z(n7687) );
  NANDN U9683 ( .A(n7664), .B(n7663), .Z(n7668) );
  NANDN U9684 ( .A(n7666), .B(n7665), .Z(n7667) );
  AND U9685 ( .A(n7668), .B(n7667), .Z(n7686) );
  XNOR U9686 ( .A(n7687), .B(n7686), .Z(n7688) );
  NANDN U9687 ( .A(n7670), .B(n7669), .Z(n7674) );
  NAND U9688 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U9689 ( .A(n7674), .B(n7673), .Z(n7689) );
  XNOR U9690 ( .A(n7688), .B(n7689), .Z(n7680) );
  XNOR U9691 ( .A(n7681), .B(n7680), .Z(n7682) );
  XNOR U9692 ( .A(n7683), .B(n7682), .Z(n7712) );
  XNOR U9693 ( .A(sreg[1113]), .B(n7712), .Z(n7714) );
  NANDN U9694 ( .A(sreg[1112]), .B(n7675), .Z(n7679) );
  NAND U9695 ( .A(n7677), .B(n7676), .Z(n7678) );
  NAND U9696 ( .A(n7679), .B(n7678), .Z(n7713) );
  XNOR U9697 ( .A(n7714), .B(n7713), .Z(c[1113]) );
  NANDN U9698 ( .A(n7681), .B(n7680), .Z(n7685) );
  NANDN U9699 ( .A(n7683), .B(n7682), .Z(n7684) );
  AND U9700 ( .A(n7685), .B(n7684), .Z(n7720) );
  NANDN U9701 ( .A(n7687), .B(n7686), .Z(n7691) );
  NANDN U9702 ( .A(n7689), .B(n7688), .Z(n7690) );
  AND U9703 ( .A(n7691), .B(n7690), .Z(n7718) );
  NAND U9704 ( .A(n42143), .B(n7692), .Z(n7694) );
  XNOR U9705 ( .A(a[92]), .B(n4085), .Z(n7729) );
  NAND U9706 ( .A(n42144), .B(n7729), .Z(n7693) );
  AND U9707 ( .A(n7694), .B(n7693), .Z(n7744) );
  XOR U9708 ( .A(a[96]), .B(n42012), .Z(n7732) );
  XNOR U9709 ( .A(n7744), .B(n7743), .Z(n7746) );
  AND U9710 ( .A(a[98]), .B(b[0]), .Z(n7696) );
  XNOR U9711 ( .A(n7696), .B(n4071), .Z(n7698) );
  NANDN U9712 ( .A(b[0]), .B(a[97]), .Z(n7697) );
  NAND U9713 ( .A(n7698), .B(n7697), .Z(n7740) );
  XOR U9714 ( .A(a[94]), .B(n42085), .Z(n7736) );
  AND U9715 ( .A(a[90]), .B(b[7]), .Z(n7737) );
  XNOR U9716 ( .A(n7738), .B(n7737), .Z(n7739) );
  XNOR U9717 ( .A(n7740), .B(n7739), .Z(n7745) );
  XOR U9718 ( .A(n7746), .B(n7745), .Z(n7724) );
  NANDN U9719 ( .A(n7701), .B(n7700), .Z(n7705) );
  NANDN U9720 ( .A(n7703), .B(n7702), .Z(n7704) );
  AND U9721 ( .A(n7705), .B(n7704), .Z(n7723) );
  XNOR U9722 ( .A(n7724), .B(n7723), .Z(n7725) );
  NANDN U9723 ( .A(n7707), .B(n7706), .Z(n7711) );
  NAND U9724 ( .A(n7709), .B(n7708), .Z(n7710) );
  NAND U9725 ( .A(n7711), .B(n7710), .Z(n7726) );
  XNOR U9726 ( .A(n7725), .B(n7726), .Z(n7717) );
  XNOR U9727 ( .A(n7718), .B(n7717), .Z(n7719) );
  XNOR U9728 ( .A(n7720), .B(n7719), .Z(n7749) );
  XNOR U9729 ( .A(sreg[1114]), .B(n7749), .Z(n7751) );
  NANDN U9730 ( .A(sreg[1113]), .B(n7712), .Z(n7716) );
  NAND U9731 ( .A(n7714), .B(n7713), .Z(n7715) );
  NAND U9732 ( .A(n7716), .B(n7715), .Z(n7750) );
  XNOR U9733 ( .A(n7751), .B(n7750), .Z(c[1114]) );
  NANDN U9734 ( .A(n7718), .B(n7717), .Z(n7722) );
  NANDN U9735 ( .A(n7720), .B(n7719), .Z(n7721) );
  AND U9736 ( .A(n7722), .B(n7721), .Z(n7757) );
  NANDN U9737 ( .A(n7724), .B(n7723), .Z(n7728) );
  NANDN U9738 ( .A(n7726), .B(n7725), .Z(n7727) );
  AND U9739 ( .A(n7728), .B(n7727), .Z(n7755) );
  NAND U9740 ( .A(n42143), .B(n7729), .Z(n7731) );
  XNOR U9741 ( .A(a[93]), .B(n4085), .Z(n7766) );
  NAND U9742 ( .A(n42144), .B(n7766), .Z(n7730) );
  AND U9743 ( .A(n7731), .B(n7730), .Z(n7781) );
  XOR U9744 ( .A(a[97]), .B(n42012), .Z(n7769) );
  XNOR U9745 ( .A(n7781), .B(n7780), .Z(n7783) );
  AND U9746 ( .A(a[99]), .B(b[0]), .Z(n7733) );
  XNOR U9747 ( .A(n7733), .B(n4071), .Z(n7735) );
  NANDN U9748 ( .A(b[0]), .B(a[98]), .Z(n7734) );
  NAND U9749 ( .A(n7735), .B(n7734), .Z(n7777) );
  XOR U9750 ( .A(a[95]), .B(n42085), .Z(n7773) );
  AND U9751 ( .A(a[91]), .B(b[7]), .Z(n7774) );
  XNOR U9752 ( .A(n7775), .B(n7774), .Z(n7776) );
  XNOR U9753 ( .A(n7777), .B(n7776), .Z(n7782) );
  XOR U9754 ( .A(n7783), .B(n7782), .Z(n7761) );
  NANDN U9755 ( .A(n7738), .B(n7737), .Z(n7742) );
  NANDN U9756 ( .A(n7740), .B(n7739), .Z(n7741) );
  AND U9757 ( .A(n7742), .B(n7741), .Z(n7760) );
  XNOR U9758 ( .A(n7761), .B(n7760), .Z(n7762) );
  NANDN U9759 ( .A(n7744), .B(n7743), .Z(n7748) );
  NAND U9760 ( .A(n7746), .B(n7745), .Z(n7747) );
  NAND U9761 ( .A(n7748), .B(n7747), .Z(n7763) );
  XNOR U9762 ( .A(n7762), .B(n7763), .Z(n7754) );
  XNOR U9763 ( .A(n7755), .B(n7754), .Z(n7756) );
  XNOR U9764 ( .A(n7757), .B(n7756), .Z(n7786) );
  XNOR U9765 ( .A(sreg[1115]), .B(n7786), .Z(n7788) );
  NANDN U9766 ( .A(sreg[1114]), .B(n7749), .Z(n7753) );
  NAND U9767 ( .A(n7751), .B(n7750), .Z(n7752) );
  NAND U9768 ( .A(n7753), .B(n7752), .Z(n7787) );
  XNOR U9769 ( .A(n7788), .B(n7787), .Z(c[1115]) );
  NANDN U9770 ( .A(n7755), .B(n7754), .Z(n7759) );
  NANDN U9771 ( .A(n7757), .B(n7756), .Z(n7758) );
  AND U9772 ( .A(n7759), .B(n7758), .Z(n7794) );
  NANDN U9773 ( .A(n7761), .B(n7760), .Z(n7765) );
  NANDN U9774 ( .A(n7763), .B(n7762), .Z(n7764) );
  AND U9775 ( .A(n7765), .B(n7764), .Z(n7792) );
  NAND U9776 ( .A(n42143), .B(n7766), .Z(n7768) );
  XNOR U9777 ( .A(a[94]), .B(n4085), .Z(n7803) );
  NAND U9778 ( .A(n42144), .B(n7803), .Z(n7767) );
  AND U9779 ( .A(n7768), .B(n7767), .Z(n7818) );
  XOR U9780 ( .A(a[98]), .B(n42012), .Z(n7806) );
  XNOR U9781 ( .A(n7818), .B(n7817), .Z(n7820) );
  AND U9782 ( .A(a[100]), .B(b[0]), .Z(n7770) );
  XNOR U9783 ( .A(n7770), .B(n4071), .Z(n7772) );
  NANDN U9784 ( .A(b[0]), .B(a[99]), .Z(n7771) );
  NAND U9785 ( .A(n7772), .B(n7771), .Z(n7814) );
  XOR U9786 ( .A(a[96]), .B(n42085), .Z(n7810) );
  AND U9787 ( .A(a[92]), .B(b[7]), .Z(n7811) );
  XNOR U9788 ( .A(n7812), .B(n7811), .Z(n7813) );
  XNOR U9789 ( .A(n7814), .B(n7813), .Z(n7819) );
  XOR U9790 ( .A(n7820), .B(n7819), .Z(n7798) );
  NANDN U9791 ( .A(n7775), .B(n7774), .Z(n7779) );
  NANDN U9792 ( .A(n7777), .B(n7776), .Z(n7778) );
  AND U9793 ( .A(n7779), .B(n7778), .Z(n7797) );
  XNOR U9794 ( .A(n7798), .B(n7797), .Z(n7799) );
  NANDN U9795 ( .A(n7781), .B(n7780), .Z(n7785) );
  NAND U9796 ( .A(n7783), .B(n7782), .Z(n7784) );
  NAND U9797 ( .A(n7785), .B(n7784), .Z(n7800) );
  XNOR U9798 ( .A(n7799), .B(n7800), .Z(n7791) );
  XNOR U9799 ( .A(n7792), .B(n7791), .Z(n7793) );
  XNOR U9800 ( .A(n7794), .B(n7793), .Z(n7823) );
  XNOR U9801 ( .A(sreg[1116]), .B(n7823), .Z(n7825) );
  NANDN U9802 ( .A(sreg[1115]), .B(n7786), .Z(n7790) );
  NAND U9803 ( .A(n7788), .B(n7787), .Z(n7789) );
  NAND U9804 ( .A(n7790), .B(n7789), .Z(n7824) );
  XNOR U9805 ( .A(n7825), .B(n7824), .Z(c[1116]) );
  NANDN U9806 ( .A(n7792), .B(n7791), .Z(n7796) );
  NANDN U9807 ( .A(n7794), .B(n7793), .Z(n7795) );
  AND U9808 ( .A(n7796), .B(n7795), .Z(n7831) );
  NANDN U9809 ( .A(n7798), .B(n7797), .Z(n7802) );
  NANDN U9810 ( .A(n7800), .B(n7799), .Z(n7801) );
  AND U9811 ( .A(n7802), .B(n7801), .Z(n7829) );
  NAND U9812 ( .A(n42143), .B(n7803), .Z(n7805) );
  XNOR U9813 ( .A(a[95]), .B(n4085), .Z(n7840) );
  NAND U9814 ( .A(n42144), .B(n7840), .Z(n7804) );
  AND U9815 ( .A(n7805), .B(n7804), .Z(n7855) );
  XOR U9816 ( .A(a[99]), .B(n42012), .Z(n7843) );
  XNOR U9817 ( .A(n7855), .B(n7854), .Z(n7857) );
  AND U9818 ( .A(a[101]), .B(b[0]), .Z(n7807) );
  XNOR U9819 ( .A(n7807), .B(n4071), .Z(n7809) );
  NANDN U9820 ( .A(b[0]), .B(a[100]), .Z(n7808) );
  NAND U9821 ( .A(n7809), .B(n7808), .Z(n7851) );
  XOR U9822 ( .A(a[97]), .B(n42085), .Z(n7847) );
  AND U9823 ( .A(a[93]), .B(b[7]), .Z(n7848) );
  XNOR U9824 ( .A(n7849), .B(n7848), .Z(n7850) );
  XNOR U9825 ( .A(n7851), .B(n7850), .Z(n7856) );
  XOR U9826 ( .A(n7857), .B(n7856), .Z(n7835) );
  NANDN U9827 ( .A(n7812), .B(n7811), .Z(n7816) );
  NANDN U9828 ( .A(n7814), .B(n7813), .Z(n7815) );
  AND U9829 ( .A(n7816), .B(n7815), .Z(n7834) );
  XNOR U9830 ( .A(n7835), .B(n7834), .Z(n7836) );
  NANDN U9831 ( .A(n7818), .B(n7817), .Z(n7822) );
  NAND U9832 ( .A(n7820), .B(n7819), .Z(n7821) );
  NAND U9833 ( .A(n7822), .B(n7821), .Z(n7837) );
  XNOR U9834 ( .A(n7836), .B(n7837), .Z(n7828) );
  XNOR U9835 ( .A(n7829), .B(n7828), .Z(n7830) );
  XNOR U9836 ( .A(n7831), .B(n7830), .Z(n7860) );
  XNOR U9837 ( .A(sreg[1117]), .B(n7860), .Z(n7862) );
  NANDN U9838 ( .A(sreg[1116]), .B(n7823), .Z(n7827) );
  NAND U9839 ( .A(n7825), .B(n7824), .Z(n7826) );
  NAND U9840 ( .A(n7827), .B(n7826), .Z(n7861) );
  XNOR U9841 ( .A(n7862), .B(n7861), .Z(c[1117]) );
  NANDN U9842 ( .A(n7829), .B(n7828), .Z(n7833) );
  NANDN U9843 ( .A(n7831), .B(n7830), .Z(n7832) );
  AND U9844 ( .A(n7833), .B(n7832), .Z(n7868) );
  NANDN U9845 ( .A(n7835), .B(n7834), .Z(n7839) );
  NANDN U9846 ( .A(n7837), .B(n7836), .Z(n7838) );
  AND U9847 ( .A(n7839), .B(n7838), .Z(n7866) );
  NAND U9848 ( .A(n42143), .B(n7840), .Z(n7842) );
  XNOR U9849 ( .A(a[96]), .B(n4085), .Z(n7877) );
  NAND U9850 ( .A(n42144), .B(n7877), .Z(n7841) );
  AND U9851 ( .A(n7842), .B(n7841), .Z(n7892) );
  XOR U9852 ( .A(a[100]), .B(n42012), .Z(n7880) );
  XNOR U9853 ( .A(n7892), .B(n7891), .Z(n7894) );
  AND U9854 ( .A(a[102]), .B(b[0]), .Z(n7844) );
  XNOR U9855 ( .A(n7844), .B(n4071), .Z(n7846) );
  NANDN U9856 ( .A(b[0]), .B(a[101]), .Z(n7845) );
  NAND U9857 ( .A(n7846), .B(n7845), .Z(n7888) );
  XOR U9858 ( .A(a[98]), .B(n42085), .Z(n7881) );
  AND U9859 ( .A(a[94]), .B(b[7]), .Z(n7885) );
  XNOR U9860 ( .A(n7886), .B(n7885), .Z(n7887) );
  XNOR U9861 ( .A(n7888), .B(n7887), .Z(n7893) );
  XOR U9862 ( .A(n7894), .B(n7893), .Z(n7872) );
  NANDN U9863 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U9864 ( .A(n7851), .B(n7850), .Z(n7852) );
  AND U9865 ( .A(n7853), .B(n7852), .Z(n7871) );
  XNOR U9866 ( .A(n7872), .B(n7871), .Z(n7873) );
  NANDN U9867 ( .A(n7855), .B(n7854), .Z(n7859) );
  NAND U9868 ( .A(n7857), .B(n7856), .Z(n7858) );
  NAND U9869 ( .A(n7859), .B(n7858), .Z(n7874) );
  XNOR U9870 ( .A(n7873), .B(n7874), .Z(n7865) );
  XNOR U9871 ( .A(n7866), .B(n7865), .Z(n7867) );
  XNOR U9872 ( .A(n7868), .B(n7867), .Z(n7897) );
  XNOR U9873 ( .A(sreg[1118]), .B(n7897), .Z(n7899) );
  NANDN U9874 ( .A(sreg[1117]), .B(n7860), .Z(n7864) );
  NAND U9875 ( .A(n7862), .B(n7861), .Z(n7863) );
  NAND U9876 ( .A(n7864), .B(n7863), .Z(n7898) );
  XNOR U9877 ( .A(n7899), .B(n7898), .Z(c[1118]) );
  NANDN U9878 ( .A(n7866), .B(n7865), .Z(n7870) );
  NANDN U9879 ( .A(n7868), .B(n7867), .Z(n7869) );
  AND U9880 ( .A(n7870), .B(n7869), .Z(n7905) );
  NANDN U9881 ( .A(n7872), .B(n7871), .Z(n7876) );
  NANDN U9882 ( .A(n7874), .B(n7873), .Z(n7875) );
  AND U9883 ( .A(n7876), .B(n7875), .Z(n7903) );
  NAND U9884 ( .A(n42143), .B(n7877), .Z(n7879) );
  XNOR U9885 ( .A(a[97]), .B(n4085), .Z(n7914) );
  NAND U9886 ( .A(n42144), .B(n7914), .Z(n7878) );
  AND U9887 ( .A(n7879), .B(n7878), .Z(n7929) );
  XOR U9888 ( .A(a[101]), .B(n42012), .Z(n7917) );
  XNOR U9889 ( .A(n7929), .B(n7928), .Z(n7931) );
  XOR U9890 ( .A(a[99]), .B(n42085), .Z(n7921) );
  AND U9891 ( .A(a[95]), .B(b[7]), .Z(n7922) );
  XNOR U9892 ( .A(n7923), .B(n7922), .Z(n7924) );
  AND U9893 ( .A(a[103]), .B(b[0]), .Z(n7882) );
  XNOR U9894 ( .A(n7882), .B(n4071), .Z(n7884) );
  NANDN U9895 ( .A(b[0]), .B(a[102]), .Z(n7883) );
  NAND U9896 ( .A(n7884), .B(n7883), .Z(n7925) );
  XNOR U9897 ( .A(n7924), .B(n7925), .Z(n7930) );
  XOR U9898 ( .A(n7931), .B(n7930), .Z(n7909) );
  NANDN U9899 ( .A(n7886), .B(n7885), .Z(n7890) );
  NANDN U9900 ( .A(n7888), .B(n7887), .Z(n7889) );
  AND U9901 ( .A(n7890), .B(n7889), .Z(n7908) );
  XNOR U9902 ( .A(n7909), .B(n7908), .Z(n7910) );
  NANDN U9903 ( .A(n7892), .B(n7891), .Z(n7896) );
  NAND U9904 ( .A(n7894), .B(n7893), .Z(n7895) );
  NAND U9905 ( .A(n7896), .B(n7895), .Z(n7911) );
  XNOR U9906 ( .A(n7910), .B(n7911), .Z(n7902) );
  XNOR U9907 ( .A(n7903), .B(n7902), .Z(n7904) );
  XNOR U9908 ( .A(n7905), .B(n7904), .Z(n7934) );
  XNOR U9909 ( .A(sreg[1119]), .B(n7934), .Z(n7936) );
  NANDN U9910 ( .A(sreg[1118]), .B(n7897), .Z(n7901) );
  NAND U9911 ( .A(n7899), .B(n7898), .Z(n7900) );
  NAND U9912 ( .A(n7901), .B(n7900), .Z(n7935) );
  XNOR U9913 ( .A(n7936), .B(n7935), .Z(c[1119]) );
  NANDN U9914 ( .A(n7903), .B(n7902), .Z(n7907) );
  NANDN U9915 ( .A(n7905), .B(n7904), .Z(n7906) );
  AND U9916 ( .A(n7907), .B(n7906), .Z(n7942) );
  NANDN U9917 ( .A(n7909), .B(n7908), .Z(n7913) );
  NANDN U9918 ( .A(n7911), .B(n7910), .Z(n7912) );
  AND U9919 ( .A(n7913), .B(n7912), .Z(n7940) );
  NAND U9920 ( .A(n42143), .B(n7914), .Z(n7916) );
  XNOR U9921 ( .A(a[98]), .B(n4085), .Z(n7951) );
  NAND U9922 ( .A(n42144), .B(n7951), .Z(n7915) );
  AND U9923 ( .A(n7916), .B(n7915), .Z(n7966) );
  XOR U9924 ( .A(a[102]), .B(n42012), .Z(n7954) );
  XNOR U9925 ( .A(n7966), .B(n7965), .Z(n7968) );
  AND U9926 ( .A(a[104]), .B(b[0]), .Z(n7918) );
  XNOR U9927 ( .A(n7918), .B(n4071), .Z(n7920) );
  NANDN U9928 ( .A(b[0]), .B(a[103]), .Z(n7919) );
  NAND U9929 ( .A(n7920), .B(n7919), .Z(n7962) );
  XOR U9930 ( .A(a[100]), .B(n42085), .Z(n7958) );
  AND U9931 ( .A(a[96]), .B(b[7]), .Z(n7959) );
  XNOR U9932 ( .A(n7960), .B(n7959), .Z(n7961) );
  XNOR U9933 ( .A(n7962), .B(n7961), .Z(n7967) );
  XOR U9934 ( .A(n7968), .B(n7967), .Z(n7946) );
  NANDN U9935 ( .A(n7923), .B(n7922), .Z(n7927) );
  NANDN U9936 ( .A(n7925), .B(n7924), .Z(n7926) );
  AND U9937 ( .A(n7927), .B(n7926), .Z(n7945) );
  XNOR U9938 ( .A(n7946), .B(n7945), .Z(n7947) );
  NANDN U9939 ( .A(n7929), .B(n7928), .Z(n7933) );
  NAND U9940 ( .A(n7931), .B(n7930), .Z(n7932) );
  NAND U9941 ( .A(n7933), .B(n7932), .Z(n7948) );
  XNOR U9942 ( .A(n7947), .B(n7948), .Z(n7939) );
  XNOR U9943 ( .A(n7940), .B(n7939), .Z(n7941) );
  XNOR U9944 ( .A(n7942), .B(n7941), .Z(n7971) );
  XNOR U9945 ( .A(sreg[1120]), .B(n7971), .Z(n7973) );
  NANDN U9946 ( .A(sreg[1119]), .B(n7934), .Z(n7938) );
  NAND U9947 ( .A(n7936), .B(n7935), .Z(n7937) );
  NAND U9948 ( .A(n7938), .B(n7937), .Z(n7972) );
  XNOR U9949 ( .A(n7973), .B(n7972), .Z(c[1120]) );
  NANDN U9950 ( .A(n7940), .B(n7939), .Z(n7944) );
  NANDN U9951 ( .A(n7942), .B(n7941), .Z(n7943) );
  AND U9952 ( .A(n7944), .B(n7943), .Z(n7979) );
  NANDN U9953 ( .A(n7946), .B(n7945), .Z(n7950) );
  NANDN U9954 ( .A(n7948), .B(n7947), .Z(n7949) );
  AND U9955 ( .A(n7950), .B(n7949), .Z(n7977) );
  NAND U9956 ( .A(n42143), .B(n7951), .Z(n7953) );
  XNOR U9957 ( .A(a[99]), .B(n4086), .Z(n7988) );
  NAND U9958 ( .A(n42144), .B(n7988), .Z(n7952) );
  AND U9959 ( .A(n7953), .B(n7952), .Z(n8003) );
  XOR U9960 ( .A(a[103]), .B(n42012), .Z(n7991) );
  XNOR U9961 ( .A(n8003), .B(n8002), .Z(n8005) );
  AND U9962 ( .A(a[105]), .B(b[0]), .Z(n7955) );
  XNOR U9963 ( .A(n7955), .B(n4071), .Z(n7957) );
  NANDN U9964 ( .A(b[0]), .B(a[104]), .Z(n7956) );
  NAND U9965 ( .A(n7957), .B(n7956), .Z(n7999) );
  XOR U9966 ( .A(a[101]), .B(n42085), .Z(n7995) );
  AND U9967 ( .A(a[97]), .B(b[7]), .Z(n7996) );
  XNOR U9968 ( .A(n7997), .B(n7996), .Z(n7998) );
  XNOR U9969 ( .A(n7999), .B(n7998), .Z(n8004) );
  XOR U9970 ( .A(n8005), .B(n8004), .Z(n7983) );
  NANDN U9971 ( .A(n7960), .B(n7959), .Z(n7964) );
  NANDN U9972 ( .A(n7962), .B(n7961), .Z(n7963) );
  AND U9973 ( .A(n7964), .B(n7963), .Z(n7982) );
  XNOR U9974 ( .A(n7983), .B(n7982), .Z(n7984) );
  NANDN U9975 ( .A(n7966), .B(n7965), .Z(n7970) );
  NAND U9976 ( .A(n7968), .B(n7967), .Z(n7969) );
  NAND U9977 ( .A(n7970), .B(n7969), .Z(n7985) );
  XNOR U9978 ( .A(n7984), .B(n7985), .Z(n7976) );
  XNOR U9979 ( .A(n7977), .B(n7976), .Z(n7978) );
  XNOR U9980 ( .A(n7979), .B(n7978), .Z(n8008) );
  XNOR U9981 ( .A(sreg[1121]), .B(n8008), .Z(n8010) );
  NANDN U9982 ( .A(sreg[1120]), .B(n7971), .Z(n7975) );
  NAND U9983 ( .A(n7973), .B(n7972), .Z(n7974) );
  NAND U9984 ( .A(n7975), .B(n7974), .Z(n8009) );
  XNOR U9985 ( .A(n8010), .B(n8009), .Z(c[1121]) );
  NANDN U9986 ( .A(n7977), .B(n7976), .Z(n7981) );
  NANDN U9987 ( .A(n7979), .B(n7978), .Z(n7980) );
  AND U9988 ( .A(n7981), .B(n7980), .Z(n8016) );
  NANDN U9989 ( .A(n7983), .B(n7982), .Z(n7987) );
  NANDN U9990 ( .A(n7985), .B(n7984), .Z(n7986) );
  AND U9991 ( .A(n7987), .B(n7986), .Z(n8014) );
  NAND U9992 ( .A(n42143), .B(n7988), .Z(n7990) );
  XNOR U9993 ( .A(a[100]), .B(n4086), .Z(n8025) );
  NAND U9994 ( .A(n42144), .B(n8025), .Z(n7989) );
  AND U9995 ( .A(n7990), .B(n7989), .Z(n8040) );
  XOR U9996 ( .A(a[104]), .B(n42012), .Z(n8028) );
  XNOR U9997 ( .A(n8040), .B(n8039), .Z(n8042) );
  NAND U9998 ( .A(a[106]), .B(b[0]), .Z(n7992) );
  XNOR U9999 ( .A(b[1]), .B(n7992), .Z(n7994) );
  NANDN U10000 ( .A(b[0]), .B(a[105]), .Z(n7993) );
  AND U10001 ( .A(n7994), .B(n7993), .Z(n8035) );
  XOR U10002 ( .A(a[102]), .B(n42085), .Z(n8032) );
  AND U10003 ( .A(a[98]), .B(b[7]), .Z(n8033) );
  XOR U10004 ( .A(n8034), .B(n8033), .Z(n8036) );
  XNOR U10005 ( .A(n8035), .B(n8036), .Z(n8041) );
  XOR U10006 ( .A(n8042), .B(n8041), .Z(n8020) );
  NANDN U10007 ( .A(n7997), .B(n7996), .Z(n8001) );
  NANDN U10008 ( .A(n7999), .B(n7998), .Z(n8000) );
  AND U10009 ( .A(n8001), .B(n8000), .Z(n8019) );
  XNOR U10010 ( .A(n8020), .B(n8019), .Z(n8021) );
  NANDN U10011 ( .A(n8003), .B(n8002), .Z(n8007) );
  NAND U10012 ( .A(n8005), .B(n8004), .Z(n8006) );
  NAND U10013 ( .A(n8007), .B(n8006), .Z(n8022) );
  XNOR U10014 ( .A(n8021), .B(n8022), .Z(n8013) );
  XNOR U10015 ( .A(n8014), .B(n8013), .Z(n8015) );
  XNOR U10016 ( .A(n8016), .B(n8015), .Z(n8045) );
  XNOR U10017 ( .A(sreg[1122]), .B(n8045), .Z(n8047) );
  NANDN U10018 ( .A(sreg[1121]), .B(n8008), .Z(n8012) );
  NAND U10019 ( .A(n8010), .B(n8009), .Z(n8011) );
  NAND U10020 ( .A(n8012), .B(n8011), .Z(n8046) );
  XNOR U10021 ( .A(n8047), .B(n8046), .Z(c[1122]) );
  NANDN U10022 ( .A(n8014), .B(n8013), .Z(n8018) );
  NANDN U10023 ( .A(n8016), .B(n8015), .Z(n8017) );
  AND U10024 ( .A(n8018), .B(n8017), .Z(n8053) );
  NANDN U10025 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U10026 ( .A(n8022), .B(n8021), .Z(n8023) );
  AND U10027 ( .A(n8024), .B(n8023), .Z(n8051) );
  NAND U10028 ( .A(n42143), .B(n8025), .Z(n8027) );
  XNOR U10029 ( .A(a[101]), .B(n4086), .Z(n8062) );
  NAND U10030 ( .A(n42144), .B(n8062), .Z(n8026) );
  AND U10031 ( .A(n8027), .B(n8026), .Z(n8077) );
  XOR U10032 ( .A(a[105]), .B(n42012), .Z(n8065) );
  XNOR U10033 ( .A(n8077), .B(n8076), .Z(n8079) );
  AND U10034 ( .A(a[107]), .B(b[0]), .Z(n8029) );
  XNOR U10035 ( .A(n8029), .B(n4071), .Z(n8031) );
  NANDN U10036 ( .A(b[0]), .B(a[106]), .Z(n8030) );
  NAND U10037 ( .A(n8031), .B(n8030), .Z(n8073) );
  XOR U10038 ( .A(a[103]), .B(n42085), .Z(n8069) );
  AND U10039 ( .A(a[99]), .B(b[7]), .Z(n8070) );
  XNOR U10040 ( .A(n8071), .B(n8070), .Z(n8072) );
  XNOR U10041 ( .A(n8073), .B(n8072), .Z(n8078) );
  XOR U10042 ( .A(n8079), .B(n8078), .Z(n8057) );
  NANDN U10043 ( .A(n8034), .B(n8033), .Z(n8038) );
  NANDN U10044 ( .A(n8036), .B(n8035), .Z(n8037) );
  AND U10045 ( .A(n8038), .B(n8037), .Z(n8056) );
  XNOR U10046 ( .A(n8057), .B(n8056), .Z(n8058) );
  NANDN U10047 ( .A(n8040), .B(n8039), .Z(n8044) );
  NAND U10048 ( .A(n8042), .B(n8041), .Z(n8043) );
  NAND U10049 ( .A(n8044), .B(n8043), .Z(n8059) );
  XNOR U10050 ( .A(n8058), .B(n8059), .Z(n8050) );
  XNOR U10051 ( .A(n8051), .B(n8050), .Z(n8052) );
  XNOR U10052 ( .A(n8053), .B(n8052), .Z(n8082) );
  XNOR U10053 ( .A(sreg[1123]), .B(n8082), .Z(n8084) );
  NANDN U10054 ( .A(sreg[1122]), .B(n8045), .Z(n8049) );
  NAND U10055 ( .A(n8047), .B(n8046), .Z(n8048) );
  NAND U10056 ( .A(n8049), .B(n8048), .Z(n8083) );
  XNOR U10057 ( .A(n8084), .B(n8083), .Z(c[1123]) );
  NANDN U10058 ( .A(n8051), .B(n8050), .Z(n8055) );
  NANDN U10059 ( .A(n8053), .B(n8052), .Z(n8054) );
  AND U10060 ( .A(n8055), .B(n8054), .Z(n8090) );
  NANDN U10061 ( .A(n8057), .B(n8056), .Z(n8061) );
  NANDN U10062 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U10063 ( .A(n8061), .B(n8060), .Z(n8088) );
  NAND U10064 ( .A(n42143), .B(n8062), .Z(n8064) );
  XNOR U10065 ( .A(a[102]), .B(n4086), .Z(n8099) );
  NAND U10066 ( .A(n42144), .B(n8099), .Z(n8063) );
  AND U10067 ( .A(n8064), .B(n8063), .Z(n8114) );
  XOR U10068 ( .A(a[106]), .B(n42012), .Z(n8102) );
  XNOR U10069 ( .A(n8114), .B(n8113), .Z(n8116) );
  AND U10070 ( .A(a[108]), .B(b[0]), .Z(n8066) );
  XNOR U10071 ( .A(n8066), .B(n4071), .Z(n8068) );
  NANDN U10072 ( .A(b[0]), .B(a[107]), .Z(n8067) );
  NAND U10073 ( .A(n8068), .B(n8067), .Z(n8110) );
  XOR U10074 ( .A(a[104]), .B(n42085), .Z(n8103) );
  AND U10075 ( .A(a[100]), .B(b[7]), .Z(n8107) );
  XNOR U10076 ( .A(n8108), .B(n8107), .Z(n8109) );
  XNOR U10077 ( .A(n8110), .B(n8109), .Z(n8115) );
  XOR U10078 ( .A(n8116), .B(n8115), .Z(n8094) );
  NANDN U10079 ( .A(n8071), .B(n8070), .Z(n8075) );
  NANDN U10080 ( .A(n8073), .B(n8072), .Z(n8074) );
  AND U10081 ( .A(n8075), .B(n8074), .Z(n8093) );
  XNOR U10082 ( .A(n8094), .B(n8093), .Z(n8095) );
  NANDN U10083 ( .A(n8077), .B(n8076), .Z(n8081) );
  NAND U10084 ( .A(n8079), .B(n8078), .Z(n8080) );
  NAND U10085 ( .A(n8081), .B(n8080), .Z(n8096) );
  XNOR U10086 ( .A(n8095), .B(n8096), .Z(n8087) );
  XNOR U10087 ( .A(n8088), .B(n8087), .Z(n8089) );
  XNOR U10088 ( .A(n8090), .B(n8089), .Z(n8119) );
  XNOR U10089 ( .A(sreg[1124]), .B(n8119), .Z(n8121) );
  NANDN U10090 ( .A(sreg[1123]), .B(n8082), .Z(n8086) );
  NAND U10091 ( .A(n8084), .B(n8083), .Z(n8085) );
  NAND U10092 ( .A(n8086), .B(n8085), .Z(n8120) );
  XNOR U10093 ( .A(n8121), .B(n8120), .Z(c[1124]) );
  NANDN U10094 ( .A(n8088), .B(n8087), .Z(n8092) );
  NANDN U10095 ( .A(n8090), .B(n8089), .Z(n8091) );
  AND U10096 ( .A(n8092), .B(n8091), .Z(n8127) );
  NANDN U10097 ( .A(n8094), .B(n8093), .Z(n8098) );
  NANDN U10098 ( .A(n8096), .B(n8095), .Z(n8097) );
  AND U10099 ( .A(n8098), .B(n8097), .Z(n8125) );
  NAND U10100 ( .A(n42143), .B(n8099), .Z(n8101) );
  XNOR U10101 ( .A(a[103]), .B(n4086), .Z(n8136) );
  NAND U10102 ( .A(n42144), .B(n8136), .Z(n8100) );
  AND U10103 ( .A(n8101), .B(n8100), .Z(n8151) );
  XOR U10104 ( .A(a[107]), .B(n42012), .Z(n8139) );
  XNOR U10105 ( .A(n8151), .B(n8150), .Z(n8153) );
  XOR U10106 ( .A(a[105]), .B(n42085), .Z(n8140) );
  AND U10107 ( .A(a[101]), .B(b[7]), .Z(n8144) );
  XNOR U10108 ( .A(n8145), .B(n8144), .Z(n8146) );
  AND U10109 ( .A(a[109]), .B(b[0]), .Z(n8104) );
  XNOR U10110 ( .A(n8104), .B(n4071), .Z(n8106) );
  NANDN U10111 ( .A(b[0]), .B(a[108]), .Z(n8105) );
  NAND U10112 ( .A(n8106), .B(n8105), .Z(n8147) );
  XNOR U10113 ( .A(n8146), .B(n8147), .Z(n8152) );
  XOR U10114 ( .A(n8153), .B(n8152), .Z(n8131) );
  NANDN U10115 ( .A(n8108), .B(n8107), .Z(n8112) );
  NANDN U10116 ( .A(n8110), .B(n8109), .Z(n8111) );
  AND U10117 ( .A(n8112), .B(n8111), .Z(n8130) );
  XNOR U10118 ( .A(n8131), .B(n8130), .Z(n8132) );
  NANDN U10119 ( .A(n8114), .B(n8113), .Z(n8118) );
  NAND U10120 ( .A(n8116), .B(n8115), .Z(n8117) );
  NAND U10121 ( .A(n8118), .B(n8117), .Z(n8133) );
  XNOR U10122 ( .A(n8132), .B(n8133), .Z(n8124) );
  XNOR U10123 ( .A(n8125), .B(n8124), .Z(n8126) );
  XNOR U10124 ( .A(n8127), .B(n8126), .Z(n8156) );
  XNOR U10125 ( .A(sreg[1125]), .B(n8156), .Z(n8158) );
  NANDN U10126 ( .A(sreg[1124]), .B(n8119), .Z(n8123) );
  NAND U10127 ( .A(n8121), .B(n8120), .Z(n8122) );
  NAND U10128 ( .A(n8123), .B(n8122), .Z(n8157) );
  XNOR U10129 ( .A(n8158), .B(n8157), .Z(c[1125]) );
  NANDN U10130 ( .A(n8125), .B(n8124), .Z(n8129) );
  NANDN U10131 ( .A(n8127), .B(n8126), .Z(n8128) );
  AND U10132 ( .A(n8129), .B(n8128), .Z(n8164) );
  NANDN U10133 ( .A(n8131), .B(n8130), .Z(n8135) );
  NANDN U10134 ( .A(n8133), .B(n8132), .Z(n8134) );
  AND U10135 ( .A(n8135), .B(n8134), .Z(n8162) );
  NAND U10136 ( .A(n42143), .B(n8136), .Z(n8138) );
  XNOR U10137 ( .A(a[104]), .B(n4086), .Z(n8173) );
  NAND U10138 ( .A(n42144), .B(n8173), .Z(n8137) );
  AND U10139 ( .A(n8138), .B(n8137), .Z(n8188) );
  XOR U10140 ( .A(a[108]), .B(n42012), .Z(n8176) );
  XNOR U10141 ( .A(n8188), .B(n8187), .Z(n8190) );
  XOR U10142 ( .A(a[106]), .B(n42085), .Z(n8177) );
  AND U10143 ( .A(a[102]), .B(b[7]), .Z(n8181) );
  XNOR U10144 ( .A(n8182), .B(n8181), .Z(n8183) );
  AND U10145 ( .A(a[110]), .B(b[0]), .Z(n8141) );
  XNOR U10146 ( .A(n8141), .B(n4071), .Z(n8143) );
  NANDN U10147 ( .A(b[0]), .B(a[109]), .Z(n8142) );
  NAND U10148 ( .A(n8143), .B(n8142), .Z(n8184) );
  XNOR U10149 ( .A(n8183), .B(n8184), .Z(n8189) );
  XOR U10150 ( .A(n8190), .B(n8189), .Z(n8168) );
  NANDN U10151 ( .A(n8145), .B(n8144), .Z(n8149) );
  NANDN U10152 ( .A(n8147), .B(n8146), .Z(n8148) );
  AND U10153 ( .A(n8149), .B(n8148), .Z(n8167) );
  XNOR U10154 ( .A(n8168), .B(n8167), .Z(n8169) );
  NANDN U10155 ( .A(n8151), .B(n8150), .Z(n8155) );
  NAND U10156 ( .A(n8153), .B(n8152), .Z(n8154) );
  NAND U10157 ( .A(n8155), .B(n8154), .Z(n8170) );
  XNOR U10158 ( .A(n8169), .B(n8170), .Z(n8161) );
  XNOR U10159 ( .A(n8162), .B(n8161), .Z(n8163) );
  XNOR U10160 ( .A(n8164), .B(n8163), .Z(n8193) );
  XNOR U10161 ( .A(sreg[1126]), .B(n8193), .Z(n8195) );
  NANDN U10162 ( .A(sreg[1125]), .B(n8156), .Z(n8160) );
  NAND U10163 ( .A(n8158), .B(n8157), .Z(n8159) );
  NAND U10164 ( .A(n8160), .B(n8159), .Z(n8194) );
  XNOR U10165 ( .A(n8195), .B(n8194), .Z(c[1126]) );
  NANDN U10166 ( .A(n8162), .B(n8161), .Z(n8166) );
  NANDN U10167 ( .A(n8164), .B(n8163), .Z(n8165) );
  AND U10168 ( .A(n8166), .B(n8165), .Z(n8201) );
  NANDN U10169 ( .A(n8168), .B(n8167), .Z(n8172) );
  NANDN U10170 ( .A(n8170), .B(n8169), .Z(n8171) );
  AND U10171 ( .A(n8172), .B(n8171), .Z(n8199) );
  NAND U10172 ( .A(n42143), .B(n8173), .Z(n8175) );
  XNOR U10173 ( .A(a[105]), .B(n4086), .Z(n8210) );
  NAND U10174 ( .A(n42144), .B(n8210), .Z(n8174) );
  AND U10175 ( .A(n8175), .B(n8174), .Z(n8225) );
  XOR U10176 ( .A(a[109]), .B(n42012), .Z(n8213) );
  XNOR U10177 ( .A(n8225), .B(n8224), .Z(n8227) );
  XOR U10178 ( .A(a[107]), .B(n42085), .Z(n8217) );
  AND U10179 ( .A(a[103]), .B(b[7]), .Z(n8218) );
  XNOR U10180 ( .A(n8219), .B(n8218), .Z(n8220) );
  AND U10181 ( .A(a[111]), .B(b[0]), .Z(n8178) );
  XNOR U10182 ( .A(n8178), .B(n4071), .Z(n8180) );
  NANDN U10183 ( .A(b[0]), .B(a[110]), .Z(n8179) );
  NAND U10184 ( .A(n8180), .B(n8179), .Z(n8221) );
  XNOR U10185 ( .A(n8220), .B(n8221), .Z(n8226) );
  XOR U10186 ( .A(n8227), .B(n8226), .Z(n8205) );
  NANDN U10187 ( .A(n8182), .B(n8181), .Z(n8186) );
  NANDN U10188 ( .A(n8184), .B(n8183), .Z(n8185) );
  AND U10189 ( .A(n8186), .B(n8185), .Z(n8204) );
  XNOR U10190 ( .A(n8205), .B(n8204), .Z(n8206) );
  NANDN U10191 ( .A(n8188), .B(n8187), .Z(n8192) );
  NAND U10192 ( .A(n8190), .B(n8189), .Z(n8191) );
  NAND U10193 ( .A(n8192), .B(n8191), .Z(n8207) );
  XNOR U10194 ( .A(n8206), .B(n8207), .Z(n8198) );
  XNOR U10195 ( .A(n8199), .B(n8198), .Z(n8200) );
  XNOR U10196 ( .A(n8201), .B(n8200), .Z(n8230) );
  XNOR U10197 ( .A(sreg[1127]), .B(n8230), .Z(n8232) );
  NANDN U10198 ( .A(sreg[1126]), .B(n8193), .Z(n8197) );
  NAND U10199 ( .A(n8195), .B(n8194), .Z(n8196) );
  NAND U10200 ( .A(n8197), .B(n8196), .Z(n8231) );
  XNOR U10201 ( .A(n8232), .B(n8231), .Z(c[1127]) );
  NANDN U10202 ( .A(n8199), .B(n8198), .Z(n8203) );
  NANDN U10203 ( .A(n8201), .B(n8200), .Z(n8202) );
  AND U10204 ( .A(n8203), .B(n8202), .Z(n8238) );
  NANDN U10205 ( .A(n8205), .B(n8204), .Z(n8209) );
  NANDN U10206 ( .A(n8207), .B(n8206), .Z(n8208) );
  AND U10207 ( .A(n8209), .B(n8208), .Z(n8236) );
  NAND U10208 ( .A(n42143), .B(n8210), .Z(n8212) );
  XNOR U10209 ( .A(a[106]), .B(n4087), .Z(n8247) );
  NAND U10210 ( .A(n42144), .B(n8247), .Z(n8211) );
  AND U10211 ( .A(n8212), .B(n8211), .Z(n8262) );
  XOR U10212 ( .A(a[110]), .B(n42012), .Z(n8250) );
  XNOR U10213 ( .A(n8262), .B(n8261), .Z(n8264) );
  AND U10214 ( .A(a[112]), .B(b[0]), .Z(n8214) );
  XNOR U10215 ( .A(n8214), .B(n4071), .Z(n8216) );
  NANDN U10216 ( .A(b[0]), .B(a[111]), .Z(n8215) );
  NAND U10217 ( .A(n8216), .B(n8215), .Z(n8258) );
  XOR U10218 ( .A(a[108]), .B(n42085), .Z(n8251) );
  AND U10219 ( .A(a[104]), .B(b[7]), .Z(n8255) );
  XNOR U10220 ( .A(n8256), .B(n8255), .Z(n8257) );
  XNOR U10221 ( .A(n8258), .B(n8257), .Z(n8263) );
  XOR U10222 ( .A(n8264), .B(n8263), .Z(n8242) );
  NANDN U10223 ( .A(n8219), .B(n8218), .Z(n8223) );
  NANDN U10224 ( .A(n8221), .B(n8220), .Z(n8222) );
  AND U10225 ( .A(n8223), .B(n8222), .Z(n8241) );
  XNOR U10226 ( .A(n8242), .B(n8241), .Z(n8243) );
  NANDN U10227 ( .A(n8225), .B(n8224), .Z(n8229) );
  NAND U10228 ( .A(n8227), .B(n8226), .Z(n8228) );
  NAND U10229 ( .A(n8229), .B(n8228), .Z(n8244) );
  XNOR U10230 ( .A(n8243), .B(n8244), .Z(n8235) );
  XNOR U10231 ( .A(n8236), .B(n8235), .Z(n8237) );
  XNOR U10232 ( .A(n8238), .B(n8237), .Z(n8267) );
  XNOR U10233 ( .A(sreg[1128]), .B(n8267), .Z(n8269) );
  NANDN U10234 ( .A(sreg[1127]), .B(n8230), .Z(n8234) );
  NAND U10235 ( .A(n8232), .B(n8231), .Z(n8233) );
  NAND U10236 ( .A(n8234), .B(n8233), .Z(n8268) );
  XNOR U10237 ( .A(n8269), .B(n8268), .Z(c[1128]) );
  NANDN U10238 ( .A(n8236), .B(n8235), .Z(n8240) );
  NANDN U10239 ( .A(n8238), .B(n8237), .Z(n8239) );
  AND U10240 ( .A(n8240), .B(n8239), .Z(n8275) );
  NANDN U10241 ( .A(n8242), .B(n8241), .Z(n8246) );
  NANDN U10242 ( .A(n8244), .B(n8243), .Z(n8245) );
  AND U10243 ( .A(n8246), .B(n8245), .Z(n8273) );
  NAND U10244 ( .A(n42143), .B(n8247), .Z(n8249) );
  XNOR U10245 ( .A(a[107]), .B(n4087), .Z(n8284) );
  NAND U10246 ( .A(n42144), .B(n8284), .Z(n8248) );
  AND U10247 ( .A(n8249), .B(n8248), .Z(n8299) );
  XOR U10248 ( .A(a[111]), .B(n42012), .Z(n8287) );
  XNOR U10249 ( .A(n8299), .B(n8298), .Z(n8301) );
  XOR U10250 ( .A(a[109]), .B(n42085), .Z(n8291) );
  AND U10251 ( .A(a[105]), .B(b[7]), .Z(n8292) );
  XNOR U10252 ( .A(n8293), .B(n8292), .Z(n8294) );
  AND U10253 ( .A(a[113]), .B(b[0]), .Z(n8252) );
  XNOR U10254 ( .A(n8252), .B(n4071), .Z(n8254) );
  NANDN U10255 ( .A(b[0]), .B(a[112]), .Z(n8253) );
  NAND U10256 ( .A(n8254), .B(n8253), .Z(n8295) );
  XNOR U10257 ( .A(n8294), .B(n8295), .Z(n8300) );
  XOR U10258 ( .A(n8301), .B(n8300), .Z(n8279) );
  NANDN U10259 ( .A(n8256), .B(n8255), .Z(n8260) );
  NANDN U10260 ( .A(n8258), .B(n8257), .Z(n8259) );
  AND U10261 ( .A(n8260), .B(n8259), .Z(n8278) );
  XNOR U10262 ( .A(n8279), .B(n8278), .Z(n8280) );
  NANDN U10263 ( .A(n8262), .B(n8261), .Z(n8266) );
  NAND U10264 ( .A(n8264), .B(n8263), .Z(n8265) );
  NAND U10265 ( .A(n8266), .B(n8265), .Z(n8281) );
  XNOR U10266 ( .A(n8280), .B(n8281), .Z(n8272) );
  XNOR U10267 ( .A(n8273), .B(n8272), .Z(n8274) );
  XNOR U10268 ( .A(n8275), .B(n8274), .Z(n8304) );
  XNOR U10269 ( .A(sreg[1129]), .B(n8304), .Z(n8306) );
  NANDN U10270 ( .A(sreg[1128]), .B(n8267), .Z(n8271) );
  NAND U10271 ( .A(n8269), .B(n8268), .Z(n8270) );
  NAND U10272 ( .A(n8271), .B(n8270), .Z(n8305) );
  XNOR U10273 ( .A(n8306), .B(n8305), .Z(c[1129]) );
  NANDN U10274 ( .A(n8273), .B(n8272), .Z(n8277) );
  NANDN U10275 ( .A(n8275), .B(n8274), .Z(n8276) );
  AND U10276 ( .A(n8277), .B(n8276), .Z(n8312) );
  NANDN U10277 ( .A(n8279), .B(n8278), .Z(n8283) );
  NANDN U10278 ( .A(n8281), .B(n8280), .Z(n8282) );
  AND U10279 ( .A(n8283), .B(n8282), .Z(n8310) );
  NAND U10280 ( .A(n42143), .B(n8284), .Z(n8286) );
  XNOR U10281 ( .A(a[108]), .B(n4087), .Z(n8321) );
  NAND U10282 ( .A(n42144), .B(n8321), .Z(n8285) );
  AND U10283 ( .A(n8286), .B(n8285), .Z(n8336) );
  XOR U10284 ( .A(a[112]), .B(n42012), .Z(n8324) );
  XNOR U10285 ( .A(n8336), .B(n8335), .Z(n8338) );
  AND U10286 ( .A(a[114]), .B(b[0]), .Z(n8288) );
  XNOR U10287 ( .A(n8288), .B(n4071), .Z(n8290) );
  NANDN U10288 ( .A(b[0]), .B(a[113]), .Z(n8289) );
  NAND U10289 ( .A(n8290), .B(n8289), .Z(n8332) );
  XOR U10290 ( .A(a[110]), .B(n42085), .Z(n8328) );
  AND U10291 ( .A(a[106]), .B(b[7]), .Z(n8329) );
  XNOR U10292 ( .A(n8330), .B(n8329), .Z(n8331) );
  XNOR U10293 ( .A(n8332), .B(n8331), .Z(n8337) );
  XOR U10294 ( .A(n8338), .B(n8337), .Z(n8316) );
  NANDN U10295 ( .A(n8293), .B(n8292), .Z(n8297) );
  NANDN U10296 ( .A(n8295), .B(n8294), .Z(n8296) );
  AND U10297 ( .A(n8297), .B(n8296), .Z(n8315) );
  XNOR U10298 ( .A(n8316), .B(n8315), .Z(n8317) );
  NANDN U10299 ( .A(n8299), .B(n8298), .Z(n8303) );
  NAND U10300 ( .A(n8301), .B(n8300), .Z(n8302) );
  NAND U10301 ( .A(n8303), .B(n8302), .Z(n8318) );
  XNOR U10302 ( .A(n8317), .B(n8318), .Z(n8309) );
  XNOR U10303 ( .A(n8310), .B(n8309), .Z(n8311) );
  XNOR U10304 ( .A(n8312), .B(n8311), .Z(n8341) );
  XNOR U10305 ( .A(sreg[1130]), .B(n8341), .Z(n8343) );
  NANDN U10306 ( .A(sreg[1129]), .B(n8304), .Z(n8308) );
  NAND U10307 ( .A(n8306), .B(n8305), .Z(n8307) );
  NAND U10308 ( .A(n8308), .B(n8307), .Z(n8342) );
  XNOR U10309 ( .A(n8343), .B(n8342), .Z(c[1130]) );
  NANDN U10310 ( .A(n8310), .B(n8309), .Z(n8314) );
  NANDN U10311 ( .A(n8312), .B(n8311), .Z(n8313) );
  AND U10312 ( .A(n8314), .B(n8313), .Z(n8349) );
  NANDN U10313 ( .A(n8316), .B(n8315), .Z(n8320) );
  NANDN U10314 ( .A(n8318), .B(n8317), .Z(n8319) );
  AND U10315 ( .A(n8320), .B(n8319), .Z(n8347) );
  NAND U10316 ( .A(n42143), .B(n8321), .Z(n8323) );
  XNOR U10317 ( .A(a[109]), .B(n4087), .Z(n8358) );
  NAND U10318 ( .A(n42144), .B(n8358), .Z(n8322) );
  AND U10319 ( .A(n8323), .B(n8322), .Z(n8373) );
  XOR U10320 ( .A(a[113]), .B(n42012), .Z(n8361) );
  XNOR U10321 ( .A(n8373), .B(n8372), .Z(n8375) );
  AND U10322 ( .A(a[115]), .B(b[0]), .Z(n8325) );
  XNOR U10323 ( .A(n8325), .B(n4071), .Z(n8327) );
  NANDN U10324 ( .A(b[0]), .B(a[114]), .Z(n8326) );
  NAND U10325 ( .A(n8327), .B(n8326), .Z(n8369) );
  XOR U10326 ( .A(a[111]), .B(n42085), .Z(n8365) );
  AND U10327 ( .A(a[107]), .B(b[7]), .Z(n8366) );
  XNOR U10328 ( .A(n8367), .B(n8366), .Z(n8368) );
  XNOR U10329 ( .A(n8369), .B(n8368), .Z(n8374) );
  XOR U10330 ( .A(n8375), .B(n8374), .Z(n8353) );
  NANDN U10331 ( .A(n8330), .B(n8329), .Z(n8334) );
  NANDN U10332 ( .A(n8332), .B(n8331), .Z(n8333) );
  AND U10333 ( .A(n8334), .B(n8333), .Z(n8352) );
  XNOR U10334 ( .A(n8353), .B(n8352), .Z(n8354) );
  NANDN U10335 ( .A(n8336), .B(n8335), .Z(n8340) );
  NAND U10336 ( .A(n8338), .B(n8337), .Z(n8339) );
  NAND U10337 ( .A(n8340), .B(n8339), .Z(n8355) );
  XNOR U10338 ( .A(n8354), .B(n8355), .Z(n8346) );
  XNOR U10339 ( .A(n8347), .B(n8346), .Z(n8348) );
  XNOR U10340 ( .A(n8349), .B(n8348), .Z(n8378) );
  XNOR U10341 ( .A(sreg[1131]), .B(n8378), .Z(n8380) );
  NANDN U10342 ( .A(sreg[1130]), .B(n8341), .Z(n8345) );
  NAND U10343 ( .A(n8343), .B(n8342), .Z(n8344) );
  NAND U10344 ( .A(n8345), .B(n8344), .Z(n8379) );
  XNOR U10345 ( .A(n8380), .B(n8379), .Z(c[1131]) );
  NANDN U10346 ( .A(n8347), .B(n8346), .Z(n8351) );
  NANDN U10347 ( .A(n8349), .B(n8348), .Z(n8350) );
  AND U10348 ( .A(n8351), .B(n8350), .Z(n8386) );
  NANDN U10349 ( .A(n8353), .B(n8352), .Z(n8357) );
  NANDN U10350 ( .A(n8355), .B(n8354), .Z(n8356) );
  AND U10351 ( .A(n8357), .B(n8356), .Z(n8384) );
  NAND U10352 ( .A(n42143), .B(n8358), .Z(n8360) );
  XNOR U10353 ( .A(a[110]), .B(n4087), .Z(n8395) );
  NAND U10354 ( .A(n42144), .B(n8395), .Z(n8359) );
  AND U10355 ( .A(n8360), .B(n8359), .Z(n8410) );
  XOR U10356 ( .A(a[114]), .B(n42012), .Z(n8398) );
  XNOR U10357 ( .A(n8410), .B(n8409), .Z(n8412) );
  AND U10358 ( .A(a[116]), .B(b[0]), .Z(n8362) );
  XNOR U10359 ( .A(n8362), .B(n4071), .Z(n8364) );
  NANDN U10360 ( .A(b[0]), .B(a[115]), .Z(n8363) );
  NAND U10361 ( .A(n8364), .B(n8363), .Z(n8406) );
  XOR U10362 ( .A(a[112]), .B(n42085), .Z(n8402) );
  AND U10363 ( .A(a[108]), .B(b[7]), .Z(n8403) );
  XNOR U10364 ( .A(n8404), .B(n8403), .Z(n8405) );
  XNOR U10365 ( .A(n8406), .B(n8405), .Z(n8411) );
  XOR U10366 ( .A(n8412), .B(n8411), .Z(n8390) );
  NANDN U10367 ( .A(n8367), .B(n8366), .Z(n8371) );
  NANDN U10368 ( .A(n8369), .B(n8368), .Z(n8370) );
  AND U10369 ( .A(n8371), .B(n8370), .Z(n8389) );
  XNOR U10370 ( .A(n8390), .B(n8389), .Z(n8391) );
  NANDN U10371 ( .A(n8373), .B(n8372), .Z(n8377) );
  NAND U10372 ( .A(n8375), .B(n8374), .Z(n8376) );
  NAND U10373 ( .A(n8377), .B(n8376), .Z(n8392) );
  XNOR U10374 ( .A(n8391), .B(n8392), .Z(n8383) );
  XNOR U10375 ( .A(n8384), .B(n8383), .Z(n8385) );
  XNOR U10376 ( .A(n8386), .B(n8385), .Z(n8415) );
  XNOR U10377 ( .A(sreg[1132]), .B(n8415), .Z(n8417) );
  NANDN U10378 ( .A(sreg[1131]), .B(n8378), .Z(n8382) );
  NAND U10379 ( .A(n8380), .B(n8379), .Z(n8381) );
  NAND U10380 ( .A(n8382), .B(n8381), .Z(n8416) );
  XNOR U10381 ( .A(n8417), .B(n8416), .Z(c[1132]) );
  NANDN U10382 ( .A(n8384), .B(n8383), .Z(n8388) );
  NANDN U10383 ( .A(n8386), .B(n8385), .Z(n8387) );
  AND U10384 ( .A(n8388), .B(n8387), .Z(n8423) );
  NANDN U10385 ( .A(n8390), .B(n8389), .Z(n8394) );
  NANDN U10386 ( .A(n8392), .B(n8391), .Z(n8393) );
  AND U10387 ( .A(n8394), .B(n8393), .Z(n8421) );
  NAND U10388 ( .A(n42143), .B(n8395), .Z(n8397) );
  XNOR U10389 ( .A(a[111]), .B(n4087), .Z(n8432) );
  NAND U10390 ( .A(n42144), .B(n8432), .Z(n8396) );
  AND U10391 ( .A(n8397), .B(n8396), .Z(n8447) );
  XOR U10392 ( .A(a[115]), .B(n42012), .Z(n8435) );
  XNOR U10393 ( .A(n8447), .B(n8446), .Z(n8449) );
  AND U10394 ( .A(a[117]), .B(b[0]), .Z(n8399) );
  XNOR U10395 ( .A(n8399), .B(n4071), .Z(n8401) );
  NANDN U10396 ( .A(b[0]), .B(a[116]), .Z(n8400) );
  NAND U10397 ( .A(n8401), .B(n8400), .Z(n8443) );
  XOR U10398 ( .A(a[113]), .B(n42085), .Z(n8439) );
  AND U10399 ( .A(a[109]), .B(b[7]), .Z(n8440) );
  XNOR U10400 ( .A(n8441), .B(n8440), .Z(n8442) );
  XNOR U10401 ( .A(n8443), .B(n8442), .Z(n8448) );
  XOR U10402 ( .A(n8449), .B(n8448), .Z(n8427) );
  NANDN U10403 ( .A(n8404), .B(n8403), .Z(n8408) );
  NANDN U10404 ( .A(n8406), .B(n8405), .Z(n8407) );
  AND U10405 ( .A(n8408), .B(n8407), .Z(n8426) );
  XNOR U10406 ( .A(n8427), .B(n8426), .Z(n8428) );
  NANDN U10407 ( .A(n8410), .B(n8409), .Z(n8414) );
  NAND U10408 ( .A(n8412), .B(n8411), .Z(n8413) );
  NAND U10409 ( .A(n8414), .B(n8413), .Z(n8429) );
  XNOR U10410 ( .A(n8428), .B(n8429), .Z(n8420) );
  XNOR U10411 ( .A(n8421), .B(n8420), .Z(n8422) );
  XNOR U10412 ( .A(n8423), .B(n8422), .Z(n8452) );
  XNOR U10413 ( .A(sreg[1133]), .B(n8452), .Z(n8454) );
  NANDN U10414 ( .A(sreg[1132]), .B(n8415), .Z(n8419) );
  NAND U10415 ( .A(n8417), .B(n8416), .Z(n8418) );
  NAND U10416 ( .A(n8419), .B(n8418), .Z(n8453) );
  XNOR U10417 ( .A(n8454), .B(n8453), .Z(c[1133]) );
  NANDN U10418 ( .A(n8421), .B(n8420), .Z(n8425) );
  NANDN U10419 ( .A(n8423), .B(n8422), .Z(n8424) );
  AND U10420 ( .A(n8425), .B(n8424), .Z(n8460) );
  NANDN U10421 ( .A(n8427), .B(n8426), .Z(n8431) );
  NANDN U10422 ( .A(n8429), .B(n8428), .Z(n8430) );
  AND U10423 ( .A(n8431), .B(n8430), .Z(n8458) );
  NAND U10424 ( .A(n42143), .B(n8432), .Z(n8434) );
  XNOR U10425 ( .A(a[112]), .B(n4087), .Z(n8469) );
  NAND U10426 ( .A(n42144), .B(n8469), .Z(n8433) );
  AND U10427 ( .A(n8434), .B(n8433), .Z(n8484) );
  XOR U10428 ( .A(a[116]), .B(n42012), .Z(n8472) );
  XNOR U10429 ( .A(n8484), .B(n8483), .Z(n8486) );
  AND U10430 ( .A(b[0]), .B(a[118]), .Z(n8436) );
  XOR U10431 ( .A(b[1]), .B(n8436), .Z(n8438) );
  NANDN U10432 ( .A(b[0]), .B(a[117]), .Z(n8437) );
  AND U10433 ( .A(n8438), .B(n8437), .Z(n8479) );
  XOR U10434 ( .A(a[114]), .B(n42085), .Z(n8476) );
  AND U10435 ( .A(a[110]), .B(b[7]), .Z(n8477) );
  XOR U10436 ( .A(n8478), .B(n8477), .Z(n8480) );
  XNOR U10437 ( .A(n8479), .B(n8480), .Z(n8485) );
  XOR U10438 ( .A(n8486), .B(n8485), .Z(n8464) );
  NANDN U10439 ( .A(n8441), .B(n8440), .Z(n8445) );
  NANDN U10440 ( .A(n8443), .B(n8442), .Z(n8444) );
  AND U10441 ( .A(n8445), .B(n8444), .Z(n8463) );
  XNOR U10442 ( .A(n8464), .B(n8463), .Z(n8465) );
  NANDN U10443 ( .A(n8447), .B(n8446), .Z(n8451) );
  NAND U10444 ( .A(n8449), .B(n8448), .Z(n8450) );
  NAND U10445 ( .A(n8451), .B(n8450), .Z(n8466) );
  XNOR U10446 ( .A(n8465), .B(n8466), .Z(n8457) );
  XNOR U10447 ( .A(n8458), .B(n8457), .Z(n8459) );
  XNOR U10448 ( .A(n8460), .B(n8459), .Z(n8489) );
  XNOR U10449 ( .A(sreg[1134]), .B(n8489), .Z(n8491) );
  NANDN U10450 ( .A(sreg[1133]), .B(n8452), .Z(n8456) );
  NAND U10451 ( .A(n8454), .B(n8453), .Z(n8455) );
  NAND U10452 ( .A(n8456), .B(n8455), .Z(n8490) );
  XNOR U10453 ( .A(n8491), .B(n8490), .Z(c[1134]) );
  NANDN U10454 ( .A(n8458), .B(n8457), .Z(n8462) );
  NANDN U10455 ( .A(n8460), .B(n8459), .Z(n8461) );
  AND U10456 ( .A(n8462), .B(n8461), .Z(n8497) );
  NANDN U10457 ( .A(n8464), .B(n8463), .Z(n8468) );
  NANDN U10458 ( .A(n8466), .B(n8465), .Z(n8467) );
  AND U10459 ( .A(n8468), .B(n8467), .Z(n8495) );
  NAND U10460 ( .A(n42143), .B(n8469), .Z(n8471) );
  XNOR U10461 ( .A(a[113]), .B(n4088), .Z(n8506) );
  NAND U10462 ( .A(n42144), .B(n8506), .Z(n8470) );
  AND U10463 ( .A(n8471), .B(n8470), .Z(n8521) );
  XOR U10464 ( .A(a[117]), .B(n42012), .Z(n8509) );
  XNOR U10465 ( .A(n8521), .B(n8520), .Z(n8523) );
  AND U10466 ( .A(a[119]), .B(b[0]), .Z(n8473) );
  XNOR U10467 ( .A(n8473), .B(n4071), .Z(n8475) );
  NANDN U10468 ( .A(b[0]), .B(a[118]), .Z(n8474) );
  NAND U10469 ( .A(n8475), .B(n8474), .Z(n8517) );
  XOR U10470 ( .A(a[115]), .B(n42085), .Z(n8513) );
  AND U10471 ( .A(a[111]), .B(b[7]), .Z(n8514) );
  XNOR U10472 ( .A(n8515), .B(n8514), .Z(n8516) );
  XNOR U10473 ( .A(n8517), .B(n8516), .Z(n8522) );
  XOR U10474 ( .A(n8523), .B(n8522), .Z(n8501) );
  NANDN U10475 ( .A(n8478), .B(n8477), .Z(n8482) );
  NANDN U10476 ( .A(n8480), .B(n8479), .Z(n8481) );
  AND U10477 ( .A(n8482), .B(n8481), .Z(n8500) );
  XNOR U10478 ( .A(n8501), .B(n8500), .Z(n8502) );
  NANDN U10479 ( .A(n8484), .B(n8483), .Z(n8488) );
  NAND U10480 ( .A(n8486), .B(n8485), .Z(n8487) );
  NAND U10481 ( .A(n8488), .B(n8487), .Z(n8503) );
  XNOR U10482 ( .A(n8502), .B(n8503), .Z(n8494) );
  XNOR U10483 ( .A(n8495), .B(n8494), .Z(n8496) );
  XNOR U10484 ( .A(n8497), .B(n8496), .Z(n8526) );
  XNOR U10485 ( .A(sreg[1135]), .B(n8526), .Z(n8528) );
  NANDN U10486 ( .A(sreg[1134]), .B(n8489), .Z(n8493) );
  NAND U10487 ( .A(n8491), .B(n8490), .Z(n8492) );
  NAND U10488 ( .A(n8493), .B(n8492), .Z(n8527) );
  XNOR U10489 ( .A(n8528), .B(n8527), .Z(c[1135]) );
  NANDN U10490 ( .A(n8495), .B(n8494), .Z(n8499) );
  NANDN U10491 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U10492 ( .A(n8499), .B(n8498), .Z(n8534) );
  NANDN U10493 ( .A(n8501), .B(n8500), .Z(n8505) );
  NANDN U10494 ( .A(n8503), .B(n8502), .Z(n8504) );
  AND U10495 ( .A(n8505), .B(n8504), .Z(n8532) );
  NAND U10496 ( .A(n42143), .B(n8506), .Z(n8508) );
  XNOR U10497 ( .A(a[114]), .B(n4088), .Z(n8543) );
  NAND U10498 ( .A(n42144), .B(n8543), .Z(n8507) );
  AND U10499 ( .A(n8508), .B(n8507), .Z(n8558) );
  XOR U10500 ( .A(a[118]), .B(n42012), .Z(n8546) );
  XNOR U10501 ( .A(n8558), .B(n8557), .Z(n8560) );
  AND U10502 ( .A(a[120]), .B(b[0]), .Z(n8510) );
  XNOR U10503 ( .A(n8510), .B(n4071), .Z(n8512) );
  NANDN U10504 ( .A(b[0]), .B(a[119]), .Z(n8511) );
  NAND U10505 ( .A(n8512), .B(n8511), .Z(n8554) );
  XOR U10506 ( .A(a[116]), .B(n42085), .Z(n8547) );
  AND U10507 ( .A(a[112]), .B(b[7]), .Z(n8551) );
  XNOR U10508 ( .A(n8552), .B(n8551), .Z(n8553) );
  XNOR U10509 ( .A(n8554), .B(n8553), .Z(n8559) );
  XOR U10510 ( .A(n8560), .B(n8559), .Z(n8538) );
  NANDN U10511 ( .A(n8515), .B(n8514), .Z(n8519) );
  NANDN U10512 ( .A(n8517), .B(n8516), .Z(n8518) );
  AND U10513 ( .A(n8519), .B(n8518), .Z(n8537) );
  XNOR U10514 ( .A(n8538), .B(n8537), .Z(n8539) );
  NANDN U10515 ( .A(n8521), .B(n8520), .Z(n8525) );
  NAND U10516 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U10517 ( .A(n8525), .B(n8524), .Z(n8540) );
  XNOR U10518 ( .A(n8539), .B(n8540), .Z(n8531) );
  XNOR U10519 ( .A(n8532), .B(n8531), .Z(n8533) );
  XNOR U10520 ( .A(n8534), .B(n8533), .Z(n8563) );
  XNOR U10521 ( .A(sreg[1136]), .B(n8563), .Z(n8565) );
  NANDN U10522 ( .A(sreg[1135]), .B(n8526), .Z(n8530) );
  NAND U10523 ( .A(n8528), .B(n8527), .Z(n8529) );
  NAND U10524 ( .A(n8530), .B(n8529), .Z(n8564) );
  XNOR U10525 ( .A(n8565), .B(n8564), .Z(c[1136]) );
  NANDN U10526 ( .A(n8532), .B(n8531), .Z(n8536) );
  NANDN U10527 ( .A(n8534), .B(n8533), .Z(n8535) );
  AND U10528 ( .A(n8536), .B(n8535), .Z(n8571) );
  NANDN U10529 ( .A(n8538), .B(n8537), .Z(n8542) );
  NANDN U10530 ( .A(n8540), .B(n8539), .Z(n8541) );
  AND U10531 ( .A(n8542), .B(n8541), .Z(n8569) );
  NAND U10532 ( .A(n42143), .B(n8543), .Z(n8545) );
  XNOR U10533 ( .A(a[115]), .B(n4088), .Z(n8580) );
  NAND U10534 ( .A(n42144), .B(n8580), .Z(n8544) );
  AND U10535 ( .A(n8545), .B(n8544), .Z(n8595) );
  XOR U10536 ( .A(a[119]), .B(n42012), .Z(n8583) );
  XNOR U10537 ( .A(n8595), .B(n8594), .Z(n8597) );
  XOR U10538 ( .A(a[117]), .B(n42085), .Z(n8587) );
  AND U10539 ( .A(a[113]), .B(b[7]), .Z(n8588) );
  XNOR U10540 ( .A(n8589), .B(n8588), .Z(n8590) );
  AND U10541 ( .A(a[121]), .B(b[0]), .Z(n8548) );
  XNOR U10542 ( .A(n8548), .B(n4071), .Z(n8550) );
  NANDN U10543 ( .A(b[0]), .B(a[120]), .Z(n8549) );
  NAND U10544 ( .A(n8550), .B(n8549), .Z(n8591) );
  XNOR U10545 ( .A(n8590), .B(n8591), .Z(n8596) );
  XOR U10546 ( .A(n8597), .B(n8596), .Z(n8575) );
  NANDN U10547 ( .A(n8552), .B(n8551), .Z(n8556) );
  NANDN U10548 ( .A(n8554), .B(n8553), .Z(n8555) );
  AND U10549 ( .A(n8556), .B(n8555), .Z(n8574) );
  XNOR U10550 ( .A(n8575), .B(n8574), .Z(n8576) );
  NANDN U10551 ( .A(n8558), .B(n8557), .Z(n8562) );
  NAND U10552 ( .A(n8560), .B(n8559), .Z(n8561) );
  NAND U10553 ( .A(n8562), .B(n8561), .Z(n8577) );
  XNOR U10554 ( .A(n8576), .B(n8577), .Z(n8568) );
  XNOR U10555 ( .A(n8569), .B(n8568), .Z(n8570) );
  XNOR U10556 ( .A(n8571), .B(n8570), .Z(n8600) );
  XNOR U10557 ( .A(sreg[1137]), .B(n8600), .Z(n8602) );
  NANDN U10558 ( .A(sreg[1136]), .B(n8563), .Z(n8567) );
  NAND U10559 ( .A(n8565), .B(n8564), .Z(n8566) );
  NAND U10560 ( .A(n8567), .B(n8566), .Z(n8601) );
  XNOR U10561 ( .A(n8602), .B(n8601), .Z(c[1137]) );
  NANDN U10562 ( .A(n8569), .B(n8568), .Z(n8573) );
  NANDN U10563 ( .A(n8571), .B(n8570), .Z(n8572) );
  AND U10564 ( .A(n8573), .B(n8572), .Z(n8608) );
  NANDN U10565 ( .A(n8575), .B(n8574), .Z(n8579) );
  NANDN U10566 ( .A(n8577), .B(n8576), .Z(n8578) );
  AND U10567 ( .A(n8579), .B(n8578), .Z(n8606) );
  NAND U10568 ( .A(n42143), .B(n8580), .Z(n8582) );
  XNOR U10569 ( .A(a[116]), .B(n4088), .Z(n8617) );
  NAND U10570 ( .A(n42144), .B(n8617), .Z(n8581) );
  AND U10571 ( .A(n8582), .B(n8581), .Z(n8632) );
  XOR U10572 ( .A(a[120]), .B(n42012), .Z(n8620) );
  XNOR U10573 ( .A(n8632), .B(n8631), .Z(n8634) );
  AND U10574 ( .A(a[122]), .B(b[0]), .Z(n8584) );
  XNOR U10575 ( .A(n8584), .B(n4071), .Z(n8586) );
  NANDN U10576 ( .A(b[0]), .B(a[121]), .Z(n8585) );
  NAND U10577 ( .A(n8586), .B(n8585), .Z(n8628) );
  XOR U10578 ( .A(a[118]), .B(n42085), .Z(n8624) );
  AND U10579 ( .A(a[114]), .B(b[7]), .Z(n8625) );
  XNOR U10580 ( .A(n8626), .B(n8625), .Z(n8627) );
  XNOR U10581 ( .A(n8628), .B(n8627), .Z(n8633) );
  XOR U10582 ( .A(n8634), .B(n8633), .Z(n8612) );
  NANDN U10583 ( .A(n8589), .B(n8588), .Z(n8593) );
  NANDN U10584 ( .A(n8591), .B(n8590), .Z(n8592) );
  AND U10585 ( .A(n8593), .B(n8592), .Z(n8611) );
  XNOR U10586 ( .A(n8612), .B(n8611), .Z(n8613) );
  NANDN U10587 ( .A(n8595), .B(n8594), .Z(n8599) );
  NAND U10588 ( .A(n8597), .B(n8596), .Z(n8598) );
  NAND U10589 ( .A(n8599), .B(n8598), .Z(n8614) );
  XNOR U10590 ( .A(n8613), .B(n8614), .Z(n8605) );
  XNOR U10591 ( .A(n8606), .B(n8605), .Z(n8607) );
  XNOR U10592 ( .A(n8608), .B(n8607), .Z(n8637) );
  XNOR U10593 ( .A(sreg[1138]), .B(n8637), .Z(n8639) );
  NANDN U10594 ( .A(sreg[1137]), .B(n8600), .Z(n8604) );
  NAND U10595 ( .A(n8602), .B(n8601), .Z(n8603) );
  NAND U10596 ( .A(n8604), .B(n8603), .Z(n8638) );
  XNOR U10597 ( .A(n8639), .B(n8638), .Z(c[1138]) );
  NANDN U10598 ( .A(n8606), .B(n8605), .Z(n8610) );
  NANDN U10599 ( .A(n8608), .B(n8607), .Z(n8609) );
  AND U10600 ( .A(n8610), .B(n8609), .Z(n8645) );
  NANDN U10601 ( .A(n8612), .B(n8611), .Z(n8616) );
  NANDN U10602 ( .A(n8614), .B(n8613), .Z(n8615) );
  AND U10603 ( .A(n8616), .B(n8615), .Z(n8643) );
  NAND U10604 ( .A(n42143), .B(n8617), .Z(n8619) );
  XNOR U10605 ( .A(a[117]), .B(n4088), .Z(n8654) );
  NAND U10606 ( .A(n42144), .B(n8654), .Z(n8618) );
  AND U10607 ( .A(n8619), .B(n8618), .Z(n8669) );
  XOR U10608 ( .A(a[121]), .B(n42012), .Z(n8657) );
  XNOR U10609 ( .A(n8669), .B(n8668), .Z(n8671) );
  AND U10610 ( .A(a[123]), .B(b[0]), .Z(n8621) );
  XNOR U10611 ( .A(n8621), .B(n4071), .Z(n8623) );
  NANDN U10612 ( .A(b[0]), .B(a[122]), .Z(n8622) );
  NAND U10613 ( .A(n8623), .B(n8622), .Z(n8665) );
  XOR U10614 ( .A(a[119]), .B(n42085), .Z(n8661) );
  AND U10615 ( .A(a[115]), .B(b[7]), .Z(n8662) );
  XNOR U10616 ( .A(n8663), .B(n8662), .Z(n8664) );
  XNOR U10617 ( .A(n8665), .B(n8664), .Z(n8670) );
  XOR U10618 ( .A(n8671), .B(n8670), .Z(n8649) );
  NANDN U10619 ( .A(n8626), .B(n8625), .Z(n8630) );
  NANDN U10620 ( .A(n8628), .B(n8627), .Z(n8629) );
  AND U10621 ( .A(n8630), .B(n8629), .Z(n8648) );
  XNOR U10622 ( .A(n8649), .B(n8648), .Z(n8650) );
  NANDN U10623 ( .A(n8632), .B(n8631), .Z(n8636) );
  NAND U10624 ( .A(n8634), .B(n8633), .Z(n8635) );
  NAND U10625 ( .A(n8636), .B(n8635), .Z(n8651) );
  XNOR U10626 ( .A(n8650), .B(n8651), .Z(n8642) );
  XNOR U10627 ( .A(n8643), .B(n8642), .Z(n8644) );
  XNOR U10628 ( .A(n8645), .B(n8644), .Z(n8674) );
  XNOR U10629 ( .A(sreg[1139]), .B(n8674), .Z(n8676) );
  NANDN U10630 ( .A(sreg[1138]), .B(n8637), .Z(n8641) );
  NAND U10631 ( .A(n8639), .B(n8638), .Z(n8640) );
  NAND U10632 ( .A(n8641), .B(n8640), .Z(n8675) );
  XNOR U10633 ( .A(n8676), .B(n8675), .Z(c[1139]) );
  NANDN U10634 ( .A(n8643), .B(n8642), .Z(n8647) );
  NANDN U10635 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U10636 ( .A(n8647), .B(n8646), .Z(n8682) );
  NANDN U10637 ( .A(n8649), .B(n8648), .Z(n8653) );
  NANDN U10638 ( .A(n8651), .B(n8650), .Z(n8652) );
  AND U10639 ( .A(n8653), .B(n8652), .Z(n8680) );
  NAND U10640 ( .A(n42143), .B(n8654), .Z(n8656) );
  XNOR U10641 ( .A(a[118]), .B(n4088), .Z(n8691) );
  NAND U10642 ( .A(n42144), .B(n8691), .Z(n8655) );
  AND U10643 ( .A(n8656), .B(n8655), .Z(n8706) );
  XOR U10644 ( .A(a[122]), .B(n42012), .Z(n8694) );
  XNOR U10645 ( .A(n8706), .B(n8705), .Z(n8708) );
  AND U10646 ( .A(a[124]), .B(b[0]), .Z(n8658) );
  XNOR U10647 ( .A(n8658), .B(n4071), .Z(n8660) );
  NANDN U10648 ( .A(b[0]), .B(a[123]), .Z(n8659) );
  NAND U10649 ( .A(n8660), .B(n8659), .Z(n8702) );
  XOR U10650 ( .A(a[120]), .B(n42085), .Z(n8695) );
  AND U10651 ( .A(a[116]), .B(b[7]), .Z(n8699) );
  XNOR U10652 ( .A(n8700), .B(n8699), .Z(n8701) );
  XNOR U10653 ( .A(n8702), .B(n8701), .Z(n8707) );
  XOR U10654 ( .A(n8708), .B(n8707), .Z(n8686) );
  NANDN U10655 ( .A(n8663), .B(n8662), .Z(n8667) );
  NANDN U10656 ( .A(n8665), .B(n8664), .Z(n8666) );
  AND U10657 ( .A(n8667), .B(n8666), .Z(n8685) );
  XNOR U10658 ( .A(n8686), .B(n8685), .Z(n8687) );
  NANDN U10659 ( .A(n8669), .B(n8668), .Z(n8673) );
  NAND U10660 ( .A(n8671), .B(n8670), .Z(n8672) );
  NAND U10661 ( .A(n8673), .B(n8672), .Z(n8688) );
  XNOR U10662 ( .A(n8687), .B(n8688), .Z(n8679) );
  XNOR U10663 ( .A(n8680), .B(n8679), .Z(n8681) );
  XNOR U10664 ( .A(n8682), .B(n8681), .Z(n8711) );
  XNOR U10665 ( .A(sreg[1140]), .B(n8711), .Z(n8713) );
  NANDN U10666 ( .A(sreg[1139]), .B(n8674), .Z(n8678) );
  NAND U10667 ( .A(n8676), .B(n8675), .Z(n8677) );
  NAND U10668 ( .A(n8678), .B(n8677), .Z(n8712) );
  XNOR U10669 ( .A(n8713), .B(n8712), .Z(c[1140]) );
  NANDN U10670 ( .A(n8680), .B(n8679), .Z(n8684) );
  NANDN U10671 ( .A(n8682), .B(n8681), .Z(n8683) );
  AND U10672 ( .A(n8684), .B(n8683), .Z(n8719) );
  NANDN U10673 ( .A(n8686), .B(n8685), .Z(n8690) );
  NANDN U10674 ( .A(n8688), .B(n8687), .Z(n8689) );
  AND U10675 ( .A(n8690), .B(n8689), .Z(n8717) );
  NAND U10676 ( .A(n42143), .B(n8691), .Z(n8693) );
  XNOR U10677 ( .A(a[119]), .B(n4088), .Z(n8728) );
  NAND U10678 ( .A(n42144), .B(n8728), .Z(n8692) );
  AND U10679 ( .A(n8693), .B(n8692), .Z(n8743) );
  XOR U10680 ( .A(a[123]), .B(n42012), .Z(n8731) );
  XNOR U10681 ( .A(n8743), .B(n8742), .Z(n8745) );
  XOR U10682 ( .A(a[121]), .B(n42085), .Z(n8732) );
  AND U10683 ( .A(a[117]), .B(b[7]), .Z(n8736) );
  XNOR U10684 ( .A(n8737), .B(n8736), .Z(n8738) );
  AND U10685 ( .A(a[125]), .B(b[0]), .Z(n8696) );
  XNOR U10686 ( .A(n8696), .B(n4071), .Z(n8698) );
  NANDN U10687 ( .A(b[0]), .B(a[124]), .Z(n8697) );
  NAND U10688 ( .A(n8698), .B(n8697), .Z(n8739) );
  XNOR U10689 ( .A(n8738), .B(n8739), .Z(n8744) );
  XOR U10690 ( .A(n8745), .B(n8744), .Z(n8723) );
  NANDN U10691 ( .A(n8700), .B(n8699), .Z(n8704) );
  NANDN U10692 ( .A(n8702), .B(n8701), .Z(n8703) );
  AND U10693 ( .A(n8704), .B(n8703), .Z(n8722) );
  XNOR U10694 ( .A(n8723), .B(n8722), .Z(n8724) );
  NANDN U10695 ( .A(n8706), .B(n8705), .Z(n8710) );
  NAND U10696 ( .A(n8708), .B(n8707), .Z(n8709) );
  NAND U10697 ( .A(n8710), .B(n8709), .Z(n8725) );
  XNOR U10698 ( .A(n8724), .B(n8725), .Z(n8716) );
  XNOR U10699 ( .A(n8717), .B(n8716), .Z(n8718) );
  XNOR U10700 ( .A(n8719), .B(n8718), .Z(n8748) );
  XNOR U10701 ( .A(sreg[1141]), .B(n8748), .Z(n8750) );
  NANDN U10702 ( .A(sreg[1140]), .B(n8711), .Z(n8715) );
  NAND U10703 ( .A(n8713), .B(n8712), .Z(n8714) );
  NAND U10704 ( .A(n8715), .B(n8714), .Z(n8749) );
  XNOR U10705 ( .A(n8750), .B(n8749), .Z(c[1141]) );
  NANDN U10706 ( .A(n8717), .B(n8716), .Z(n8721) );
  NANDN U10707 ( .A(n8719), .B(n8718), .Z(n8720) );
  AND U10708 ( .A(n8721), .B(n8720), .Z(n8756) );
  NANDN U10709 ( .A(n8723), .B(n8722), .Z(n8727) );
  NANDN U10710 ( .A(n8725), .B(n8724), .Z(n8726) );
  AND U10711 ( .A(n8727), .B(n8726), .Z(n8754) );
  NAND U10712 ( .A(n42143), .B(n8728), .Z(n8730) );
  XNOR U10713 ( .A(a[120]), .B(n4089), .Z(n8765) );
  NAND U10714 ( .A(n42144), .B(n8765), .Z(n8729) );
  AND U10715 ( .A(n8730), .B(n8729), .Z(n8780) );
  XOR U10716 ( .A(a[124]), .B(n42012), .Z(n8768) );
  XNOR U10717 ( .A(n8780), .B(n8779), .Z(n8782) );
  XOR U10718 ( .A(a[122]), .B(n42085), .Z(n8772) );
  AND U10719 ( .A(a[118]), .B(b[7]), .Z(n8773) );
  XNOR U10720 ( .A(n8774), .B(n8773), .Z(n8775) );
  AND U10721 ( .A(a[126]), .B(b[0]), .Z(n8733) );
  XNOR U10722 ( .A(n8733), .B(n4071), .Z(n8735) );
  NANDN U10723 ( .A(b[0]), .B(a[125]), .Z(n8734) );
  NAND U10724 ( .A(n8735), .B(n8734), .Z(n8776) );
  XNOR U10725 ( .A(n8775), .B(n8776), .Z(n8781) );
  XOR U10726 ( .A(n8782), .B(n8781), .Z(n8760) );
  NANDN U10727 ( .A(n8737), .B(n8736), .Z(n8741) );
  NANDN U10728 ( .A(n8739), .B(n8738), .Z(n8740) );
  AND U10729 ( .A(n8741), .B(n8740), .Z(n8759) );
  XNOR U10730 ( .A(n8760), .B(n8759), .Z(n8761) );
  NANDN U10731 ( .A(n8743), .B(n8742), .Z(n8747) );
  NAND U10732 ( .A(n8745), .B(n8744), .Z(n8746) );
  NAND U10733 ( .A(n8747), .B(n8746), .Z(n8762) );
  XNOR U10734 ( .A(n8761), .B(n8762), .Z(n8753) );
  XNOR U10735 ( .A(n8754), .B(n8753), .Z(n8755) );
  XNOR U10736 ( .A(n8756), .B(n8755), .Z(n8785) );
  XNOR U10737 ( .A(sreg[1142]), .B(n8785), .Z(n8787) );
  NANDN U10738 ( .A(sreg[1141]), .B(n8748), .Z(n8752) );
  NAND U10739 ( .A(n8750), .B(n8749), .Z(n8751) );
  NAND U10740 ( .A(n8752), .B(n8751), .Z(n8786) );
  XNOR U10741 ( .A(n8787), .B(n8786), .Z(c[1142]) );
  NANDN U10742 ( .A(n8754), .B(n8753), .Z(n8758) );
  NANDN U10743 ( .A(n8756), .B(n8755), .Z(n8757) );
  AND U10744 ( .A(n8758), .B(n8757), .Z(n8793) );
  NANDN U10745 ( .A(n8760), .B(n8759), .Z(n8764) );
  NANDN U10746 ( .A(n8762), .B(n8761), .Z(n8763) );
  AND U10747 ( .A(n8764), .B(n8763), .Z(n8791) );
  NAND U10748 ( .A(n42143), .B(n8765), .Z(n8767) );
  XNOR U10749 ( .A(a[121]), .B(n4089), .Z(n8802) );
  NAND U10750 ( .A(n42144), .B(n8802), .Z(n8766) );
  AND U10751 ( .A(n8767), .B(n8766), .Z(n8817) );
  XOR U10752 ( .A(a[125]), .B(n42012), .Z(n8805) );
  XNOR U10753 ( .A(n8817), .B(n8816), .Z(n8819) );
  AND U10754 ( .A(a[127]), .B(b[0]), .Z(n8769) );
  XNOR U10755 ( .A(n8769), .B(n4071), .Z(n8771) );
  NANDN U10756 ( .A(b[0]), .B(a[126]), .Z(n8770) );
  NAND U10757 ( .A(n8771), .B(n8770), .Z(n8813) );
  XOR U10758 ( .A(a[123]), .B(n42085), .Z(n8806) );
  AND U10759 ( .A(a[119]), .B(b[7]), .Z(n8810) );
  XNOR U10760 ( .A(n8811), .B(n8810), .Z(n8812) );
  XNOR U10761 ( .A(n8813), .B(n8812), .Z(n8818) );
  XOR U10762 ( .A(n8819), .B(n8818), .Z(n8797) );
  NANDN U10763 ( .A(n8774), .B(n8773), .Z(n8778) );
  NANDN U10764 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U10765 ( .A(n8778), .B(n8777), .Z(n8796) );
  XNOR U10766 ( .A(n8797), .B(n8796), .Z(n8798) );
  NANDN U10767 ( .A(n8780), .B(n8779), .Z(n8784) );
  NAND U10768 ( .A(n8782), .B(n8781), .Z(n8783) );
  NAND U10769 ( .A(n8784), .B(n8783), .Z(n8799) );
  XNOR U10770 ( .A(n8798), .B(n8799), .Z(n8790) );
  XNOR U10771 ( .A(n8791), .B(n8790), .Z(n8792) );
  XNOR U10772 ( .A(n8793), .B(n8792), .Z(n8822) );
  XNOR U10773 ( .A(sreg[1143]), .B(n8822), .Z(n8824) );
  NANDN U10774 ( .A(sreg[1142]), .B(n8785), .Z(n8789) );
  NAND U10775 ( .A(n8787), .B(n8786), .Z(n8788) );
  NAND U10776 ( .A(n8789), .B(n8788), .Z(n8823) );
  XNOR U10777 ( .A(n8824), .B(n8823), .Z(c[1143]) );
  NANDN U10778 ( .A(n8791), .B(n8790), .Z(n8795) );
  NANDN U10779 ( .A(n8793), .B(n8792), .Z(n8794) );
  AND U10780 ( .A(n8795), .B(n8794), .Z(n8830) );
  NANDN U10781 ( .A(n8797), .B(n8796), .Z(n8801) );
  NANDN U10782 ( .A(n8799), .B(n8798), .Z(n8800) );
  AND U10783 ( .A(n8801), .B(n8800), .Z(n8828) );
  NAND U10784 ( .A(n42143), .B(n8802), .Z(n8804) );
  XNOR U10785 ( .A(a[122]), .B(n4089), .Z(n8839) );
  NAND U10786 ( .A(n42144), .B(n8839), .Z(n8803) );
  AND U10787 ( .A(n8804), .B(n8803), .Z(n8854) );
  XOR U10788 ( .A(a[126]), .B(n42012), .Z(n8842) );
  XNOR U10789 ( .A(n8854), .B(n8853), .Z(n8856) );
  XOR U10790 ( .A(a[124]), .B(n42085), .Z(n8843) );
  AND U10791 ( .A(a[120]), .B(b[7]), .Z(n8847) );
  XNOR U10792 ( .A(n8848), .B(n8847), .Z(n8849) );
  AND U10793 ( .A(a[128]), .B(b[0]), .Z(n8807) );
  XNOR U10794 ( .A(n8807), .B(n4071), .Z(n8809) );
  NANDN U10795 ( .A(b[0]), .B(a[127]), .Z(n8808) );
  NAND U10796 ( .A(n8809), .B(n8808), .Z(n8850) );
  XNOR U10797 ( .A(n8849), .B(n8850), .Z(n8855) );
  XOR U10798 ( .A(n8856), .B(n8855), .Z(n8834) );
  NANDN U10799 ( .A(n8811), .B(n8810), .Z(n8815) );
  NANDN U10800 ( .A(n8813), .B(n8812), .Z(n8814) );
  AND U10801 ( .A(n8815), .B(n8814), .Z(n8833) );
  XNOR U10802 ( .A(n8834), .B(n8833), .Z(n8835) );
  NANDN U10803 ( .A(n8817), .B(n8816), .Z(n8821) );
  NAND U10804 ( .A(n8819), .B(n8818), .Z(n8820) );
  NAND U10805 ( .A(n8821), .B(n8820), .Z(n8836) );
  XNOR U10806 ( .A(n8835), .B(n8836), .Z(n8827) );
  XNOR U10807 ( .A(n8828), .B(n8827), .Z(n8829) );
  XNOR U10808 ( .A(n8830), .B(n8829), .Z(n8859) );
  XNOR U10809 ( .A(sreg[1144]), .B(n8859), .Z(n8861) );
  NANDN U10810 ( .A(sreg[1143]), .B(n8822), .Z(n8826) );
  NAND U10811 ( .A(n8824), .B(n8823), .Z(n8825) );
  NAND U10812 ( .A(n8826), .B(n8825), .Z(n8860) );
  XNOR U10813 ( .A(n8861), .B(n8860), .Z(c[1144]) );
  NANDN U10814 ( .A(n8828), .B(n8827), .Z(n8832) );
  NANDN U10815 ( .A(n8830), .B(n8829), .Z(n8831) );
  AND U10816 ( .A(n8832), .B(n8831), .Z(n8867) );
  NANDN U10817 ( .A(n8834), .B(n8833), .Z(n8838) );
  NANDN U10818 ( .A(n8836), .B(n8835), .Z(n8837) );
  AND U10819 ( .A(n8838), .B(n8837), .Z(n8865) );
  NAND U10820 ( .A(n42143), .B(n8839), .Z(n8841) );
  XNOR U10821 ( .A(a[123]), .B(n4089), .Z(n8876) );
  NAND U10822 ( .A(n42144), .B(n8876), .Z(n8840) );
  AND U10823 ( .A(n8841), .B(n8840), .Z(n8891) );
  XOR U10824 ( .A(a[127]), .B(n42012), .Z(n8879) );
  XNOR U10825 ( .A(n8891), .B(n8890), .Z(n8893) );
  XOR U10826 ( .A(a[125]), .B(n42085), .Z(n8883) );
  AND U10827 ( .A(a[121]), .B(b[7]), .Z(n8884) );
  XNOR U10828 ( .A(n8885), .B(n8884), .Z(n8886) );
  AND U10829 ( .A(a[129]), .B(b[0]), .Z(n8844) );
  XNOR U10830 ( .A(n8844), .B(n4071), .Z(n8846) );
  NANDN U10831 ( .A(b[0]), .B(a[128]), .Z(n8845) );
  NAND U10832 ( .A(n8846), .B(n8845), .Z(n8887) );
  XNOR U10833 ( .A(n8886), .B(n8887), .Z(n8892) );
  XOR U10834 ( .A(n8893), .B(n8892), .Z(n8871) );
  NANDN U10835 ( .A(n8848), .B(n8847), .Z(n8852) );
  NANDN U10836 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U10837 ( .A(n8852), .B(n8851), .Z(n8870) );
  XNOR U10838 ( .A(n8871), .B(n8870), .Z(n8872) );
  NANDN U10839 ( .A(n8854), .B(n8853), .Z(n8858) );
  NAND U10840 ( .A(n8856), .B(n8855), .Z(n8857) );
  NAND U10841 ( .A(n8858), .B(n8857), .Z(n8873) );
  XNOR U10842 ( .A(n8872), .B(n8873), .Z(n8864) );
  XNOR U10843 ( .A(n8865), .B(n8864), .Z(n8866) );
  XNOR U10844 ( .A(n8867), .B(n8866), .Z(n8896) );
  XNOR U10845 ( .A(sreg[1145]), .B(n8896), .Z(n8898) );
  NANDN U10846 ( .A(sreg[1144]), .B(n8859), .Z(n8863) );
  NAND U10847 ( .A(n8861), .B(n8860), .Z(n8862) );
  NAND U10848 ( .A(n8863), .B(n8862), .Z(n8897) );
  XNOR U10849 ( .A(n8898), .B(n8897), .Z(c[1145]) );
  NANDN U10850 ( .A(n8865), .B(n8864), .Z(n8869) );
  NANDN U10851 ( .A(n8867), .B(n8866), .Z(n8868) );
  AND U10852 ( .A(n8869), .B(n8868), .Z(n8904) );
  NANDN U10853 ( .A(n8871), .B(n8870), .Z(n8875) );
  NANDN U10854 ( .A(n8873), .B(n8872), .Z(n8874) );
  AND U10855 ( .A(n8875), .B(n8874), .Z(n8902) );
  NAND U10856 ( .A(n42143), .B(n8876), .Z(n8878) );
  XNOR U10857 ( .A(a[124]), .B(n4089), .Z(n8913) );
  NAND U10858 ( .A(n42144), .B(n8913), .Z(n8877) );
  AND U10859 ( .A(n8878), .B(n8877), .Z(n8928) );
  XOR U10860 ( .A(a[128]), .B(n42012), .Z(n8916) );
  XNOR U10861 ( .A(n8928), .B(n8927), .Z(n8930) );
  AND U10862 ( .A(a[130]), .B(b[0]), .Z(n8880) );
  XNOR U10863 ( .A(n8880), .B(n4071), .Z(n8882) );
  NANDN U10864 ( .A(b[0]), .B(a[129]), .Z(n8881) );
  NAND U10865 ( .A(n8882), .B(n8881), .Z(n8924) );
  XOR U10866 ( .A(a[126]), .B(n42085), .Z(n8920) );
  AND U10867 ( .A(a[122]), .B(b[7]), .Z(n8921) );
  XNOR U10868 ( .A(n8922), .B(n8921), .Z(n8923) );
  XNOR U10869 ( .A(n8924), .B(n8923), .Z(n8929) );
  XOR U10870 ( .A(n8930), .B(n8929), .Z(n8908) );
  NANDN U10871 ( .A(n8885), .B(n8884), .Z(n8889) );
  NANDN U10872 ( .A(n8887), .B(n8886), .Z(n8888) );
  AND U10873 ( .A(n8889), .B(n8888), .Z(n8907) );
  XNOR U10874 ( .A(n8908), .B(n8907), .Z(n8909) );
  NANDN U10875 ( .A(n8891), .B(n8890), .Z(n8895) );
  NAND U10876 ( .A(n8893), .B(n8892), .Z(n8894) );
  NAND U10877 ( .A(n8895), .B(n8894), .Z(n8910) );
  XNOR U10878 ( .A(n8909), .B(n8910), .Z(n8901) );
  XNOR U10879 ( .A(n8902), .B(n8901), .Z(n8903) );
  XNOR U10880 ( .A(n8904), .B(n8903), .Z(n8933) );
  XNOR U10881 ( .A(sreg[1146]), .B(n8933), .Z(n8935) );
  NANDN U10882 ( .A(sreg[1145]), .B(n8896), .Z(n8900) );
  NAND U10883 ( .A(n8898), .B(n8897), .Z(n8899) );
  NAND U10884 ( .A(n8900), .B(n8899), .Z(n8934) );
  XNOR U10885 ( .A(n8935), .B(n8934), .Z(c[1146]) );
  NANDN U10886 ( .A(n8902), .B(n8901), .Z(n8906) );
  NANDN U10887 ( .A(n8904), .B(n8903), .Z(n8905) );
  AND U10888 ( .A(n8906), .B(n8905), .Z(n8941) );
  NANDN U10889 ( .A(n8908), .B(n8907), .Z(n8912) );
  NANDN U10890 ( .A(n8910), .B(n8909), .Z(n8911) );
  AND U10891 ( .A(n8912), .B(n8911), .Z(n8939) );
  NAND U10892 ( .A(n42143), .B(n8913), .Z(n8915) );
  XNOR U10893 ( .A(a[125]), .B(n4089), .Z(n8950) );
  NAND U10894 ( .A(n42144), .B(n8950), .Z(n8914) );
  AND U10895 ( .A(n8915), .B(n8914), .Z(n8965) );
  XOR U10896 ( .A(a[129]), .B(n42012), .Z(n8953) );
  XNOR U10897 ( .A(n8965), .B(n8964), .Z(n8967) );
  AND U10898 ( .A(a[131]), .B(b[0]), .Z(n8917) );
  XNOR U10899 ( .A(n8917), .B(n4071), .Z(n8919) );
  NANDN U10900 ( .A(b[0]), .B(a[130]), .Z(n8918) );
  NAND U10901 ( .A(n8919), .B(n8918), .Z(n8961) );
  XOR U10902 ( .A(a[127]), .B(n42085), .Z(n8957) );
  AND U10903 ( .A(a[123]), .B(b[7]), .Z(n8958) );
  XNOR U10904 ( .A(n8959), .B(n8958), .Z(n8960) );
  XNOR U10905 ( .A(n8961), .B(n8960), .Z(n8966) );
  XOR U10906 ( .A(n8967), .B(n8966), .Z(n8945) );
  NANDN U10907 ( .A(n8922), .B(n8921), .Z(n8926) );
  NANDN U10908 ( .A(n8924), .B(n8923), .Z(n8925) );
  AND U10909 ( .A(n8926), .B(n8925), .Z(n8944) );
  XNOR U10910 ( .A(n8945), .B(n8944), .Z(n8946) );
  NANDN U10911 ( .A(n8928), .B(n8927), .Z(n8932) );
  NAND U10912 ( .A(n8930), .B(n8929), .Z(n8931) );
  NAND U10913 ( .A(n8932), .B(n8931), .Z(n8947) );
  XNOR U10914 ( .A(n8946), .B(n8947), .Z(n8938) );
  XNOR U10915 ( .A(n8939), .B(n8938), .Z(n8940) );
  XNOR U10916 ( .A(n8941), .B(n8940), .Z(n8970) );
  XNOR U10917 ( .A(sreg[1147]), .B(n8970), .Z(n8972) );
  NANDN U10918 ( .A(sreg[1146]), .B(n8933), .Z(n8937) );
  NAND U10919 ( .A(n8935), .B(n8934), .Z(n8936) );
  NAND U10920 ( .A(n8937), .B(n8936), .Z(n8971) );
  XNOR U10921 ( .A(n8972), .B(n8971), .Z(c[1147]) );
  NANDN U10922 ( .A(n8939), .B(n8938), .Z(n8943) );
  NANDN U10923 ( .A(n8941), .B(n8940), .Z(n8942) );
  AND U10924 ( .A(n8943), .B(n8942), .Z(n8978) );
  NANDN U10925 ( .A(n8945), .B(n8944), .Z(n8949) );
  NANDN U10926 ( .A(n8947), .B(n8946), .Z(n8948) );
  AND U10927 ( .A(n8949), .B(n8948), .Z(n8976) );
  NAND U10928 ( .A(n42143), .B(n8950), .Z(n8952) );
  XNOR U10929 ( .A(a[126]), .B(n4089), .Z(n8987) );
  NAND U10930 ( .A(n42144), .B(n8987), .Z(n8951) );
  AND U10931 ( .A(n8952), .B(n8951), .Z(n9002) );
  XOR U10932 ( .A(a[130]), .B(n42012), .Z(n8990) );
  XNOR U10933 ( .A(n9002), .B(n9001), .Z(n9004) );
  AND U10934 ( .A(a[132]), .B(b[0]), .Z(n8954) );
  XNOR U10935 ( .A(n8954), .B(n4071), .Z(n8956) );
  NANDN U10936 ( .A(b[0]), .B(a[131]), .Z(n8955) );
  NAND U10937 ( .A(n8956), .B(n8955), .Z(n8998) );
  XOR U10938 ( .A(a[128]), .B(n42085), .Z(n8994) );
  AND U10939 ( .A(a[124]), .B(b[7]), .Z(n8995) );
  XNOR U10940 ( .A(n8996), .B(n8995), .Z(n8997) );
  XNOR U10941 ( .A(n8998), .B(n8997), .Z(n9003) );
  XOR U10942 ( .A(n9004), .B(n9003), .Z(n8982) );
  NANDN U10943 ( .A(n8959), .B(n8958), .Z(n8963) );
  NANDN U10944 ( .A(n8961), .B(n8960), .Z(n8962) );
  AND U10945 ( .A(n8963), .B(n8962), .Z(n8981) );
  XNOR U10946 ( .A(n8982), .B(n8981), .Z(n8983) );
  NANDN U10947 ( .A(n8965), .B(n8964), .Z(n8969) );
  NAND U10948 ( .A(n8967), .B(n8966), .Z(n8968) );
  NAND U10949 ( .A(n8969), .B(n8968), .Z(n8984) );
  XNOR U10950 ( .A(n8983), .B(n8984), .Z(n8975) );
  XNOR U10951 ( .A(n8976), .B(n8975), .Z(n8977) );
  XNOR U10952 ( .A(n8978), .B(n8977), .Z(n9007) );
  XNOR U10953 ( .A(sreg[1148]), .B(n9007), .Z(n9009) );
  NANDN U10954 ( .A(sreg[1147]), .B(n8970), .Z(n8974) );
  NAND U10955 ( .A(n8972), .B(n8971), .Z(n8973) );
  NAND U10956 ( .A(n8974), .B(n8973), .Z(n9008) );
  XNOR U10957 ( .A(n9009), .B(n9008), .Z(c[1148]) );
  NANDN U10958 ( .A(n8976), .B(n8975), .Z(n8980) );
  NANDN U10959 ( .A(n8978), .B(n8977), .Z(n8979) );
  AND U10960 ( .A(n8980), .B(n8979), .Z(n9019) );
  NANDN U10961 ( .A(n8982), .B(n8981), .Z(n8986) );
  NANDN U10962 ( .A(n8984), .B(n8983), .Z(n8985) );
  AND U10963 ( .A(n8986), .B(n8985), .Z(n9018) );
  NAND U10964 ( .A(n42143), .B(n8987), .Z(n8989) );
  XNOR U10965 ( .A(a[127]), .B(n4090), .Z(n9029) );
  NAND U10966 ( .A(n42144), .B(n9029), .Z(n8988) );
  AND U10967 ( .A(n8989), .B(n8988), .Z(n9044) );
  XOR U10968 ( .A(a[131]), .B(n42012), .Z(n9032) );
  XNOR U10969 ( .A(n9044), .B(n9043), .Z(n9046) );
  AND U10970 ( .A(a[133]), .B(b[0]), .Z(n8991) );
  XNOR U10971 ( .A(n8991), .B(n4071), .Z(n8993) );
  NANDN U10972 ( .A(b[0]), .B(a[132]), .Z(n8992) );
  NAND U10973 ( .A(n8993), .B(n8992), .Z(n9040) );
  XOR U10974 ( .A(a[129]), .B(n42085), .Z(n9033) );
  AND U10975 ( .A(a[125]), .B(b[7]), .Z(n9037) );
  XNOR U10976 ( .A(n9038), .B(n9037), .Z(n9039) );
  XNOR U10977 ( .A(n9040), .B(n9039), .Z(n9045) );
  XOR U10978 ( .A(n9046), .B(n9045), .Z(n9024) );
  NANDN U10979 ( .A(n8996), .B(n8995), .Z(n9000) );
  NANDN U10980 ( .A(n8998), .B(n8997), .Z(n8999) );
  AND U10981 ( .A(n9000), .B(n8999), .Z(n9023) );
  XNOR U10982 ( .A(n9024), .B(n9023), .Z(n9025) );
  NANDN U10983 ( .A(n9002), .B(n9001), .Z(n9006) );
  NAND U10984 ( .A(n9004), .B(n9003), .Z(n9005) );
  NAND U10985 ( .A(n9006), .B(n9005), .Z(n9026) );
  XNOR U10986 ( .A(n9025), .B(n9026), .Z(n9017) );
  XOR U10987 ( .A(n9018), .B(n9017), .Z(n9020) );
  XOR U10988 ( .A(n9019), .B(n9020), .Z(n9012) );
  XNOR U10989 ( .A(n9012), .B(sreg[1149]), .Z(n9014) );
  NANDN U10990 ( .A(sreg[1148]), .B(n9007), .Z(n9011) );
  NAND U10991 ( .A(n9009), .B(n9008), .Z(n9010) );
  AND U10992 ( .A(n9011), .B(n9010), .Z(n9013) );
  XOR U10993 ( .A(n9014), .B(n9013), .Z(c[1149]) );
  NANDN U10994 ( .A(n9012), .B(sreg[1149]), .Z(n9016) );
  NAND U10995 ( .A(n9014), .B(n9013), .Z(n9015) );
  AND U10996 ( .A(n9016), .B(n9015), .Z(n9083) );
  NANDN U10997 ( .A(n9018), .B(n9017), .Z(n9022) );
  OR U10998 ( .A(n9020), .B(n9019), .Z(n9021) );
  AND U10999 ( .A(n9022), .B(n9021), .Z(n9052) );
  NANDN U11000 ( .A(n9024), .B(n9023), .Z(n9028) );
  NANDN U11001 ( .A(n9026), .B(n9025), .Z(n9027) );
  AND U11002 ( .A(n9028), .B(n9027), .Z(n9050) );
  NAND U11003 ( .A(n42143), .B(n9029), .Z(n9031) );
  XNOR U11004 ( .A(a[128]), .B(n4090), .Z(n9061) );
  NAND U11005 ( .A(n42144), .B(n9061), .Z(n9030) );
  AND U11006 ( .A(n9031), .B(n9030), .Z(n9076) );
  XOR U11007 ( .A(a[132]), .B(n42012), .Z(n9064) );
  XNOR U11008 ( .A(n9076), .B(n9075), .Z(n9078) );
  XOR U11009 ( .A(a[130]), .B(n42085), .Z(n9068) );
  AND U11010 ( .A(a[126]), .B(b[7]), .Z(n9069) );
  XNOR U11011 ( .A(n9070), .B(n9069), .Z(n9071) );
  AND U11012 ( .A(a[134]), .B(b[0]), .Z(n9034) );
  XNOR U11013 ( .A(n9034), .B(n4071), .Z(n9036) );
  NANDN U11014 ( .A(b[0]), .B(a[133]), .Z(n9035) );
  NAND U11015 ( .A(n9036), .B(n9035), .Z(n9072) );
  XNOR U11016 ( .A(n9071), .B(n9072), .Z(n9077) );
  XOR U11017 ( .A(n9078), .B(n9077), .Z(n9056) );
  NANDN U11018 ( .A(n9038), .B(n9037), .Z(n9042) );
  NANDN U11019 ( .A(n9040), .B(n9039), .Z(n9041) );
  AND U11020 ( .A(n9042), .B(n9041), .Z(n9055) );
  XNOR U11021 ( .A(n9056), .B(n9055), .Z(n9057) );
  NANDN U11022 ( .A(n9044), .B(n9043), .Z(n9048) );
  NAND U11023 ( .A(n9046), .B(n9045), .Z(n9047) );
  NAND U11024 ( .A(n9048), .B(n9047), .Z(n9058) );
  XNOR U11025 ( .A(n9057), .B(n9058), .Z(n9049) );
  XNOR U11026 ( .A(n9050), .B(n9049), .Z(n9051) );
  XNOR U11027 ( .A(n9052), .B(n9051), .Z(n9081) );
  XNOR U11028 ( .A(sreg[1150]), .B(n9081), .Z(n9082) );
  XNOR U11029 ( .A(n9083), .B(n9082), .Z(c[1150]) );
  NANDN U11030 ( .A(n9050), .B(n9049), .Z(n9054) );
  NANDN U11031 ( .A(n9052), .B(n9051), .Z(n9053) );
  AND U11032 ( .A(n9054), .B(n9053), .Z(n9089) );
  NANDN U11033 ( .A(n9056), .B(n9055), .Z(n9060) );
  NANDN U11034 ( .A(n9058), .B(n9057), .Z(n9059) );
  AND U11035 ( .A(n9060), .B(n9059), .Z(n9087) );
  NAND U11036 ( .A(n42143), .B(n9061), .Z(n9063) );
  XNOR U11037 ( .A(a[129]), .B(n4090), .Z(n9098) );
  NAND U11038 ( .A(n42144), .B(n9098), .Z(n9062) );
  AND U11039 ( .A(n9063), .B(n9062), .Z(n9113) );
  XOR U11040 ( .A(a[133]), .B(n42012), .Z(n9101) );
  XNOR U11041 ( .A(n9113), .B(n9112), .Z(n9115) );
  AND U11042 ( .A(a[135]), .B(b[0]), .Z(n9065) );
  XNOR U11043 ( .A(n9065), .B(n4071), .Z(n9067) );
  NANDN U11044 ( .A(b[0]), .B(a[134]), .Z(n9066) );
  NAND U11045 ( .A(n9067), .B(n9066), .Z(n9109) );
  XOR U11046 ( .A(a[131]), .B(n42085), .Z(n9105) );
  AND U11047 ( .A(a[127]), .B(b[7]), .Z(n9106) );
  XNOR U11048 ( .A(n9107), .B(n9106), .Z(n9108) );
  XNOR U11049 ( .A(n9109), .B(n9108), .Z(n9114) );
  XOR U11050 ( .A(n9115), .B(n9114), .Z(n9093) );
  NANDN U11051 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U11052 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U11053 ( .A(n9074), .B(n9073), .Z(n9092) );
  XNOR U11054 ( .A(n9093), .B(n9092), .Z(n9094) );
  NANDN U11055 ( .A(n9076), .B(n9075), .Z(n9080) );
  NAND U11056 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U11057 ( .A(n9080), .B(n9079), .Z(n9095) );
  XNOR U11058 ( .A(n9094), .B(n9095), .Z(n9086) );
  XNOR U11059 ( .A(n9087), .B(n9086), .Z(n9088) );
  XNOR U11060 ( .A(n9089), .B(n9088), .Z(n9118) );
  XNOR U11061 ( .A(sreg[1151]), .B(n9118), .Z(n9120) );
  NANDN U11062 ( .A(sreg[1150]), .B(n9081), .Z(n9085) );
  NAND U11063 ( .A(n9083), .B(n9082), .Z(n9084) );
  NAND U11064 ( .A(n9085), .B(n9084), .Z(n9119) );
  XNOR U11065 ( .A(n9120), .B(n9119), .Z(c[1151]) );
  NANDN U11066 ( .A(n9087), .B(n9086), .Z(n9091) );
  NANDN U11067 ( .A(n9089), .B(n9088), .Z(n9090) );
  AND U11068 ( .A(n9091), .B(n9090), .Z(n9126) );
  NANDN U11069 ( .A(n9093), .B(n9092), .Z(n9097) );
  NANDN U11070 ( .A(n9095), .B(n9094), .Z(n9096) );
  AND U11071 ( .A(n9097), .B(n9096), .Z(n9124) );
  NAND U11072 ( .A(n42143), .B(n9098), .Z(n9100) );
  XNOR U11073 ( .A(a[130]), .B(n4090), .Z(n9135) );
  NAND U11074 ( .A(n42144), .B(n9135), .Z(n9099) );
  AND U11075 ( .A(n9100), .B(n9099), .Z(n9150) );
  XOR U11076 ( .A(a[134]), .B(n42012), .Z(n9138) );
  XNOR U11077 ( .A(n9150), .B(n9149), .Z(n9152) );
  AND U11078 ( .A(a[136]), .B(b[0]), .Z(n9102) );
  XNOR U11079 ( .A(n9102), .B(n4071), .Z(n9104) );
  NANDN U11080 ( .A(b[0]), .B(a[135]), .Z(n9103) );
  NAND U11081 ( .A(n9104), .B(n9103), .Z(n9146) );
  XOR U11082 ( .A(a[132]), .B(n42085), .Z(n9142) );
  AND U11083 ( .A(a[128]), .B(b[7]), .Z(n9143) );
  XNOR U11084 ( .A(n9144), .B(n9143), .Z(n9145) );
  XNOR U11085 ( .A(n9146), .B(n9145), .Z(n9151) );
  XOR U11086 ( .A(n9152), .B(n9151), .Z(n9130) );
  NANDN U11087 ( .A(n9107), .B(n9106), .Z(n9111) );
  NANDN U11088 ( .A(n9109), .B(n9108), .Z(n9110) );
  AND U11089 ( .A(n9111), .B(n9110), .Z(n9129) );
  XNOR U11090 ( .A(n9130), .B(n9129), .Z(n9131) );
  NANDN U11091 ( .A(n9113), .B(n9112), .Z(n9117) );
  NAND U11092 ( .A(n9115), .B(n9114), .Z(n9116) );
  NAND U11093 ( .A(n9117), .B(n9116), .Z(n9132) );
  XNOR U11094 ( .A(n9131), .B(n9132), .Z(n9123) );
  XNOR U11095 ( .A(n9124), .B(n9123), .Z(n9125) );
  XNOR U11096 ( .A(n9126), .B(n9125), .Z(n9155) );
  XNOR U11097 ( .A(sreg[1152]), .B(n9155), .Z(n9157) );
  NANDN U11098 ( .A(sreg[1151]), .B(n9118), .Z(n9122) );
  NAND U11099 ( .A(n9120), .B(n9119), .Z(n9121) );
  NAND U11100 ( .A(n9122), .B(n9121), .Z(n9156) );
  XNOR U11101 ( .A(n9157), .B(n9156), .Z(c[1152]) );
  NANDN U11102 ( .A(n9124), .B(n9123), .Z(n9128) );
  NANDN U11103 ( .A(n9126), .B(n9125), .Z(n9127) );
  AND U11104 ( .A(n9128), .B(n9127), .Z(n9163) );
  NANDN U11105 ( .A(n9130), .B(n9129), .Z(n9134) );
  NANDN U11106 ( .A(n9132), .B(n9131), .Z(n9133) );
  AND U11107 ( .A(n9134), .B(n9133), .Z(n9161) );
  NAND U11108 ( .A(n42143), .B(n9135), .Z(n9137) );
  XNOR U11109 ( .A(a[131]), .B(n4090), .Z(n9172) );
  NAND U11110 ( .A(n42144), .B(n9172), .Z(n9136) );
  AND U11111 ( .A(n9137), .B(n9136), .Z(n9187) );
  XOR U11112 ( .A(a[135]), .B(n42012), .Z(n9175) );
  XNOR U11113 ( .A(n9187), .B(n9186), .Z(n9189) );
  AND U11114 ( .A(a[137]), .B(b[0]), .Z(n9139) );
  XNOR U11115 ( .A(n9139), .B(n4071), .Z(n9141) );
  NANDN U11116 ( .A(b[0]), .B(a[136]), .Z(n9140) );
  NAND U11117 ( .A(n9141), .B(n9140), .Z(n9183) );
  XOR U11118 ( .A(a[133]), .B(n42085), .Z(n9179) );
  AND U11119 ( .A(a[129]), .B(b[7]), .Z(n9180) );
  XNOR U11120 ( .A(n9181), .B(n9180), .Z(n9182) );
  XNOR U11121 ( .A(n9183), .B(n9182), .Z(n9188) );
  XOR U11122 ( .A(n9189), .B(n9188), .Z(n9167) );
  NANDN U11123 ( .A(n9144), .B(n9143), .Z(n9148) );
  NANDN U11124 ( .A(n9146), .B(n9145), .Z(n9147) );
  AND U11125 ( .A(n9148), .B(n9147), .Z(n9166) );
  XNOR U11126 ( .A(n9167), .B(n9166), .Z(n9168) );
  NANDN U11127 ( .A(n9150), .B(n9149), .Z(n9154) );
  NAND U11128 ( .A(n9152), .B(n9151), .Z(n9153) );
  NAND U11129 ( .A(n9154), .B(n9153), .Z(n9169) );
  XNOR U11130 ( .A(n9168), .B(n9169), .Z(n9160) );
  XNOR U11131 ( .A(n9161), .B(n9160), .Z(n9162) );
  XNOR U11132 ( .A(n9163), .B(n9162), .Z(n9192) );
  XNOR U11133 ( .A(sreg[1153]), .B(n9192), .Z(n9194) );
  NANDN U11134 ( .A(sreg[1152]), .B(n9155), .Z(n9159) );
  NAND U11135 ( .A(n9157), .B(n9156), .Z(n9158) );
  NAND U11136 ( .A(n9159), .B(n9158), .Z(n9193) );
  XNOR U11137 ( .A(n9194), .B(n9193), .Z(c[1153]) );
  NANDN U11138 ( .A(n9161), .B(n9160), .Z(n9165) );
  NANDN U11139 ( .A(n9163), .B(n9162), .Z(n9164) );
  AND U11140 ( .A(n9165), .B(n9164), .Z(n9200) );
  NANDN U11141 ( .A(n9167), .B(n9166), .Z(n9171) );
  NANDN U11142 ( .A(n9169), .B(n9168), .Z(n9170) );
  AND U11143 ( .A(n9171), .B(n9170), .Z(n9198) );
  NAND U11144 ( .A(n42143), .B(n9172), .Z(n9174) );
  XNOR U11145 ( .A(a[132]), .B(n4090), .Z(n9209) );
  NAND U11146 ( .A(n42144), .B(n9209), .Z(n9173) );
  AND U11147 ( .A(n9174), .B(n9173), .Z(n9224) );
  XOR U11148 ( .A(a[136]), .B(n42012), .Z(n9212) );
  XNOR U11149 ( .A(n9224), .B(n9223), .Z(n9226) );
  AND U11150 ( .A(a[138]), .B(b[0]), .Z(n9176) );
  XNOR U11151 ( .A(n9176), .B(n4071), .Z(n9178) );
  NANDN U11152 ( .A(b[0]), .B(a[137]), .Z(n9177) );
  NAND U11153 ( .A(n9178), .B(n9177), .Z(n9220) );
  XOR U11154 ( .A(a[134]), .B(n42085), .Z(n9216) );
  AND U11155 ( .A(a[130]), .B(b[7]), .Z(n9217) );
  XNOR U11156 ( .A(n9218), .B(n9217), .Z(n9219) );
  XNOR U11157 ( .A(n9220), .B(n9219), .Z(n9225) );
  XOR U11158 ( .A(n9226), .B(n9225), .Z(n9204) );
  NANDN U11159 ( .A(n9181), .B(n9180), .Z(n9185) );
  NANDN U11160 ( .A(n9183), .B(n9182), .Z(n9184) );
  AND U11161 ( .A(n9185), .B(n9184), .Z(n9203) );
  XNOR U11162 ( .A(n9204), .B(n9203), .Z(n9205) );
  NANDN U11163 ( .A(n9187), .B(n9186), .Z(n9191) );
  NAND U11164 ( .A(n9189), .B(n9188), .Z(n9190) );
  NAND U11165 ( .A(n9191), .B(n9190), .Z(n9206) );
  XNOR U11166 ( .A(n9205), .B(n9206), .Z(n9197) );
  XNOR U11167 ( .A(n9198), .B(n9197), .Z(n9199) );
  XNOR U11168 ( .A(n9200), .B(n9199), .Z(n9229) );
  XNOR U11169 ( .A(sreg[1154]), .B(n9229), .Z(n9231) );
  NANDN U11170 ( .A(sreg[1153]), .B(n9192), .Z(n9196) );
  NAND U11171 ( .A(n9194), .B(n9193), .Z(n9195) );
  NAND U11172 ( .A(n9196), .B(n9195), .Z(n9230) );
  XNOR U11173 ( .A(n9231), .B(n9230), .Z(c[1154]) );
  NANDN U11174 ( .A(n9198), .B(n9197), .Z(n9202) );
  NANDN U11175 ( .A(n9200), .B(n9199), .Z(n9201) );
  AND U11176 ( .A(n9202), .B(n9201), .Z(n9237) );
  NANDN U11177 ( .A(n9204), .B(n9203), .Z(n9208) );
  NANDN U11178 ( .A(n9206), .B(n9205), .Z(n9207) );
  AND U11179 ( .A(n9208), .B(n9207), .Z(n9235) );
  NAND U11180 ( .A(n42143), .B(n9209), .Z(n9211) );
  XNOR U11181 ( .A(a[133]), .B(n4090), .Z(n9246) );
  NAND U11182 ( .A(n42144), .B(n9246), .Z(n9210) );
  AND U11183 ( .A(n9211), .B(n9210), .Z(n9261) );
  XOR U11184 ( .A(a[137]), .B(n42012), .Z(n9249) );
  XNOR U11185 ( .A(n9261), .B(n9260), .Z(n9263) );
  AND U11186 ( .A(a[139]), .B(b[0]), .Z(n9213) );
  XNOR U11187 ( .A(n9213), .B(n4071), .Z(n9215) );
  NANDN U11188 ( .A(b[0]), .B(a[138]), .Z(n9214) );
  NAND U11189 ( .A(n9215), .B(n9214), .Z(n9257) );
  XOR U11190 ( .A(a[135]), .B(n42085), .Z(n9253) );
  AND U11191 ( .A(a[131]), .B(b[7]), .Z(n9254) );
  XNOR U11192 ( .A(n9255), .B(n9254), .Z(n9256) );
  XNOR U11193 ( .A(n9257), .B(n9256), .Z(n9262) );
  XOR U11194 ( .A(n9263), .B(n9262), .Z(n9241) );
  NANDN U11195 ( .A(n9218), .B(n9217), .Z(n9222) );
  NANDN U11196 ( .A(n9220), .B(n9219), .Z(n9221) );
  AND U11197 ( .A(n9222), .B(n9221), .Z(n9240) );
  XNOR U11198 ( .A(n9241), .B(n9240), .Z(n9242) );
  NANDN U11199 ( .A(n9224), .B(n9223), .Z(n9228) );
  NAND U11200 ( .A(n9226), .B(n9225), .Z(n9227) );
  NAND U11201 ( .A(n9228), .B(n9227), .Z(n9243) );
  XNOR U11202 ( .A(n9242), .B(n9243), .Z(n9234) );
  XNOR U11203 ( .A(n9235), .B(n9234), .Z(n9236) );
  XNOR U11204 ( .A(n9237), .B(n9236), .Z(n9266) );
  XNOR U11205 ( .A(sreg[1155]), .B(n9266), .Z(n9268) );
  NANDN U11206 ( .A(sreg[1154]), .B(n9229), .Z(n9233) );
  NAND U11207 ( .A(n9231), .B(n9230), .Z(n9232) );
  NAND U11208 ( .A(n9233), .B(n9232), .Z(n9267) );
  XNOR U11209 ( .A(n9268), .B(n9267), .Z(c[1155]) );
  NANDN U11210 ( .A(n9235), .B(n9234), .Z(n9239) );
  NANDN U11211 ( .A(n9237), .B(n9236), .Z(n9238) );
  AND U11212 ( .A(n9239), .B(n9238), .Z(n9274) );
  NANDN U11213 ( .A(n9241), .B(n9240), .Z(n9245) );
  NANDN U11214 ( .A(n9243), .B(n9242), .Z(n9244) );
  AND U11215 ( .A(n9245), .B(n9244), .Z(n9272) );
  NAND U11216 ( .A(n42143), .B(n9246), .Z(n9248) );
  XNOR U11217 ( .A(a[134]), .B(n4091), .Z(n9283) );
  NAND U11218 ( .A(n42144), .B(n9283), .Z(n9247) );
  AND U11219 ( .A(n9248), .B(n9247), .Z(n9298) );
  XOR U11220 ( .A(a[138]), .B(n42012), .Z(n9286) );
  XNOR U11221 ( .A(n9298), .B(n9297), .Z(n9300) );
  AND U11222 ( .A(a[140]), .B(b[0]), .Z(n9250) );
  XNOR U11223 ( .A(n9250), .B(n4071), .Z(n9252) );
  NANDN U11224 ( .A(b[0]), .B(a[139]), .Z(n9251) );
  NAND U11225 ( .A(n9252), .B(n9251), .Z(n9294) );
  XOR U11226 ( .A(a[136]), .B(n42085), .Z(n9290) );
  AND U11227 ( .A(a[132]), .B(b[7]), .Z(n9291) );
  XNOR U11228 ( .A(n9292), .B(n9291), .Z(n9293) );
  XNOR U11229 ( .A(n9294), .B(n9293), .Z(n9299) );
  XOR U11230 ( .A(n9300), .B(n9299), .Z(n9278) );
  NANDN U11231 ( .A(n9255), .B(n9254), .Z(n9259) );
  NANDN U11232 ( .A(n9257), .B(n9256), .Z(n9258) );
  AND U11233 ( .A(n9259), .B(n9258), .Z(n9277) );
  XNOR U11234 ( .A(n9278), .B(n9277), .Z(n9279) );
  NANDN U11235 ( .A(n9261), .B(n9260), .Z(n9265) );
  NAND U11236 ( .A(n9263), .B(n9262), .Z(n9264) );
  NAND U11237 ( .A(n9265), .B(n9264), .Z(n9280) );
  XNOR U11238 ( .A(n9279), .B(n9280), .Z(n9271) );
  XNOR U11239 ( .A(n9272), .B(n9271), .Z(n9273) );
  XNOR U11240 ( .A(n9274), .B(n9273), .Z(n9303) );
  XNOR U11241 ( .A(sreg[1156]), .B(n9303), .Z(n9305) );
  NANDN U11242 ( .A(sreg[1155]), .B(n9266), .Z(n9270) );
  NAND U11243 ( .A(n9268), .B(n9267), .Z(n9269) );
  NAND U11244 ( .A(n9270), .B(n9269), .Z(n9304) );
  XNOR U11245 ( .A(n9305), .B(n9304), .Z(c[1156]) );
  NANDN U11246 ( .A(n9272), .B(n9271), .Z(n9276) );
  NANDN U11247 ( .A(n9274), .B(n9273), .Z(n9275) );
  AND U11248 ( .A(n9276), .B(n9275), .Z(n9311) );
  NANDN U11249 ( .A(n9278), .B(n9277), .Z(n9282) );
  NANDN U11250 ( .A(n9280), .B(n9279), .Z(n9281) );
  AND U11251 ( .A(n9282), .B(n9281), .Z(n9309) );
  NAND U11252 ( .A(n42143), .B(n9283), .Z(n9285) );
  XNOR U11253 ( .A(a[135]), .B(n4091), .Z(n9320) );
  NAND U11254 ( .A(n42144), .B(n9320), .Z(n9284) );
  AND U11255 ( .A(n9285), .B(n9284), .Z(n9335) );
  XOR U11256 ( .A(a[139]), .B(n42012), .Z(n9323) );
  XNOR U11257 ( .A(n9335), .B(n9334), .Z(n9337) );
  AND U11258 ( .A(a[141]), .B(b[0]), .Z(n9287) );
  XNOR U11259 ( .A(n9287), .B(n4071), .Z(n9289) );
  NANDN U11260 ( .A(b[0]), .B(a[140]), .Z(n9288) );
  NAND U11261 ( .A(n9289), .B(n9288), .Z(n9331) );
  XOR U11262 ( .A(a[137]), .B(n42085), .Z(n9327) );
  AND U11263 ( .A(a[133]), .B(b[7]), .Z(n9328) );
  XNOR U11264 ( .A(n9329), .B(n9328), .Z(n9330) );
  XNOR U11265 ( .A(n9331), .B(n9330), .Z(n9336) );
  XOR U11266 ( .A(n9337), .B(n9336), .Z(n9315) );
  NANDN U11267 ( .A(n9292), .B(n9291), .Z(n9296) );
  NANDN U11268 ( .A(n9294), .B(n9293), .Z(n9295) );
  AND U11269 ( .A(n9296), .B(n9295), .Z(n9314) );
  XNOR U11270 ( .A(n9315), .B(n9314), .Z(n9316) );
  NANDN U11271 ( .A(n9298), .B(n9297), .Z(n9302) );
  NAND U11272 ( .A(n9300), .B(n9299), .Z(n9301) );
  NAND U11273 ( .A(n9302), .B(n9301), .Z(n9317) );
  XNOR U11274 ( .A(n9316), .B(n9317), .Z(n9308) );
  XNOR U11275 ( .A(n9309), .B(n9308), .Z(n9310) );
  XNOR U11276 ( .A(n9311), .B(n9310), .Z(n9340) );
  XNOR U11277 ( .A(sreg[1157]), .B(n9340), .Z(n9342) );
  NANDN U11278 ( .A(sreg[1156]), .B(n9303), .Z(n9307) );
  NAND U11279 ( .A(n9305), .B(n9304), .Z(n9306) );
  NAND U11280 ( .A(n9307), .B(n9306), .Z(n9341) );
  XNOR U11281 ( .A(n9342), .B(n9341), .Z(c[1157]) );
  NANDN U11282 ( .A(n9309), .B(n9308), .Z(n9313) );
  NANDN U11283 ( .A(n9311), .B(n9310), .Z(n9312) );
  AND U11284 ( .A(n9313), .B(n9312), .Z(n9348) );
  NANDN U11285 ( .A(n9315), .B(n9314), .Z(n9319) );
  NANDN U11286 ( .A(n9317), .B(n9316), .Z(n9318) );
  AND U11287 ( .A(n9319), .B(n9318), .Z(n9346) );
  NAND U11288 ( .A(n42143), .B(n9320), .Z(n9322) );
  XNOR U11289 ( .A(a[136]), .B(n4091), .Z(n9357) );
  NAND U11290 ( .A(n42144), .B(n9357), .Z(n9321) );
  AND U11291 ( .A(n9322), .B(n9321), .Z(n9372) );
  XOR U11292 ( .A(a[140]), .B(n42012), .Z(n9360) );
  XNOR U11293 ( .A(n9372), .B(n9371), .Z(n9374) );
  AND U11294 ( .A(a[142]), .B(b[0]), .Z(n9324) );
  XNOR U11295 ( .A(n9324), .B(n4071), .Z(n9326) );
  NANDN U11296 ( .A(b[0]), .B(a[141]), .Z(n9325) );
  NAND U11297 ( .A(n9326), .B(n9325), .Z(n9368) );
  XOR U11298 ( .A(a[138]), .B(n42085), .Z(n9364) );
  AND U11299 ( .A(a[134]), .B(b[7]), .Z(n9365) );
  XNOR U11300 ( .A(n9366), .B(n9365), .Z(n9367) );
  XNOR U11301 ( .A(n9368), .B(n9367), .Z(n9373) );
  XOR U11302 ( .A(n9374), .B(n9373), .Z(n9352) );
  NANDN U11303 ( .A(n9329), .B(n9328), .Z(n9333) );
  NANDN U11304 ( .A(n9331), .B(n9330), .Z(n9332) );
  AND U11305 ( .A(n9333), .B(n9332), .Z(n9351) );
  XNOR U11306 ( .A(n9352), .B(n9351), .Z(n9353) );
  NANDN U11307 ( .A(n9335), .B(n9334), .Z(n9339) );
  NAND U11308 ( .A(n9337), .B(n9336), .Z(n9338) );
  NAND U11309 ( .A(n9339), .B(n9338), .Z(n9354) );
  XNOR U11310 ( .A(n9353), .B(n9354), .Z(n9345) );
  XNOR U11311 ( .A(n9346), .B(n9345), .Z(n9347) );
  XNOR U11312 ( .A(n9348), .B(n9347), .Z(n9377) );
  XNOR U11313 ( .A(sreg[1158]), .B(n9377), .Z(n9379) );
  NANDN U11314 ( .A(sreg[1157]), .B(n9340), .Z(n9344) );
  NAND U11315 ( .A(n9342), .B(n9341), .Z(n9343) );
  NAND U11316 ( .A(n9344), .B(n9343), .Z(n9378) );
  XNOR U11317 ( .A(n9379), .B(n9378), .Z(c[1158]) );
  NANDN U11318 ( .A(n9346), .B(n9345), .Z(n9350) );
  NANDN U11319 ( .A(n9348), .B(n9347), .Z(n9349) );
  AND U11320 ( .A(n9350), .B(n9349), .Z(n9385) );
  NANDN U11321 ( .A(n9352), .B(n9351), .Z(n9356) );
  NANDN U11322 ( .A(n9354), .B(n9353), .Z(n9355) );
  AND U11323 ( .A(n9356), .B(n9355), .Z(n9383) );
  NAND U11324 ( .A(n42143), .B(n9357), .Z(n9359) );
  XNOR U11325 ( .A(a[137]), .B(n4091), .Z(n9394) );
  NAND U11326 ( .A(n42144), .B(n9394), .Z(n9358) );
  AND U11327 ( .A(n9359), .B(n9358), .Z(n9409) );
  XOR U11328 ( .A(a[141]), .B(n42012), .Z(n9397) );
  XNOR U11329 ( .A(n9409), .B(n9408), .Z(n9411) );
  AND U11330 ( .A(a[143]), .B(b[0]), .Z(n9361) );
  XNOR U11331 ( .A(n9361), .B(n4071), .Z(n9363) );
  NANDN U11332 ( .A(b[0]), .B(a[142]), .Z(n9362) );
  NAND U11333 ( .A(n9363), .B(n9362), .Z(n9405) );
  XOR U11334 ( .A(a[139]), .B(n42085), .Z(n9398) );
  AND U11335 ( .A(a[135]), .B(b[7]), .Z(n9402) );
  XNOR U11336 ( .A(n9403), .B(n9402), .Z(n9404) );
  XNOR U11337 ( .A(n9405), .B(n9404), .Z(n9410) );
  XOR U11338 ( .A(n9411), .B(n9410), .Z(n9389) );
  NANDN U11339 ( .A(n9366), .B(n9365), .Z(n9370) );
  NANDN U11340 ( .A(n9368), .B(n9367), .Z(n9369) );
  AND U11341 ( .A(n9370), .B(n9369), .Z(n9388) );
  XNOR U11342 ( .A(n9389), .B(n9388), .Z(n9390) );
  NANDN U11343 ( .A(n9372), .B(n9371), .Z(n9376) );
  NAND U11344 ( .A(n9374), .B(n9373), .Z(n9375) );
  NAND U11345 ( .A(n9376), .B(n9375), .Z(n9391) );
  XNOR U11346 ( .A(n9390), .B(n9391), .Z(n9382) );
  XNOR U11347 ( .A(n9383), .B(n9382), .Z(n9384) );
  XNOR U11348 ( .A(n9385), .B(n9384), .Z(n9414) );
  XNOR U11349 ( .A(sreg[1159]), .B(n9414), .Z(n9416) );
  NANDN U11350 ( .A(sreg[1158]), .B(n9377), .Z(n9381) );
  NAND U11351 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U11352 ( .A(n9381), .B(n9380), .Z(n9415) );
  XNOR U11353 ( .A(n9416), .B(n9415), .Z(c[1159]) );
  NANDN U11354 ( .A(n9383), .B(n9382), .Z(n9387) );
  NANDN U11355 ( .A(n9385), .B(n9384), .Z(n9386) );
  AND U11356 ( .A(n9387), .B(n9386), .Z(n9422) );
  NANDN U11357 ( .A(n9389), .B(n9388), .Z(n9393) );
  NANDN U11358 ( .A(n9391), .B(n9390), .Z(n9392) );
  AND U11359 ( .A(n9393), .B(n9392), .Z(n9420) );
  NAND U11360 ( .A(n42143), .B(n9394), .Z(n9396) );
  XNOR U11361 ( .A(a[138]), .B(n4091), .Z(n9431) );
  NAND U11362 ( .A(n42144), .B(n9431), .Z(n9395) );
  AND U11363 ( .A(n9396), .B(n9395), .Z(n9446) );
  XOR U11364 ( .A(a[142]), .B(n42012), .Z(n9434) );
  XNOR U11365 ( .A(n9446), .B(n9445), .Z(n9448) );
  XOR U11366 ( .A(a[140]), .B(n42085), .Z(n9435) );
  AND U11367 ( .A(a[136]), .B(b[7]), .Z(n9439) );
  XNOR U11368 ( .A(n9440), .B(n9439), .Z(n9441) );
  AND U11369 ( .A(a[144]), .B(b[0]), .Z(n9399) );
  XNOR U11370 ( .A(n9399), .B(n4071), .Z(n9401) );
  NANDN U11371 ( .A(b[0]), .B(a[143]), .Z(n9400) );
  NAND U11372 ( .A(n9401), .B(n9400), .Z(n9442) );
  XNOR U11373 ( .A(n9441), .B(n9442), .Z(n9447) );
  XOR U11374 ( .A(n9448), .B(n9447), .Z(n9426) );
  NANDN U11375 ( .A(n9403), .B(n9402), .Z(n9407) );
  NANDN U11376 ( .A(n9405), .B(n9404), .Z(n9406) );
  AND U11377 ( .A(n9407), .B(n9406), .Z(n9425) );
  XNOR U11378 ( .A(n9426), .B(n9425), .Z(n9427) );
  NANDN U11379 ( .A(n9409), .B(n9408), .Z(n9413) );
  NAND U11380 ( .A(n9411), .B(n9410), .Z(n9412) );
  NAND U11381 ( .A(n9413), .B(n9412), .Z(n9428) );
  XNOR U11382 ( .A(n9427), .B(n9428), .Z(n9419) );
  XNOR U11383 ( .A(n9420), .B(n9419), .Z(n9421) );
  XNOR U11384 ( .A(n9422), .B(n9421), .Z(n9451) );
  XNOR U11385 ( .A(sreg[1160]), .B(n9451), .Z(n9453) );
  NANDN U11386 ( .A(sreg[1159]), .B(n9414), .Z(n9418) );
  NAND U11387 ( .A(n9416), .B(n9415), .Z(n9417) );
  NAND U11388 ( .A(n9418), .B(n9417), .Z(n9452) );
  XNOR U11389 ( .A(n9453), .B(n9452), .Z(c[1160]) );
  NANDN U11390 ( .A(n9420), .B(n9419), .Z(n9424) );
  NANDN U11391 ( .A(n9422), .B(n9421), .Z(n9423) );
  AND U11392 ( .A(n9424), .B(n9423), .Z(n9459) );
  NANDN U11393 ( .A(n9426), .B(n9425), .Z(n9430) );
  NANDN U11394 ( .A(n9428), .B(n9427), .Z(n9429) );
  AND U11395 ( .A(n9430), .B(n9429), .Z(n9457) );
  NAND U11396 ( .A(n42143), .B(n9431), .Z(n9433) );
  XNOR U11397 ( .A(a[139]), .B(n4091), .Z(n9468) );
  NAND U11398 ( .A(n42144), .B(n9468), .Z(n9432) );
  AND U11399 ( .A(n9433), .B(n9432), .Z(n9483) );
  XOR U11400 ( .A(a[143]), .B(n42012), .Z(n9471) );
  XNOR U11401 ( .A(n9483), .B(n9482), .Z(n9485) );
  XOR U11402 ( .A(a[141]), .B(n42085), .Z(n9475) );
  AND U11403 ( .A(a[137]), .B(b[7]), .Z(n9476) );
  XNOR U11404 ( .A(n9477), .B(n9476), .Z(n9478) );
  AND U11405 ( .A(a[145]), .B(b[0]), .Z(n9436) );
  XNOR U11406 ( .A(n9436), .B(n4071), .Z(n9438) );
  NANDN U11407 ( .A(b[0]), .B(a[144]), .Z(n9437) );
  NAND U11408 ( .A(n9438), .B(n9437), .Z(n9479) );
  XNOR U11409 ( .A(n9478), .B(n9479), .Z(n9484) );
  XOR U11410 ( .A(n9485), .B(n9484), .Z(n9463) );
  NANDN U11411 ( .A(n9440), .B(n9439), .Z(n9444) );
  NANDN U11412 ( .A(n9442), .B(n9441), .Z(n9443) );
  AND U11413 ( .A(n9444), .B(n9443), .Z(n9462) );
  XNOR U11414 ( .A(n9463), .B(n9462), .Z(n9464) );
  NANDN U11415 ( .A(n9446), .B(n9445), .Z(n9450) );
  NAND U11416 ( .A(n9448), .B(n9447), .Z(n9449) );
  NAND U11417 ( .A(n9450), .B(n9449), .Z(n9465) );
  XNOR U11418 ( .A(n9464), .B(n9465), .Z(n9456) );
  XNOR U11419 ( .A(n9457), .B(n9456), .Z(n9458) );
  XNOR U11420 ( .A(n9459), .B(n9458), .Z(n9488) );
  XNOR U11421 ( .A(sreg[1161]), .B(n9488), .Z(n9490) );
  NANDN U11422 ( .A(sreg[1160]), .B(n9451), .Z(n9455) );
  NAND U11423 ( .A(n9453), .B(n9452), .Z(n9454) );
  NAND U11424 ( .A(n9455), .B(n9454), .Z(n9489) );
  XNOR U11425 ( .A(n9490), .B(n9489), .Z(c[1161]) );
  NANDN U11426 ( .A(n9457), .B(n9456), .Z(n9461) );
  NANDN U11427 ( .A(n9459), .B(n9458), .Z(n9460) );
  AND U11428 ( .A(n9461), .B(n9460), .Z(n9496) );
  NANDN U11429 ( .A(n9463), .B(n9462), .Z(n9467) );
  NANDN U11430 ( .A(n9465), .B(n9464), .Z(n9466) );
  AND U11431 ( .A(n9467), .B(n9466), .Z(n9494) );
  NAND U11432 ( .A(n42143), .B(n9468), .Z(n9470) );
  XNOR U11433 ( .A(a[140]), .B(n4091), .Z(n9505) );
  NAND U11434 ( .A(n42144), .B(n9505), .Z(n9469) );
  AND U11435 ( .A(n9470), .B(n9469), .Z(n9520) );
  XOR U11436 ( .A(a[144]), .B(n42012), .Z(n9508) );
  XNOR U11437 ( .A(n9520), .B(n9519), .Z(n9522) );
  AND U11438 ( .A(a[146]), .B(b[0]), .Z(n9472) );
  XNOR U11439 ( .A(n9472), .B(n4071), .Z(n9474) );
  NANDN U11440 ( .A(b[0]), .B(a[145]), .Z(n9473) );
  NAND U11441 ( .A(n9474), .B(n9473), .Z(n9516) );
  XOR U11442 ( .A(a[142]), .B(n42085), .Z(n9509) );
  AND U11443 ( .A(a[138]), .B(b[7]), .Z(n9513) );
  XNOR U11444 ( .A(n9514), .B(n9513), .Z(n9515) );
  XNOR U11445 ( .A(n9516), .B(n9515), .Z(n9521) );
  XOR U11446 ( .A(n9522), .B(n9521), .Z(n9500) );
  NANDN U11447 ( .A(n9477), .B(n9476), .Z(n9481) );
  NANDN U11448 ( .A(n9479), .B(n9478), .Z(n9480) );
  AND U11449 ( .A(n9481), .B(n9480), .Z(n9499) );
  XNOR U11450 ( .A(n9500), .B(n9499), .Z(n9501) );
  NANDN U11451 ( .A(n9483), .B(n9482), .Z(n9487) );
  NAND U11452 ( .A(n9485), .B(n9484), .Z(n9486) );
  NAND U11453 ( .A(n9487), .B(n9486), .Z(n9502) );
  XNOR U11454 ( .A(n9501), .B(n9502), .Z(n9493) );
  XNOR U11455 ( .A(n9494), .B(n9493), .Z(n9495) );
  XNOR U11456 ( .A(n9496), .B(n9495), .Z(n9525) );
  XNOR U11457 ( .A(sreg[1162]), .B(n9525), .Z(n9527) );
  NANDN U11458 ( .A(sreg[1161]), .B(n9488), .Z(n9492) );
  NAND U11459 ( .A(n9490), .B(n9489), .Z(n9491) );
  NAND U11460 ( .A(n9492), .B(n9491), .Z(n9526) );
  XNOR U11461 ( .A(n9527), .B(n9526), .Z(c[1162]) );
  NANDN U11462 ( .A(n9494), .B(n9493), .Z(n9498) );
  NANDN U11463 ( .A(n9496), .B(n9495), .Z(n9497) );
  AND U11464 ( .A(n9498), .B(n9497), .Z(n9533) );
  NANDN U11465 ( .A(n9500), .B(n9499), .Z(n9504) );
  NANDN U11466 ( .A(n9502), .B(n9501), .Z(n9503) );
  AND U11467 ( .A(n9504), .B(n9503), .Z(n9531) );
  NAND U11468 ( .A(n42143), .B(n9505), .Z(n9507) );
  XNOR U11469 ( .A(a[141]), .B(n4092), .Z(n9542) );
  NAND U11470 ( .A(n42144), .B(n9542), .Z(n9506) );
  AND U11471 ( .A(n9507), .B(n9506), .Z(n9557) );
  XOR U11472 ( .A(a[145]), .B(n42012), .Z(n9545) );
  XNOR U11473 ( .A(n9557), .B(n9556), .Z(n9559) );
  XOR U11474 ( .A(a[143]), .B(n42085), .Z(n9546) );
  AND U11475 ( .A(a[139]), .B(b[7]), .Z(n9550) );
  XNOR U11476 ( .A(n9551), .B(n9550), .Z(n9552) );
  AND U11477 ( .A(a[147]), .B(b[0]), .Z(n9510) );
  XNOR U11478 ( .A(n9510), .B(n4071), .Z(n9512) );
  NANDN U11479 ( .A(b[0]), .B(a[146]), .Z(n9511) );
  NAND U11480 ( .A(n9512), .B(n9511), .Z(n9553) );
  XNOR U11481 ( .A(n9552), .B(n9553), .Z(n9558) );
  XOR U11482 ( .A(n9559), .B(n9558), .Z(n9537) );
  NANDN U11483 ( .A(n9514), .B(n9513), .Z(n9518) );
  NANDN U11484 ( .A(n9516), .B(n9515), .Z(n9517) );
  AND U11485 ( .A(n9518), .B(n9517), .Z(n9536) );
  XNOR U11486 ( .A(n9537), .B(n9536), .Z(n9538) );
  NANDN U11487 ( .A(n9520), .B(n9519), .Z(n9524) );
  NAND U11488 ( .A(n9522), .B(n9521), .Z(n9523) );
  NAND U11489 ( .A(n9524), .B(n9523), .Z(n9539) );
  XNOR U11490 ( .A(n9538), .B(n9539), .Z(n9530) );
  XNOR U11491 ( .A(n9531), .B(n9530), .Z(n9532) );
  XNOR U11492 ( .A(n9533), .B(n9532), .Z(n9562) );
  XNOR U11493 ( .A(sreg[1163]), .B(n9562), .Z(n9564) );
  NANDN U11494 ( .A(sreg[1162]), .B(n9525), .Z(n9529) );
  NAND U11495 ( .A(n9527), .B(n9526), .Z(n9528) );
  NAND U11496 ( .A(n9529), .B(n9528), .Z(n9563) );
  XNOR U11497 ( .A(n9564), .B(n9563), .Z(c[1163]) );
  NANDN U11498 ( .A(n9531), .B(n9530), .Z(n9535) );
  NANDN U11499 ( .A(n9533), .B(n9532), .Z(n9534) );
  AND U11500 ( .A(n9535), .B(n9534), .Z(n9570) );
  NANDN U11501 ( .A(n9537), .B(n9536), .Z(n9541) );
  NANDN U11502 ( .A(n9539), .B(n9538), .Z(n9540) );
  AND U11503 ( .A(n9541), .B(n9540), .Z(n9568) );
  NAND U11504 ( .A(n42143), .B(n9542), .Z(n9544) );
  XNOR U11505 ( .A(a[142]), .B(n4092), .Z(n9579) );
  NAND U11506 ( .A(n42144), .B(n9579), .Z(n9543) );
  AND U11507 ( .A(n9544), .B(n9543), .Z(n9594) );
  XOR U11508 ( .A(a[146]), .B(n42012), .Z(n9582) );
  XNOR U11509 ( .A(n9594), .B(n9593), .Z(n9596) );
  XOR U11510 ( .A(a[144]), .B(n42085), .Z(n9586) );
  AND U11511 ( .A(a[140]), .B(b[7]), .Z(n9587) );
  XNOR U11512 ( .A(n9588), .B(n9587), .Z(n9589) );
  AND U11513 ( .A(a[148]), .B(b[0]), .Z(n9547) );
  XNOR U11514 ( .A(n9547), .B(n4071), .Z(n9549) );
  NANDN U11515 ( .A(b[0]), .B(a[147]), .Z(n9548) );
  NAND U11516 ( .A(n9549), .B(n9548), .Z(n9590) );
  XNOR U11517 ( .A(n9589), .B(n9590), .Z(n9595) );
  XOR U11518 ( .A(n9596), .B(n9595), .Z(n9574) );
  NANDN U11519 ( .A(n9551), .B(n9550), .Z(n9555) );
  NANDN U11520 ( .A(n9553), .B(n9552), .Z(n9554) );
  AND U11521 ( .A(n9555), .B(n9554), .Z(n9573) );
  XNOR U11522 ( .A(n9574), .B(n9573), .Z(n9575) );
  NANDN U11523 ( .A(n9557), .B(n9556), .Z(n9561) );
  NAND U11524 ( .A(n9559), .B(n9558), .Z(n9560) );
  NAND U11525 ( .A(n9561), .B(n9560), .Z(n9576) );
  XNOR U11526 ( .A(n9575), .B(n9576), .Z(n9567) );
  XNOR U11527 ( .A(n9568), .B(n9567), .Z(n9569) );
  XNOR U11528 ( .A(n9570), .B(n9569), .Z(n9599) );
  XNOR U11529 ( .A(sreg[1164]), .B(n9599), .Z(n9601) );
  NANDN U11530 ( .A(sreg[1163]), .B(n9562), .Z(n9566) );
  NAND U11531 ( .A(n9564), .B(n9563), .Z(n9565) );
  NAND U11532 ( .A(n9566), .B(n9565), .Z(n9600) );
  XNOR U11533 ( .A(n9601), .B(n9600), .Z(c[1164]) );
  NANDN U11534 ( .A(n9568), .B(n9567), .Z(n9572) );
  NANDN U11535 ( .A(n9570), .B(n9569), .Z(n9571) );
  AND U11536 ( .A(n9572), .B(n9571), .Z(n9607) );
  NANDN U11537 ( .A(n9574), .B(n9573), .Z(n9578) );
  NANDN U11538 ( .A(n9576), .B(n9575), .Z(n9577) );
  AND U11539 ( .A(n9578), .B(n9577), .Z(n9605) );
  NAND U11540 ( .A(n42143), .B(n9579), .Z(n9581) );
  XNOR U11541 ( .A(a[143]), .B(n4092), .Z(n9616) );
  NAND U11542 ( .A(n42144), .B(n9616), .Z(n9580) );
  AND U11543 ( .A(n9581), .B(n9580), .Z(n9631) );
  XOR U11544 ( .A(a[147]), .B(n42012), .Z(n9619) );
  XNOR U11545 ( .A(n9631), .B(n9630), .Z(n9633) );
  AND U11546 ( .A(a[149]), .B(b[0]), .Z(n9583) );
  XNOR U11547 ( .A(n9583), .B(n4071), .Z(n9585) );
  NANDN U11548 ( .A(b[0]), .B(a[148]), .Z(n9584) );
  NAND U11549 ( .A(n9585), .B(n9584), .Z(n9627) );
  XOR U11550 ( .A(a[145]), .B(n42085), .Z(n9623) );
  AND U11551 ( .A(a[141]), .B(b[7]), .Z(n9624) );
  XNOR U11552 ( .A(n9625), .B(n9624), .Z(n9626) );
  XNOR U11553 ( .A(n9627), .B(n9626), .Z(n9632) );
  XOR U11554 ( .A(n9633), .B(n9632), .Z(n9611) );
  NANDN U11555 ( .A(n9588), .B(n9587), .Z(n9592) );
  NANDN U11556 ( .A(n9590), .B(n9589), .Z(n9591) );
  AND U11557 ( .A(n9592), .B(n9591), .Z(n9610) );
  XNOR U11558 ( .A(n9611), .B(n9610), .Z(n9612) );
  NANDN U11559 ( .A(n9594), .B(n9593), .Z(n9598) );
  NAND U11560 ( .A(n9596), .B(n9595), .Z(n9597) );
  NAND U11561 ( .A(n9598), .B(n9597), .Z(n9613) );
  XNOR U11562 ( .A(n9612), .B(n9613), .Z(n9604) );
  XNOR U11563 ( .A(n9605), .B(n9604), .Z(n9606) );
  XNOR U11564 ( .A(n9607), .B(n9606), .Z(n9636) );
  XNOR U11565 ( .A(sreg[1165]), .B(n9636), .Z(n9638) );
  NANDN U11566 ( .A(sreg[1164]), .B(n9599), .Z(n9603) );
  NAND U11567 ( .A(n9601), .B(n9600), .Z(n9602) );
  NAND U11568 ( .A(n9603), .B(n9602), .Z(n9637) );
  XNOR U11569 ( .A(n9638), .B(n9637), .Z(c[1165]) );
  NANDN U11570 ( .A(n9605), .B(n9604), .Z(n9609) );
  NANDN U11571 ( .A(n9607), .B(n9606), .Z(n9608) );
  AND U11572 ( .A(n9609), .B(n9608), .Z(n9644) );
  NANDN U11573 ( .A(n9611), .B(n9610), .Z(n9615) );
  NANDN U11574 ( .A(n9613), .B(n9612), .Z(n9614) );
  AND U11575 ( .A(n9615), .B(n9614), .Z(n9642) );
  NAND U11576 ( .A(n42143), .B(n9616), .Z(n9618) );
  XNOR U11577 ( .A(a[144]), .B(n4092), .Z(n9653) );
  NAND U11578 ( .A(n42144), .B(n9653), .Z(n9617) );
  AND U11579 ( .A(n9618), .B(n9617), .Z(n9668) );
  XOR U11580 ( .A(a[148]), .B(n42012), .Z(n9656) );
  XNOR U11581 ( .A(n9668), .B(n9667), .Z(n9670) );
  AND U11582 ( .A(a[150]), .B(b[0]), .Z(n9620) );
  XNOR U11583 ( .A(n9620), .B(n4071), .Z(n9622) );
  NANDN U11584 ( .A(b[0]), .B(a[149]), .Z(n9621) );
  NAND U11585 ( .A(n9622), .B(n9621), .Z(n9664) );
  XOR U11586 ( .A(a[146]), .B(n42085), .Z(n9657) );
  AND U11587 ( .A(a[142]), .B(b[7]), .Z(n9661) );
  XNOR U11588 ( .A(n9662), .B(n9661), .Z(n9663) );
  XNOR U11589 ( .A(n9664), .B(n9663), .Z(n9669) );
  XOR U11590 ( .A(n9670), .B(n9669), .Z(n9648) );
  NANDN U11591 ( .A(n9625), .B(n9624), .Z(n9629) );
  NANDN U11592 ( .A(n9627), .B(n9626), .Z(n9628) );
  AND U11593 ( .A(n9629), .B(n9628), .Z(n9647) );
  XNOR U11594 ( .A(n9648), .B(n9647), .Z(n9649) );
  NANDN U11595 ( .A(n9631), .B(n9630), .Z(n9635) );
  NAND U11596 ( .A(n9633), .B(n9632), .Z(n9634) );
  NAND U11597 ( .A(n9635), .B(n9634), .Z(n9650) );
  XNOR U11598 ( .A(n9649), .B(n9650), .Z(n9641) );
  XNOR U11599 ( .A(n9642), .B(n9641), .Z(n9643) );
  XNOR U11600 ( .A(n9644), .B(n9643), .Z(n9673) );
  XNOR U11601 ( .A(sreg[1166]), .B(n9673), .Z(n9675) );
  NANDN U11602 ( .A(sreg[1165]), .B(n9636), .Z(n9640) );
  NAND U11603 ( .A(n9638), .B(n9637), .Z(n9639) );
  NAND U11604 ( .A(n9640), .B(n9639), .Z(n9674) );
  XNOR U11605 ( .A(n9675), .B(n9674), .Z(c[1166]) );
  NANDN U11606 ( .A(n9642), .B(n9641), .Z(n9646) );
  NANDN U11607 ( .A(n9644), .B(n9643), .Z(n9645) );
  AND U11608 ( .A(n9646), .B(n9645), .Z(n9685) );
  NANDN U11609 ( .A(n9648), .B(n9647), .Z(n9652) );
  NANDN U11610 ( .A(n9650), .B(n9649), .Z(n9651) );
  AND U11611 ( .A(n9652), .B(n9651), .Z(n9684) );
  NAND U11612 ( .A(n42143), .B(n9653), .Z(n9655) );
  XNOR U11613 ( .A(a[145]), .B(n4092), .Z(n9695) );
  NAND U11614 ( .A(n42144), .B(n9695), .Z(n9654) );
  AND U11615 ( .A(n9655), .B(n9654), .Z(n9710) );
  XOR U11616 ( .A(a[149]), .B(n42012), .Z(n9698) );
  XNOR U11617 ( .A(n9710), .B(n9709), .Z(n9712) );
  XOR U11618 ( .A(a[147]), .B(n42085), .Z(n9702) );
  AND U11619 ( .A(a[143]), .B(b[7]), .Z(n9703) );
  XNOR U11620 ( .A(n9704), .B(n9703), .Z(n9705) );
  AND U11621 ( .A(a[151]), .B(b[0]), .Z(n9658) );
  XNOR U11622 ( .A(n9658), .B(n4071), .Z(n9660) );
  NANDN U11623 ( .A(b[0]), .B(a[150]), .Z(n9659) );
  NAND U11624 ( .A(n9660), .B(n9659), .Z(n9706) );
  XNOR U11625 ( .A(n9705), .B(n9706), .Z(n9711) );
  XOR U11626 ( .A(n9712), .B(n9711), .Z(n9690) );
  NANDN U11627 ( .A(n9662), .B(n9661), .Z(n9666) );
  NANDN U11628 ( .A(n9664), .B(n9663), .Z(n9665) );
  AND U11629 ( .A(n9666), .B(n9665), .Z(n9689) );
  XNOR U11630 ( .A(n9690), .B(n9689), .Z(n9691) );
  NANDN U11631 ( .A(n9668), .B(n9667), .Z(n9672) );
  NAND U11632 ( .A(n9670), .B(n9669), .Z(n9671) );
  NAND U11633 ( .A(n9672), .B(n9671), .Z(n9692) );
  XNOR U11634 ( .A(n9691), .B(n9692), .Z(n9683) );
  XOR U11635 ( .A(n9684), .B(n9683), .Z(n9686) );
  XOR U11636 ( .A(n9685), .B(n9686), .Z(n9678) );
  XNOR U11637 ( .A(n9678), .B(sreg[1167]), .Z(n9680) );
  NANDN U11638 ( .A(sreg[1166]), .B(n9673), .Z(n9677) );
  NAND U11639 ( .A(n9675), .B(n9674), .Z(n9676) );
  AND U11640 ( .A(n9677), .B(n9676), .Z(n9679) );
  XOR U11641 ( .A(n9680), .B(n9679), .Z(c[1167]) );
  NANDN U11642 ( .A(n9678), .B(sreg[1167]), .Z(n9682) );
  NAND U11643 ( .A(n9680), .B(n9679), .Z(n9681) );
  AND U11644 ( .A(n9682), .B(n9681), .Z(n9749) );
  NANDN U11645 ( .A(n9684), .B(n9683), .Z(n9688) );
  OR U11646 ( .A(n9686), .B(n9685), .Z(n9687) );
  AND U11647 ( .A(n9688), .B(n9687), .Z(n9718) );
  NANDN U11648 ( .A(n9690), .B(n9689), .Z(n9694) );
  NANDN U11649 ( .A(n9692), .B(n9691), .Z(n9693) );
  AND U11650 ( .A(n9694), .B(n9693), .Z(n9716) );
  NAND U11651 ( .A(n42143), .B(n9695), .Z(n9697) );
  XNOR U11652 ( .A(a[146]), .B(n4092), .Z(n9727) );
  NAND U11653 ( .A(n42144), .B(n9727), .Z(n9696) );
  AND U11654 ( .A(n9697), .B(n9696), .Z(n9742) );
  XOR U11655 ( .A(a[150]), .B(n42012), .Z(n9730) );
  XNOR U11656 ( .A(n9742), .B(n9741), .Z(n9744) );
  AND U11657 ( .A(a[152]), .B(b[0]), .Z(n9699) );
  XNOR U11658 ( .A(n9699), .B(n4071), .Z(n9701) );
  NANDN U11659 ( .A(b[0]), .B(a[151]), .Z(n9700) );
  NAND U11660 ( .A(n9701), .B(n9700), .Z(n9738) );
  XOR U11661 ( .A(a[148]), .B(n42085), .Z(n9734) );
  AND U11662 ( .A(a[144]), .B(b[7]), .Z(n9735) );
  XNOR U11663 ( .A(n9736), .B(n9735), .Z(n9737) );
  XNOR U11664 ( .A(n9738), .B(n9737), .Z(n9743) );
  XOR U11665 ( .A(n9744), .B(n9743), .Z(n9722) );
  NANDN U11666 ( .A(n9704), .B(n9703), .Z(n9708) );
  NANDN U11667 ( .A(n9706), .B(n9705), .Z(n9707) );
  AND U11668 ( .A(n9708), .B(n9707), .Z(n9721) );
  XNOR U11669 ( .A(n9722), .B(n9721), .Z(n9723) );
  NANDN U11670 ( .A(n9710), .B(n9709), .Z(n9714) );
  NAND U11671 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U11672 ( .A(n9714), .B(n9713), .Z(n9724) );
  XNOR U11673 ( .A(n9723), .B(n9724), .Z(n9715) );
  XNOR U11674 ( .A(n9716), .B(n9715), .Z(n9717) );
  XNOR U11675 ( .A(n9718), .B(n9717), .Z(n9747) );
  XNOR U11676 ( .A(sreg[1168]), .B(n9747), .Z(n9748) );
  XNOR U11677 ( .A(n9749), .B(n9748), .Z(c[1168]) );
  NANDN U11678 ( .A(n9716), .B(n9715), .Z(n9720) );
  NANDN U11679 ( .A(n9718), .B(n9717), .Z(n9719) );
  AND U11680 ( .A(n9720), .B(n9719), .Z(n9755) );
  NANDN U11681 ( .A(n9722), .B(n9721), .Z(n9726) );
  NANDN U11682 ( .A(n9724), .B(n9723), .Z(n9725) );
  AND U11683 ( .A(n9726), .B(n9725), .Z(n9753) );
  NAND U11684 ( .A(n42143), .B(n9727), .Z(n9729) );
  XNOR U11685 ( .A(a[147]), .B(n4092), .Z(n9764) );
  NAND U11686 ( .A(n42144), .B(n9764), .Z(n9728) );
  AND U11687 ( .A(n9729), .B(n9728), .Z(n9779) );
  XOR U11688 ( .A(a[151]), .B(n42012), .Z(n9767) );
  XNOR U11689 ( .A(n9779), .B(n9778), .Z(n9781) );
  AND U11690 ( .A(a[153]), .B(b[0]), .Z(n9731) );
  XNOR U11691 ( .A(n9731), .B(n4071), .Z(n9733) );
  NANDN U11692 ( .A(b[0]), .B(a[152]), .Z(n9732) );
  NAND U11693 ( .A(n9733), .B(n9732), .Z(n9775) );
  XOR U11694 ( .A(a[149]), .B(n42085), .Z(n9771) );
  AND U11695 ( .A(a[145]), .B(b[7]), .Z(n9772) );
  XNOR U11696 ( .A(n9773), .B(n9772), .Z(n9774) );
  XNOR U11697 ( .A(n9775), .B(n9774), .Z(n9780) );
  XOR U11698 ( .A(n9781), .B(n9780), .Z(n9759) );
  NANDN U11699 ( .A(n9736), .B(n9735), .Z(n9740) );
  NANDN U11700 ( .A(n9738), .B(n9737), .Z(n9739) );
  AND U11701 ( .A(n9740), .B(n9739), .Z(n9758) );
  XNOR U11702 ( .A(n9759), .B(n9758), .Z(n9760) );
  NANDN U11703 ( .A(n9742), .B(n9741), .Z(n9746) );
  NAND U11704 ( .A(n9744), .B(n9743), .Z(n9745) );
  NAND U11705 ( .A(n9746), .B(n9745), .Z(n9761) );
  XNOR U11706 ( .A(n9760), .B(n9761), .Z(n9752) );
  XNOR U11707 ( .A(n9753), .B(n9752), .Z(n9754) );
  XNOR U11708 ( .A(n9755), .B(n9754), .Z(n9784) );
  XNOR U11709 ( .A(sreg[1169]), .B(n9784), .Z(n9786) );
  NANDN U11710 ( .A(sreg[1168]), .B(n9747), .Z(n9751) );
  NAND U11711 ( .A(n9749), .B(n9748), .Z(n9750) );
  NAND U11712 ( .A(n9751), .B(n9750), .Z(n9785) );
  XNOR U11713 ( .A(n9786), .B(n9785), .Z(c[1169]) );
  NANDN U11714 ( .A(n9753), .B(n9752), .Z(n9757) );
  NANDN U11715 ( .A(n9755), .B(n9754), .Z(n9756) );
  AND U11716 ( .A(n9757), .B(n9756), .Z(n9792) );
  NANDN U11717 ( .A(n9759), .B(n9758), .Z(n9763) );
  NANDN U11718 ( .A(n9761), .B(n9760), .Z(n9762) );
  AND U11719 ( .A(n9763), .B(n9762), .Z(n9790) );
  NAND U11720 ( .A(n42143), .B(n9764), .Z(n9766) );
  XNOR U11721 ( .A(a[148]), .B(n4093), .Z(n9801) );
  NAND U11722 ( .A(n42144), .B(n9801), .Z(n9765) );
  AND U11723 ( .A(n9766), .B(n9765), .Z(n9816) );
  XOR U11724 ( .A(a[152]), .B(n42012), .Z(n9804) );
  XNOR U11725 ( .A(n9816), .B(n9815), .Z(n9818) );
  AND U11726 ( .A(a[154]), .B(b[0]), .Z(n9768) );
  XNOR U11727 ( .A(n9768), .B(n4071), .Z(n9770) );
  NANDN U11728 ( .A(b[0]), .B(a[153]), .Z(n9769) );
  NAND U11729 ( .A(n9770), .B(n9769), .Z(n9812) );
  XOR U11730 ( .A(a[150]), .B(n42085), .Z(n9808) );
  AND U11731 ( .A(a[146]), .B(b[7]), .Z(n9809) );
  XNOR U11732 ( .A(n9810), .B(n9809), .Z(n9811) );
  XNOR U11733 ( .A(n9812), .B(n9811), .Z(n9817) );
  XOR U11734 ( .A(n9818), .B(n9817), .Z(n9796) );
  NANDN U11735 ( .A(n9773), .B(n9772), .Z(n9777) );
  NANDN U11736 ( .A(n9775), .B(n9774), .Z(n9776) );
  AND U11737 ( .A(n9777), .B(n9776), .Z(n9795) );
  XNOR U11738 ( .A(n9796), .B(n9795), .Z(n9797) );
  NANDN U11739 ( .A(n9779), .B(n9778), .Z(n9783) );
  NAND U11740 ( .A(n9781), .B(n9780), .Z(n9782) );
  NAND U11741 ( .A(n9783), .B(n9782), .Z(n9798) );
  XNOR U11742 ( .A(n9797), .B(n9798), .Z(n9789) );
  XNOR U11743 ( .A(n9790), .B(n9789), .Z(n9791) );
  XNOR U11744 ( .A(n9792), .B(n9791), .Z(n9821) );
  XNOR U11745 ( .A(sreg[1170]), .B(n9821), .Z(n9823) );
  NANDN U11746 ( .A(sreg[1169]), .B(n9784), .Z(n9788) );
  NAND U11747 ( .A(n9786), .B(n9785), .Z(n9787) );
  NAND U11748 ( .A(n9788), .B(n9787), .Z(n9822) );
  XNOR U11749 ( .A(n9823), .B(n9822), .Z(c[1170]) );
  NANDN U11750 ( .A(n9790), .B(n9789), .Z(n9794) );
  NANDN U11751 ( .A(n9792), .B(n9791), .Z(n9793) );
  AND U11752 ( .A(n9794), .B(n9793), .Z(n9829) );
  NANDN U11753 ( .A(n9796), .B(n9795), .Z(n9800) );
  NANDN U11754 ( .A(n9798), .B(n9797), .Z(n9799) );
  AND U11755 ( .A(n9800), .B(n9799), .Z(n9827) );
  NAND U11756 ( .A(n42143), .B(n9801), .Z(n9803) );
  XNOR U11757 ( .A(a[149]), .B(n4093), .Z(n9838) );
  NAND U11758 ( .A(n42144), .B(n9838), .Z(n9802) );
  AND U11759 ( .A(n9803), .B(n9802), .Z(n9853) );
  XOR U11760 ( .A(a[153]), .B(n42012), .Z(n9841) );
  XNOR U11761 ( .A(n9853), .B(n9852), .Z(n9855) );
  AND U11762 ( .A(a[155]), .B(b[0]), .Z(n9805) );
  XNOR U11763 ( .A(n9805), .B(n4071), .Z(n9807) );
  NANDN U11764 ( .A(b[0]), .B(a[154]), .Z(n9806) );
  NAND U11765 ( .A(n9807), .B(n9806), .Z(n9849) );
  XOR U11766 ( .A(a[151]), .B(n42085), .Z(n9842) );
  AND U11767 ( .A(a[147]), .B(b[7]), .Z(n9846) );
  XNOR U11768 ( .A(n9847), .B(n9846), .Z(n9848) );
  XNOR U11769 ( .A(n9849), .B(n9848), .Z(n9854) );
  XOR U11770 ( .A(n9855), .B(n9854), .Z(n9833) );
  NANDN U11771 ( .A(n9810), .B(n9809), .Z(n9814) );
  NANDN U11772 ( .A(n9812), .B(n9811), .Z(n9813) );
  AND U11773 ( .A(n9814), .B(n9813), .Z(n9832) );
  XNOR U11774 ( .A(n9833), .B(n9832), .Z(n9834) );
  NANDN U11775 ( .A(n9816), .B(n9815), .Z(n9820) );
  NAND U11776 ( .A(n9818), .B(n9817), .Z(n9819) );
  NAND U11777 ( .A(n9820), .B(n9819), .Z(n9835) );
  XNOR U11778 ( .A(n9834), .B(n9835), .Z(n9826) );
  XNOR U11779 ( .A(n9827), .B(n9826), .Z(n9828) );
  XNOR U11780 ( .A(n9829), .B(n9828), .Z(n9858) );
  XNOR U11781 ( .A(sreg[1171]), .B(n9858), .Z(n9860) );
  NANDN U11782 ( .A(sreg[1170]), .B(n9821), .Z(n9825) );
  NAND U11783 ( .A(n9823), .B(n9822), .Z(n9824) );
  NAND U11784 ( .A(n9825), .B(n9824), .Z(n9859) );
  XNOR U11785 ( .A(n9860), .B(n9859), .Z(c[1171]) );
  NANDN U11786 ( .A(n9827), .B(n9826), .Z(n9831) );
  NANDN U11787 ( .A(n9829), .B(n9828), .Z(n9830) );
  AND U11788 ( .A(n9831), .B(n9830), .Z(n9866) );
  NANDN U11789 ( .A(n9833), .B(n9832), .Z(n9837) );
  NANDN U11790 ( .A(n9835), .B(n9834), .Z(n9836) );
  AND U11791 ( .A(n9837), .B(n9836), .Z(n9864) );
  NAND U11792 ( .A(n42143), .B(n9838), .Z(n9840) );
  XNOR U11793 ( .A(a[150]), .B(n4093), .Z(n9875) );
  NAND U11794 ( .A(n42144), .B(n9875), .Z(n9839) );
  AND U11795 ( .A(n9840), .B(n9839), .Z(n9890) );
  XOR U11796 ( .A(a[154]), .B(n42012), .Z(n9878) );
  XNOR U11797 ( .A(n9890), .B(n9889), .Z(n9892) );
  XOR U11798 ( .A(a[152]), .B(n42085), .Z(n9882) );
  AND U11799 ( .A(a[148]), .B(b[7]), .Z(n9883) );
  XNOR U11800 ( .A(n9884), .B(n9883), .Z(n9885) );
  AND U11801 ( .A(a[156]), .B(b[0]), .Z(n9843) );
  XNOR U11802 ( .A(n9843), .B(n4071), .Z(n9845) );
  NANDN U11803 ( .A(b[0]), .B(a[155]), .Z(n9844) );
  NAND U11804 ( .A(n9845), .B(n9844), .Z(n9886) );
  XNOR U11805 ( .A(n9885), .B(n9886), .Z(n9891) );
  XOR U11806 ( .A(n9892), .B(n9891), .Z(n9870) );
  NANDN U11807 ( .A(n9847), .B(n9846), .Z(n9851) );
  NANDN U11808 ( .A(n9849), .B(n9848), .Z(n9850) );
  AND U11809 ( .A(n9851), .B(n9850), .Z(n9869) );
  XNOR U11810 ( .A(n9870), .B(n9869), .Z(n9871) );
  NANDN U11811 ( .A(n9853), .B(n9852), .Z(n9857) );
  NAND U11812 ( .A(n9855), .B(n9854), .Z(n9856) );
  NAND U11813 ( .A(n9857), .B(n9856), .Z(n9872) );
  XNOR U11814 ( .A(n9871), .B(n9872), .Z(n9863) );
  XNOR U11815 ( .A(n9864), .B(n9863), .Z(n9865) );
  XNOR U11816 ( .A(n9866), .B(n9865), .Z(n9895) );
  XNOR U11817 ( .A(sreg[1172]), .B(n9895), .Z(n9897) );
  NANDN U11818 ( .A(sreg[1171]), .B(n9858), .Z(n9862) );
  NAND U11819 ( .A(n9860), .B(n9859), .Z(n9861) );
  NAND U11820 ( .A(n9862), .B(n9861), .Z(n9896) );
  XNOR U11821 ( .A(n9897), .B(n9896), .Z(c[1172]) );
  NANDN U11822 ( .A(n9864), .B(n9863), .Z(n9868) );
  NANDN U11823 ( .A(n9866), .B(n9865), .Z(n9867) );
  AND U11824 ( .A(n9868), .B(n9867), .Z(n9903) );
  NANDN U11825 ( .A(n9870), .B(n9869), .Z(n9874) );
  NANDN U11826 ( .A(n9872), .B(n9871), .Z(n9873) );
  AND U11827 ( .A(n9874), .B(n9873), .Z(n9901) );
  NAND U11828 ( .A(n42143), .B(n9875), .Z(n9877) );
  XNOR U11829 ( .A(a[151]), .B(n4093), .Z(n9912) );
  NAND U11830 ( .A(n42144), .B(n9912), .Z(n9876) );
  AND U11831 ( .A(n9877), .B(n9876), .Z(n9927) );
  XOR U11832 ( .A(a[155]), .B(n42012), .Z(n9915) );
  XNOR U11833 ( .A(n9927), .B(n9926), .Z(n9929) );
  AND U11834 ( .A(a[157]), .B(b[0]), .Z(n9879) );
  XNOR U11835 ( .A(n9879), .B(n4071), .Z(n9881) );
  NANDN U11836 ( .A(b[0]), .B(a[156]), .Z(n9880) );
  NAND U11837 ( .A(n9881), .B(n9880), .Z(n9923) );
  XOR U11838 ( .A(a[153]), .B(n42085), .Z(n9919) );
  AND U11839 ( .A(a[149]), .B(b[7]), .Z(n9920) );
  XNOR U11840 ( .A(n9921), .B(n9920), .Z(n9922) );
  XNOR U11841 ( .A(n9923), .B(n9922), .Z(n9928) );
  XOR U11842 ( .A(n9929), .B(n9928), .Z(n9907) );
  NANDN U11843 ( .A(n9884), .B(n9883), .Z(n9888) );
  NANDN U11844 ( .A(n9886), .B(n9885), .Z(n9887) );
  AND U11845 ( .A(n9888), .B(n9887), .Z(n9906) );
  XNOR U11846 ( .A(n9907), .B(n9906), .Z(n9908) );
  NANDN U11847 ( .A(n9890), .B(n9889), .Z(n9894) );
  NAND U11848 ( .A(n9892), .B(n9891), .Z(n9893) );
  NAND U11849 ( .A(n9894), .B(n9893), .Z(n9909) );
  XNOR U11850 ( .A(n9908), .B(n9909), .Z(n9900) );
  XNOR U11851 ( .A(n9901), .B(n9900), .Z(n9902) );
  XNOR U11852 ( .A(n9903), .B(n9902), .Z(n9932) );
  XNOR U11853 ( .A(sreg[1173]), .B(n9932), .Z(n9934) );
  NANDN U11854 ( .A(sreg[1172]), .B(n9895), .Z(n9899) );
  NAND U11855 ( .A(n9897), .B(n9896), .Z(n9898) );
  NAND U11856 ( .A(n9899), .B(n9898), .Z(n9933) );
  XNOR U11857 ( .A(n9934), .B(n9933), .Z(c[1173]) );
  NANDN U11858 ( .A(n9901), .B(n9900), .Z(n9905) );
  NANDN U11859 ( .A(n9903), .B(n9902), .Z(n9904) );
  AND U11860 ( .A(n9905), .B(n9904), .Z(n9940) );
  NANDN U11861 ( .A(n9907), .B(n9906), .Z(n9911) );
  NANDN U11862 ( .A(n9909), .B(n9908), .Z(n9910) );
  AND U11863 ( .A(n9911), .B(n9910), .Z(n9938) );
  NAND U11864 ( .A(n42143), .B(n9912), .Z(n9914) );
  XNOR U11865 ( .A(a[152]), .B(n4093), .Z(n9949) );
  NAND U11866 ( .A(n42144), .B(n9949), .Z(n9913) );
  AND U11867 ( .A(n9914), .B(n9913), .Z(n9964) );
  XOR U11868 ( .A(a[156]), .B(n42012), .Z(n9952) );
  XNOR U11869 ( .A(n9964), .B(n9963), .Z(n9966) );
  AND U11870 ( .A(a[158]), .B(b[0]), .Z(n9916) );
  XNOR U11871 ( .A(n9916), .B(n4071), .Z(n9918) );
  NANDN U11872 ( .A(b[0]), .B(a[157]), .Z(n9917) );
  NAND U11873 ( .A(n9918), .B(n9917), .Z(n9960) );
  XOR U11874 ( .A(a[154]), .B(n42085), .Z(n9956) );
  AND U11875 ( .A(a[150]), .B(b[7]), .Z(n9957) );
  XNOR U11876 ( .A(n9958), .B(n9957), .Z(n9959) );
  XNOR U11877 ( .A(n9960), .B(n9959), .Z(n9965) );
  XOR U11878 ( .A(n9966), .B(n9965), .Z(n9944) );
  NANDN U11879 ( .A(n9921), .B(n9920), .Z(n9925) );
  NANDN U11880 ( .A(n9923), .B(n9922), .Z(n9924) );
  AND U11881 ( .A(n9925), .B(n9924), .Z(n9943) );
  XNOR U11882 ( .A(n9944), .B(n9943), .Z(n9945) );
  NANDN U11883 ( .A(n9927), .B(n9926), .Z(n9931) );
  NAND U11884 ( .A(n9929), .B(n9928), .Z(n9930) );
  NAND U11885 ( .A(n9931), .B(n9930), .Z(n9946) );
  XNOR U11886 ( .A(n9945), .B(n9946), .Z(n9937) );
  XNOR U11887 ( .A(n9938), .B(n9937), .Z(n9939) );
  XNOR U11888 ( .A(n9940), .B(n9939), .Z(n9969) );
  XNOR U11889 ( .A(sreg[1174]), .B(n9969), .Z(n9971) );
  NANDN U11890 ( .A(sreg[1173]), .B(n9932), .Z(n9936) );
  NAND U11891 ( .A(n9934), .B(n9933), .Z(n9935) );
  NAND U11892 ( .A(n9936), .B(n9935), .Z(n9970) );
  XNOR U11893 ( .A(n9971), .B(n9970), .Z(c[1174]) );
  NANDN U11894 ( .A(n9938), .B(n9937), .Z(n9942) );
  NANDN U11895 ( .A(n9940), .B(n9939), .Z(n9941) );
  AND U11896 ( .A(n9942), .B(n9941), .Z(n9977) );
  NANDN U11897 ( .A(n9944), .B(n9943), .Z(n9948) );
  NANDN U11898 ( .A(n9946), .B(n9945), .Z(n9947) );
  AND U11899 ( .A(n9948), .B(n9947), .Z(n9975) );
  NAND U11900 ( .A(n42143), .B(n9949), .Z(n9951) );
  XNOR U11901 ( .A(a[153]), .B(n4093), .Z(n9986) );
  NAND U11902 ( .A(n42144), .B(n9986), .Z(n9950) );
  AND U11903 ( .A(n9951), .B(n9950), .Z(n10001) );
  XOR U11904 ( .A(a[157]), .B(n42012), .Z(n9989) );
  XNOR U11905 ( .A(n10001), .B(n10000), .Z(n10003) );
  AND U11906 ( .A(a[159]), .B(b[0]), .Z(n9953) );
  XNOR U11907 ( .A(n9953), .B(n4071), .Z(n9955) );
  NANDN U11908 ( .A(b[0]), .B(a[158]), .Z(n9954) );
  NAND U11909 ( .A(n9955), .B(n9954), .Z(n9997) );
  XOR U11910 ( .A(a[155]), .B(n42085), .Z(n9993) );
  AND U11911 ( .A(a[151]), .B(b[7]), .Z(n9994) );
  XNOR U11912 ( .A(n9995), .B(n9994), .Z(n9996) );
  XNOR U11913 ( .A(n9997), .B(n9996), .Z(n10002) );
  XOR U11914 ( .A(n10003), .B(n10002), .Z(n9981) );
  NANDN U11915 ( .A(n9958), .B(n9957), .Z(n9962) );
  NANDN U11916 ( .A(n9960), .B(n9959), .Z(n9961) );
  AND U11917 ( .A(n9962), .B(n9961), .Z(n9980) );
  XNOR U11918 ( .A(n9981), .B(n9980), .Z(n9982) );
  NANDN U11919 ( .A(n9964), .B(n9963), .Z(n9968) );
  NAND U11920 ( .A(n9966), .B(n9965), .Z(n9967) );
  NAND U11921 ( .A(n9968), .B(n9967), .Z(n9983) );
  XNOR U11922 ( .A(n9982), .B(n9983), .Z(n9974) );
  XNOR U11923 ( .A(n9975), .B(n9974), .Z(n9976) );
  XNOR U11924 ( .A(n9977), .B(n9976), .Z(n10006) );
  XNOR U11925 ( .A(sreg[1175]), .B(n10006), .Z(n10008) );
  NANDN U11926 ( .A(sreg[1174]), .B(n9969), .Z(n9973) );
  NAND U11927 ( .A(n9971), .B(n9970), .Z(n9972) );
  NAND U11928 ( .A(n9973), .B(n9972), .Z(n10007) );
  XNOR U11929 ( .A(n10008), .B(n10007), .Z(c[1175]) );
  NANDN U11930 ( .A(n9975), .B(n9974), .Z(n9979) );
  NANDN U11931 ( .A(n9977), .B(n9976), .Z(n9978) );
  AND U11932 ( .A(n9979), .B(n9978), .Z(n10014) );
  NANDN U11933 ( .A(n9981), .B(n9980), .Z(n9985) );
  NANDN U11934 ( .A(n9983), .B(n9982), .Z(n9984) );
  AND U11935 ( .A(n9985), .B(n9984), .Z(n10012) );
  NAND U11936 ( .A(n42143), .B(n9986), .Z(n9988) );
  XNOR U11937 ( .A(a[154]), .B(n4093), .Z(n10023) );
  NAND U11938 ( .A(n42144), .B(n10023), .Z(n9987) );
  AND U11939 ( .A(n9988), .B(n9987), .Z(n10038) );
  XOR U11940 ( .A(a[158]), .B(n42012), .Z(n10026) );
  XNOR U11941 ( .A(n10038), .B(n10037), .Z(n10040) );
  AND U11942 ( .A(a[160]), .B(b[0]), .Z(n9990) );
  XNOR U11943 ( .A(n9990), .B(n4071), .Z(n9992) );
  NANDN U11944 ( .A(b[0]), .B(a[159]), .Z(n9991) );
  NAND U11945 ( .A(n9992), .B(n9991), .Z(n10034) );
  XOR U11946 ( .A(a[156]), .B(n42085), .Z(n10030) );
  AND U11947 ( .A(a[152]), .B(b[7]), .Z(n10031) );
  XNOR U11948 ( .A(n10032), .B(n10031), .Z(n10033) );
  XNOR U11949 ( .A(n10034), .B(n10033), .Z(n10039) );
  XOR U11950 ( .A(n10040), .B(n10039), .Z(n10018) );
  NANDN U11951 ( .A(n9995), .B(n9994), .Z(n9999) );
  NANDN U11952 ( .A(n9997), .B(n9996), .Z(n9998) );
  AND U11953 ( .A(n9999), .B(n9998), .Z(n10017) );
  XNOR U11954 ( .A(n10018), .B(n10017), .Z(n10019) );
  NANDN U11955 ( .A(n10001), .B(n10000), .Z(n10005) );
  NAND U11956 ( .A(n10003), .B(n10002), .Z(n10004) );
  NAND U11957 ( .A(n10005), .B(n10004), .Z(n10020) );
  XNOR U11958 ( .A(n10019), .B(n10020), .Z(n10011) );
  XNOR U11959 ( .A(n10012), .B(n10011), .Z(n10013) );
  XNOR U11960 ( .A(n10014), .B(n10013), .Z(n10043) );
  XNOR U11961 ( .A(sreg[1176]), .B(n10043), .Z(n10045) );
  NANDN U11962 ( .A(sreg[1175]), .B(n10006), .Z(n10010) );
  NAND U11963 ( .A(n10008), .B(n10007), .Z(n10009) );
  NAND U11964 ( .A(n10010), .B(n10009), .Z(n10044) );
  XNOR U11965 ( .A(n10045), .B(n10044), .Z(c[1176]) );
  NANDN U11966 ( .A(n10012), .B(n10011), .Z(n10016) );
  NANDN U11967 ( .A(n10014), .B(n10013), .Z(n10015) );
  AND U11968 ( .A(n10016), .B(n10015), .Z(n10051) );
  NANDN U11969 ( .A(n10018), .B(n10017), .Z(n10022) );
  NANDN U11970 ( .A(n10020), .B(n10019), .Z(n10021) );
  AND U11971 ( .A(n10022), .B(n10021), .Z(n10049) );
  NAND U11972 ( .A(n42143), .B(n10023), .Z(n10025) );
  XNOR U11973 ( .A(a[155]), .B(n4094), .Z(n10060) );
  NAND U11974 ( .A(n42144), .B(n10060), .Z(n10024) );
  AND U11975 ( .A(n10025), .B(n10024), .Z(n10075) );
  XOR U11976 ( .A(a[159]), .B(n42012), .Z(n10063) );
  XNOR U11977 ( .A(n10075), .B(n10074), .Z(n10077) );
  AND U11978 ( .A(a[161]), .B(b[0]), .Z(n10027) );
  XNOR U11979 ( .A(n10027), .B(n4071), .Z(n10029) );
  NANDN U11980 ( .A(b[0]), .B(a[160]), .Z(n10028) );
  NAND U11981 ( .A(n10029), .B(n10028), .Z(n10071) );
  XOR U11982 ( .A(a[157]), .B(n42085), .Z(n10067) );
  AND U11983 ( .A(a[153]), .B(b[7]), .Z(n10068) );
  XNOR U11984 ( .A(n10069), .B(n10068), .Z(n10070) );
  XNOR U11985 ( .A(n10071), .B(n10070), .Z(n10076) );
  XOR U11986 ( .A(n10077), .B(n10076), .Z(n10055) );
  NANDN U11987 ( .A(n10032), .B(n10031), .Z(n10036) );
  NANDN U11988 ( .A(n10034), .B(n10033), .Z(n10035) );
  AND U11989 ( .A(n10036), .B(n10035), .Z(n10054) );
  XNOR U11990 ( .A(n10055), .B(n10054), .Z(n10056) );
  NANDN U11991 ( .A(n10038), .B(n10037), .Z(n10042) );
  NAND U11992 ( .A(n10040), .B(n10039), .Z(n10041) );
  NAND U11993 ( .A(n10042), .B(n10041), .Z(n10057) );
  XNOR U11994 ( .A(n10056), .B(n10057), .Z(n10048) );
  XNOR U11995 ( .A(n10049), .B(n10048), .Z(n10050) );
  XNOR U11996 ( .A(n10051), .B(n10050), .Z(n10080) );
  XNOR U11997 ( .A(sreg[1177]), .B(n10080), .Z(n10082) );
  NANDN U11998 ( .A(sreg[1176]), .B(n10043), .Z(n10047) );
  NAND U11999 ( .A(n10045), .B(n10044), .Z(n10046) );
  NAND U12000 ( .A(n10047), .B(n10046), .Z(n10081) );
  XNOR U12001 ( .A(n10082), .B(n10081), .Z(c[1177]) );
  NANDN U12002 ( .A(n10049), .B(n10048), .Z(n10053) );
  NANDN U12003 ( .A(n10051), .B(n10050), .Z(n10052) );
  AND U12004 ( .A(n10053), .B(n10052), .Z(n10088) );
  NANDN U12005 ( .A(n10055), .B(n10054), .Z(n10059) );
  NANDN U12006 ( .A(n10057), .B(n10056), .Z(n10058) );
  AND U12007 ( .A(n10059), .B(n10058), .Z(n10086) );
  NAND U12008 ( .A(n42143), .B(n10060), .Z(n10062) );
  XNOR U12009 ( .A(a[156]), .B(n4094), .Z(n10097) );
  NAND U12010 ( .A(n42144), .B(n10097), .Z(n10061) );
  AND U12011 ( .A(n10062), .B(n10061), .Z(n10112) );
  XOR U12012 ( .A(a[160]), .B(n42012), .Z(n10100) );
  XNOR U12013 ( .A(n10112), .B(n10111), .Z(n10114) );
  AND U12014 ( .A(a[162]), .B(b[0]), .Z(n10064) );
  XNOR U12015 ( .A(n10064), .B(n4071), .Z(n10066) );
  NANDN U12016 ( .A(b[0]), .B(a[161]), .Z(n10065) );
  NAND U12017 ( .A(n10066), .B(n10065), .Z(n10108) );
  XOR U12018 ( .A(a[158]), .B(n42085), .Z(n10104) );
  AND U12019 ( .A(a[154]), .B(b[7]), .Z(n10105) );
  XNOR U12020 ( .A(n10106), .B(n10105), .Z(n10107) );
  XNOR U12021 ( .A(n10108), .B(n10107), .Z(n10113) );
  XOR U12022 ( .A(n10114), .B(n10113), .Z(n10092) );
  NANDN U12023 ( .A(n10069), .B(n10068), .Z(n10073) );
  NANDN U12024 ( .A(n10071), .B(n10070), .Z(n10072) );
  AND U12025 ( .A(n10073), .B(n10072), .Z(n10091) );
  XNOR U12026 ( .A(n10092), .B(n10091), .Z(n10093) );
  NANDN U12027 ( .A(n10075), .B(n10074), .Z(n10079) );
  NAND U12028 ( .A(n10077), .B(n10076), .Z(n10078) );
  NAND U12029 ( .A(n10079), .B(n10078), .Z(n10094) );
  XNOR U12030 ( .A(n10093), .B(n10094), .Z(n10085) );
  XNOR U12031 ( .A(n10086), .B(n10085), .Z(n10087) );
  XNOR U12032 ( .A(n10088), .B(n10087), .Z(n10117) );
  XNOR U12033 ( .A(sreg[1178]), .B(n10117), .Z(n10119) );
  NANDN U12034 ( .A(sreg[1177]), .B(n10080), .Z(n10084) );
  NAND U12035 ( .A(n10082), .B(n10081), .Z(n10083) );
  NAND U12036 ( .A(n10084), .B(n10083), .Z(n10118) );
  XNOR U12037 ( .A(n10119), .B(n10118), .Z(c[1178]) );
  NANDN U12038 ( .A(n10086), .B(n10085), .Z(n10090) );
  NANDN U12039 ( .A(n10088), .B(n10087), .Z(n10089) );
  AND U12040 ( .A(n10090), .B(n10089), .Z(n10125) );
  NANDN U12041 ( .A(n10092), .B(n10091), .Z(n10096) );
  NANDN U12042 ( .A(n10094), .B(n10093), .Z(n10095) );
  AND U12043 ( .A(n10096), .B(n10095), .Z(n10123) );
  NAND U12044 ( .A(n42143), .B(n10097), .Z(n10099) );
  XNOR U12045 ( .A(a[157]), .B(n4094), .Z(n10134) );
  NAND U12046 ( .A(n42144), .B(n10134), .Z(n10098) );
  AND U12047 ( .A(n10099), .B(n10098), .Z(n10149) );
  XOR U12048 ( .A(a[161]), .B(n42012), .Z(n10137) );
  XNOR U12049 ( .A(n10149), .B(n10148), .Z(n10151) );
  AND U12050 ( .A(a[163]), .B(b[0]), .Z(n10101) );
  XNOR U12051 ( .A(n10101), .B(n4071), .Z(n10103) );
  NANDN U12052 ( .A(b[0]), .B(a[162]), .Z(n10102) );
  NAND U12053 ( .A(n10103), .B(n10102), .Z(n10145) );
  XOR U12054 ( .A(a[159]), .B(n42085), .Z(n10138) );
  AND U12055 ( .A(a[155]), .B(b[7]), .Z(n10142) );
  XNOR U12056 ( .A(n10143), .B(n10142), .Z(n10144) );
  XNOR U12057 ( .A(n10145), .B(n10144), .Z(n10150) );
  XOR U12058 ( .A(n10151), .B(n10150), .Z(n10129) );
  NANDN U12059 ( .A(n10106), .B(n10105), .Z(n10110) );
  NANDN U12060 ( .A(n10108), .B(n10107), .Z(n10109) );
  AND U12061 ( .A(n10110), .B(n10109), .Z(n10128) );
  XNOR U12062 ( .A(n10129), .B(n10128), .Z(n10130) );
  NANDN U12063 ( .A(n10112), .B(n10111), .Z(n10116) );
  NAND U12064 ( .A(n10114), .B(n10113), .Z(n10115) );
  NAND U12065 ( .A(n10116), .B(n10115), .Z(n10131) );
  XNOR U12066 ( .A(n10130), .B(n10131), .Z(n10122) );
  XNOR U12067 ( .A(n10123), .B(n10122), .Z(n10124) );
  XNOR U12068 ( .A(n10125), .B(n10124), .Z(n10154) );
  XNOR U12069 ( .A(sreg[1179]), .B(n10154), .Z(n10156) );
  NANDN U12070 ( .A(sreg[1178]), .B(n10117), .Z(n10121) );
  NAND U12071 ( .A(n10119), .B(n10118), .Z(n10120) );
  NAND U12072 ( .A(n10121), .B(n10120), .Z(n10155) );
  XNOR U12073 ( .A(n10156), .B(n10155), .Z(c[1179]) );
  NANDN U12074 ( .A(n10123), .B(n10122), .Z(n10127) );
  NANDN U12075 ( .A(n10125), .B(n10124), .Z(n10126) );
  AND U12076 ( .A(n10127), .B(n10126), .Z(n10162) );
  NANDN U12077 ( .A(n10129), .B(n10128), .Z(n10133) );
  NANDN U12078 ( .A(n10131), .B(n10130), .Z(n10132) );
  AND U12079 ( .A(n10133), .B(n10132), .Z(n10160) );
  NAND U12080 ( .A(n42143), .B(n10134), .Z(n10136) );
  XNOR U12081 ( .A(a[158]), .B(n4094), .Z(n10171) );
  NAND U12082 ( .A(n42144), .B(n10171), .Z(n10135) );
  AND U12083 ( .A(n10136), .B(n10135), .Z(n10186) );
  XOR U12084 ( .A(a[162]), .B(n42012), .Z(n10174) );
  XNOR U12085 ( .A(n10186), .B(n10185), .Z(n10188) );
  XOR U12086 ( .A(a[160]), .B(n42085), .Z(n10175) );
  AND U12087 ( .A(a[156]), .B(b[7]), .Z(n10179) );
  XNOR U12088 ( .A(n10180), .B(n10179), .Z(n10181) );
  AND U12089 ( .A(a[164]), .B(b[0]), .Z(n10139) );
  XNOR U12090 ( .A(n10139), .B(n4071), .Z(n10141) );
  NANDN U12091 ( .A(b[0]), .B(a[163]), .Z(n10140) );
  NAND U12092 ( .A(n10141), .B(n10140), .Z(n10182) );
  XNOR U12093 ( .A(n10181), .B(n10182), .Z(n10187) );
  XOR U12094 ( .A(n10188), .B(n10187), .Z(n10166) );
  NANDN U12095 ( .A(n10143), .B(n10142), .Z(n10147) );
  NANDN U12096 ( .A(n10145), .B(n10144), .Z(n10146) );
  AND U12097 ( .A(n10147), .B(n10146), .Z(n10165) );
  XNOR U12098 ( .A(n10166), .B(n10165), .Z(n10167) );
  NANDN U12099 ( .A(n10149), .B(n10148), .Z(n10153) );
  NAND U12100 ( .A(n10151), .B(n10150), .Z(n10152) );
  NAND U12101 ( .A(n10153), .B(n10152), .Z(n10168) );
  XNOR U12102 ( .A(n10167), .B(n10168), .Z(n10159) );
  XNOR U12103 ( .A(n10160), .B(n10159), .Z(n10161) );
  XNOR U12104 ( .A(n10162), .B(n10161), .Z(n10191) );
  XNOR U12105 ( .A(sreg[1180]), .B(n10191), .Z(n10193) );
  NANDN U12106 ( .A(sreg[1179]), .B(n10154), .Z(n10158) );
  NAND U12107 ( .A(n10156), .B(n10155), .Z(n10157) );
  NAND U12108 ( .A(n10158), .B(n10157), .Z(n10192) );
  XNOR U12109 ( .A(n10193), .B(n10192), .Z(c[1180]) );
  NANDN U12110 ( .A(n10160), .B(n10159), .Z(n10164) );
  NANDN U12111 ( .A(n10162), .B(n10161), .Z(n10163) );
  AND U12112 ( .A(n10164), .B(n10163), .Z(n10199) );
  NANDN U12113 ( .A(n10166), .B(n10165), .Z(n10170) );
  NANDN U12114 ( .A(n10168), .B(n10167), .Z(n10169) );
  AND U12115 ( .A(n10170), .B(n10169), .Z(n10197) );
  NAND U12116 ( .A(n42143), .B(n10171), .Z(n10173) );
  XNOR U12117 ( .A(a[159]), .B(n4094), .Z(n10208) );
  NAND U12118 ( .A(n42144), .B(n10208), .Z(n10172) );
  AND U12119 ( .A(n10173), .B(n10172), .Z(n10223) );
  XOR U12120 ( .A(a[163]), .B(n42012), .Z(n10211) );
  XNOR U12121 ( .A(n10223), .B(n10222), .Z(n10225) );
  XOR U12122 ( .A(a[161]), .B(n42085), .Z(n10215) );
  AND U12123 ( .A(a[157]), .B(b[7]), .Z(n10216) );
  XNOR U12124 ( .A(n10217), .B(n10216), .Z(n10218) );
  AND U12125 ( .A(a[165]), .B(b[0]), .Z(n10176) );
  XNOR U12126 ( .A(n10176), .B(n4071), .Z(n10178) );
  NANDN U12127 ( .A(b[0]), .B(a[164]), .Z(n10177) );
  NAND U12128 ( .A(n10178), .B(n10177), .Z(n10219) );
  XNOR U12129 ( .A(n10218), .B(n10219), .Z(n10224) );
  XOR U12130 ( .A(n10225), .B(n10224), .Z(n10203) );
  NANDN U12131 ( .A(n10180), .B(n10179), .Z(n10184) );
  NANDN U12132 ( .A(n10182), .B(n10181), .Z(n10183) );
  AND U12133 ( .A(n10184), .B(n10183), .Z(n10202) );
  XNOR U12134 ( .A(n10203), .B(n10202), .Z(n10204) );
  NANDN U12135 ( .A(n10186), .B(n10185), .Z(n10190) );
  NAND U12136 ( .A(n10188), .B(n10187), .Z(n10189) );
  NAND U12137 ( .A(n10190), .B(n10189), .Z(n10205) );
  XNOR U12138 ( .A(n10204), .B(n10205), .Z(n10196) );
  XNOR U12139 ( .A(n10197), .B(n10196), .Z(n10198) );
  XNOR U12140 ( .A(n10199), .B(n10198), .Z(n10228) );
  XNOR U12141 ( .A(sreg[1181]), .B(n10228), .Z(n10230) );
  NANDN U12142 ( .A(sreg[1180]), .B(n10191), .Z(n10195) );
  NAND U12143 ( .A(n10193), .B(n10192), .Z(n10194) );
  NAND U12144 ( .A(n10195), .B(n10194), .Z(n10229) );
  XNOR U12145 ( .A(n10230), .B(n10229), .Z(c[1181]) );
  NANDN U12146 ( .A(n10197), .B(n10196), .Z(n10201) );
  NANDN U12147 ( .A(n10199), .B(n10198), .Z(n10200) );
  AND U12148 ( .A(n10201), .B(n10200), .Z(n10236) );
  NANDN U12149 ( .A(n10203), .B(n10202), .Z(n10207) );
  NANDN U12150 ( .A(n10205), .B(n10204), .Z(n10206) );
  AND U12151 ( .A(n10207), .B(n10206), .Z(n10234) );
  NAND U12152 ( .A(n42143), .B(n10208), .Z(n10210) );
  XNOR U12153 ( .A(a[160]), .B(n4094), .Z(n10245) );
  NAND U12154 ( .A(n42144), .B(n10245), .Z(n10209) );
  AND U12155 ( .A(n10210), .B(n10209), .Z(n10260) );
  XOR U12156 ( .A(a[164]), .B(n42012), .Z(n10248) );
  XNOR U12157 ( .A(n10260), .B(n10259), .Z(n10262) );
  AND U12158 ( .A(a[166]), .B(b[0]), .Z(n10212) );
  XNOR U12159 ( .A(n10212), .B(n4071), .Z(n10214) );
  NANDN U12160 ( .A(b[0]), .B(a[165]), .Z(n10213) );
  NAND U12161 ( .A(n10214), .B(n10213), .Z(n10256) );
  XOR U12162 ( .A(a[162]), .B(n42085), .Z(n10252) );
  AND U12163 ( .A(a[158]), .B(b[7]), .Z(n10253) );
  XNOR U12164 ( .A(n10254), .B(n10253), .Z(n10255) );
  XNOR U12165 ( .A(n10256), .B(n10255), .Z(n10261) );
  XOR U12166 ( .A(n10262), .B(n10261), .Z(n10240) );
  NANDN U12167 ( .A(n10217), .B(n10216), .Z(n10221) );
  NANDN U12168 ( .A(n10219), .B(n10218), .Z(n10220) );
  AND U12169 ( .A(n10221), .B(n10220), .Z(n10239) );
  XNOR U12170 ( .A(n10240), .B(n10239), .Z(n10241) );
  NANDN U12171 ( .A(n10223), .B(n10222), .Z(n10227) );
  NAND U12172 ( .A(n10225), .B(n10224), .Z(n10226) );
  NAND U12173 ( .A(n10227), .B(n10226), .Z(n10242) );
  XNOR U12174 ( .A(n10241), .B(n10242), .Z(n10233) );
  XNOR U12175 ( .A(n10234), .B(n10233), .Z(n10235) );
  XNOR U12176 ( .A(n10236), .B(n10235), .Z(n10265) );
  XNOR U12177 ( .A(sreg[1182]), .B(n10265), .Z(n10267) );
  NANDN U12178 ( .A(sreg[1181]), .B(n10228), .Z(n10232) );
  NAND U12179 ( .A(n10230), .B(n10229), .Z(n10231) );
  NAND U12180 ( .A(n10232), .B(n10231), .Z(n10266) );
  XNOR U12181 ( .A(n10267), .B(n10266), .Z(c[1182]) );
  NANDN U12182 ( .A(n10234), .B(n10233), .Z(n10238) );
  NANDN U12183 ( .A(n10236), .B(n10235), .Z(n10237) );
  AND U12184 ( .A(n10238), .B(n10237), .Z(n10273) );
  NANDN U12185 ( .A(n10240), .B(n10239), .Z(n10244) );
  NANDN U12186 ( .A(n10242), .B(n10241), .Z(n10243) );
  AND U12187 ( .A(n10244), .B(n10243), .Z(n10271) );
  NAND U12188 ( .A(n42143), .B(n10245), .Z(n10247) );
  XNOR U12189 ( .A(a[161]), .B(n4094), .Z(n10282) );
  NAND U12190 ( .A(n42144), .B(n10282), .Z(n10246) );
  AND U12191 ( .A(n10247), .B(n10246), .Z(n10297) );
  XOR U12192 ( .A(a[165]), .B(n42012), .Z(n10285) );
  XNOR U12193 ( .A(n10297), .B(n10296), .Z(n10299) );
  AND U12194 ( .A(a[167]), .B(b[0]), .Z(n10249) );
  XNOR U12195 ( .A(n10249), .B(n4071), .Z(n10251) );
  NANDN U12196 ( .A(b[0]), .B(a[166]), .Z(n10250) );
  NAND U12197 ( .A(n10251), .B(n10250), .Z(n10293) );
  XOR U12198 ( .A(a[163]), .B(n42085), .Z(n10289) );
  AND U12199 ( .A(a[159]), .B(b[7]), .Z(n10290) );
  XNOR U12200 ( .A(n10291), .B(n10290), .Z(n10292) );
  XNOR U12201 ( .A(n10293), .B(n10292), .Z(n10298) );
  XOR U12202 ( .A(n10299), .B(n10298), .Z(n10277) );
  NANDN U12203 ( .A(n10254), .B(n10253), .Z(n10258) );
  NANDN U12204 ( .A(n10256), .B(n10255), .Z(n10257) );
  AND U12205 ( .A(n10258), .B(n10257), .Z(n10276) );
  XNOR U12206 ( .A(n10277), .B(n10276), .Z(n10278) );
  NANDN U12207 ( .A(n10260), .B(n10259), .Z(n10264) );
  NAND U12208 ( .A(n10262), .B(n10261), .Z(n10263) );
  NAND U12209 ( .A(n10264), .B(n10263), .Z(n10279) );
  XNOR U12210 ( .A(n10278), .B(n10279), .Z(n10270) );
  XNOR U12211 ( .A(n10271), .B(n10270), .Z(n10272) );
  XNOR U12212 ( .A(n10273), .B(n10272), .Z(n10302) );
  XNOR U12213 ( .A(sreg[1183]), .B(n10302), .Z(n10304) );
  NANDN U12214 ( .A(sreg[1182]), .B(n10265), .Z(n10269) );
  NAND U12215 ( .A(n10267), .B(n10266), .Z(n10268) );
  NAND U12216 ( .A(n10269), .B(n10268), .Z(n10303) );
  XNOR U12217 ( .A(n10304), .B(n10303), .Z(c[1183]) );
  NANDN U12218 ( .A(n10271), .B(n10270), .Z(n10275) );
  NANDN U12219 ( .A(n10273), .B(n10272), .Z(n10274) );
  AND U12220 ( .A(n10275), .B(n10274), .Z(n10310) );
  NANDN U12221 ( .A(n10277), .B(n10276), .Z(n10281) );
  NANDN U12222 ( .A(n10279), .B(n10278), .Z(n10280) );
  AND U12223 ( .A(n10281), .B(n10280), .Z(n10308) );
  NAND U12224 ( .A(n42143), .B(n10282), .Z(n10284) );
  XNOR U12225 ( .A(a[162]), .B(n4095), .Z(n10319) );
  NAND U12226 ( .A(n42144), .B(n10319), .Z(n10283) );
  AND U12227 ( .A(n10284), .B(n10283), .Z(n10334) );
  XOR U12228 ( .A(a[166]), .B(n42012), .Z(n10322) );
  XNOR U12229 ( .A(n10334), .B(n10333), .Z(n10336) );
  AND U12230 ( .A(a[168]), .B(b[0]), .Z(n10286) );
  XNOR U12231 ( .A(n10286), .B(n4071), .Z(n10288) );
  NANDN U12232 ( .A(b[0]), .B(a[167]), .Z(n10287) );
  NAND U12233 ( .A(n10288), .B(n10287), .Z(n10330) );
  XOR U12234 ( .A(a[164]), .B(n42085), .Z(n10326) );
  AND U12235 ( .A(a[160]), .B(b[7]), .Z(n10327) );
  XNOR U12236 ( .A(n10328), .B(n10327), .Z(n10329) );
  XNOR U12237 ( .A(n10330), .B(n10329), .Z(n10335) );
  XOR U12238 ( .A(n10336), .B(n10335), .Z(n10314) );
  NANDN U12239 ( .A(n10291), .B(n10290), .Z(n10295) );
  NANDN U12240 ( .A(n10293), .B(n10292), .Z(n10294) );
  AND U12241 ( .A(n10295), .B(n10294), .Z(n10313) );
  XNOR U12242 ( .A(n10314), .B(n10313), .Z(n10315) );
  NANDN U12243 ( .A(n10297), .B(n10296), .Z(n10301) );
  NAND U12244 ( .A(n10299), .B(n10298), .Z(n10300) );
  NAND U12245 ( .A(n10301), .B(n10300), .Z(n10316) );
  XNOR U12246 ( .A(n10315), .B(n10316), .Z(n10307) );
  XNOR U12247 ( .A(n10308), .B(n10307), .Z(n10309) );
  XNOR U12248 ( .A(n10310), .B(n10309), .Z(n10339) );
  XNOR U12249 ( .A(sreg[1184]), .B(n10339), .Z(n10341) );
  NANDN U12250 ( .A(sreg[1183]), .B(n10302), .Z(n10306) );
  NAND U12251 ( .A(n10304), .B(n10303), .Z(n10305) );
  NAND U12252 ( .A(n10306), .B(n10305), .Z(n10340) );
  XNOR U12253 ( .A(n10341), .B(n10340), .Z(c[1184]) );
  NANDN U12254 ( .A(n10308), .B(n10307), .Z(n10312) );
  NANDN U12255 ( .A(n10310), .B(n10309), .Z(n10311) );
  AND U12256 ( .A(n10312), .B(n10311), .Z(n10347) );
  NANDN U12257 ( .A(n10314), .B(n10313), .Z(n10318) );
  NANDN U12258 ( .A(n10316), .B(n10315), .Z(n10317) );
  AND U12259 ( .A(n10318), .B(n10317), .Z(n10345) );
  NAND U12260 ( .A(n42143), .B(n10319), .Z(n10321) );
  XNOR U12261 ( .A(a[163]), .B(n4095), .Z(n10356) );
  NAND U12262 ( .A(n42144), .B(n10356), .Z(n10320) );
  AND U12263 ( .A(n10321), .B(n10320), .Z(n10371) );
  XOR U12264 ( .A(a[167]), .B(n42012), .Z(n10359) );
  XNOR U12265 ( .A(n10371), .B(n10370), .Z(n10373) );
  AND U12266 ( .A(a[169]), .B(b[0]), .Z(n10323) );
  XNOR U12267 ( .A(n10323), .B(n4071), .Z(n10325) );
  NANDN U12268 ( .A(b[0]), .B(a[168]), .Z(n10324) );
  NAND U12269 ( .A(n10325), .B(n10324), .Z(n10367) );
  XOR U12270 ( .A(a[165]), .B(n42085), .Z(n10363) );
  AND U12271 ( .A(a[161]), .B(b[7]), .Z(n10364) );
  XNOR U12272 ( .A(n10365), .B(n10364), .Z(n10366) );
  XNOR U12273 ( .A(n10367), .B(n10366), .Z(n10372) );
  XOR U12274 ( .A(n10373), .B(n10372), .Z(n10351) );
  NANDN U12275 ( .A(n10328), .B(n10327), .Z(n10332) );
  NANDN U12276 ( .A(n10330), .B(n10329), .Z(n10331) );
  AND U12277 ( .A(n10332), .B(n10331), .Z(n10350) );
  XNOR U12278 ( .A(n10351), .B(n10350), .Z(n10352) );
  NANDN U12279 ( .A(n10334), .B(n10333), .Z(n10338) );
  NAND U12280 ( .A(n10336), .B(n10335), .Z(n10337) );
  NAND U12281 ( .A(n10338), .B(n10337), .Z(n10353) );
  XNOR U12282 ( .A(n10352), .B(n10353), .Z(n10344) );
  XNOR U12283 ( .A(n10345), .B(n10344), .Z(n10346) );
  XNOR U12284 ( .A(n10347), .B(n10346), .Z(n10376) );
  XNOR U12285 ( .A(sreg[1185]), .B(n10376), .Z(n10378) );
  NANDN U12286 ( .A(sreg[1184]), .B(n10339), .Z(n10343) );
  NAND U12287 ( .A(n10341), .B(n10340), .Z(n10342) );
  NAND U12288 ( .A(n10343), .B(n10342), .Z(n10377) );
  XNOR U12289 ( .A(n10378), .B(n10377), .Z(c[1185]) );
  NANDN U12290 ( .A(n10345), .B(n10344), .Z(n10349) );
  NANDN U12291 ( .A(n10347), .B(n10346), .Z(n10348) );
  AND U12292 ( .A(n10349), .B(n10348), .Z(n10384) );
  NANDN U12293 ( .A(n10351), .B(n10350), .Z(n10355) );
  NANDN U12294 ( .A(n10353), .B(n10352), .Z(n10354) );
  AND U12295 ( .A(n10355), .B(n10354), .Z(n10382) );
  NAND U12296 ( .A(n42143), .B(n10356), .Z(n10358) );
  XNOR U12297 ( .A(a[164]), .B(n4095), .Z(n10393) );
  NAND U12298 ( .A(n42144), .B(n10393), .Z(n10357) );
  AND U12299 ( .A(n10358), .B(n10357), .Z(n10408) );
  XOR U12300 ( .A(a[168]), .B(n42012), .Z(n10396) );
  XNOR U12301 ( .A(n10408), .B(n10407), .Z(n10410) );
  AND U12302 ( .A(a[170]), .B(b[0]), .Z(n10360) );
  XNOR U12303 ( .A(n10360), .B(n4071), .Z(n10362) );
  NANDN U12304 ( .A(b[0]), .B(a[169]), .Z(n10361) );
  NAND U12305 ( .A(n10362), .B(n10361), .Z(n10404) );
  XOR U12306 ( .A(a[166]), .B(n42085), .Z(n10400) );
  AND U12307 ( .A(a[162]), .B(b[7]), .Z(n10401) );
  XNOR U12308 ( .A(n10402), .B(n10401), .Z(n10403) );
  XNOR U12309 ( .A(n10404), .B(n10403), .Z(n10409) );
  XOR U12310 ( .A(n10410), .B(n10409), .Z(n10388) );
  NANDN U12311 ( .A(n10365), .B(n10364), .Z(n10369) );
  NANDN U12312 ( .A(n10367), .B(n10366), .Z(n10368) );
  AND U12313 ( .A(n10369), .B(n10368), .Z(n10387) );
  XNOR U12314 ( .A(n10388), .B(n10387), .Z(n10389) );
  NANDN U12315 ( .A(n10371), .B(n10370), .Z(n10375) );
  NAND U12316 ( .A(n10373), .B(n10372), .Z(n10374) );
  NAND U12317 ( .A(n10375), .B(n10374), .Z(n10390) );
  XNOR U12318 ( .A(n10389), .B(n10390), .Z(n10381) );
  XNOR U12319 ( .A(n10382), .B(n10381), .Z(n10383) );
  XNOR U12320 ( .A(n10384), .B(n10383), .Z(n10413) );
  XNOR U12321 ( .A(sreg[1186]), .B(n10413), .Z(n10415) );
  NANDN U12322 ( .A(sreg[1185]), .B(n10376), .Z(n10380) );
  NAND U12323 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND U12324 ( .A(n10380), .B(n10379), .Z(n10414) );
  XNOR U12325 ( .A(n10415), .B(n10414), .Z(c[1186]) );
  NANDN U12326 ( .A(n10382), .B(n10381), .Z(n10386) );
  NANDN U12327 ( .A(n10384), .B(n10383), .Z(n10385) );
  AND U12328 ( .A(n10386), .B(n10385), .Z(n10421) );
  NANDN U12329 ( .A(n10388), .B(n10387), .Z(n10392) );
  NANDN U12330 ( .A(n10390), .B(n10389), .Z(n10391) );
  AND U12331 ( .A(n10392), .B(n10391), .Z(n10419) );
  NAND U12332 ( .A(n42143), .B(n10393), .Z(n10395) );
  XNOR U12333 ( .A(a[165]), .B(n4095), .Z(n10430) );
  NAND U12334 ( .A(n42144), .B(n10430), .Z(n10394) );
  AND U12335 ( .A(n10395), .B(n10394), .Z(n10445) );
  XOR U12336 ( .A(a[169]), .B(n42012), .Z(n10433) );
  XNOR U12337 ( .A(n10445), .B(n10444), .Z(n10447) );
  AND U12338 ( .A(a[171]), .B(b[0]), .Z(n10397) );
  XNOR U12339 ( .A(n10397), .B(n4071), .Z(n10399) );
  NANDN U12340 ( .A(b[0]), .B(a[170]), .Z(n10398) );
  NAND U12341 ( .A(n10399), .B(n10398), .Z(n10441) );
  XOR U12342 ( .A(a[167]), .B(n42085), .Z(n10437) );
  AND U12343 ( .A(a[163]), .B(b[7]), .Z(n10438) );
  XNOR U12344 ( .A(n10439), .B(n10438), .Z(n10440) );
  XNOR U12345 ( .A(n10441), .B(n10440), .Z(n10446) );
  XOR U12346 ( .A(n10447), .B(n10446), .Z(n10425) );
  NANDN U12347 ( .A(n10402), .B(n10401), .Z(n10406) );
  NANDN U12348 ( .A(n10404), .B(n10403), .Z(n10405) );
  AND U12349 ( .A(n10406), .B(n10405), .Z(n10424) );
  XNOR U12350 ( .A(n10425), .B(n10424), .Z(n10426) );
  NANDN U12351 ( .A(n10408), .B(n10407), .Z(n10412) );
  NAND U12352 ( .A(n10410), .B(n10409), .Z(n10411) );
  NAND U12353 ( .A(n10412), .B(n10411), .Z(n10427) );
  XNOR U12354 ( .A(n10426), .B(n10427), .Z(n10418) );
  XNOR U12355 ( .A(n10419), .B(n10418), .Z(n10420) );
  XNOR U12356 ( .A(n10421), .B(n10420), .Z(n10450) );
  XNOR U12357 ( .A(sreg[1187]), .B(n10450), .Z(n10452) );
  NANDN U12358 ( .A(sreg[1186]), .B(n10413), .Z(n10417) );
  NAND U12359 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U12360 ( .A(n10417), .B(n10416), .Z(n10451) );
  XNOR U12361 ( .A(n10452), .B(n10451), .Z(c[1187]) );
  NANDN U12362 ( .A(n10419), .B(n10418), .Z(n10423) );
  NANDN U12363 ( .A(n10421), .B(n10420), .Z(n10422) );
  AND U12364 ( .A(n10423), .B(n10422), .Z(n10458) );
  NANDN U12365 ( .A(n10425), .B(n10424), .Z(n10429) );
  NANDN U12366 ( .A(n10427), .B(n10426), .Z(n10428) );
  AND U12367 ( .A(n10429), .B(n10428), .Z(n10456) );
  NAND U12368 ( .A(n42143), .B(n10430), .Z(n10432) );
  XNOR U12369 ( .A(a[166]), .B(n4095), .Z(n10467) );
  NAND U12370 ( .A(n42144), .B(n10467), .Z(n10431) );
  AND U12371 ( .A(n10432), .B(n10431), .Z(n10482) );
  XOR U12372 ( .A(a[170]), .B(n42012), .Z(n10470) );
  XNOR U12373 ( .A(n10482), .B(n10481), .Z(n10484) );
  AND U12374 ( .A(a[172]), .B(b[0]), .Z(n10434) );
  XNOR U12375 ( .A(n10434), .B(n4071), .Z(n10436) );
  NANDN U12376 ( .A(b[0]), .B(a[171]), .Z(n10435) );
  NAND U12377 ( .A(n10436), .B(n10435), .Z(n10478) );
  XOR U12378 ( .A(a[168]), .B(n42085), .Z(n10474) );
  AND U12379 ( .A(a[164]), .B(b[7]), .Z(n10475) );
  XNOR U12380 ( .A(n10476), .B(n10475), .Z(n10477) );
  XNOR U12381 ( .A(n10478), .B(n10477), .Z(n10483) );
  XOR U12382 ( .A(n10484), .B(n10483), .Z(n10462) );
  NANDN U12383 ( .A(n10439), .B(n10438), .Z(n10443) );
  NANDN U12384 ( .A(n10441), .B(n10440), .Z(n10442) );
  AND U12385 ( .A(n10443), .B(n10442), .Z(n10461) );
  XNOR U12386 ( .A(n10462), .B(n10461), .Z(n10463) );
  NANDN U12387 ( .A(n10445), .B(n10444), .Z(n10449) );
  NAND U12388 ( .A(n10447), .B(n10446), .Z(n10448) );
  NAND U12389 ( .A(n10449), .B(n10448), .Z(n10464) );
  XNOR U12390 ( .A(n10463), .B(n10464), .Z(n10455) );
  XNOR U12391 ( .A(n10456), .B(n10455), .Z(n10457) );
  XNOR U12392 ( .A(n10458), .B(n10457), .Z(n10487) );
  XNOR U12393 ( .A(sreg[1188]), .B(n10487), .Z(n10489) );
  NANDN U12394 ( .A(sreg[1187]), .B(n10450), .Z(n10454) );
  NAND U12395 ( .A(n10452), .B(n10451), .Z(n10453) );
  NAND U12396 ( .A(n10454), .B(n10453), .Z(n10488) );
  XNOR U12397 ( .A(n10489), .B(n10488), .Z(c[1188]) );
  NANDN U12398 ( .A(n10456), .B(n10455), .Z(n10460) );
  NANDN U12399 ( .A(n10458), .B(n10457), .Z(n10459) );
  AND U12400 ( .A(n10460), .B(n10459), .Z(n10495) );
  NANDN U12401 ( .A(n10462), .B(n10461), .Z(n10466) );
  NANDN U12402 ( .A(n10464), .B(n10463), .Z(n10465) );
  AND U12403 ( .A(n10466), .B(n10465), .Z(n10493) );
  NAND U12404 ( .A(n42143), .B(n10467), .Z(n10469) );
  XNOR U12405 ( .A(a[167]), .B(n4095), .Z(n10504) );
  NAND U12406 ( .A(n42144), .B(n10504), .Z(n10468) );
  AND U12407 ( .A(n10469), .B(n10468), .Z(n10519) );
  XOR U12408 ( .A(a[171]), .B(n42012), .Z(n10507) );
  XNOR U12409 ( .A(n10519), .B(n10518), .Z(n10521) );
  AND U12410 ( .A(a[173]), .B(b[0]), .Z(n10471) );
  XNOR U12411 ( .A(n10471), .B(n4071), .Z(n10473) );
  NANDN U12412 ( .A(b[0]), .B(a[172]), .Z(n10472) );
  NAND U12413 ( .A(n10473), .B(n10472), .Z(n10515) );
  XOR U12414 ( .A(a[169]), .B(n42085), .Z(n10511) );
  AND U12415 ( .A(a[165]), .B(b[7]), .Z(n10512) );
  XNOR U12416 ( .A(n10513), .B(n10512), .Z(n10514) );
  XNOR U12417 ( .A(n10515), .B(n10514), .Z(n10520) );
  XOR U12418 ( .A(n10521), .B(n10520), .Z(n10499) );
  NANDN U12419 ( .A(n10476), .B(n10475), .Z(n10480) );
  NANDN U12420 ( .A(n10478), .B(n10477), .Z(n10479) );
  AND U12421 ( .A(n10480), .B(n10479), .Z(n10498) );
  XNOR U12422 ( .A(n10499), .B(n10498), .Z(n10500) );
  NANDN U12423 ( .A(n10482), .B(n10481), .Z(n10486) );
  NAND U12424 ( .A(n10484), .B(n10483), .Z(n10485) );
  NAND U12425 ( .A(n10486), .B(n10485), .Z(n10501) );
  XNOR U12426 ( .A(n10500), .B(n10501), .Z(n10492) );
  XNOR U12427 ( .A(n10493), .B(n10492), .Z(n10494) );
  XNOR U12428 ( .A(n10495), .B(n10494), .Z(n10524) );
  XNOR U12429 ( .A(sreg[1189]), .B(n10524), .Z(n10526) );
  NANDN U12430 ( .A(sreg[1188]), .B(n10487), .Z(n10491) );
  NAND U12431 ( .A(n10489), .B(n10488), .Z(n10490) );
  NAND U12432 ( .A(n10491), .B(n10490), .Z(n10525) );
  XNOR U12433 ( .A(n10526), .B(n10525), .Z(c[1189]) );
  NANDN U12434 ( .A(n10493), .B(n10492), .Z(n10497) );
  NANDN U12435 ( .A(n10495), .B(n10494), .Z(n10496) );
  AND U12436 ( .A(n10497), .B(n10496), .Z(n10532) );
  NANDN U12437 ( .A(n10499), .B(n10498), .Z(n10503) );
  NANDN U12438 ( .A(n10501), .B(n10500), .Z(n10502) );
  AND U12439 ( .A(n10503), .B(n10502), .Z(n10530) );
  NAND U12440 ( .A(n42143), .B(n10504), .Z(n10506) );
  XNOR U12441 ( .A(a[168]), .B(n4095), .Z(n10541) );
  NAND U12442 ( .A(n42144), .B(n10541), .Z(n10505) );
  AND U12443 ( .A(n10506), .B(n10505), .Z(n10556) );
  XOR U12444 ( .A(a[172]), .B(n42012), .Z(n10544) );
  XNOR U12445 ( .A(n10556), .B(n10555), .Z(n10558) );
  AND U12446 ( .A(a[174]), .B(b[0]), .Z(n10508) );
  XNOR U12447 ( .A(n10508), .B(n4071), .Z(n10510) );
  NANDN U12448 ( .A(b[0]), .B(a[173]), .Z(n10509) );
  NAND U12449 ( .A(n10510), .B(n10509), .Z(n10552) );
  XOR U12450 ( .A(a[170]), .B(n42085), .Z(n10548) );
  AND U12451 ( .A(a[166]), .B(b[7]), .Z(n10549) );
  XNOR U12452 ( .A(n10550), .B(n10549), .Z(n10551) );
  XNOR U12453 ( .A(n10552), .B(n10551), .Z(n10557) );
  XOR U12454 ( .A(n10558), .B(n10557), .Z(n10536) );
  NANDN U12455 ( .A(n10513), .B(n10512), .Z(n10517) );
  NANDN U12456 ( .A(n10515), .B(n10514), .Z(n10516) );
  AND U12457 ( .A(n10517), .B(n10516), .Z(n10535) );
  XNOR U12458 ( .A(n10536), .B(n10535), .Z(n10537) );
  NANDN U12459 ( .A(n10519), .B(n10518), .Z(n10523) );
  NAND U12460 ( .A(n10521), .B(n10520), .Z(n10522) );
  NAND U12461 ( .A(n10523), .B(n10522), .Z(n10538) );
  XNOR U12462 ( .A(n10537), .B(n10538), .Z(n10529) );
  XNOR U12463 ( .A(n10530), .B(n10529), .Z(n10531) );
  XNOR U12464 ( .A(n10532), .B(n10531), .Z(n10561) );
  XNOR U12465 ( .A(sreg[1190]), .B(n10561), .Z(n10563) );
  NANDN U12466 ( .A(sreg[1189]), .B(n10524), .Z(n10528) );
  NAND U12467 ( .A(n10526), .B(n10525), .Z(n10527) );
  NAND U12468 ( .A(n10528), .B(n10527), .Z(n10562) );
  XNOR U12469 ( .A(n10563), .B(n10562), .Z(c[1190]) );
  NANDN U12470 ( .A(n10530), .B(n10529), .Z(n10534) );
  NANDN U12471 ( .A(n10532), .B(n10531), .Z(n10533) );
  AND U12472 ( .A(n10534), .B(n10533), .Z(n10569) );
  NANDN U12473 ( .A(n10536), .B(n10535), .Z(n10540) );
  NANDN U12474 ( .A(n10538), .B(n10537), .Z(n10539) );
  AND U12475 ( .A(n10540), .B(n10539), .Z(n10567) );
  NAND U12476 ( .A(n42143), .B(n10541), .Z(n10543) );
  XNOR U12477 ( .A(a[169]), .B(n4096), .Z(n10578) );
  NAND U12478 ( .A(n42144), .B(n10578), .Z(n10542) );
  AND U12479 ( .A(n10543), .B(n10542), .Z(n10593) );
  XOR U12480 ( .A(a[173]), .B(n42012), .Z(n10581) );
  XNOR U12481 ( .A(n10593), .B(n10592), .Z(n10595) );
  AND U12482 ( .A(a[175]), .B(b[0]), .Z(n10545) );
  XNOR U12483 ( .A(n10545), .B(n4071), .Z(n10547) );
  NANDN U12484 ( .A(b[0]), .B(a[174]), .Z(n10546) );
  NAND U12485 ( .A(n10547), .B(n10546), .Z(n10589) );
  XOR U12486 ( .A(a[171]), .B(n42085), .Z(n10585) );
  AND U12487 ( .A(a[167]), .B(b[7]), .Z(n10586) );
  XNOR U12488 ( .A(n10587), .B(n10586), .Z(n10588) );
  XNOR U12489 ( .A(n10589), .B(n10588), .Z(n10594) );
  XOR U12490 ( .A(n10595), .B(n10594), .Z(n10573) );
  NANDN U12491 ( .A(n10550), .B(n10549), .Z(n10554) );
  NANDN U12492 ( .A(n10552), .B(n10551), .Z(n10553) );
  AND U12493 ( .A(n10554), .B(n10553), .Z(n10572) );
  XNOR U12494 ( .A(n10573), .B(n10572), .Z(n10574) );
  NANDN U12495 ( .A(n10556), .B(n10555), .Z(n10560) );
  NAND U12496 ( .A(n10558), .B(n10557), .Z(n10559) );
  NAND U12497 ( .A(n10560), .B(n10559), .Z(n10575) );
  XNOR U12498 ( .A(n10574), .B(n10575), .Z(n10566) );
  XNOR U12499 ( .A(n10567), .B(n10566), .Z(n10568) );
  XNOR U12500 ( .A(n10569), .B(n10568), .Z(n10598) );
  XNOR U12501 ( .A(sreg[1191]), .B(n10598), .Z(n10600) );
  NANDN U12502 ( .A(sreg[1190]), .B(n10561), .Z(n10565) );
  NAND U12503 ( .A(n10563), .B(n10562), .Z(n10564) );
  NAND U12504 ( .A(n10565), .B(n10564), .Z(n10599) );
  XNOR U12505 ( .A(n10600), .B(n10599), .Z(c[1191]) );
  NANDN U12506 ( .A(n10567), .B(n10566), .Z(n10571) );
  NANDN U12507 ( .A(n10569), .B(n10568), .Z(n10570) );
  AND U12508 ( .A(n10571), .B(n10570), .Z(n10606) );
  NANDN U12509 ( .A(n10573), .B(n10572), .Z(n10577) );
  NANDN U12510 ( .A(n10575), .B(n10574), .Z(n10576) );
  AND U12511 ( .A(n10577), .B(n10576), .Z(n10604) );
  NAND U12512 ( .A(n42143), .B(n10578), .Z(n10580) );
  XNOR U12513 ( .A(a[170]), .B(n4096), .Z(n10615) );
  NAND U12514 ( .A(n42144), .B(n10615), .Z(n10579) );
  AND U12515 ( .A(n10580), .B(n10579), .Z(n10630) );
  XOR U12516 ( .A(a[174]), .B(n42012), .Z(n10618) );
  XNOR U12517 ( .A(n10630), .B(n10629), .Z(n10632) );
  AND U12518 ( .A(a[176]), .B(b[0]), .Z(n10582) );
  XNOR U12519 ( .A(n10582), .B(n4071), .Z(n10584) );
  NANDN U12520 ( .A(b[0]), .B(a[175]), .Z(n10583) );
  NAND U12521 ( .A(n10584), .B(n10583), .Z(n10626) );
  XOR U12522 ( .A(a[172]), .B(n42085), .Z(n10619) );
  AND U12523 ( .A(a[168]), .B(b[7]), .Z(n10623) );
  XNOR U12524 ( .A(n10624), .B(n10623), .Z(n10625) );
  XNOR U12525 ( .A(n10626), .B(n10625), .Z(n10631) );
  XOR U12526 ( .A(n10632), .B(n10631), .Z(n10610) );
  NANDN U12527 ( .A(n10587), .B(n10586), .Z(n10591) );
  NANDN U12528 ( .A(n10589), .B(n10588), .Z(n10590) );
  AND U12529 ( .A(n10591), .B(n10590), .Z(n10609) );
  XNOR U12530 ( .A(n10610), .B(n10609), .Z(n10611) );
  NANDN U12531 ( .A(n10593), .B(n10592), .Z(n10597) );
  NAND U12532 ( .A(n10595), .B(n10594), .Z(n10596) );
  NAND U12533 ( .A(n10597), .B(n10596), .Z(n10612) );
  XNOR U12534 ( .A(n10611), .B(n10612), .Z(n10603) );
  XNOR U12535 ( .A(n10604), .B(n10603), .Z(n10605) );
  XNOR U12536 ( .A(n10606), .B(n10605), .Z(n10635) );
  XNOR U12537 ( .A(sreg[1192]), .B(n10635), .Z(n10637) );
  NANDN U12538 ( .A(sreg[1191]), .B(n10598), .Z(n10602) );
  NAND U12539 ( .A(n10600), .B(n10599), .Z(n10601) );
  NAND U12540 ( .A(n10602), .B(n10601), .Z(n10636) );
  XNOR U12541 ( .A(n10637), .B(n10636), .Z(c[1192]) );
  NANDN U12542 ( .A(n10604), .B(n10603), .Z(n10608) );
  NANDN U12543 ( .A(n10606), .B(n10605), .Z(n10607) );
  AND U12544 ( .A(n10608), .B(n10607), .Z(n10643) );
  NANDN U12545 ( .A(n10610), .B(n10609), .Z(n10614) );
  NANDN U12546 ( .A(n10612), .B(n10611), .Z(n10613) );
  AND U12547 ( .A(n10614), .B(n10613), .Z(n10641) );
  NAND U12548 ( .A(n42143), .B(n10615), .Z(n10617) );
  XNOR U12549 ( .A(a[171]), .B(n4096), .Z(n10652) );
  NAND U12550 ( .A(n42144), .B(n10652), .Z(n10616) );
  AND U12551 ( .A(n10617), .B(n10616), .Z(n10667) );
  XOR U12552 ( .A(a[175]), .B(n42012), .Z(n10655) );
  XNOR U12553 ( .A(n10667), .B(n10666), .Z(n10669) );
  XOR U12554 ( .A(a[173]), .B(n42085), .Z(n10656) );
  AND U12555 ( .A(a[169]), .B(b[7]), .Z(n10660) );
  XNOR U12556 ( .A(n10661), .B(n10660), .Z(n10662) );
  AND U12557 ( .A(a[177]), .B(b[0]), .Z(n10620) );
  XNOR U12558 ( .A(n10620), .B(n4071), .Z(n10622) );
  NANDN U12559 ( .A(b[0]), .B(a[176]), .Z(n10621) );
  NAND U12560 ( .A(n10622), .B(n10621), .Z(n10663) );
  XNOR U12561 ( .A(n10662), .B(n10663), .Z(n10668) );
  XOR U12562 ( .A(n10669), .B(n10668), .Z(n10647) );
  NANDN U12563 ( .A(n10624), .B(n10623), .Z(n10628) );
  NANDN U12564 ( .A(n10626), .B(n10625), .Z(n10627) );
  AND U12565 ( .A(n10628), .B(n10627), .Z(n10646) );
  XNOR U12566 ( .A(n10647), .B(n10646), .Z(n10648) );
  NANDN U12567 ( .A(n10630), .B(n10629), .Z(n10634) );
  NAND U12568 ( .A(n10632), .B(n10631), .Z(n10633) );
  NAND U12569 ( .A(n10634), .B(n10633), .Z(n10649) );
  XNOR U12570 ( .A(n10648), .B(n10649), .Z(n10640) );
  XNOR U12571 ( .A(n10641), .B(n10640), .Z(n10642) );
  XNOR U12572 ( .A(n10643), .B(n10642), .Z(n10672) );
  XNOR U12573 ( .A(sreg[1193]), .B(n10672), .Z(n10674) );
  NANDN U12574 ( .A(sreg[1192]), .B(n10635), .Z(n10639) );
  NAND U12575 ( .A(n10637), .B(n10636), .Z(n10638) );
  NAND U12576 ( .A(n10639), .B(n10638), .Z(n10673) );
  XNOR U12577 ( .A(n10674), .B(n10673), .Z(c[1193]) );
  NANDN U12578 ( .A(n10641), .B(n10640), .Z(n10645) );
  NANDN U12579 ( .A(n10643), .B(n10642), .Z(n10644) );
  AND U12580 ( .A(n10645), .B(n10644), .Z(n10680) );
  NANDN U12581 ( .A(n10647), .B(n10646), .Z(n10651) );
  NANDN U12582 ( .A(n10649), .B(n10648), .Z(n10650) );
  AND U12583 ( .A(n10651), .B(n10650), .Z(n10678) );
  NAND U12584 ( .A(n42143), .B(n10652), .Z(n10654) );
  XNOR U12585 ( .A(a[172]), .B(n4096), .Z(n10689) );
  NAND U12586 ( .A(n42144), .B(n10689), .Z(n10653) );
  AND U12587 ( .A(n10654), .B(n10653), .Z(n10704) );
  XOR U12588 ( .A(a[176]), .B(n42012), .Z(n10692) );
  XNOR U12589 ( .A(n10704), .B(n10703), .Z(n10706) );
  XOR U12590 ( .A(a[174]), .B(n42085), .Z(n10696) );
  AND U12591 ( .A(a[170]), .B(b[7]), .Z(n10697) );
  XNOR U12592 ( .A(n10698), .B(n10697), .Z(n10699) );
  AND U12593 ( .A(a[178]), .B(b[0]), .Z(n10657) );
  XNOR U12594 ( .A(n10657), .B(n4071), .Z(n10659) );
  NANDN U12595 ( .A(b[0]), .B(a[177]), .Z(n10658) );
  NAND U12596 ( .A(n10659), .B(n10658), .Z(n10700) );
  XNOR U12597 ( .A(n10699), .B(n10700), .Z(n10705) );
  XOR U12598 ( .A(n10706), .B(n10705), .Z(n10684) );
  NANDN U12599 ( .A(n10661), .B(n10660), .Z(n10665) );
  NANDN U12600 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U12601 ( .A(n10665), .B(n10664), .Z(n10683) );
  XNOR U12602 ( .A(n10684), .B(n10683), .Z(n10685) );
  NANDN U12603 ( .A(n10667), .B(n10666), .Z(n10671) );
  NAND U12604 ( .A(n10669), .B(n10668), .Z(n10670) );
  NAND U12605 ( .A(n10671), .B(n10670), .Z(n10686) );
  XNOR U12606 ( .A(n10685), .B(n10686), .Z(n10677) );
  XNOR U12607 ( .A(n10678), .B(n10677), .Z(n10679) );
  XNOR U12608 ( .A(n10680), .B(n10679), .Z(n10709) );
  XNOR U12609 ( .A(sreg[1194]), .B(n10709), .Z(n10711) );
  NANDN U12610 ( .A(sreg[1193]), .B(n10672), .Z(n10676) );
  NAND U12611 ( .A(n10674), .B(n10673), .Z(n10675) );
  NAND U12612 ( .A(n10676), .B(n10675), .Z(n10710) );
  XNOR U12613 ( .A(n10711), .B(n10710), .Z(c[1194]) );
  NANDN U12614 ( .A(n10678), .B(n10677), .Z(n10682) );
  NANDN U12615 ( .A(n10680), .B(n10679), .Z(n10681) );
  AND U12616 ( .A(n10682), .B(n10681), .Z(n10717) );
  NANDN U12617 ( .A(n10684), .B(n10683), .Z(n10688) );
  NANDN U12618 ( .A(n10686), .B(n10685), .Z(n10687) );
  AND U12619 ( .A(n10688), .B(n10687), .Z(n10715) );
  NAND U12620 ( .A(n42143), .B(n10689), .Z(n10691) );
  XNOR U12621 ( .A(a[173]), .B(n4096), .Z(n10726) );
  NAND U12622 ( .A(n42144), .B(n10726), .Z(n10690) );
  AND U12623 ( .A(n10691), .B(n10690), .Z(n10741) );
  XOR U12624 ( .A(a[177]), .B(n42012), .Z(n10729) );
  XNOR U12625 ( .A(n10741), .B(n10740), .Z(n10743) );
  AND U12626 ( .A(a[179]), .B(b[0]), .Z(n10693) );
  XNOR U12627 ( .A(n10693), .B(n4071), .Z(n10695) );
  NANDN U12628 ( .A(b[0]), .B(a[178]), .Z(n10694) );
  NAND U12629 ( .A(n10695), .B(n10694), .Z(n10737) );
  XOR U12630 ( .A(a[175]), .B(n42085), .Z(n10730) );
  AND U12631 ( .A(a[171]), .B(b[7]), .Z(n10734) );
  XNOR U12632 ( .A(n10735), .B(n10734), .Z(n10736) );
  XNOR U12633 ( .A(n10737), .B(n10736), .Z(n10742) );
  XOR U12634 ( .A(n10743), .B(n10742), .Z(n10721) );
  NANDN U12635 ( .A(n10698), .B(n10697), .Z(n10702) );
  NANDN U12636 ( .A(n10700), .B(n10699), .Z(n10701) );
  AND U12637 ( .A(n10702), .B(n10701), .Z(n10720) );
  XNOR U12638 ( .A(n10721), .B(n10720), .Z(n10722) );
  NANDN U12639 ( .A(n10704), .B(n10703), .Z(n10708) );
  NAND U12640 ( .A(n10706), .B(n10705), .Z(n10707) );
  NAND U12641 ( .A(n10708), .B(n10707), .Z(n10723) );
  XNOR U12642 ( .A(n10722), .B(n10723), .Z(n10714) );
  XNOR U12643 ( .A(n10715), .B(n10714), .Z(n10716) );
  XNOR U12644 ( .A(n10717), .B(n10716), .Z(n10746) );
  XNOR U12645 ( .A(sreg[1195]), .B(n10746), .Z(n10748) );
  NANDN U12646 ( .A(sreg[1194]), .B(n10709), .Z(n10713) );
  NAND U12647 ( .A(n10711), .B(n10710), .Z(n10712) );
  NAND U12648 ( .A(n10713), .B(n10712), .Z(n10747) );
  XNOR U12649 ( .A(n10748), .B(n10747), .Z(c[1195]) );
  NANDN U12650 ( .A(n10715), .B(n10714), .Z(n10719) );
  NANDN U12651 ( .A(n10717), .B(n10716), .Z(n10718) );
  AND U12652 ( .A(n10719), .B(n10718), .Z(n10754) );
  NANDN U12653 ( .A(n10721), .B(n10720), .Z(n10725) );
  NANDN U12654 ( .A(n10723), .B(n10722), .Z(n10724) );
  AND U12655 ( .A(n10725), .B(n10724), .Z(n10752) );
  NAND U12656 ( .A(n42143), .B(n10726), .Z(n10728) );
  XNOR U12657 ( .A(a[174]), .B(n4096), .Z(n10763) );
  NAND U12658 ( .A(n42144), .B(n10763), .Z(n10727) );
  AND U12659 ( .A(n10728), .B(n10727), .Z(n10778) );
  XOR U12660 ( .A(a[178]), .B(n42012), .Z(n10766) );
  XNOR U12661 ( .A(n10778), .B(n10777), .Z(n10780) );
  XOR U12662 ( .A(a[176]), .B(n42085), .Z(n10770) );
  AND U12663 ( .A(a[172]), .B(b[7]), .Z(n10771) );
  XNOR U12664 ( .A(n10772), .B(n10771), .Z(n10773) );
  AND U12665 ( .A(a[180]), .B(b[0]), .Z(n10731) );
  XNOR U12666 ( .A(n10731), .B(n4071), .Z(n10733) );
  NANDN U12667 ( .A(b[0]), .B(a[179]), .Z(n10732) );
  NAND U12668 ( .A(n10733), .B(n10732), .Z(n10774) );
  XNOR U12669 ( .A(n10773), .B(n10774), .Z(n10779) );
  XOR U12670 ( .A(n10780), .B(n10779), .Z(n10758) );
  NANDN U12671 ( .A(n10735), .B(n10734), .Z(n10739) );
  NANDN U12672 ( .A(n10737), .B(n10736), .Z(n10738) );
  AND U12673 ( .A(n10739), .B(n10738), .Z(n10757) );
  XNOR U12674 ( .A(n10758), .B(n10757), .Z(n10759) );
  NANDN U12675 ( .A(n10741), .B(n10740), .Z(n10745) );
  NAND U12676 ( .A(n10743), .B(n10742), .Z(n10744) );
  NAND U12677 ( .A(n10745), .B(n10744), .Z(n10760) );
  XNOR U12678 ( .A(n10759), .B(n10760), .Z(n10751) );
  XNOR U12679 ( .A(n10752), .B(n10751), .Z(n10753) );
  XNOR U12680 ( .A(n10754), .B(n10753), .Z(n10783) );
  XNOR U12681 ( .A(sreg[1196]), .B(n10783), .Z(n10785) );
  NANDN U12682 ( .A(sreg[1195]), .B(n10746), .Z(n10750) );
  NAND U12683 ( .A(n10748), .B(n10747), .Z(n10749) );
  NAND U12684 ( .A(n10750), .B(n10749), .Z(n10784) );
  XNOR U12685 ( .A(n10785), .B(n10784), .Z(c[1196]) );
  NANDN U12686 ( .A(n10752), .B(n10751), .Z(n10756) );
  NANDN U12687 ( .A(n10754), .B(n10753), .Z(n10755) );
  AND U12688 ( .A(n10756), .B(n10755), .Z(n10791) );
  NANDN U12689 ( .A(n10758), .B(n10757), .Z(n10762) );
  NANDN U12690 ( .A(n10760), .B(n10759), .Z(n10761) );
  AND U12691 ( .A(n10762), .B(n10761), .Z(n10789) );
  NAND U12692 ( .A(n42143), .B(n10763), .Z(n10765) );
  XNOR U12693 ( .A(a[175]), .B(n4096), .Z(n10800) );
  NAND U12694 ( .A(n42144), .B(n10800), .Z(n10764) );
  AND U12695 ( .A(n10765), .B(n10764), .Z(n10815) );
  XOR U12696 ( .A(a[179]), .B(n42012), .Z(n10803) );
  XNOR U12697 ( .A(n10815), .B(n10814), .Z(n10817) );
  AND U12698 ( .A(a[181]), .B(b[0]), .Z(n10767) );
  XNOR U12699 ( .A(n10767), .B(n4071), .Z(n10769) );
  NANDN U12700 ( .A(b[0]), .B(a[180]), .Z(n10768) );
  NAND U12701 ( .A(n10769), .B(n10768), .Z(n10811) );
  XOR U12702 ( .A(a[177]), .B(n42085), .Z(n10807) );
  AND U12703 ( .A(a[173]), .B(b[7]), .Z(n10808) );
  XNOR U12704 ( .A(n10809), .B(n10808), .Z(n10810) );
  XNOR U12705 ( .A(n10811), .B(n10810), .Z(n10816) );
  XOR U12706 ( .A(n10817), .B(n10816), .Z(n10795) );
  NANDN U12707 ( .A(n10772), .B(n10771), .Z(n10776) );
  NANDN U12708 ( .A(n10774), .B(n10773), .Z(n10775) );
  AND U12709 ( .A(n10776), .B(n10775), .Z(n10794) );
  XNOR U12710 ( .A(n10795), .B(n10794), .Z(n10796) );
  NANDN U12711 ( .A(n10778), .B(n10777), .Z(n10782) );
  NAND U12712 ( .A(n10780), .B(n10779), .Z(n10781) );
  NAND U12713 ( .A(n10782), .B(n10781), .Z(n10797) );
  XNOR U12714 ( .A(n10796), .B(n10797), .Z(n10788) );
  XNOR U12715 ( .A(n10789), .B(n10788), .Z(n10790) );
  XNOR U12716 ( .A(n10791), .B(n10790), .Z(n10820) );
  XNOR U12717 ( .A(sreg[1197]), .B(n10820), .Z(n10822) );
  NANDN U12718 ( .A(sreg[1196]), .B(n10783), .Z(n10787) );
  NAND U12719 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U12720 ( .A(n10787), .B(n10786), .Z(n10821) );
  XNOR U12721 ( .A(n10822), .B(n10821), .Z(c[1197]) );
  NANDN U12722 ( .A(n10789), .B(n10788), .Z(n10793) );
  NANDN U12723 ( .A(n10791), .B(n10790), .Z(n10792) );
  AND U12724 ( .A(n10793), .B(n10792), .Z(n10828) );
  NANDN U12725 ( .A(n10795), .B(n10794), .Z(n10799) );
  NANDN U12726 ( .A(n10797), .B(n10796), .Z(n10798) );
  AND U12727 ( .A(n10799), .B(n10798), .Z(n10826) );
  NAND U12728 ( .A(n42143), .B(n10800), .Z(n10802) );
  XNOR U12729 ( .A(a[176]), .B(n4097), .Z(n10837) );
  NAND U12730 ( .A(n42144), .B(n10837), .Z(n10801) );
  AND U12731 ( .A(n10802), .B(n10801), .Z(n10852) );
  XOR U12732 ( .A(a[180]), .B(n42012), .Z(n10840) );
  XNOR U12733 ( .A(n10852), .B(n10851), .Z(n10854) );
  AND U12734 ( .A(a[182]), .B(b[0]), .Z(n10804) );
  XNOR U12735 ( .A(n10804), .B(n4071), .Z(n10806) );
  NANDN U12736 ( .A(b[0]), .B(a[181]), .Z(n10805) );
  NAND U12737 ( .A(n10806), .B(n10805), .Z(n10848) );
  XOR U12738 ( .A(a[178]), .B(n42085), .Z(n10844) );
  AND U12739 ( .A(a[174]), .B(b[7]), .Z(n10845) );
  XNOR U12740 ( .A(n10846), .B(n10845), .Z(n10847) );
  XNOR U12741 ( .A(n10848), .B(n10847), .Z(n10853) );
  XOR U12742 ( .A(n10854), .B(n10853), .Z(n10832) );
  NANDN U12743 ( .A(n10809), .B(n10808), .Z(n10813) );
  NANDN U12744 ( .A(n10811), .B(n10810), .Z(n10812) );
  AND U12745 ( .A(n10813), .B(n10812), .Z(n10831) );
  XNOR U12746 ( .A(n10832), .B(n10831), .Z(n10833) );
  NANDN U12747 ( .A(n10815), .B(n10814), .Z(n10819) );
  NAND U12748 ( .A(n10817), .B(n10816), .Z(n10818) );
  NAND U12749 ( .A(n10819), .B(n10818), .Z(n10834) );
  XNOR U12750 ( .A(n10833), .B(n10834), .Z(n10825) );
  XNOR U12751 ( .A(n10826), .B(n10825), .Z(n10827) );
  XNOR U12752 ( .A(n10828), .B(n10827), .Z(n10857) );
  XNOR U12753 ( .A(sreg[1198]), .B(n10857), .Z(n10859) );
  NANDN U12754 ( .A(sreg[1197]), .B(n10820), .Z(n10824) );
  NAND U12755 ( .A(n10822), .B(n10821), .Z(n10823) );
  NAND U12756 ( .A(n10824), .B(n10823), .Z(n10858) );
  XNOR U12757 ( .A(n10859), .B(n10858), .Z(c[1198]) );
  NANDN U12758 ( .A(n10826), .B(n10825), .Z(n10830) );
  NANDN U12759 ( .A(n10828), .B(n10827), .Z(n10829) );
  AND U12760 ( .A(n10830), .B(n10829), .Z(n10865) );
  NANDN U12761 ( .A(n10832), .B(n10831), .Z(n10836) );
  NANDN U12762 ( .A(n10834), .B(n10833), .Z(n10835) );
  AND U12763 ( .A(n10836), .B(n10835), .Z(n10863) );
  NAND U12764 ( .A(n42143), .B(n10837), .Z(n10839) );
  XNOR U12765 ( .A(a[177]), .B(n4097), .Z(n10874) );
  NAND U12766 ( .A(n42144), .B(n10874), .Z(n10838) );
  AND U12767 ( .A(n10839), .B(n10838), .Z(n10889) );
  XOR U12768 ( .A(a[181]), .B(n42012), .Z(n10877) );
  XNOR U12769 ( .A(n10889), .B(n10888), .Z(n10891) );
  AND U12770 ( .A(b[0]), .B(a[183]), .Z(n10841) );
  XOR U12771 ( .A(b[1]), .B(n10841), .Z(n10843) );
  NANDN U12772 ( .A(b[0]), .B(a[182]), .Z(n10842) );
  AND U12773 ( .A(n10843), .B(n10842), .Z(n10884) );
  XOR U12774 ( .A(a[179]), .B(n42085), .Z(n10881) );
  AND U12775 ( .A(a[175]), .B(b[7]), .Z(n10882) );
  XOR U12776 ( .A(n10883), .B(n10882), .Z(n10885) );
  XNOR U12777 ( .A(n10884), .B(n10885), .Z(n10890) );
  XOR U12778 ( .A(n10891), .B(n10890), .Z(n10869) );
  NANDN U12779 ( .A(n10846), .B(n10845), .Z(n10850) );
  NANDN U12780 ( .A(n10848), .B(n10847), .Z(n10849) );
  AND U12781 ( .A(n10850), .B(n10849), .Z(n10868) );
  XNOR U12782 ( .A(n10869), .B(n10868), .Z(n10870) );
  NANDN U12783 ( .A(n10852), .B(n10851), .Z(n10856) );
  NAND U12784 ( .A(n10854), .B(n10853), .Z(n10855) );
  NAND U12785 ( .A(n10856), .B(n10855), .Z(n10871) );
  XNOR U12786 ( .A(n10870), .B(n10871), .Z(n10862) );
  XNOR U12787 ( .A(n10863), .B(n10862), .Z(n10864) );
  XNOR U12788 ( .A(n10865), .B(n10864), .Z(n10894) );
  XNOR U12789 ( .A(sreg[1199]), .B(n10894), .Z(n10896) );
  NANDN U12790 ( .A(sreg[1198]), .B(n10857), .Z(n10861) );
  NAND U12791 ( .A(n10859), .B(n10858), .Z(n10860) );
  NAND U12792 ( .A(n10861), .B(n10860), .Z(n10895) );
  XNOR U12793 ( .A(n10896), .B(n10895), .Z(c[1199]) );
  NANDN U12794 ( .A(n10863), .B(n10862), .Z(n10867) );
  NANDN U12795 ( .A(n10865), .B(n10864), .Z(n10866) );
  AND U12796 ( .A(n10867), .B(n10866), .Z(n10902) );
  NANDN U12797 ( .A(n10869), .B(n10868), .Z(n10873) );
  NANDN U12798 ( .A(n10871), .B(n10870), .Z(n10872) );
  AND U12799 ( .A(n10873), .B(n10872), .Z(n10900) );
  NAND U12800 ( .A(n42143), .B(n10874), .Z(n10876) );
  XNOR U12801 ( .A(a[178]), .B(n4097), .Z(n10911) );
  NAND U12802 ( .A(n42144), .B(n10911), .Z(n10875) );
  AND U12803 ( .A(n10876), .B(n10875), .Z(n10926) );
  XOR U12804 ( .A(a[182]), .B(n42012), .Z(n10914) );
  XNOR U12805 ( .A(n10926), .B(n10925), .Z(n10928) );
  AND U12806 ( .A(a[184]), .B(b[0]), .Z(n10878) );
  XNOR U12807 ( .A(n10878), .B(n4071), .Z(n10880) );
  NANDN U12808 ( .A(b[0]), .B(a[183]), .Z(n10879) );
  NAND U12809 ( .A(n10880), .B(n10879), .Z(n10922) );
  XOR U12810 ( .A(a[180]), .B(n42085), .Z(n10918) );
  AND U12811 ( .A(a[176]), .B(b[7]), .Z(n10919) );
  XNOR U12812 ( .A(n10920), .B(n10919), .Z(n10921) );
  XNOR U12813 ( .A(n10922), .B(n10921), .Z(n10927) );
  XOR U12814 ( .A(n10928), .B(n10927), .Z(n10906) );
  NANDN U12815 ( .A(n10883), .B(n10882), .Z(n10887) );
  NANDN U12816 ( .A(n10885), .B(n10884), .Z(n10886) );
  AND U12817 ( .A(n10887), .B(n10886), .Z(n10905) );
  XNOR U12818 ( .A(n10906), .B(n10905), .Z(n10907) );
  NANDN U12819 ( .A(n10889), .B(n10888), .Z(n10893) );
  NAND U12820 ( .A(n10891), .B(n10890), .Z(n10892) );
  NAND U12821 ( .A(n10893), .B(n10892), .Z(n10908) );
  XNOR U12822 ( .A(n10907), .B(n10908), .Z(n10899) );
  XNOR U12823 ( .A(n10900), .B(n10899), .Z(n10901) );
  XNOR U12824 ( .A(n10902), .B(n10901), .Z(n10931) );
  XNOR U12825 ( .A(sreg[1200]), .B(n10931), .Z(n10933) );
  NANDN U12826 ( .A(sreg[1199]), .B(n10894), .Z(n10898) );
  NAND U12827 ( .A(n10896), .B(n10895), .Z(n10897) );
  NAND U12828 ( .A(n10898), .B(n10897), .Z(n10932) );
  XNOR U12829 ( .A(n10933), .B(n10932), .Z(c[1200]) );
  NANDN U12830 ( .A(n10900), .B(n10899), .Z(n10904) );
  NANDN U12831 ( .A(n10902), .B(n10901), .Z(n10903) );
  AND U12832 ( .A(n10904), .B(n10903), .Z(n10939) );
  NANDN U12833 ( .A(n10906), .B(n10905), .Z(n10910) );
  NANDN U12834 ( .A(n10908), .B(n10907), .Z(n10909) );
  AND U12835 ( .A(n10910), .B(n10909), .Z(n10937) );
  NAND U12836 ( .A(n42143), .B(n10911), .Z(n10913) );
  XNOR U12837 ( .A(a[179]), .B(n4097), .Z(n10948) );
  NAND U12838 ( .A(n42144), .B(n10948), .Z(n10912) );
  AND U12839 ( .A(n10913), .B(n10912), .Z(n10963) );
  XOR U12840 ( .A(a[183]), .B(n42012), .Z(n10951) );
  XNOR U12841 ( .A(n10963), .B(n10962), .Z(n10965) );
  AND U12842 ( .A(a[185]), .B(b[0]), .Z(n10915) );
  XNOR U12843 ( .A(n10915), .B(n4071), .Z(n10917) );
  NANDN U12844 ( .A(b[0]), .B(a[184]), .Z(n10916) );
  NAND U12845 ( .A(n10917), .B(n10916), .Z(n10959) );
  XOR U12846 ( .A(a[181]), .B(n42085), .Z(n10955) );
  AND U12847 ( .A(a[177]), .B(b[7]), .Z(n10956) );
  XNOR U12848 ( .A(n10957), .B(n10956), .Z(n10958) );
  XNOR U12849 ( .A(n10959), .B(n10958), .Z(n10964) );
  XOR U12850 ( .A(n10965), .B(n10964), .Z(n10943) );
  NANDN U12851 ( .A(n10920), .B(n10919), .Z(n10924) );
  NANDN U12852 ( .A(n10922), .B(n10921), .Z(n10923) );
  AND U12853 ( .A(n10924), .B(n10923), .Z(n10942) );
  XNOR U12854 ( .A(n10943), .B(n10942), .Z(n10944) );
  NANDN U12855 ( .A(n10926), .B(n10925), .Z(n10930) );
  NAND U12856 ( .A(n10928), .B(n10927), .Z(n10929) );
  NAND U12857 ( .A(n10930), .B(n10929), .Z(n10945) );
  XNOR U12858 ( .A(n10944), .B(n10945), .Z(n10936) );
  XNOR U12859 ( .A(n10937), .B(n10936), .Z(n10938) );
  XNOR U12860 ( .A(n10939), .B(n10938), .Z(n10968) );
  XNOR U12861 ( .A(sreg[1201]), .B(n10968), .Z(n10970) );
  NANDN U12862 ( .A(sreg[1200]), .B(n10931), .Z(n10935) );
  NAND U12863 ( .A(n10933), .B(n10932), .Z(n10934) );
  NAND U12864 ( .A(n10935), .B(n10934), .Z(n10969) );
  XNOR U12865 ( .A(n10970), .B(n10969), .Z(c[1201]) );
  NANDN U12866 ( .A(n10937), .B(n10936), .Z(n10941) );
  NANDN U12867 ( .A(n10939), .B(n10938), .Z(n10940) );
  AND U12868 ( .A(n10941), .B(n10940), .Z(n10976) );
  NANDN U12869 ( .A(n10943), .B(n10942), .Z(n10947) );
  NANDN U12870 ( .A(n10945), .B(n10944), .Z(n10946) );
  AND U12871 ( .A(n10947), .B(n10946), .Z(n10974) );
  NAND U12872 ( .A(n42143), .B(n10948), .Z(n10950) );
  XNOR U12873 ( .A(a[180]), .B(n4097), .Z(n10985) );
  NAND U12874 ( .A(n42144), .B(n10985), .Z(n10949) );
  AND U12875 ( .A(n10950), .B(n10949), .Z(n11000) );
  XOR U12876 ( .A(a[184]), .B(n42012), .Z(n10988) );
  XNOR U12877 ( .A(n11000), .B(n10999), .Z(n11002) );
  AND U12878 ( .A(a[186]), .B(b[0]), .Z(n10952) );
  XNOR U12879 ( .A(n10952), .B(n4071), .Z(n10954) );
  NANDN U12880 ( .A(b[0]), .B(a[185]), .Z(n10953) );
  NAND U12881 ( .A(n10954), .B(n10953), .Z(n10996) );
  XOR U12882 ( .A(a[182]), .B(n42085), .Z(n10992) );
  AND U12883 ( .A(a[178]), .B(b[7]), .Z(n10993) );
  XNOR U12884 ( .A(n10994), .B(n10993), .Z(n10995) );
  XNOR U12885 ( .A(n10996), .B(n10995), .Z(n11001) );
  XOR U12886 ( .A(n11002), .B(n11001), .Z(n10980) );
  NANDN U12887 ( .A(n10957), .B(n10956), .Z(n10961) );
  NANDN U12888 ( .A(n10959), .B(n10958), .Z(n10960) );
  AND U12889 ( .A(n10961), .B(n10960), .Z(n10979) );
  XNOR U12890 ( .A(n10980), .B(n10979), .Z(n10981) );
  NANDN U12891 ( .A(n10963), .B(n10962), .Z(n10967) );
  NAND U12892 ( .A(n10965), .B(n10964), .Z(n10966) );
  NAND U12893 ( .A(n10967), .B(n10966), .Z(n10982) );
  XNOR U12894 ( .A(n10981), .B(n10982), .Z(n10973) );
  XNOR U12895 ( .A(n10974), .B(n10973), .Z(n10975) );
  XNOR U12896 ( .A(n10976), .B(n10975), .Z(n11005) );
  XNOR U12897 ( .A(sreg[1202]), .B(n11005), .Z(n11007) );
  NANDN U12898 ( .A(sreg[1201]), .B(n10968), .Z(n10972) );
  NAND U12899 ( .A(n10970), .B(n10969), .Z(n10971) );
  NAND U12900 ( .A(n10972), .B(n10971), .Z(n11006) );
  XNOR U12901 ( .A(n11007), .B(n11006), .Z(c[1202]) );
  NANDN U12902 ( .A(n10974), .B(n10973), .Z(n10978) );
  NANDN U12903 ( .A(n10976), .B(n10975), .Z(n10977) );
  AND U12904 ( .A(n10978), .B(n10977), .Z(n11013) );
  NANDN U12905 ( .A(n10980), .B(n10979), .Z(n10984) );
  NANDN U12906 ( .A(n10982), .B(n10981), .Z(n10983) );
  AND U12907 ( .A(n10984), .B(n10983), .Z(n11011) );
  NAND U12908 ( .A(n42143), .B(n10985), .Z(n10987) );
  XNOR U12909 ( .A(a[181]), .B(n4097), .Z(n11022) );
  NAND U12910 ( .A(n42144), .B(n11022), .Z(n10986) );
  AND U12911 ( .A(n10987), .B(n10986), .Z(n11037) );
  XOR U12912 ( .A(a[185]), .B(n42012), .Z(n11025) );
  XNOR U12913 ( .A(n11037), .B(n11036), .Z(n11039) );
  AND U12914 ( .A(a[187]), .B(b[0]), .Z(n10989) );
  XNOR U12915 ( .A(n10989), .B(n4071), .Z(n10991) );
  NANDN U12916 ( .A(b[0]), .B(a[186]), .Z(n10990) );
  NAND U12917 ( .A(n10991), .B(n10990), .Z(n11033) );
  XOR U12918 ( .A(a[183]), .B(n42085), .Z(n11026) );
  AND U12919 ( .A(a[179]), .B(b[7]), .Z(n11030) );
  XNOR U12920 ( .A(n11031), .B(n11030), .Z(n11032) );
  XNOR U12921 ( .A(n11033), .B(n11032), .Z(n11038) );
  XOR U12922 ( .A(n11039), .B(n11038), .Z(n11017) );
  NANDN U12923 ( .A(n10994), .B(n10993), .Z(n10998) );
  NANDN U12924 ( .A(n10996), .B(n10995), .Z(n10997) );
  AND U12925 ( .A(n10998), .B(n10997), .Z(n11016) );
  XNOR U12926 ( .A(n11017), .B(n11016), .Z(n11018) );
  NANDN U12927 ( .A(n11000), .B(n10999), .Z(n11004) );
  NAND U12928 ( .A(n11002), .B(n11001), .Z(n11003) );
  NAND U12929 ( .A(n11004), .B(n11003), .Z(n11019) );
  XNOR U12930 ( .A(n11018), .B(n11019), .Z(n11010) );
  XNOR U12931 ( .A(n11011), .B(n11010), .Z(n11012) );
  XNOR U12932 ( .A(n11013), .B(n11012), .Z(n11042) );
  XNOR U12933 ( .A(sreg[1203]), .B(n11042), .Z(n11044) );
  NANDN U12934 ( .A(sreg[1202]), .B(n11005), .Z(n11009) );
  NAND U12935 ( .A(n11007), .B(n11006), .Z(n11008) );
  NAND U12936 ( .A(n11009), .B(n11008), .Z(n11043) );
  XNOR U12937 ( .A(n11044), .B(n11043), .Z(c[1203]) );
  NANDN U12938 ( .A(n11011), .B(n11010), .Z(n11015) );
  NANDN U12939 ( .A(n11013), .B(n11012), .Z(n11014) );
  AND U12940 ( .A(n11015), .B(n11014), .Z(n11050) );
  NANDN U12941 ( .A(n11017), .B(n11016), .Z(n11021) );
  NANDN U12942 ( .A(n11019), .B(n11018), .Z(n11020) );
  AND U12943 ( .A(n11021), .B(n11020), .Z(n11048) );
  NAND U12944 ( .A(n42143), .B(n11022), .Z(n11024) );
  XNOR U12945 ( .A(a[182]), .B(n4097), .Z(n11059) );
  NAND U12946 ( .A(n42144), .B(n11059), .Z(n11023) );
  AND U12947 ( .A(n11024), .B(n11023), .Z(n11074) );
  XOR U12948 ( .A(a[186]), .B(n42012), .Z(n11062) );
  XNOR U12949 ( .A(n11074), .B(n11073), .Z(n11076) );
  XOR U12950 ( .A(a[184]), .B(n42085), .Z(n11066) );
  AND U12951 ( .A(a[180]), .B(b[7]), .Z(n11067) );
  XNOR U12952 ( .A(n11068), .B(n11067), .Z(n11069) );
  AND U12953 ( .A(a[188]), .B(b[0]), .Z(n11027) );
  XNOR U12954 ( .A(n11027), .B(n4071), .Z(n11029) );
  NANDN U12955 ( .A(b[0]), .B(a[187]), .Z(n11028) );
  NAND U12956 ( .A(n11029), .B(n11028), .Z(n11070) );
  XNOR U12957 ( .A(n11069), .B(n11070), .Z(n11075) );
  XOR U12958 ( .A(n11076), .B(n11075), .Z(n11054) );
  NANDN U12959 ( .A(n11031), .B(n11030), .Z(n11035) );
  NANDN U12960 ( .A(n11033), .B(n11032), .Z(n11034) );
  AND U12961 ( .A(n11035), .B(n11034), .Z(n11053) );
  XNOR U12962 ( .A(n11054), .B(n11053), .Z(n11055) );
  NANDN U12963 ( .A(n11037), .B(n11036), .Z(n11041) );
  NAND U12964 ( .A(n11039), .B(n11038), .Z(n11040) );
  NAND U12965 ( .A(n11041), .B(n11040), .Z(n11056) );
  XNOR U12966 ( .A(n11055), .B(n11056), .Z(n11047) );
  XNOR U12967 ( .A(n11048), .B(n11047), .Z(n11049) );
  XNOR U12968 ( .A(n11050), .B(n11049), .Z(n11079) );
  XNOR U12969 ( .A(sreg[1204]), .B(n11079), .Z(n11081) );
  NANDN U12970 ( .A(sreg[1203]), .B(n11042), .Z(n11046) );
  NAND U12971 ( .A(n11044), .B(n11043), .Z(n11045) );
  NAND U12972 ( .A(n11046), .B(n11045), .Z(n11080) );
  XNOR U12973 ( .A(n11081), .B(n11080), .Z(c[1204]) );
  NANDN U12974 ( .A(n11048), .B(n11047), .Z(n11052) );
  NANDN U12975 ( .A(n11050), .B(n11049), .Z(n11051) );
  AND U12976 ( .A(n11052), .B(n11051), .Z(n11087) );
  NANDN U12977 ( .A(n11054), .B(n11053), .Z(n11058) );
  NANDN U12978 ( .A(n11056), .B(n11055), .Z(n11057) );
  AND U12979 ( .A(n11058), .B(n11057), .Z(n11085) );
  NAND U12980 ( .A(n42143), .B(n11059), .Z(n11061) );
  XNOR U12981 ( .A(a[183]), .B(n4098), .Z(n11096) );
  NAND U12982 ( .A(n42144), .B(n11096), .Z(n11060) );
  AND U12983 ( .A(n11061), .B(n11060), .Z(n11111) );
  XOR U12984 ( .A(a[187]), .B(n42012), .Z(n11099) );
  XNOR U12985 ( .A(n11111), .B(n11110), .Z(n11113) );
  AND U12986 ( .A(a[189]), .B(b[0]), .Z(n11063) );
  XNOR U12987 ( .A(n11063), .B(n4071), .Z(n11065) );
  NANDN U12988 ( .A(b[0]), .B(a[188]), .Z(n11064) );
  NAND U12989 ( .A(n11065), .B(n11064), .Z(n11107) );
  XOR U12990 ( .A(a[185]), .B(n42085), .Z(n11100) );
  AND U12991 ( .A(a[181]), .B(b[7]), .Z(n11104) );
  XNOR U12992 ( .A(n11105), .B(n11104), .Z(n11106) );
  XNOR U12993 ( .A(n11107), .B(n11106), .Z(n11112) );
  XOR U12994 ( .A(n11113), .B(n11112), .Z(n11091) );
  NANDN U12995 ( .A(n11068), .B(n11067), .Z(n11072) );
  NANDN U12996 ( .A(n11070), .B(n11069), .Z(n11071) );
  AND U12997 ( .A(n11072), .B(n11071), .Z(n11090) );
  XNOR U12998 ( .A(n11091), .B(n11090), .Z(n11092) );
  NANDN U12999 ( .A(n11074), .B(n11073), .Z(n11078) );
  NAND U13000 ( .A(n11076), .B(n11075), .Z(n11077) );
  NAND U13001 ( .A(n11078), .B(n11077), .Z(n11093) );
  XNOR U13002 ( .A(n11092), .B(n11093), .Z(n11084) );
  XNOR U13003 ( .A(n11085), .B(n11084), .Z(n11086) );
  XNOR U13004 ( .A(n11087), .B(n11086), .Z(n11116) );
  XNOR U13005 ( .A(sreg[1205]), .B(n11116), .Z(n11118) );
  NANDN U13006 ( .A(sreg[1204]), .B(n11079), .Z(n11083) );
  NAND U13007 ( .A(n11081), .B(n11080), .Z(n11082) );
  NAND U13008 ( .A(n11083), .B(n11082), .Z(n11117) );
  XNOR U13009 ( .A(n11118), .B(n11117), .Z(c[1205]) );
  NANDN U13010 ( .A(n11085), .B(n11084), .Z(n11089) );
  NANDN U13011 ( .A(n11087), .B(n11086), .Z(n11088) );
  AND U13012 ( .A(n11089), .B(n11088), .Z(n11124) );
  NANDN U13013 ( .A(n11091), .B(n11090), .Z(n11095) );
  NANDN U13014 ( .A(n11093), .B(n11092), .Z(n11094) );
  AND U13015 ( .A(n11095), .B(n11094), .Z(n11122) );
  NAND U13016 ( .A(n42143), .B(n11096), .Z(n11098) );
  XNOR U13017 ( .A(a[184]), .B(n4098), .Z(n11133) );
  NAND U13018 ( .A(n42144), .B(n11133), .Z(n11097) );
  AND U13019 ( .A(n11098), .B(n11097), .Z(n11148) );
  XOR U13020 ( .A(a[188]), .B(n42012), .Z(n11136) );
  XNOR U13021 ( .A(n11148), .B(n11147), .Z(n11150) );
  XOR U13022 ( .A(a[186]), .B(n42085), .Z(n11137) );
  AND U13023 ( .A(a[182]), .B(b[7]), .Z(n11141) );
  XNOR U13024 ( .A(n11142), .B(n11141), .Z(n11143) );
  AND U13025 ( .A(a[190]), .B(b[0]), .Z(n11101) );
  XNOR U13026 ( .A(n11101), .B(n4071), .Z(n11103) );
  NANDN U13027 ( .A(b[0]), .B(a[189]), .Z(n11102) );
  NAND U13028 ( .A(n11103), .B(n11102), .Z(n11144) );
  XNOR U13029 ( .A(n11143), .B(n11144), .Z(n11149) );
  XOR U13030 ( .A(n11150), .B(n11149), .Z(n11128) );
  NANDN U13031 ( .A(n11105), .B(n11104), .Z(n11109) );
  NANDN U13032 ( .A(n11107), .B(n11106), .Z(n11108) );
  AND U13033 ( .A(n11109), .B(n11108), .Z(n11127) );
  XNOR U13034 ( .A(n11128), .B(n11127), .Z(n11129) );
  NANDN U13035 ( .A(n11111), .B(n11110), .Z(n11115) );
  NAND U13036 ( .A(n11113), .B(n11112), .Z(n11114) );
  NAND U13037 ( .A(n11115), .B(n11114), .Z(n11130) );
  XNOR U13038 ( .A(n11129), .B(n11130), .Z(n11121) );
  XNOR U13039 ( .A(n11122), .B(n11121), .Z(n11123) );
  XNOR U13040 ( .A(n11124), .B(n11123), .Z(n11153) );
  XNOR U13041 ( .A(sreg[1206]), .B(n11153), .Z(n11155) );
  NANDN U13042 ( .A(sreg[1205]), .B(n11116), .Z(n11120) );
  NAND U13043 ( .A(n11118), .B(n11117), .Z(n11119) );
  NAND U13044 ( .A(n11120), .B(n11119), .Z(n11154) );
  XNOR U13045 ( .A(n11155), .B(n11154), .Z(c[1206]) );
  NANDN U13046 ( .A(n11122), .B(n11121), .Z(n11126) );
  NANDN U13047 ( .A(n11124), .B(n11123), .Z(n11125) );
  AND U13048 ( .A(n11126), .B(n11125), .Z(n11161) );
  NANDN U13049 ( .A(n11128), .B(n11127), .Z(n11132) );
  NANDN U13050 ( .A(n11130), .B(n11129), .Z(n11131) );
  AND U13051 ( .A(n11132), .B(n11131), .Z(n11159) );
  NAND U13052 ( .A(n42143), .B(n11133), .Z(n11135) );
  XNOR U13053 ( .A(a[185]), .B(n4098), .Z(n11170) );
  NAND U13054 ( .A(n42144), .B(n11170), .Z(n11134) );
  AND U13055 ( .A(n11135), .B(n11134), .Z(n11185) );
  XOR U13056 ( .A(a[189]), .B(n42012), .Z(n11173) );
  XNOR U13057 ( .A(n11185), .B(n11184), .Z(n11187) );
  XOR U13058 ( .A(a[187]), .B(n42085), .Z(n11177) );
  AND U13059 ( .A(a[183]), .B(b[7]), .Z(n11178) );
  XNOR U13060 ( .A(n11179), .B(n11178), .Z(n11180) );
  AND U13061 ( .A(a[191]), .B(b[0]), .Z(n11138) );
  XNOR U13062 ( .A(n11138), .B(n4071), .Z(n11140) );
  NANDN U13063 ( .A(b[0]), .B(a[190]), .Z(n11139) );
  NAND U13064 ( .A(n11140), .B(n11139), .Z(n11181) );
  XNOR U13065 ( .A(n11180), .B(n11181), .Z(n11186) );
  XOR U13066 ( .A(n11187), .B(n11186), .Z(n11165) );
  NANDN U13067 ( .A(n11142), .B(n11141), .Z(n11146) );
  NANDN U13068 ( .A(n11144), .B(n11143), .Z(n11145) );
  AND U13069 ( .A(n11146), .B(n11145), .Z(n11164) );
  XNOR U13070 ( .A(n11165), .B(n11164), .Z(n11166) );
  NANDN U13071 ( .A(n11148), .B(n11147), .Z(n11152) );
  NAND U13072 ( .A(n11150), .B(n11149), .Z(n11151) );
  NAND U13073 ( .A(n11152), .B(n11151), .Z(n11167) );
  XNOR U13074 ( .A(n11166), .B(n11167), .Z(n11158) );
  XNOR U13075 ( .A(n11159), .B(n11158), .Z(n11160) );
  XNOR U13076 ( .A(n11161), .B(n11160), .Z(n11190) );
  XNOR U13077 ( .A(sreg[1207]), .B(n11190), .Z(n11192) );
  NANDN U13078 ( .A(sreg[1206]), .B(n11153), .Z(n11157) );
  NAND U13079 ( .A(n11155), .B(n11154), .Z(n11156) );
  NAND U13080 ( .A(n11157), .B(n11156), .Z(n11191) );
  XNOR U13081 ( .A(n11192), .B(n11191), .Z(c[1207]) );
  NANDN U13082 ( .A(n11159), .B(n11158), .Z(n11163) );
  NANDN U13083 ( .A(n11161), .B(n11160), .Z(n11162) );
  AND U13084 ( .A(n11163), .B(n11162), .Z(n11198) );
  NANDN U13085 ( .A(n11165), .B(n11164), .Z(n11169) );
  NANDN U13086 ( .A(n11167), .B(n11166), .Z(n11168) );
  AND U13087 ( .A(n11169), .B(n11168), .Z(n11196) );
  NAND U13088 ( .A(n42143), .B(n11170), .Z(n11172) );
  XNOR U13089 ( .A(a[186]), .B(n4098), .Z(n11207) );
  NAND U13090 ( .A(n42144), .B(n11207), .Z(n11171) );
  AND U13091 ( .A(n11172), .B(n11171), .Z(n11222) );
  XOR U13092 ( .A(a[190]), .B(n42012), .Z(n11210) );
  XNOR U13093 ( .A(n11222), .B(n11221), .Z(n11224) );
  AND U13094 ( .A(a[192]), .B(b[0]), .Z(n11174) );
  XNOR U13095 ( .A(n11174), .B(n4071), .Z(n11176) );
  NANDN U13096 ( .A(b[0]), .B(a[191]), .Z(n11175) );
  NAND U13097 ( .A(n11176), .B(n11175), .Z(n11218) );
  XOR U13098 ( .A(a[188]), .B(n42085), .Z(n11214) );
  AND U13099 ( .A(a[184]), .B(b[7]), .Z(n11215) );
  XNOR U13100 ( .A(n11216), .B(n11215), .Z(n11217) );
  XNOR U13101 ( .A(n11218), .B(n11217), .Z(n11223) );
  XOR U13102 ( .A(n11224), .B(n11223), .Z(n11202) );
  NANDN U13103 ( .A(n11179), .B(n11178), .Z(n11183) );
  NANDN U13104 ( .A(n11181), .B(n11180), .Z(n11182) );
  AND U13105 ( .A(n11183), .B(n11182), .Z(n11201) );
  XNOR U13106 ( .A(n11202), .B(n11201), .Z(n11203) );
  NANDN U13107 ( .A(n11185), .B(n11184), .Z(n11189) );
  NAND U13108 ( .A(n11187), .B(n11186), .Z(n11188) );
  NAND U13109 ( .A(n11189), .B(n11188), .Z(n11204) );
  XNOR U13110 ( .A(n11203), .B(n11204), .Z(n11195) );
  XNOR U13111 ( .A(n11196), .B(n11195), .Z(n11197) );
  XNOR U13112 ( .A(n11198), .B(n11197), .Z(n11227) );
  XNOR U13113 ( .A(sreg[1208]), .B(n11227), .Z(n11229) );
  NANDN U13114 ( .A(sreg[1207]), .B(n11190), .Z(n11194) );
  NAND U13115 ( .A(n11192), .B(n11191), .Z(n11193) );
  NAND U13116 ( .A(n11194), .B(n11193), .Z(n11228) );
  XNOR U13117 ( .A(n11229), .B(n11228), .Z(c[1208]) );
  NANDN U13118 ( .A(n11196), .B(n11195), .Z(n11200) );
  NANDN U13119 ( .A(n11198), .B(n11197), .Z(n11199) );
  AND U13120 ( .A(n11200), .B(n11199), .Z(n11235) );
  NANDN U13121 ( .A(n11202), .B(n11201), .Z(n11206) );
  NANDN U13122 ( .A(n11204), .B(n11203), .Z(n11205) );
  AND U13123 ( .A(n11206), .B(n11205), .Z(n11233) );
  NAND U13124 ( .A(n42143), .B(n11207), .Z(n11209) );
  XNOR U13125 ( .A(a[187]), .B(n4098), .Z(n11244) );
  NAND U13126 ( .A(n42144), .B(n11244), .Z(n11208) );
  AND U13127 ( .A(n11209), .B(n11208), .Z(n11259) );
  XOR U13128 ( .A(a[191]), .B(n42012), .Z(n11247) );
  XNOR U13129 ( .A(n11259), .B(n11258), .Z(n11261) );
  AND U13130 ( .A(a[193]), .B(b[0]), .Z(n11211) );
  XNOR U13131 ( .A(n11211), .B(n4071), .Z(n11213) );
  NANDN U13132 ( .A(b[0]), .B(a[192]), .Z(n11212) );
  NAND U13133 ( .A(n11213), .B(n11212), .Z(n11255) );
  XOR U13134 ( .A(a[189]), .B(n42085), .Z(n11251) );
  AND U13135 ( .A(a[185]), .B(b[7]), .Z(n11252) );
  XNOR U13136 ( .A(n11253), .B(n11252), .Z(n11254) );
  XNOR U13137 ( .A(n11255), .B(n11254), .Z(n11260) );
  XOR U13138 ( .A(n11261), .B(n11260), .Z(n11239) );
  NANDN U13139 ( .A(n11216), .B(n11215), .Z(n11220) );
  NANDN U13140 ( .A(n11218), .B(n11217), .Z(n11219) );
  AND U13141 ( .A(n11220), .B(n11219), .Z(n11238) );
  XNOR U13142 ( .A(n11239), .B(n11238), .Z(n11240) );
  NANDN U13143 ( .A(n11222), .B(n11221), .Z(n11226) );
  NAND U13144 ( .A(n11224), .B(n11223), .Z(n11225) );
  NAND U13145 ( .A(n11226), .B(n11225), .Z(n11241) );
  XNOR U13146 ( .A(n11240), .B(n11241), .Z(n11232) );
  XNOR U13147 ( .A(n11233), .B(n11232), .Z(n11234) );
  XNOR U13148 ( .A(n11235), .B(n11234), .Z(n11264) );
  XNOR U13149 ( .A(sreg[1209]), .B(n11264), .Z(n11266) );
  NANDN U13150 ( .A(sreg[1208]), .B(n11227), .Z(n11231) );
  NAND U13151 ( .A(n11229), .B(n11228), .Z(n11230) );
  NAND U13152 ( .A(n11231), .B(n11230), .Z(n11265) );
  XNOR U13153 ( .A(n11266), .B(n11265), .Z(c[1209]) );
  NANDN U13154 ( .A(n11233), .B(n11232), .Z(n11237) );
  NANDN U13155 ( .A(n11235), .B(n11234), .Z(n11236) );
  AND U13156 ( .A(n11237), .B(n11236), .Z(n11272) );
  NANDN U13157 ( .A(n11239), .B(n11238), .Z(n11243) );
  NANDN U13158 ( .A(n11241), .B(n11240), .Z(n11242) );
  AND U13159 ( .A(n11243), .B(n11242), .Z(n11270) );
  NAND U13160 ( .A(n42143), .B(n11244), .Z(n11246) );
  XNOR U13161 ( .A(a[188]), .B(n4098), .Z(n11281) );
  NAND U13162 ( .A(n42144), .B(n11281), .Z(n11245) );
  AND U13163 ( .A(n11246), .B(n11245), .Z(n11296) );
  XOR U13164 ( .A(a[192]), .B(n42012), .Z(n11284) );
  XNOR U13165 ( .A(n11296), .B(n11295), .Z(n11298) );
  AND U13166 ( .A(a[194]), .B(b[0]), .Z(n11248) );
  XNOR U13167 ( .A(n11248), .B(n4071), .Z(n11250) );
  NANDN U13168 ( .A(b[0]), .B(a[193]), .Z(n11249) );
  NAND U13169 ( .A(n11250), .B(n11249), .Z(n11292) );
  XOR U13170 ( .A(a[190]), .B(n42085), .Z(n11285) );
  AND U13171 ( .A(a[186]), .B(b[7]), .Z(n11289) );
  XNOR U13172 ( .A(n11290), .B(n11289), .Z(n11291) );
  XNOR U13173 ( .A(n11292), .B(n11291), .Z(n11297) );
  XOR U13174 ( .A(n11298), .B(n11297), .Z(n11276) );
  NANDN U13175 ( .A(n11253), .B(n11252), .Z(n11257) );
  NANDN U13176 ( .A(n11255), .B(n11254), .Z(n11256) );
  AND U13177 ( .A(n11257), .B(n11256), .Z(n11275) );
  XNOR U13178 ( .A(n11276), .B(n11275), .Z(n11277) );
  NANDN U13179 ( .A(n11259), .B(n11258), .Z(n11263) );
  NAND U13180 ( .A(n11261), .B(n11260), .Z(n11262) );
  NAND U13181 ( .A(n11263), .B(n11262), .Z(n11278) );
  XNOR U13182 ( .A(n11277), .B(n11278), .Z(n11269) );
  XNOR U13183 ( .A(n11270), .B(n11269), .Z(n11271) );
  XNOR U13184 ( .A(n11272), .B(n11271), .Z(n11301) );
  XNOR U13185 ( .A(sreg[1210]), .B(n11301), .Z(n11303) );
  NANDN U13186 ( .A(sreg[1209]), .B(n11264), .Z(n11268) );
  NAND U13187 ( .A(n11266), .B(n11265), .Z(n11267) );
  NAND U13188 ( .A(n11268), .B(n11267), .Z(n11302) );
  XNOR U13189 ( .A(n11303), .B(n11302), .Z(c[1210]) );
  NANDN U13190 ( .A(n11270), .B(n11269), .Z(n11274) );
  NANDN U13191 ( .A(n11272), .B(n11271), .Z(n11273) );
  AND U13192 ( .A(n11274), .B(n11273), .Z(n11309) );
  NANDN U13193 ( .A(n11276), .B(n11275), .Z(n11280) );
  NANDN U13194 ( .A(n11278), .B(n11277), .Z(n11279) );
  AND U13195 ( .A(n11280), .B(n11279), .Z(n11307) );
  NAND U13196 ( .A(n42143), .B(n11281), .Z(n11283) );
  XNOR U13197 ( .A(a[189]), .B(n4098), .Z(n11318) );
  NAND U13198 ( .A(n42144), .B(n11318), .Z(n11282) );
  AND U13199 ( .A(n11283), .B(n11282), .Z(n11333) );
  XOR U13200 ( .A(a[193]), .B(n42012), .Z(n11321) );
  XNOR U13201 ( .A(n11333), .B(n11332), .Z(n11335) );
  XOR U13202 ( .A(a[191]), .B(n42085), .Z(n11322) );
  AND U13203 ( .A(a[187]), .B(b[7]), .Z(n11326) );
  XNOR U13204 ( .A(n11327), .B(n11326), .Z(n11328) );
  AND U13205 ( .A(a[195]), .B(b[0]), .Z(n11286) );
  XNOR U13206 ( .A(n11286), .B(n4071), .Z(n11288) );
  NANDN U13207 ( .A(b[0]), .B(a[194]), .Z(n11287) );
  NAND U13208 ( .A(n11288), .B(n11287), .Z(n11329) );
  XNOR U13209 ( .A(n11328), .B(n11329), .Z(n11334) );
  XOR U13210 ( .A(n11335), .B(n11334), .Z(n11313) );
  NANDN U13211 ( .A(n11290), .B(n11289), .Z(n11294) );
  NANDN U13212 ( .A(n11292), .B(n11291), .Z(n11293) );
  AND U13213 ( .A(n11294), .B(n11293), .Z(n11312) );
  XNOR U13214 ( .A(n11313), .B(n11312), .Z(n11314) );
  NANDN U13215 ( .A(n11296), .B(n11295), .Z(n11300) );
  NAND U13216 ( .A(n11298), .B(n11297), .Z(n11299) );
  NAND U13217 ( .A(n11300), .B(n11299), .Z(n11315) );
  XNOR U13218 ( .A(n11314), .B(n11315), .Z(n11306) );
  XNOR U13219 ( .A(n11307), .B(n11306), .Z(n11308) );
  XNOR U13220 ( .A(n11309), .B(n11308), .Z(n11338) );
  XNOR U13221 ( .A(sreg[1211]), .B(n11338), .Z(n11340) );
  NANDN U13222 ( .A(sreg[1210]), .B(n11301), .Z(n11305) );
  NAND U13223 ( .A(n11303), .B(n11302), .Z(n11304) );
  NAND U13224 ( .A(n11305), .B(n11304), .Z(n11339) );
  XNOR U13225 ( .A(n11340), .B(n11339), .Z(c[1211]) );
  NANDN U13226 ( .A(n11307), .B(n11306), .Z(n11311) );
  NANDN U13227 ( .A(n11309), .B(n11308), .Z(n11310) );
  AND U13228 ( .A(n11311), .B(n11310), .Z(n11346) );
  NANDN U13229 ( .A(n11313), .B(n11312), .Z(n11317) );
  NANDN U13230 ( .A(n11315), .B(n11314), .Z(n11316) );
  AND U13231 ( .A(n11317), .B(n11316), .Z(n11344) );
  NAND U13232 ( .A(n42143), .B(n11318), .Z(n11320) );
  XNOR U13233 ( .A(a[190]), .B(n4099), .Z(n11355) );
  NAND U13234 ( .A(n42144), .B(n11355), .Z(n11319) );
  AND U13235 ( .A(n11320), .B(n11319), .Z(n11370) );
  XOR U13236 ( .A(a[194]), .B(n42012), .Z(n11358) );
  XNOR U13237 ( .A(n11370), .B(n11369), .Z(n11372) );
  XOR U13238 ( .A(a[192]), .B(n42085), .Z(n11362) );
  AND U13239 ( .A(a[188]), .B(b[7]), .Z(n11363) );
  XNOR U13240 ( .A(n11364), .B(n11363), .Z(n11365) );
  AND U13241 ( .A(a[196]), .B(b[0]), .Z(n11323) );
  XNOR U13242 ( .A(n11323), .B(n4071), .Z(n11325) );
  NANDN U13243 ( .A(b[0]), .B(a[195]), .Z(n11324) );
  NAND U13244 ( .A(n11325), .B(n11324), .Z(n11366) );
  XNOR U13245 ( .A(n11365), .B(n11366), .Z(n11371) );
  XOR U13246 ( .A(n11372), .B(n11371), .Z(n11350) );
  NANDN U13247 ( .A(n11327), .B(n11326), .Z(n11331) );
  NANDN U13248 ( .A(n11329), .B(n11328), .Z(n11330) );
  AND U13249 ( .A(n11331), .B(n11330), .Z(n11349) );
  XNOR U13250 ( .A(n11350), .B(n11349), .Z(n11351) );
  NANDN U13251 ( .A(n11333), .B(n11332), .Z(n11337) );
  NAND U13252 ( .A(n11335), .B(n11334), .Z(n11336) );
  NAND U13253 ( .A(n11337), .B(n11336), .Z(n11352) );
  XNOR U13254 ( .A(n11351), .B(n11352), .Z(n11343) );
  XNOR U13255 ( .A(n11344), .B(n11343), .Z(n11345) );
  XNOR U13256 ( .A(n11346), .B(n11345), .Z(n11375) );
  XNOR U13257 ( .A(sreg[1212]), .B(n11375), .Z(n11377) );
  NANDN U13258 ( .A(sreg[1211]), .B(n11338), .Z(n11342) );
  NAND U13259 ( .A(n11340), .B(n11339), .Z(n11341) );
  NAND U13260 ( .A(n11342), .B(n11341), .Z(n11376) );
  XNOR U13261 ( .A(n11377), .B(n11376), .Z(c[1212]) );
  NANDN U13262 ( .A(n11344), .B(n11343), .Z(n11348) );
  NANDN U13263 ( .A(n11346), .B(n11345), .Z(n11347) );
  AND U13264 ( .A(n11348), .B(n11347), .Z(n11383) );
  NANDN U13265 ( .A(n11350), .B(n11349), .Z(n11354) );
  NANDN U13266 ( .A(n11352), .B(n11351), .Z(n11353) );
  AND U13267 ( .A(n11354), .B(n11353), .Z(n11381) );
  NAND U13268 ( .A(n42143), .B(n11355), .Z(n11357) );
  XNOR U13269 ( .A(a[191]), .B(n4099), .Z(n11392) );
  NAND U13270 ( .A(n42144), .B(n11392), .Z(n11356) );
  AND U13271 ( .A(n11357), .B(n11356), .Z(n11407) );
  XOR U13272 ( .A(a[195]), .B(n42012), .Z(n11395) );
  XNOR U13273 ( .A(n11407), .B(n11406), .Z(n11409) );
  AND U13274 ( .A(a[197]), .B(b[0]), .Z(n11359) );
  XNOR U13275 ( .A(n11359), .B(n4071), .Z(n11361) );
  NANDN U13276 ( .A(b[0]), .B(a[196]), .Z(n11360) );
  NAND U13277 ( .A(n11361), .B(n11360), .Z(n11403) );
  XOR U13278 ( .A(a[193]), .B(n42085), .Z(n11396) );
  AND U13279 ( .A(a[189]), .B(b[7]), .Z(n11400) );
  XNOR U13280 ( .A(n11401), .B(n11400), .Z(n11402) );
  XNOR U13281 ( .A(n11403), .B(n11402), .Z(n11408) );
  XOR U13282 ( .A(n11409), .B(n11408), .Z(n11387) );
  NANDN U13283 ( .A(n11364), .B(n11363), .Z(n11368) );
  NANDN U13284 ( .A(n11366), .B(n11365), .Z(n11367) );
  AND U13285 ( .A(n11368), .B(n11367), .Z(n11386) );
  XNOR U13286 ( .A(n11387), .B(n11386), .Z(n11388) );
  NANDN U13287 ( .A(n11370), .B(n11369), .Z(n11374) );
  NAND U13288 ( .A(n11372), .B(n11371), .Z(n11373) );
  NAND U13289 ( .A(n11374), .B(n11373), .Z(n11389) );
  XNOR U13290 ( .A(n11388), .B(n11389), .Z(n11380) );
  XNOR U13291 ( .A(n11381), .B(n11380), .Z(n11382) );
  XNOR U13292 ( .A(n11383), .B(n11382), .Z(n11412) );
  XNOR U13293 ( .A(sreg[1213]), .B(n11412), .Z(n11414) );
  NANDN U13294 ( .A(sreg[1212]), .B(n11375), .Z(n11379) );
  NAND U13295 ( .A(n11377), .B(n11376), .Z(n11378) );
  NAND U13296 ( .A(n11379), .B(n11378), .Z(n11413) );
  XNOR U13297 ( .A(n11414), .B(n11413), .Z(c[1213]) );
  NANDN U13298 ( .A(n11381), .B(n11380), .Z(n11385) );
  NANDN U13299 ( .A(n11383), .B(n11382), .Z(n11384) );
  AND U13300 ( .A(n11385), .B(n11384), .Z(n11420) );
  NANDN U13301 ( .A(n11387), .B(n11386), .Z(n11391) );
  NANDN U13302 ( .A(n11389), .B(n11388), .Z(n11390) );
  AND U13303 ( .A(n11391), .B(n11390), .Z(n11418) );
  NAND U13304 ( .A(n42143), .B(n11392), .Z(n11394) );
  XNOR U13305 ( .A(a[192]), .B(n4099), .Z(n11429) );
  NAND U13306 ( .A(n42144), .B(n11429), .Z(n11393) );
  AND U13307 ( .A(n11394), .B(n11393), .Z(n11444) );
  XOR U13308 ( .A(a[196]), .B(n42012), .Z(n11432) );
  XNOR U13309 ( .A(n11444), .B(n11443), .Z(n11446) );
  XOR U13310 ( .A(a[194]), .B(n42085), .Z(n11433) );
  AND U13311 ( .A(a[190]), .B(b[7]), .Z(n11437) );
  XNOR U13312 ( .A(n11438), .B(n11437), .Z(n11439) );
  AND U13313 ( .A(a[198]), .B(b[0]), .Z(n11397) );
  XNOR U13314 ( .A(n11397), .B(n4071), .Z(n11399) );
  NANDN U13315 ( .A(b[0]), .B(a[197]), .Z(n11398) );
  NAND U13316 ( .A(n11399), .B(n11398), .Z(n11440) );
  XNOR U13317 ( .A(n11439), .B(n11440), .Z(n11445) );
  XOR U13318 ( .A(n11446), .B(n11445), .Z(n11424) );
  NANDN U13319 ( .A(n11401), .B(n11400), .Z(n11405) );
  NANDN U13320 ( .A(n11403), .B(n11402), .Z(n11404) );
  AND U13321 ( .A(n11405), .B(n11404), .Z(n11423) );
  XNOR U13322 ( .A(n11424), .B(n11423), .Z(n11425) );
  NANDN U13323 ( .A(n11407), .B(n11406), .Z(n11411) );
  NAND U13324 ( .A(n11409), .B(n11408), .Z(n11410) );
  NAND U13325 ( .A(n11411), .B(n11410), .Z(n11426) );
  XNOR U13326 ( .A(n11425), .B(n11426), .Z(n11417) );
  XNOR U13327 ( .A(n11418), .B(n11417), .Z(n11419) );
  XNOR U13328 ( .A(n11420), .B(n11419), .Z(n11449) );
  XNOR U13329 ( .A(sreg[1214]), .B(n11449), .Z(n11451) );
  NANDN U13330 ( .A(sreg[1213]), .B(n11412), .Z(n11416) );
  NAND U13331 ( .A(n11414), .B(n11413), .Z(n11415) );
  NAND U13332 ( .A(n11416), .B(n11415), .Z(n11450) );
  XNOR U13333 ( .A(n11451), .B(n11450), .Z(c[1214]) );
  NANDN U13334 ( .A(n11418), .B(n11417), .Z(n11422) );
  NANDN U13335 ( .A(n11420), .B(n11419), .Z(n11421) );
  AND U13336 ( .A(n11422), .B(n11421), .Z(n11457) );
  NANDN U13337 ( .A(n11424), .B(n11423), .Z(n11428) );
  NANDN U13338 ( .A(n11426), .B(n11425), .Z(n11427) );
  AND U13339 ( .A(n11428), .B(n11427), .Z(n11455) );
  NAND U13340 ( .A(n42143), .B(n11429), .Z(n11431) );
  XNOR U13341 ( .A(a[193]), .B(n4099), .Z(n11466) );
  NAND U13342 ( .A(n42144), .B(n11466), .Z(n11430) );
  AND U13343 ( .A(n11431), .B(n11430), .Z(n11481) );
  XOR U13344 ( .A(a[197]), .B(n42012), .Z(n11469) );
  XNOR U13345 ( .A(n11481), .B(n11480), .Z(n11483) );
  XOR U13346 ( .A(a[195]), .B(n42085), .Z(n11473) );
  AND U13347 ( .A(a[191]), .B(b[7]), .Z(n11474) );
  XNOR U13348 ( .A(n11475), .B(n11474), .Z(n11476) );
  AND U13349 ( .A(a[199]), .B(b[0]), .Z(n11434) );
  XNOR U13350 ( .A(n11434), .B(n4071), .Z(n11436) );
  NANDN U13351 ( .A(b[0]), .B(a[198]), .Z(n11435) );
  NAND U13352 ( .A(n11436), .B(n11435), .Z(n11477) );
  XNOR U13353 ( .A(n11476), .B(n11477), .Z(n11482) );
  XOR U13354 ( .A(n11483), .B(n11482), .Z(n11461) );
  NANDN U13355 ( .A(n11438), .B(n11437), .Z(n11442) );
  NANDN U13356 ( .A(n11440), .B(n11439), .Z(n11441) );
  AND U13357 ( .A(n11442), .B(n11441), .Z(n11460) );
  XNOR U13358 ( .A(n11461), .B(n11460), .Z(n11462) );
  NANDN U13359 ( .A(n11444), .B(n11443), .Z(n11448) );
  NAND U13360 ( .A(n11446), .B(n11445), .Z(n11447) );
  NAND U13361 ( .A(n11448), .B(n11447), .Z(n11463) );
  XNOR U13362 ( .A(n11462), .B(n11463), .Z(n11454) );
  XNOR U13363 ( .A(n11455), .B(n11454), .Z(n11456) );
  XNOR U13364 ( .A(n11457), .B(n11456), .Z(n11486) );
  XNOR U13365 ( .A(sreg[1215]), .B(n11486), .Z(n11488) );
  NANDN U13366 ( .A(sreg[1214]), .B(n11449), .Z(n11453) );
  NAND U13367 ( .A(n11451), .B(n11450), .Z(n11452) );
  NAND U13368 ( .A(n11453), .B(n11452), .Z(n11487) );
  XNOR U13369 ( .A(n11488), .B(n11487), .Z(c[1215]) );
  NANDN U13370 ( .A(n11455), .B(n11454), .Z(n11459) );
  NANDN U13371 ( .A(n11457), .B(n11456), .Z(n11458) );
  AND U13372 ( .A(n11459), .B(n11458), .Z(n11494) );
  NANDN U13373 ( .A(n11461), .B(n11460), .Z(n11465) );
  NANDN U13374 ( .A(n11463), .B(n11462), .Z(n11464) );
  AND U13375 ( .A(n11465), .B(n11464), .Z(n11492) );
  NAND U13376 ( .A(n42143), .B(n11466), .Z(n11468) );
  XNOR U13377 ( .A(a[194]), .B(n4099), .Z(n11503) );
  NAND U13378 ( .A(n42144), .B(n11503), .Z(n11467) );
  AND U13379 ( .A(n11468), .B(n11467), .Z(n11518) );
  XOR U13380 ( .A(a[198]), .B(n42012), .Z(n11506) );
  XNOR U13381 ( .A(n11518), .B(n11517), .Z(n11520) );
  AND U13382 ( .A(a[200]), .B(b[0]), .Z(n11470) );
  XNOR U13383 ( .A(n11470), .B(n4071), .Z(n11472) );
  NANDN U13384 ( .A(b[0]), .B(a[199]), .Z(n11471) );
  NAND U13385 ( .A(n11472), .B(n11471), .Z(n11514) );
  XOR U13386 ( .A(a[196]), .B(n42085), .Z(n11510) );
  AND U13387 ( .A(a[192]), .B(b[7]), .Z(n11511) );
  XNOR U13388 ( .A(n11512), .B(n11511), .Z(n11513) );
  XNOR U13389 ( .A(n11514), .B(n11513), .Z(n11519) );
  XOR U13390 ( .A(n11520), .B(n11519), .Z(n11498) );
  NANDN U13391 ( .A(n11475), .B(n11474), .Z(n11479) );
  NANDN U13392 ( .A(n11477), .B(n11476), .Z(n11478) );
  AND U13393 ( .A(n11479), .B(n11478), .Z(n11497) );
  XNOR U13394 ( .A(n11498), .B(n11497), .Z(n11499) );
  NANDN U13395 ( .A(n11481), .B(n11480), .Z(n11485) );
  NAND U13396 ( .A(n11483), .B(n11482), .Z(n11484) );
  NAND U13397 ( .A(n11485), .B(n11484), .Z(n11500) );
  XNOR U13398 ( .A(n11499), .B(n11500), .Z(n11491) );
  XNOR U13399 ( .A(n11492), .B(n11491), .Z(n11493) );
  XNOR U13400 ( .A(n11494), .B(n11493), .Z(n11523) );
  XNOR U13401 ( .A(sreg[1216]), .B(n11523), .Z(n11525) );
  NANDN U13402 ( .A(sreg[1215]), .B(n11486), .Z(n11490) );
  NAND U13403 ( .A(n11488), .B(n11487), .Z(n11489) );
  NAND U13404 ( .A(n11490), .B(n11489), .Z(n11524) );
  XNOR U13405 ( .A(n11525), .B(n11524), .Z(c[1216]) );
  NANDN U13406 ( .A(n11492), .B(n11491), .Z(n11496) );
  NANDN U13407 ( .A(n11494), .B(n11493), .Z(n11495) );
  AND U13408 ( .A(n11496), .B(n11495), .Z(n11531) );
  NANDN U13409 ( .A(n11498), .B(n11497), .Z(n11502) );
  NANDN U13410 ( .A(n11500), .B(n11499), .Z(n11501) );
  AND U13411 ( .A(n11502), .B(n11501), .Z(n11529) );
  NAND U13412 ( .A(n42143), .B(n11503), .Z(n11505) );
  XNOR U13413 ( .A(a[195]), .B(n4099), .Z(n11540) );
  NAND U13414 ( .A(n42144), .B(n11540), .Z(n11504) );
  AND U13415 ( .A(n11505), .B(n11504), .Z(n11555) );
  XOR U13416 ( .A(a[199]), .B(n42012), .Z(n11543) );
  XNOR U13417 ( .A(n11555), .B(n11554), .Z(n11557) );
  AND U13418 ( .A(a[201]), .B(b[0]), .Z(n11507) );
  XNOR U13419 ( .A(n11507), .B(n4071), .Z(n11509) );
  NANDN U13420 ( .A(b[0]), .B(a[200]), .Z(n11508) );
  NAND U13421 ( .A(n11509), .B(n11508), .Z(n11551) );
  XOR U13422 ( .A(a[197]), .B(n42085), .Z(n11547) );
  AND U13423 ( .A(a[193]), .B(b[7]), .Z(n11548) );
  XNOR U13424 ( .A(n11549), .B(n11548), .Z(n11550) );
  XNOR U13425 ( .A(n11551), .B(n11550), .Z(n11556) );
  XOR U13426 ( .A(n11557), .B(n11556), .Z(n11535) );
  NANDN U13427 ( .A(n11512), .B(n11511), .Z(n11516) );
  NANDN U13428 ( .A(n11514), .B(n11513), .Z(n11515) );
  AND U13429 ( .A(n11516), .B(n11515), .Z(n11534) );
  XNOR U13430 ( .A(n11535), .B(n11534), .Z(n11536) );
  NANDN U13431 ( .A(n11518), .B(n11517), .Z(n11522) );
  NAND U13432 ( .A(n11520), .B(n11519), .Z(n11521) );
  NAND U13433 ( .A(n11522), .B(n11521), .Z(n11537) );
  XNOR U13434 ( .A(n11536), .B(n11537), .Z(n11528) );
  XNOR U13435 ( .A(n11529), .B(n11528), .Z(n11530) );
  XNOR U13436 ( .A(n11531), .B(n11530), .Z(n11560) );
  XNOR U13437 ( .A(sreg[1217]), .B(n11560), .Z(n11562) );
  NANDN U13438 ( .A(sreg[1216]), .B(n11523), .Z(n11527) );
  NAND U13439 ( .A(n11525), .B(n11524), .Z(n11526) );
  NAND U13440 ( .A(n11527), .B(n11526), .Z(n11561) );
  XNOR U13441 ( .A(n11562), .B(n11561), .Z(c[1217]) );
  NANDN U13442 ( .A(n11529), .B(n11528), .Z(n11533) );
  NANDN U13443 ( .A(n11531), .B(n11530), .Z(n11532) );
  AND U13444 ( .A(n11533), .B(n11532), .Z(n11568) );
  NANDN U13445 ( .A(n11535), .B(n11534), .Z(n11539) );
  NANDN U13446 ( .A(n11537), .B(n11536), .Z(n11538) );
  AND U13447 ( .A(n11539), .B(n11538), .Z(n11566) );
  NAND U13448 ( .A(n42143), .B(n11540), .Z(n11542) );
  XNOR U13449 ( .A(a[196]), .B(n4099), .Z(n11577) );
  NAND U13450 ( .A(n42144), .B(n11577), .Z(n11541) );
  AND U13451 ( .A(n11542), .B(n11541), .Z(n11592) );
  XOR U13452 ( .A(a[200]), .B(n42012), .Z(n11580) );
  XNOR U13453 ( .A(n11592), .B(n11591), .Z(n11594) );
  AND U13454 ( .A(a[202]), .B(b[0]), .Z(n11544) );
  XNOR U13455 ( .A(n11544), .B(n4071), .Z(n11546) );
  NANDN U13456 ( .A(b[0]), .B(a[201]), .Z(n11545) );
  NAND U13457 ( .A(n11546), .B(n11545), .Z(n11588) );
  XOR U13458 ( .A(a[198]), .B(n42085), .Z(n11581) );
  AND U13459 ( .A(a[194]), .B(b[7]), .Z(n11585) );
  XNOR U13460 ( .A(n11586), .B(n11585), .Z(n11587) );
  XNOR U13461 ( .A(n11588), .B(n11587), .Z(n11593) );
  XOR U13462 ( .A(n11594), .B(n11593), .Z(n11572) );
  NANDN U13463 ( .A(n11549), .B(n11548), .Z(n11553) );
  NANDN U13464 ( .A(n11551), .B(n11550), .Z(n11552) );
  AND U13465 ( .A(n11553), .B(n11552), .Z(n11571) );
  XNOR U13466 ( .A(n11572), .B(n11571), .Z(n11573) );
  NANDN U13467 ( .A(n11555), .B(n11554), .Z(n11559) );
  NAND U13468 ( .A(n11557), .B(n11556), .Z(n11558) );
  NAND U13469 ( .A(n11559), .B(n11558), .Z(n11574) );
  XNOR U13470 ( .A(n11573), .B(n11574), .Z(n11565) );
  XNOR U13471 ( .A(n11566), .B(n11565), .Z(n11567) );
  XNOR U13472 ( .A(n11568), .B(n11567), .Z(n11597) );
  XNOR U13473 ( .A(sreg[1218]), .B(n11597), .Z(n11599) );
  NANDN U13474 ( .A(sreg[1217]), .B(n11560), .Z(n11564) );
  NAND U13475 ( .A(n11562), .B(n11561), .Z(n11563) );
  NAND U13476 ( .A(n11564), .B(n11563), .Z(n11598) );
  XNOR U13477 ( .A(n11599), .B(n11598), .Z(c[1218]) );
  NANDN U13478 ( .A(n11566), .B(n11565), .Z(n11570) );
  NANDN U13479 ( .A(n11568), .B(n11567), .Z(n11569) );
  AND U13480 ( .A(n11570), .B(n11569), .Z(n11605) );
  NANDN U13481 ( .A(n11572), .B(n11571), .Z(n11576) );
  NANDN U13482 ( .A(n11574), .B(n11573), .Z(n11575) );
  AND U13483 ( .A(n11576), .B(n11575), .Z(n11603) );
  NAND U13484 ( .A(n42143), .B(n11577), .Z(n11579) );
  XNOR U13485 ( .A(a[197]), .B(n4100), .Z(n11614) );
  NAND U13486 ( .A(n42144), .B(n11614), .Z(n11578) );
  AND U13487 ( .A(n11579), .B(n11578), .Z(n11629) );
  XOR U13488 ( .A(a[201]), .B(n42012), .Z(n11617) );
  XNOR U13489 ( .A(n11629), .B(n11628), .Z(n11631) );
  XOR U13490 ( .A(a[199]), .B(n42085), .Z(n11621) );
  AND U13491 ( .A(a[195]), .B(b[7]), .Z(n11622) );
  XNOR U13492 ( .A(n11623), .B(n11622), .Z(n11624) );
  AND U13493 ( .A(a[203]), .B(b[0]), .Z(n11582) );
  XNOR U13494 ( .A(n11582), .B(n4071), .Z(n11584) );
  NANDN U13495 ( .A(b[0]), .B(a[202]), .Z(n11583) );
  NAND U13496 ( .A(n11584), .B(n11583), .Z(n11625) );
  XNOR U13497 ( .A(n11624), .B(n11625), .Z(n11630) );
  XOR U13498 ( .A(n11631), .B(n11630), .Z(n11609) );
  NANDN U13499 ( .A(n11586), .B(n11585), .Z(n11590) );
  NANDN U13500 ( .A(n11588), .B(n11587), .Z(n11589) );
  AND U13501 ( .A(n11590), .B(n11589), .Z(n11608) );
  XNOR U13502 ( .A(n11609), .B(n11608), .Z(n11610) );
  NANDN U13503 ( .A(n11592), .B(n11591), .Z(n11596) );
  NAND U13504 ( .A(n11594), .B(n11593), .Z(n11595) );
  NAND U13505 ( .A(n11596), .B(n11595), .Z(n11611) );
  XNOR U13506 ( .A(n11610), .B(n11611), .Z(n11602) );
  XNOR U13507 ( .A(n11603), .B(n11602), .Z(n11604) );
  XNOR U13508 ( .A(n11605), .B(n11604), .Z(n11634) );
  XNOR U13509 ( .A(sreg[1219]), .B(n11634), .Z(n11636) );
  NANDN U13510 ( .A(sreg[1218]), .B(n11597), .Z(n11601) );
  NAND U13511 ( .A(n11599), .B(n11598), .Z(n11600) );
  NAND U13512 ( .A(n11601), .B(n11600), .Z(n11635) );
  XNOR U13513 ( .A(n11636), .B(n11635), .Z(c[1219]) );
  NANDN U13514 ( .A(n11603), .B(n11602), .Z(n11607) );
  NANDN U13515 ( .A(n11605), .B(n11604), .Z(n11606) );
  AND U13516 ( .A(n11607), .B(n11606), .Z(n11642) );
  NANDN U13517 ( .A(n11609), .B(n11608), .Z(n11613) );
  NANDN U13518 ( .A(n11611), .B(n11610), .Z(n11612) );
  AND U13519 ( .A(n11613), .B(n11612), .Z(n11640) );
  NAND U13520 ( .A(n42143), .B(n11614), .Z(n11616) );
  XNOR U13521 ( .A(a[198]), .B(n4100), .Z(n11651) );
  NAND U13522 ( .A(n42144), .B(n11651), .Z(n11615) );
  AND U13523 ( .A(n11616), .B(n11615), .Z(n11666) );
  XOR U13524 ( .A(a[202]), .B(n42012), .Z(n11654) );
  XNOR U13525 ( .A(n11666), .B(n11665), .Z(n11668) );
  AND U13526 ( .A(a[204]), .B(b[0]), .Z(n11618) );
  XNOR U13527 ( .A(n11618), .B(n4071), .Z(n11620) );
  NANDN U13528 ( .A(b[0]), .B(a[203]), .Z(n11619) );
  NAND U13529 ( .A(n11620), .B(n11619), .Z(n11662) );
  XOR U13530 ( .A(a[200]), .B(n42085), .Z(n11655) );
  AND U13531 ( .A(a[196]), .B(b[7]), .Z(n11659) );
  XNOR U13532 ( .A(n11660), .B(n11659), .Z(n11661) );
  XNOR U13533 ( .A(n11662), .B(n11661), .Z(n11667) );
  XOR U13534 ( .A(n11668), .B(n11667), .Z(n11646) );
  NANDN U13535 ( .A(n11623), .B(n11622), .Z(n11627) );
  NANDN U13536 ( .A(n11625), .B(n11624), .Z(n11626) );
  AND U13537 ( .A(n11627), .B(n11626), .Z(n11645) );
  XNOR U13538 ( .A(n11646), .B(n11645), .Z(n11647) );
  NANDN U13539 ( .A(n11629), .B(n11628), .Z(n11633) );
  NAND U13540 ( .A(n11631), .B(n11630), .Z(n11632) );
  NAND U13541 ( .A(n11633), .B(n11632), .Z(n11648) );
  XNOR U13542 ( .A(n11647), .B(n11648), .Z(n11639) );
  XNOR U13543 ( .A(n11640), .B(n11639), .Z(n11641) );
  XNOR U13544 ( .A(n11642), .B(n11641), .Z(n11671) );
  XNOR U13545 ( .A(sreg[1220]), .B(n11671), .Z(n11673) );
  NANDN U13546 ( .A(sreg[1219]), .B(n11634), .Z(n11638) );
  NAND U13547 ( .A(n11636), .B(n11635), .Z(n11637) );
  NAND U13548 ( .A(n11638), .B(n11637), .Z(n11672) );
  XNOR U13549 ( .A(n11673), .B(n11672), .Z(c[1220]) );
  NANDN U13550 ( .A(n11640), .B(n11639), .Z(n11644) );
  NANDN U13551 ( .A(n11642), .B(n11641), .Z(n11643) );
  AND U13552 ( .A(n11644), .B(n11643), .Z(n11679) );
  NANDN U13553 ( .A(n11646), .B(n11645), .Z(n11650) );
  NANDN U13554 ( .A(n11648), .B(n11647), .Z(n11649) );
  AND U13555 ( .A(n11650), .B(n11649), .Z(n11677) );
  NAND U13556 ( .A(n42143), .B(n11651), .Z(n11653) );
  XNOR U13557 ( .A(a[199]), .B(n4100), .Z(n11688) );
  NAND U13558 ( .A(n42144), .B(n11688), .Z(n11652) );
  AND U13559 ( .A(n11653), .B(n11652), .Z(n11703) );
  XOR U13560 ( .A(a[203]), .B(n42012), .Z(n11691) );
  XNOR U13561 ( .A(n11703), .B(n11702), .Z(n11705) );
  XOR U13562 ( .A(a[201]), .B(n42085), .Z(n11695) );
  AND U13563 ( .A(a[197]), .B(b[7]), .Z(n11696) );
  XNOR U13564 ( .A(n11697), .B(n11696), .Z(n11698) );
  AND U13565 ( .A(a[205]), .B(b[0]), .Z(n11656) );
  XNOR U13566 ( .A(n11656), .B(n4071), .Z(n11658) );
  NANDN U13567 ( .A(b[0]), .B(a[204]), .Z(n11657) );
  NAND U13568 ( .A(n11658), .B(n11657), .Z(n11699) );
  XNOR U13569 ( .A(n11698), .B(n11699), .Z(n11704) );
  XOR U13570 ( .A(n11705), .B(n11704), .Z(n11683) );
  NANDN U13571 ( .A(n11660), .B(n11659), .Z(n11664) );
  NANDN U13572 ( .A(n11662), .B(n11661), .Z(n11663) );
  AND U13573 ( .A(n11664), .B(n11663), .Z(n11682) );
  XNOR U13574 ( .A(n11683), .B(n11682), .Z(n11684) );
  NANDN U13575 ( .A(n11666), .B(n11665), .Z(n11670) );
  NAND U13576 ( .A(n11668), .B(n11667), .Z(n11669) );
  NAND U13577 ( .A(n11670), .B(n11669), .Z(n11685) );
  XNOR U13578 ( .A(n11684), .B(n11685), .Z(n11676) );
  XNOR U13579 ( .A(n11677), .B(n11676), .Z(n11678) );
  XNOR U13580 ( .A(n11679), .B(n11678), .Z(n11708) );
  XNOR U13581 ( .A(sreg[1221]), .B(n11708), .Z(n11710) );
  NANDN U13582 ( .A(sreg[1220]), .B(n11671), .Z(n11675) );
  NAND U13583 ( .A(n11673), .B(n11672), .Z(n11674) );
  NAND U13584 ( .A(n11675), .B(n11674), .Z(n11709) );
  XNOR U13585 ( .A(n11710), .B(n11709), .Z(c[1221]) );
  NANDN U13586 ( .A(n11677), .B(n11676), .Z(n11681) );
  NANDN U13587 ( .A(n11679), .B(n11678), .Z(n11680) );
  AND U13588 ( .A(n11681), .B(n11680), .Z(n11716) );
  NANDN U13589 ( .A(n11683), .B(n11682), .Z(n11687) );
  NANDN U13590 ( .A(n11685), .B(n11684), .Z(n11686) );
  AND U13591 ( .A(n11687), .B(n11686), .Z(n11714) );
  NAND U13592 ( .A(n42143), .B(n11688), .Z(n11690) );
  XNOR U13593 ( .A(a[200]), .B(n4100), .Z(n11725) );
  NAND U13594 ( .A(n42144), .B(n11725), .Z(n11689) );
  AND U13595 ( .A(n11690), .B(n11689), .Z(n11740) );
  XOR U13596 ( .A(a[204]), .B(n42012), .Z(n11728) );
  XNOR U13597 ( .A(n11740), .B(n11739), .Z(n11742) );
  AND U13598 ( .A(b[0]), .B(a[206]), .Z(n11692) );
  XOR U13599 ( .A(b[1]), .B(n11692), .Z(n11694) );
  NANDN U13600 ( .A(b[0]), .B(a[205]), .Z(n11693) );
  AND U13601 ( .A(n11694), .B(n11693), .Z(n11735) );
  XOR U13602 ( .A(a[202]), .B(n42085), .Z(n11732) );
  AND U13603 ( .A(a[198]), .B(b[7]), .Z(n11733) );
  XOR U13604 ( .A(n11734), .B(n11733), .Z(n11736) );
  XNOR U13605 ( .A(n11735), .B(n11736), .Z(n11741) );
  XOR U13606 ( .A(n11742), .B(n11741), .Z(n11720) );
  NANDN U13607 ( .A(n11697), .B(n11696), .Z(n11701) );
  NANDN U13608 ( .A(n11699), .B(n11698), .Z(n11700) );
  AND U13609 ( .A(n11701), .B(n11700), .Z(n11719) );
  XNOR U13610 ( .A(n11720), .B(n11719), .Z(n11721) );
  NANDN U13611 ( .A(n11703), .B(n11702), .Z(n11707) );
  NAND U13612 ( .A(n11705), .B(n11704), .Z(n11706) );
  NAND U13613 ( .A(n11707), .B(n11706), .Z(n11722) );
  XNOR U13614 ( .A(n11721), .B(n11722), .Z(n11713) );
  XNOR U13615 ( .A(n11714), .B(n11713), .Z(n11715) );
  XNOR U13616 ( .A(n11716), .B(n11715), .Z(n11745) );
  XNOR U13617 ( .A(sreg[1222]), .B(n11745), .Z(n11747) );
  NANDN U13618 ( .A(sreg[1221]), .B(n11708), .Z(n11712) );
  NAND U13619 ( .A(n11710), .B(n11709), .Z(n11711) );
  NAND U13620 ( .A(n11712), .B(n11711), .Z(n11746) );
  XNOR U13621 ( .A(n11747), .B(n11746), .Z(c[1222]) );
  NANDN U13622 ( .A(n11714), .B(n11713), .Z(n11718) );
  NANDN U13623 ( .A(n11716), .B(n11715), .Z(n11717) );
  AND U13624 ( .A(n11718), .B(n11717), .Z(n11753) );
  NANDN U13625 ( .A(n11720), .B(n11719), .Z(n11724) );
  NANDN U13626 ( .A(n11722), .B(n11721), .Z(n11723) );
  AND U13627 ( .A(n11724), .B(n11723), .Z(n11751) );
  NAND U13628 ( .A(n42143), .B(n11725), .Z(n11727) );
  XNOR U13629 ( .A(a[201]), .B(n4100), .Z(n11762) );
  NAND U13630 ( .A(n42144), .B(n11762), .Z(n11726) );
  AND U13631 ( .A(n11727), .B(n11726), .Z(n11777) );
  XOR U13632 ( .A(a[205]), .B(n42012), .Z(n11765) );
  XNOR U13633 ( .A(n11777), .B(n11776), .Z(n11779) );
  AND U13634 ( .A(a[207]), .B(b[0]), .Z(n11729) );
  XNOR U13635 ( .A(n11729), .B(n4071), .Z(n11731) );
  NANDN U13636 ( .A(b[0]), .B(a[206]), .Z(n11730) );
  NAND U13637 ( .A(n11731), .B(n11730), .Z(n11773) );
  XOR U13638 ( .A(a[203]), .B(n42085), .Z(n11769) );
  AND U13639 ( .A(a[199]), .B(b[7]), .Z(n11770) );
  XNOR U13640 ( .A(n11771), .B(n11770), .Z(n11772) );
  XNOR U13641 ( .A(n11773), .B(n11772), .Z(n11778) );
  XOR U13642 ( .A(n11779), .B(n11778), .Z(n11757) );
  NANDN U13643 ( .A(n11734), .B(n11733), .Z(n11738) );
  NANDN U13644 ( .A(n11736), .B(n11735), .Z(n11737) );
  AND U13645 ( .A(n11738), .B(n11737), .Z(n11756) );
  XNOR U13646 ( .A(n11757), .B(n11756), .Z(n11758) );
  NANDN U13647 ( .A(n11740), .B(n11739), .Z(n11744) );
  NAND U13648 ( .A(n11742), .B(n11741), .Z(n11743) );
  NAND U13649 ( .A(n11744), .B(n11743), .Z(n11759) );
  XNOR U13650 ( .A(n11758), .B(n11759), .Z(n11750) );
  XNOR U13651 ( .A(n11751), .B(n11750), .Z(n11752) );
  XNOR U13652 ( .A(n11753), .B(n11752), .Z(n11782) );
  XNOR U13653 ( .A(sreg[1223]), .B(n11782), .Z(n11784) );
  NANDN U13654 ( .A(sreg[1222]), .B(n11745), .Z(n11749) );
  NAND U13655 ( .A(n11747), .B(n11746), .Z(n11748) );
  NAND U13656 ( .A(n11749), .B(n11748), .Z(n11783) );
  XNOR U13657 ( .A(n11784), .B(n11783), .Z(c[1223]) );
  NANDN U13658 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U13659 ( .A(n11753), .B(n11752), .Z(n11754) );
  AND U13660 ( .A(n11755), .B(n11754), .Z(n11790) );
  NANDN U13661 ( .A(n11757), .B(n11756), .Z(n11761) );
  NANDN U13662 ( .A(n11759), .B(n11758), .Z(n11760) );
  AND U13663 ( .A(n11761), .B(n11760), .Z(n11788) );
  NAND U13664 ( .A(n42143), .B(n11762), .Z(n11764) );
  XNOR U13665 ( .A(a[202]), .B(n4100), .Z(n11799) );
  NAND U13666 ( .A(n42144), .B(n11799), .Z(n11763) );
  AND U13667 ( .A(n11764), .B(n11763), .Z(n11814) );
  XOR U13668 ( .A(a[206]), .B(n42012), .Z(n11802) );
  XNOR U13669 ( .A(n11814), .B(n11813), .Z(n11816) );
  AND U13670 ( .A(a[208]), .B(b[0]), .Z(n11766) );
  XNOR U13671 ( .A(n11766), .B(n4071), .Z(n11768) );
  NANDN U13672 ( .A(b[0]), .B(a[207]), .Z(n11767) );
  NAND U13673 ( .A(n11768), .B(n11767), .Z(n11810) );
  XOR U13674 ( .A(a[204]), .B(n42085), .Z(n11803) );
  AND U13675 ( .A(a[200]), .B(b[7]), .Z(n11807) );
  XNOR U13676 ( .A(n11808), .B(n11807), .Z(n11809) );
  XNOR U13677 ( .A(n11810), .B(n11809), .Z(n11815) );
  XOR U13678 ( .A(n11816), .B(n11815), .Z(n11794) );
  NANDN U13679 ( .A(n11771), .B(n11770), .Z(n11775) );
  NANDN U13680 ( .A(n11773), .B(n11772), .Z(n11774) );
  AND U13681 ( .A(n11775), .B(n11774), .Z(n11793) );
  XNOR U13682 ( .A(n11794), .B(n11793), .Z(n11795) );
  NANDN U13683 ( .A(n11777), .B(n11776), .Z(n11781) );
  NAND U13684 ( .A(n11779), .B(n11778), .Z(n11780) );
  NAND U13685 ( .A(n11781), .B(n11780), .Z(n11796) );
  XNOR U13686 ( .A(n11795), .B(n11796), .Z(n11787) );
  XNOR U13687 ( .A(n11788), .B(n11787), .Z(n11789) );
  XNOR U13688 ( .A(n11790), .B(n11789), .Z(n11819) );
  XNOR U13689 ( .A(sreg[1224]), .B(n11819), .Z(n11821) );
  NANDN U13690 ( .A(sreg[1223]), .B(n11782), .Z(n11786) );
  NAND U13691 ( .A(n11784), .B(n11783), .Z(n11785) );
  NAND U13692 ( .A(n11786), .B(n11785), .Z(n11820) );
  XNOR U13693 ( .A(n11821), .B(n11820), .Z(c[1224]) );
  NANDN U13694 ( .A(n11788), .B(n11787), .Z(n11792) );
  NANDN U13695 ( .A(n11790), .B(n11789), .Z(n11791) );
  AND U13696 ( .A(n11792), .B(n11791), .Z(n11827) );
  NANDN U13697 ( .A(n11794), .B(n11793), .Z(n11798) );
  NANDN U13698 ( .A(n11796), .B(n11795), .Z(n11797) );
  AND U13699 ( .A(n11798), .B(n11797), .Z(n11825) );
  NAND U13700 ( .A(n42143), .B(n11799), .Z(n11801) );
  XNOR U13701 ( .A(a[203]), .B(n4100), .Z(n11836) );
  NAND U13702 ( .A(n42144), .B(n11836), .Z(n11800) );
  AND U13703 ( .A(n11801), .B(n11800), .Z(n11851) );
  XOR U13704 ( .A(a[207]), .B(n42012), .Z(n11839) );
  XNOR U13705 ( .A(n11851), .B(n11850), .Z(n11853) );
  XOR U13706 ( .A(a[205]), .B(n42085), .Z(n11843) );
  AND U13707 ( .A(a[201]), .B(b[7]), .Z(n11844) );
  XNOR U13708 ( .A(n11845), .B(n11844), .Z(n11846) );
  AND U13709 ( .A(a[209]), .B(b[0]), .Z(n11804) );
  XNOR U13710 ( .A(n11804), .B(n4071), .Z(n11806) );
  NANDN U13711 ( .A(b[0]), .B(a[208]), .Z(n11805) );
  NAND U13712 ( .A(n11806), .B(n11805), .Z(n11847) );
  XNOR U13713 ( .A(n11846), .B(n11847), .Z(n11852) );
  XOR U13714 ( .A(n11853), .B(n11852), .Z(n11831) );
  NANDN U13715 ( .A(n11808), .B(n11807), .Z(n11812) );
  NANDN U13716 ( .A(n11810), .B(n11809), .Z(n11811) );
  AND U13717 ( .A(n11812), .B(n11811), .Z(n11830) );
  XNOR U13718 ( .A(n11831), .B(n11830), .Z(n11832) );
  NANDN U13719 ( .A(n11814), .B(n11813), .Z(n11818) );
  NAND U13720 ( .A(n11816), .B(n11815), .Z(n11817) );
  NAND U13721 ( .A(n11818), .B(n11817), .Z(n11833) );
  XNOR U13722 ( .A(n11832), .B(n11833), .Z(n11824) );
  XNOR U13723 ( .A(n11825), .B(n11824), .Z(n11826) );
  XNOR U13724 ( .A(n11827), .B(n11826), .Z(n11856) );
  XNOR U13725 ( .A(sreg[1225]), .B(n11856), .Z(n11858) );
  NANDN U13726 ( .A(sreg[1224]), .B(n11819), .Z(n11823) );
  NAND U13727 ( .A(n11821), .B(n11820), .Z(n11822) );
  NAND U13728 ( .A(n11823), .B(n11822), .Z(n11857) );
  XNOR U13729 ( .A(n11858), .B(n11857), .Z(c[1225]) );
  NANDN U13730 ( .A(n11825), .B(n11824), .Z(n11829) );
  NANDN U13731 ( .A(n11827), .B(n11826), .Z(n11828) );
  AND U13732 ( .A(n11829), .B(n11828), .Z(n11864) );
  NANDN U13733 ( .A(n11831), .B(n11830), .Z(n11835) );
  NANDN U13734 ( .A(n11833), .B(n11832), .Z(n11834) );
  AND U13735 ( .A(n11835), .B(n11834), .Z(n11862) );
  NAND U13736 ( .A(n42143), .B(n11836), .Z(n11838) );
  XNOR U13737 ( .A(a[204]), .B(n4101), .Z(n11873) );
  NAND U13738 ( .A(n42144), .B(n11873), .Z(n11837) );
  AND U13739 ( .A(n11838), .B(n11837), .Z(n11888) );
  XOR U13740 ( .A(a[208]), .B(n42012), .Z(n11876) );
  XNOR U13741 ( .A(n11888), .B(n11887), .Z(n11890) );
  AND U13742 ( .A(a[210]), .B(b[0]), .Z(n11840) );
  XNOR U13743 ( .A(n11840), .B(n4071), .Z(n11842) );
  NANDN U13744 ( .A(b[0]), .B(a[209]), .Z(n11841) );
  NAND U13745 ( .A(n11842), .B(n11841), .Z(n11884) );
  XOR U13746 ( .A(a[206]), .B(n42085), .Z(n11880) );
  AND U13747 ( .A(a[202]), .B(b[7]), .Z(n11881) );
  XNOR U13748 ( .A(n11882), .B(n11881), .Z(n11883) );
  XNOR U13749 ( .A(n11884), .B(n11883), .Z(n11889) );
  XOR U13750 ( .A(n11890), .B(n11889), .Z(n11868) );
  NANDN U13751 ( .A(n11845), .B(n11844), .Z(n11849) );
  NANDN U13752 ( .A(n11847), .B(n11846), .Z(n11848) );
  AND U13753 ( .A(n11849), .B(n11848), .Z(n11867) );
  XNOR U13754 ( .A(n11868), .B(n11867), .Z(n11869) );
  NANDN U13755 ( .A(n11851), .B(n11850), .Z(n11855) );
  NAND U13756 ( .A(n11853), .B(n11852), .Z(n11854) );
  NAND U13757 ( .A(n11855), .B(n11854), .Z(n11870) );
  XNOR U13758 ( .A(n11869), .B(n11870), .Z(n11861) );
  XNOR U13759 ( .A(n11862), .B(n11861), .Z(n11863) );
  XNOR U13760 ( .A(n11864), .B(n11863), .Z(n11893) );
  XNOR U13761 ( .A(sreg[1226]), .B(n11893), .Z(n11895) );
  NANDN U13762 ( .A(sreg[1225]), .B(n11856), .Z(n11860) );
  NAND U13763 ( .A(n11858), .B(n11857), .Z(n11859) );
  NAND U13764 ( .A(n11860), .B(n11859), .Z(n11894) );
  XNOR U13765 ( .A(n11895), .B(n11894), .Z(c[1226]) );
  NANDN U13766 ( .A(n11862), .B(n11861), .Z(n11866) );
  NANDN U13767 ( .A(n11864), .B(n11863), .Z(n11865) );
  AND U13768 ( .A(n11866), .B(n11865), .Z(n11901) );
  NANDN U13769 ( .A(n11868), .B(n11867), .Z(n11872) );
  NANDN U13770 ( .A(n11870), .B(n11869), .Z(n11871) );
  AND U13771 ( .A(n11872), .B(n11871), .Z(n11899) );
  NAND U13772 ( .A(n42143), .B(n11873), .Z(n11875) );
  XNOR U13773 ( .A(a[205]), .B(n4101), .Z(n11910) );
  NAND U13774 ( .A(n42144), .B(n11910), .Z(n11874) );
  AND U13775 ( .A(n11875), .B(n11874), .Z(n11925) );
  XOR U13776 ( .A(a[209]), .B(n42012), .Z(n11913) );
  XNOR U13777 ( .A(n11925), .B(n11924), .Z(n11927) );
  AND U13778 ( .A(a[211]), .B(b[0]), .Z(n11877) );
  XNOR U13779 ( .A(n11877), .B(n4071), .Z(n11879) );
  NANDN U13780 ( .A(b[0]), .B(a[210]), .Z(n11878) );
  NAND U13781 ( .A(n11879), .B(n11878), .Z(n11921) );
  XOR U13782 ( .A(a[207]), .B(n42085), .Z(n11917) );
  AND U13783 ( .A(a[203]), .B(b[7]), .Z(n11918) );
  XNOR U13784 ( .A(n11919), .B(n11918), .Z(n11920) );
  XNOR U13785 ( .A(n11921), .B(n11920), .Z(n11926) );
  XOR U13786 ( .A(n11927), .B(n11926), .Z(n11905) );
  NANDN U13787 ( .A(n11882), .B(n11881), .Z(n11886) );
  NANDN U13788 ( .A(n11884), .B(n11883), .Z(n11885) );
  AND U13789 ( .A(n11886), .B(n11885), .Z(n11904) );
  XNOR U13790 ( .A(n11905), .B(n11904), .Z(n11906) );
  NANDN U13791 ( .A(n11888), .B(n11887), .Z(n11892) );
  NAND U13792 ( .A(n11890), .B(n11889), .Z(n11891) );
  NAND U13793 ( .A(n11892), .B(n11891), .Z(n11907) );
  XNOR U13794 ( .A(n11906), .B(n11907), .Z(n11898) );
  XNOR U13795 ( .A(n11899), .B(n11898), .Z(n11900) );
  XNOR U13796 ( .A(n11901), .B(n11900), .Z(n11930) );
  XNOR U13797 ( .A(sreg[1227]), .B(n11930), .Z(n11932) );
  NANDN U13798 ( .A(sreg[1226]), .B(n11893), .Z(n11897) );
  NAND U13799 ( .A(n11895), .B(n11894), .Z(n11896) );
  NAND U13800 ( .A(n11897), .B(n11896), .Z(n11931) );
  XNOR U13801 ( .A(n11932), .B(n11931), .Z(c[1227]) );
  NANDN U13802 ( .A(n11899), .B(n11898), .Z(n11903) );
  NANDN U13803 ( .A(n11901), .B(n11900), .Z(n11902) );
  AND U13804 ( .A(n11903), .B(n11902), .Z(n11938) );
  NANDN U13805 ( .A(n11905), .B(n11904), .Z(n11909) );
  NANDN U13806 ( .A(n11907), .B(n11906), .Z(n11908) );
  AND U13807 ( .A(n11909), .B(n11908), .Z(n11936) );
  NAND U13808 ( .A(n42143), .B(n11910), .Z(n11912) );
  XNOR U13809 ( .A(a[206]), .B(n4101), .Z(n11947) );
  NAND U13810 ( .A(n42144), .B(n11947), .Z(n11911) );
  AND U13811 ( .A(n11912), .B(n11911), .Z(n11962) );
  XOR U13812 ( .A(a[210]), .B(n42012), .Z(n11950) );
  XNOR U13813 ( .A(n11962), .B(n11961), .Z(n11964) );
  AND U13814 ( .A(a[212]), .B(b[0]), .Z(n11914) );
  XNOR U13815 ( .A(n11914), .B(n4071), .Z(n11916) );
  NANDN U13816 ( .A(b[0]), .B(a[211]), .Z(n11915) );
  NAND U13817 ( .A(n11916), .B(n11915), .Z(n11958) );
  XOR U13818 ( .A(a[208]), .B(n42085), .Z(n11954) );
  AND U13819 ( .A(a[204]), .B(b[7]), .Z(n11955) );
  XNOR U13820 ( .A(n11956), .B(n11955), .Z(n11957) );
  XNOR U13821 ( .A(n11958), .B(n11957), .Z(n11963) );
  XOR U13822 ( .A(n11964), .B(n11963), .Z(n11942) );
  NANDN U13823 ( .A(n11919), .B(n11918), .Z(n11923) );
  NANDN U13824 ( .A(n11921), .B(n11920), .Z(n11922) );
  AND U13825 ( .A(n11923), .B(n11922), .Z(n11941) );
  XNOR U13826 ( .A(n11942), .B(n11941), .Z(n11943) );
  NANDN U13827 ( .A(n11925), .B(n11924), .Z(n11929) );
  NAND U13828 ( .A(n11927), .B(n11926), .Z(n11928) );
  NAND U13829 ( .A(n11929), .B(n11928), .Z(n11944) );
  XNOR U13830 ( .A(n11943), .B(n11944), .Z(n11935) );
  XNOR U13831 ( .A(n11936), .B(n11935), .Z(n11937) );
  XNOR U13832 ( .A(n11938), .B(n11937), .Z(n11967) );
  XNOR U13833 ( .A(sreg[1228]), .B(n11967), .Z(n11969) );
  NANDN U13834 ( .A(sreg[1227]), .B(n11930), .Z(n11934) );
  NAND U13835 ( .A(n11932), .B(n11931), .Z(n11933) );
  NAND U13836 ( .A(n11934), .B(n11933), .Z(n11968) );
  XNOR U13837 ( .A(n11969), .B(n11968), .Z(c[1228]) );
  NANDN U13838 ( .A(n11936), .B(n11935), .Z(n11940) );
  NANDN U13839 ( .A(n11938), .B(n11937), .Z(n11939) );
  AND U13840 ( .A(n11940), .B(n11939), .Z(n11975) );
  NANDN U13841 ( .A(n11942), .B(n11941), .Z(n11946) );
  NANDN U13842 ( .A(n11944), .B(n11943), .Z(n11945) );
  AND U13843 ( .A(n11946), .B(n11945), .Z(n11973) );
  NAND U13844 ( .A(n42143), .B(n11947), .Z(n11949) );
  XNOR U13845 ( .A(a[207]), .B(n4101), .Z(n11984) );
  NAND U13846 ( .A(n42144), .B(n11984), .Z(n11948) );
  AND U13847 ( .A(n11949), .B(n11948), .Z(n11999) );
  XOR U13848 ( .A(a[211]), .B(n42012), .Z(n11987) );
  XNOR U13849 ( .A(n11999), .B(n11998), .Z(n12001) );
  AND U13850 ( .A(a[213]), .B(b[0]), .Z(n11951) );
  XNOR U13851 ( .A(n11951), .B(n4071), .Z(n11953) );
  NANDN U13852 ( .A(b[0]), .B(a[212]), .Z(n11952) );
  NAND U13853 ( .A(n11953), .B(n11952), .Z(n11995) );
  XOR U13854 ( .A(a[209]), .B(n42085), .Z(n11991) );
  AND U13855 ( .A(a[205]), .B(b[7]), .Z(n11992) );
  XNOR U13856 ( .A(n11993), .B(n11992), .Z(n11994) );
  XNOR U13857 ( .A(n11995), .B(n11994), .Z(n12000) );
  XOR U13858 ( .A(n12001), .B(n12000), .Z(n11979) );
  NANDN U13859 ( .A(n11956), .B(n11955), .Z(n11960) );
  NANDN U13860 ( .A(n11958), .B(n11957), .Z(n11959) );
  AND U13861 ( .A(n11960), .B(n11959), .Z(n11978) );
  XNOR U13862 ( .A(n11979), .B(n11978), .Z(n11980) );
  NANDN U13863 ( .A(n11962), .B(n11961), .Z(n11966) );
  NAND U13864 ( .A(n11964), .B(n11963), .Z(n11965) );
  NAND U13865 ( .A(n11966), .B(n11965), .Z(n11981) );
  XNOR U13866 ( .A(n11980), .B(n11981), .Z(n11972) );
  XNOR U13867 ( .A(n11973), .B(n11972), .Z(n11974) );
  XNOR U13868 ( .A(n11975), .B(n11974), .Z(n12004) );
  XNOR U13869 ( .A(sreg[1229]), .B(n12004), .Z(n12006) );
  NANDN U13870 ( .A(sreg[1228]), .B(n11967), .Z(n11971) );
  NAND U13871 ( .A(n11969), .B(n11968), .Z(n11970) );
  NAND U13872 ( .A(n11971), .B(n11970), .Z(n12005) );
  XNOR U13873 ( .A(n12006), .B(n12005), .Z(c[1229]) );
  NANDN U13874 ( .A(n11973), .B(n11972), .Z(n11977) );
  NANDN U13875 ( .A(n11975), .B(n11974), .Z(n11976) );
  AND U13876 ( .A(n11977), .B(n11976), .Z(n12012) );
  NANDN U13877 ( .A(n11979), .B(n11978), .Z(n11983) );
  NANDN U13878 ( .A(n11981), .B(n11980), .Z(n11982) );
  AND U13879 ( .A(n11983), .B(n11982), .Z(n12010) );
  NAND U13880 ( .A(n42143), .B(n11984), .Z(n11986) );
  XNOR U13881 ( .A(a[208]), .B(n4101), .Z(n12021) );
  NAND U13882 ( .A(n42144), .B(n12021), .Z(n11985) );
  AND U13883 ( .A(n11986), .B(n11985), .Z(n12036) );
  XOR U13884 ( .A(a[212]), .B(n42012), .Z(n12024) );
  XNOR U13885 ( .A(n12036), .B(n12035), .Z(n12038) );
  AND U13886 ( .A(a[214]), .B(b[0]), .Z(n11988) );
  XNOR U13887 ( .A(n11988), .B(n4071), .Z(n11990) );
  NANDN U13888 ( .A(b[0]), .B(a[213]), .Z(n11989) );
  NAND U13889 ( .A(n11990), .B(n11989), .Z(n12032) );
  XOR U13890 ( .A(a[210]), .B(n42085), .Z(n12025) );
  AND U13891 ( .A(a[206]), .B(b[7]), .Z(n12029) );
  XNOR U13892 ( .A(n12030), .B(n12029), .Z(n12031) );
  XNOR U13893 ( .A(n12032), .B(n12031), .Z(n12037) );
  XOR U13894 ( .A(n12038), .B(n12037), .Z(n12016) );
  NANDN U13895 ( .A(n11993), .B(n11992), .Z(n11997) );
  NANDN U13896 ( .A(n11995), .B(n11994), .Z(n11996) );
  AND U13897 ( .A(n11997), .B(n11996), .Z(n12015) );
  XNOR U13898 ( .A(n12016), .B(n12015), .Z(n12017) );
  NANDN U13899 ( .A(n11999), .B(n11998), .Z(n12003) );
  NAND U13900 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U13901 ( .A(n12003), .B(n12002), .Z(n12018) );
  XNOR U13902 ( .A(n12017), .B(n12018), .Z(n12009) );
  XNOR U13903 ( .A(n12010), .B(n12009), .Z(n12011) );
  XNOR U13904 ( .A(n12012), .B(n12011), .Z(n12041) );
  XNOR U13905 ( .A(sreg[1230]), .B(n12041), .Z(n12043) );
  NANDN U13906 ( .A(sreg[1229]), .B(n12004), .Z(n12008) );
  NAND U13907 ( .A(n12006), .B(n12005), .Z(n12007) );
  NAND U13908 ( .A(n12008), .B(n12007), .Z(n12042) );
  XNOR U13909 ( .A(n12043), .B(n12042), .Z(c[1230]) );
  NANDN U13910 ( .A(n12010), .B(n12009), .Z(n12014) );
  NANDN U13911 ( .A(n12012), .B(n12011), .Z(n12013) );
  AND U13912 ( .A(n12014), .B(n12013), .Z(n12049) );
  NANDN U13913 ( .A(n12016), .B(n12015), .Z(n12020) );
  NANDN U13914 ( .A(n12018), .B(n12017), .Z(n12019) );
  AND U13915 ( .A(n12020), .B(n12019), .Z(n12047) );
  NAND U13916 ( .A(n42143), .B(n12021), .Z(n12023) );
  XNOR U13917 ( .A(a[209]), .B(n4101), .Z(n12058) );
  NAND U13918 ( .A(n42144), .B(n12058), .Z(n12022) );
  AND U13919 ( .A(n12023), .B(n12022), .Z(n12073) );
  XOR U13920 ( .A(a[213]), .B(n42012), .Z(n12061) );
  XNOR U13921 ( .A(n12073), .B(n12072), .Z(n12075) );
  XOR U13922 ( .A(a[211]), .B(n42085), .Z(n12065) );
  AND U13923 ( .A(a[207]), .B(b[7]), .Z(n12066) );
  XNOR U13924 ( .A(n12067), .B(n12066), .Z(n12068) );
  AND U13925 ( .A(a[215]), .B(b[0]), .Z(n12026) );
  XNOR U13926 ( .A(n12026), .B(n4071), .Z(n12028) );
  NANDN U13927 ( .A(b[0]), .B(a[214]), .Z(n12027) );
  NAND U13928 ( .A(n12028), .B(n12027), .Z(n12069) );
  XNOR U13929 ( .A(n12068), .B(n12069), .Z(n12074) );
  XOR U13930 ( .A(n12075), .B(n12074), .Z(n12053) );
  NANDN U13931 ( .A(n12030), .B(n12029), .Z(n12034) );
  NANDN U13932 ( .A(n12032), .B(n12031), .Z(n12033) );
  AND U13933 ( .A(n12034), .B(n12033), .Z(n12052) );
  XNOR U13934 ( .A(n12053), .B(n12052), .Z(n12054) );
  NANDN U13935 ( .A(n12036), .B(n12035), .Z(n12040) );
  NAND U13936 ( .A(n12038), .B(n12037), .Z(n12039) );
  NAND U13937 ( .A(n12040), .B(n12039), .Z(n12055) );
  XNOR U13938 ( .A(n12054), .B(n12055), .Z(n12046) );
  XNOR U13939 ( .A(n12047), .B(n12046), .Z(n12048) );
  XNOR U13940 ( .A(n12049), .B(n12048), .Z(n12078) );
  XNOR U13941 ( .A(sreg[1231]), .B(n12078), .Z(n12080) );
  NANDN U13942 ( .A(sreg[1230]), .B(n12041), .Z(n12045) );
  NAND U13943 ( .A(n12043), .B(n12042), .Z(n12044) );
  NAND U13944 ( .A(n12045), .B(n12044), .Z(n12079) );
  XNOR U13945 ( .A(n12080), .B(n12079), .Z(c[1231]) );
  NANDN U13946 ( .A(n12047), .B(n12046), .Z(n12051) );
  NANDN U13947 ( .A(n12049), .B(n12048), .Z(n12050) );
  AND U13948 ( .A(n12051), .B(n12050), .Z(n12086) );
  NANDN U13949 ( .A(n12053), .B(n12052), .Z(n12057) );
  NANDN U13950 ( .A(n12055), .B(n12054), .Z(n12056) );
  AND U13951 ( .A(n12057), .B(n12056), .Z(n12084) );
  NAND U13952 ( .A(n42143), .B(n12058), .Z(n12060) );
  XNOR U13953 ( .A(a[210]), .B(n4101), .Z(n12095) );
  NAND U13954 ( .A(n42144), .B(n12095), .Z(n12059) );
  AND U13955 ( .A(n12060), .B(n12059), .Z(n12110) );
  XOR U13956 ( .A(a[214]), .B(n42012), .Z(n12098) );
  XNOR U13957 ( .A(n12110), .B(n12109), .Z(n12112) );
  AND U13958 ( .A(a[216]), .B(b[0]), .Z(n12062) );
  XNOR U13959 ( .A(n12062), .B(n4071), .Z(n12064) );
  NANDN U13960 ( .A(b[0]), .B(a[215]), .Z(n12063) );
  NAND U13961 ( .A(n12064), .B(n12063), .Z(n12106) );
  XOR U13962 ( .A(a[212]), .B(n42085), .Z(n12099) );
  AND U13963 ( .A(a[208]), .B(b[7]), .Z(n12103) );
  XNOR U13964 ( .A(n12104), .B(n12103), .Z(n12105) );
  XNOR U13965 ( .A(n12106), .B(n12105), .Z(n12111) );
  XOR U13966 ( .A(n12112), .B(n12111), .Z(n12090) );
  NANDN U13967 ( .A(n12067), .B(n12066), .Z(n12071) );
  NANDN U13968 ( .A(n12069), .B(n12068), .Z(n12070) );
  AND U13969 ( .A(n12071), .B(n12070), .Z(n12089) );
  XNOR U13970 ( .A(n12090), .B(n12089), .Z(n12091) );
  NANDN U13971 ( .A(n12073), .B(n12072), .Z(n12077) );
  NAND U13972 ( .A(n12075), .B(n12074), .Z(n12076) );
  NAND U13973 ( .A(n12077), .B(n12076), .Z(n12092) );
  XNOR U13974 ( .A(n12091), .B(n12092), .Z(n12083) );
  XNOR U13975 ( .A(n12084), .B(n12083), .Z(n12085) );
  XNOR U13976 ( .A(n12086), .B(n12085), .Z(n12115) );
  XNOR U13977 ( .A(sreg[1232]), .B(n12115), .Z(n12117) );
  NANDN U13978 ( .A(sreg[1231]), .B(n12078), .Z(n12082) );
  NAND U13979 ( .A(n12080), .B(n12079), .Z(n12081) );
  NAND U13980 ( .A(n12082), .B(n12081), .Z(n12116) );
  XNOR U13981 ( .A(n12117), .B(n12116), .Z(c[1232]) );
  NANDN U13982 ( .A(n12084), .B(n12083), .Z(n12088) );
  NANDN U13983 ( .A(n12086), .B(n12085), .Z(n12087) );
  AND U13984 ( .A(n12088), .B(n12087), .Z(n12123) );
  NANDN U13985 ( .A(n12090), .B(n12089), .Z(n12094) );
  NANDN U13986 ( .A(n12092), .B(n12091), .Z(n12093) );
  AND U13987 ( .A(n12094), .B(n12093), .Z(n12121) );
  NAND U13988 ( .A(n42143), .B(n12095), .Z(n12097) );
  XNOR U13989 ( .A(a[211]), .B(n4102), .Z(n12132) );
  NAND U13990 ( .A(n42144), .B(n12132), .Z(n12096) );
  AND U13991 ( .A(n12097), .B(n12096), .Z(n12147) );
  XOR U13992 ( .A(a[215]), .B(n42012), .Z(n12135) );
  XNOR U13993 ( .A(n12147), .B(n12146), .Z(n12149) );
  XOR U13994 ( .A(a[213]), .B(n42085), .Z(n12139) );
  AND U13995 ( .A(a[209]), .B(b[7]), .Z(n12140) );
  XNOR U13996 ( .A(n12141), .B(n12140), .Z(n12142) );
  AND U13997 ( .A(a[217]), .B(b[0]), .Z(n12100) );
  XNOR U13998 ( .A(n12100), .B(n4071), .Z(n12102) );
  NANDN U13999 ( .A(b[0]), .B(a[216]), .Z(n12101) );
  NAND U14000 ( .A(n12102), .B(n12101), .Z(n12143) );
  XNOR U14001 ( .A(n12142), .B(n12143), .Z(n12148) );
  XOR U14002 ( .A(n12149), .B(n12148), .Z(n12127) );
  NANDN U14003 ( .A(n12104), .B(n12103), .Z(n12108) );
  NANDN U14004 ( .A(n12106), .B(n12105), .Z(n12107) );
  AND U14005 ( .A(n12108), .B(n12107), .Z(n12126) );
  XNOR U14006 ( .A(n12127), .B(n12126), .Z(n12128) );
  NANDN U14007 ( .A(n12110), .B(n12109), .Z(n12114) );
  NAND U14008 ( .A(n12112), .B(n12111), .Z(n12113) );
  NAND U14009 ( .A(n12114), .B(n12113), .Z(n12129) );
  XNOR U14010 ( .A(n12128), .B(n12129), .Z(n12120) );
  XNOR U14011 ( .A(n12121), .B(n12120), .Z(n12122) );
  XNOR U14012 ( .A(n12123), .B(n12122), .Z(n12152) );
  XNOR U14013 ( .A(sreg[1233]), .B(n12152), .Z(n12154) );
  NANDN U14014 ( .A(sreg[1232]), .B(n12115), .Z(n12119) );
  NAND U14015 ( .A(n12117), .B(n12116), .Z(n12118) );
  NAND U14016 ( .A(n12119), .B(n12118), .Z(n12153) );
  XNOR U14017 ( .A(n12154), .B(n12153), .Z(c[1233]) );
  NANDN U14018 ( .A(n12121), .B(n12120), .Z(n12125) );
  NANDN U14019 ( .A(n12123), .B(n12122), .Z(n12124) );
  AND U14020 ( .A(n12125), .B(n12124), .Z(n12160) );
  NANDN U14021 ( .A(n12127), .B(n12126), .Z(n12131) );
  NANDN U14022 ( .A(n12129), .B(n12128), .Z(n12130) );
  AND U14023 ( .A(n12131), .B(n12130), .Z(n12158) );
  NAND U14024 ( .A(n42143), .B(n12132), .Z(n12134) );
  XNOR U14025 ( .A(a[212]), .B(n4102), .Z(n12169) );
  NAND U14026 ( .A(n42144), .B(n12169), .Z(n12133) );
  AND U14027 ( .A(n12134), .B(n12133), .Z(n12184) );
  XOR U14028 ( .A(a[216]), .B(n42012), .Z(n12172) );
  XNOR U14029 ( .A(n12184), .B(n12183), .Z(n12186) );
  AND U14030 ( .A(a[218]), .B(b[0]), .Z(n12136) );
  XNOR U14031 ( .A(n12136), .B(n4071), .Z(n12138) );
  NANDN U14032 ( .A(b[0]), .B(a[217]), .Z(n12137) );
  NAND U14033 ( .A(n12138), .B(n12137), .Z(n12180) );
  XOR U14034 ( .A(a[214]), .B(n42085), .Z(n12176) );
  AND U14035 ( .A(a[210]), .B(b[7]), .Z(n12177) );
  XNOR U14036 ( .A(n12178), .B(n12177), .Z(n12179) );
  XNOR U14037 ( .A(n12180), .B(n12179), .Z(n12185) );
  XOR U14038 ( .A(n12186), .B(n12185), .Z(n12164) );
  NANDN U14039 ( .A(n12141), .B(n12140), .Z(n12145) );
  NANDN U14040 ( .A(n12143), .B(n12142), .Z(n12144) );
  AND U14041 ( .A(n12145), .B(n12144), .Z(n12163) );
  XNOR U14042 ( .A(n12164), .B(n12163), .Z(n12165) );
  NANDN U14043 ( .A(n12147), .B(n12146), .Z(n12151) );
  NAND U14044 ( .A(n12149), .B(n12148), .Z(n12150) );
  NAND U14045 ( .A(n12151), .B(n12150), .Z(n12166) );
  XNOR U14046 ( .A(n12165), .B(n12166), .Z(n12157) );
  XNOR U14047 ( .A(n12158), .B(n12157), .Z(n12159) );
  XNOR U14048 ( .A(n12160), .B(n12159), .Z(n12189) );
  XNOR U14049 ( .A(sreg[1234]), .B(n12189), .Z(n12191) );
  NANDN U14050 ( .A(sreg[1233]), .B(n12152), .Z(n12156) );
  NAND U14051 ( .A(n12154), .B(n12153), .Z(n12155) );
  NAND U14052 ( .A(n12156), .B(n12155), .Z(n12190) );
  XNOR U14053 ( .A(n12191), .B(n12190), .Z(c[1234]) );
  NANDN U14054 ( .A(n12158), .B(n12157), .Z(n12162) );
  NANDN U14055 ( .A(n12160), .B(n12159), .Z(n12161) );
  AND U14056 ( .A(n12162), .B(n12161), .Z(n12197) );
  NANDN U14057 ( .A(n12164), .B(n12163), .Z(n12168) );
  NANDN U14058 ( .A(n12166), .B(n12165), .Z(n12167) );
  AND U14059 ( .A(n12168), .B(n12167), .Z(n12195) );
  NAND U14060 ( .A(n42143), .B(n12169), .Z(n12171) );
  XNOR U14061 ( .A(a[213]), .B(n4102), .Z(n12206) );
  NAND U14062 ( .A(n42144), .B(n12206), .Z(n12170) );
  AND U14063 ( .A(n12171), .B(n12170), .Z(n12221) );
  XOR U14064 ( .A(a[217]), .B(n42012), .Z(n12209) );
  XNOR U14065 ( .A(n12221), .B(n12220), .Z(n12223) );
  AND U14066 ( .A(a[219]), .B(b[0]), .Z(n12173) );
  XNOR U14067 ( .A(n12173), .B(n4071), .Z(n12175) );
  NANDN U14068 ( .A(b[0]), .B(a[218]), .Z(n12174) );
  NAND U14069 ( .A(n12175), .B(n12174), .Z(n12217) );
  XOR U14070 ( .A(a[215]), .B(n42085), .Z(n12213) );
  AND U14071 ( .A(a[211]), .B(b[7]), .Z(n12214) );
  XNOR U14072 ( .A(n12215), .B(n12214), .Z(n12216) );
  XNOR U14073 ( .A(n12217), .B(n12216), .Z(n12222) );
  XOR U14074 ( .A(n12223), .B(n12222), .Z(n12201) );
  NANDN U14075 ( .A(n12178), .B(n12177), .Z(n12182) );
  NANDN U14076 ( .A(n12180), .B(n12179), .Z(n12181) );
  AND U14077 ( .A(n12182), .B(n12181), .Z(n12200) );
  XNOR U14078 ( .A(n12201), .B(n12200), .Z(n12202) );
  NANDN U14079 ( .A(n12184), .B(n12183), .Z(n12188) );
  NAND U14080 ( .A(n12186), .B(n12185), .Z(n12187) );
  NAND U14081 ( .A(n12188), .B(n12187), .Z(n12203) );
  XNOR U14082 ( .A(n12202), .B(n12203), .Z(n12194) );
  XNOR U14083 ( .A(n12195), .B(n12194), .Z(n12196) );
  XNOR U14084 ( .A(n12197), .B(n12196), .Z(n12226) );
  XNOR U14085 ( .A(sreg[1235]), .B(n12226), .Z(n12228) );
  NANDN U14086 ( .A(sreg[1234]), .B(n12189), .Z(n12193) );
  NAND U14087 ( .A(n12191), .B(n12190), .Z(n12192) );
  NAND U14088 ( .A(n12193), .B(n12192), .Z(n12227) );
  XNOR U14089 ( .A(n12228), .B(n12227), .Z(c[1235]) );
  NANDN U14090 ( .A(n12195), .B(n12194), .Z(n12199) );
  NANDN U14091 ( .A(n12197), .B(n12196), .Z(n12198) );
  AND U14092 ( .A(n12199), .B(n12198), .Z(n12234) );
  NANDN U14093 ( .A(n12201), .B(n12200), .Z(n12205) );
  NANDN U14094 ( .A(n12203), .B(n12202), .Z(n12204) );
  AND U14095 ( .A(n12205), .B(n12204), .Z(n12232) );
  NAND U14096 ( .A(n42143), .B(n12206), .Z(n12208) );
  XNOR U14097 ( .A(a[214]), .B(n4102), .Z(n12243) );
  NAND U14098 ( .A(n42144), .B(n12243), .Z(n12207) );
  AND U14099 ( .A(n12208), .B(n12207), .Z(n12258) );
  XOR U14100 ( .A(a[218]), .B(n42012), .Z(n12246) );
  XNOR U14101 ( .A(n12258), .B(n12257), .Z(n12260) );
  AND U14102 ( .A(a[220]), .B(b[0]), .Z(n12210) );
  XNOR U14103 ( .A(n12210), .B(n4071), .Z(n12212) );
  NANDN U14104 ( .A(b[0]), .B(a[219]), .Z(n12211) );
  NAND U14105 ( .A(n12212), .B(n12211), .Z(n12254) );
  XOR U14106 ( .A(a[216]), .B(n42085), .Z(n12250) );
  AND U14107 ( .A(a[212]), .B(b[7]), .Z(n12251) );
  XNOR U14108 ( .A(n12252), .B(n12251), .Z(n12253) );
  XNOR U14109 ( .A(n12254), .B(n12253), .Z(n12259) );
  XOR U14110 ( .A(n12260), .B(n12259), .Z(n12238) );
  NANDN U14111 ( .A(n12215), .B(n12214), .Z(n12219) );
  NANDN U14112 ( .A(n12217), .B(n12216), .Z(n12218) );
  AND U14113 ( .A(n12219), .B(n12218), .Z(n12237) );
  XNOR U14114 ( .A(n12238), .B(n12237), .Z(n12239) );
  NANDN U14115 ( .A(n12221), .B(n12220), .Z(n12225) );
  NAND U14116 ( .A(n12223), .B(n12222), .Z(n12224) );
  NAND U14117 ( .A(n12225), .B(n12224), .Z(n12240) );
  XNOR U14118 ( .A(n12239), .B(n12240), .Z(n12231) );
  XNOR U14119 ( .A(n12232), .B(n12231), .Z(n12233) );
  XNOR U14120 ( .A(n12234), .B(n12233), .Z(n12263) );
  XNOR U14121 ( .A(sreg[1236]), .B(n12263), .Z(n12265) );
  NANDN U14122 ( .A(sreg[1235]), .B(n12226), .Z(n12230) );
  NAND U14123 ( .A(n12228), .B(n12227), .Z(n12229) );
  NAND U14124 ( .A(n12230), .B(n12229), .Z(n12264) );
  XNOR U14125 ( .A(n12265), .B(n12264), .Z(c[1236]) );
  NANDN U14126 ( .A(n12232), .B(n12231), .Z(n12236) );
  NANDN U14127 ( .A(n12234), .B(n12233), .Z(n12235) );
  AND U14128 ( .A(n12236), .B(n12235), .Z(n12271) );
  NANDN U14129 ( .A(n12238), .B(n12237), .Z(n12242) );
  NANDN U14130 ( .A(n12240), .B(n12239), .Z(n12241) );
  AND U14131 ( .A(n12242), .B(n12241), .Z(n12269) );
  NAND U14132 ( .A(n42143), .B(n12243), .Z(n12245) );
  XNOR U14133 ( .A(a[215]), .B(n4102), .Z(n12280) );
  NAND U14134 ( .A(n42144), .B(n12280), .Z(n12244) );
  AND U14135 ( .A(n12245), .B(n12244), .Z(n12295) );
  XOR U14136 ( .A(a[219]), .B(n42012), .Z(n12283) );
  XNOR U14137 ( .A(n12295), .B(n12294), .Z(n12297) );
  AND U14138 ( .A(a[221]), .B(b[0]), .Z(n12247) );
  XNOR U14139 ( .A(n12247), .B(n4071), .Z(n12249) );
  NANDN U14140 ( .A(b[0]), .B(a[220]), .Z(n12248) );
  NAND U14141 ( .A(n12249), .B(n12248), .Z(n12291) );
  XOR U14142 ( .A(a[217]), .B(n42085), .Z(n12284) );
  AND U14143 ( .A(a[213]), .B(b[7]), .Z(n12288) );
  XNOR U14144 ( .A(n12289), .B(n12288), .Z(n12290) );
  XNOR U14145 ( .A(n12291), .B(n12290), .Z(n12296) );
  XOR U14146 ( .A(n12297), .B(n12296), .Z(n12275) );
  NANDN U14147 ( .A(n12252), .B(n12251), .Z(n12256) );
  NANDN U14148 ( .A(n12254), .B(n12253), .Z(n12255) );
  AND U14149 ( .A(n12256), .B(n12255), .Z(n12274) );
  XNOR U14150 ( .A(n12275), .B(n12274), .Z(n12276) );
  NANDN U14151 ( .A(n12258), .B(n12257), .Z(n12262) );
  NAND U14152 ( .A(n12260), .B(n12259), .Z(n12261) );
  NAND U14153 ( .A(n12262), .B(n12261), .Z(n12277) );
  XNOR U14154 ( .A(n12276), .B(n12277), .Z(n12268) );
  XNOR U14155 ( .A(n12269), .B(n12268), .Z(n12270) );
  XNOR U14156 ( .A(n12271), .B(n12270), .Z(n12300) );
  XNOR U14157 ( .A(sreg[1237]), .B(n12300), .Z(n12302) );
  NANDN U14158 ( .A(sreg[1236]), .B(n12263), .Z(n12267) );
  NAND U14159 ( .A(n12265), .B(n12264), .Z(n12266) );
  NAND U14160 ( .A(n12267), .B(n12266), .Z(n12301) );
  XNOR U14161 ( .A(n12302), .B(n12301), .Z(c[1237]) );
  NANDN U14162 ( .A(n12269), .B(n12268), .Z(n12273) );
  NANDN U14163 ( .A(n12271), .B(n12270), .Z(n12272) );
  AND U14164 ( .A(n12273), .B(n12272), .Z(n12308) );
  NANDN U14165 ( .A(n12275), .B(n12274), .Z(n12279) );
  NANDN U14166 ( .A(n12277), .B(n12276), .Z(n12278) );
  AND U14167 ( .A(n12279), .B(n12278), .Z(n12306) );
  NAND U14168 ( .A(n42143), .B(n12280), .Z(n12282) );
  XNOR U14169 ( .A(a[216]), .B(n4102), .Z(n12317) );
  NAND U14170 ( .A(n42144), .B(n12317), .Z(n12281) );
  AND U14171 ( .A(n12282), .B(n12281), .Z(n12332) );
  XOR U14172 ( .A(a[220]), .B(n42012), .Z(n12320) );
  XNOR U14173 ( .A(n12332), .B(n12331), .Z(n12334) );
  XOR U14174 ( .A(a[218]), .B(n42085), .Z(n12324) );
  AND U14175 ( .A(a[214]), .B(b[7]), .Z(n12325) );
  XNOR U14176 ( .A(n12326), .B(n12325), .Z(n12327) );
  AND U14177 ( .A(a[222]), .B(b[0]), .Z(n12285) );
  XNOR U14178 ( .A(n12285), .B(n4071), .Z(n12287) );
  NANDN U14179 ( .A(b[0]), .B(a[221]), .Z(n12286) );
  NAND U14180 ( .A(n12287), .B(n12286), .Z(n12328) );
  XNOR U14181 ( .A(n12327), .B(n12328), .Z(n12333) );
  XOR U14182 ( .A(n12334), .B(n12333), .Z(n12312) );
  NANDN U14183 ( .A(n12289), .B(n12288), .Z(n12293) );
  NANDN U14184 ( .A(n12291), .B(n12290), .Z(n12292) );
  AND U14185 ( .A(n12293), .B(n12292), .Z(n12311) );
  XNOR U14186 ( .A(n12312), .B(n12311), .Z(n12313) );
  NANDN U14187 ( .A(n12295), .B(n12294), .Z(n12299) );
  NAND U14188 ( .A(n12297), .B(n12296), .Z(n12298) );
  NAND U14189 ( .A(n12299), .B(n12298), .Z(n12314) );
  XNOR U14190 ( .A(n12313), .B(n12314), .Z(n12305) );
  XNOR U14191 ( .A(n12306), .B(n12305), .Z(n12307) );
  XNOR U14192 ( .A(n12308), .B(n12307), .Z(n12337) );
  XNOR U14193 ( .A(sreg[1238]), .B(n12337), .Z(n12339) );
  NANDN U14194 ( .A(sreg[1237]), .B(n12300), .Z(n12304) );
  NAND U14195 ( .A(n12302), .B(n12301), .Z(n12303) );
  NAND U14196 ( .A(n12304), .B(n12303), .Z(n12338) );
  XNOR U14197 ( .A(n12339), .B(n12338), .Z(c[1238]) );
  NANDN U14198 ( .A(n12306), .B(n12305), .Z(n12310) );
  NANDN U14199 ( .A(n12308), .B(n12307), .Z(n12309) );
  AND U14200 ( .A(n12310), .B(n12309), .Z(n12345) );
  NANDN U14201 ( .A(n12312), .B(n12311), .Z(n12316) );
  NANDN U14202 ( .A(n12314), .B(n12313), .Z(n12315) );
  AND U14203 ( .A(n12316), .B(n12315), .Z(n12343) );
  NAND U14204 ( .A(n42143), .B(n12317), .Z(n12319) );
  XNOR U14205 ( .A(a[217]), .B(n4102), .Z(n12354) );
  NAND U14206 ( .A(n42144), .B(n12354), .Z(n12318) );
  AND U14207 ( .A(n12319), .B(n12318), .Z(n12369) );
  XOR U14208 ( .A(a[221]), .B(n42012), .Z(n12357) );
  XNOR U14209 ( .A(n12369), .B(n12368), .Z(n12371) );
  AND U14210 ( .A(a[223]), .B(b[0]), .Z(n12321) );
  XNOR U14211 ( .A(n12321), .B(n4071), .Z(n12323) );
  NANDN U14212 ( .A(b[0]), .B(a[222]), .Z(n12322) );
  NAND U14213 ( .A(n12323), .B(n12322), .Z(n12365) );
  XOR U14214 ( .A(a[219]), .B(n42085), .Z(n12361) );
  AND U14215 ( .A(a[215]), .B(b[7]), .Z(n12362) );
  XNOR U14216 ( .A(n12363), .B(n12362), .Z(n12364) );
  XNOR U14217 ( .A(n12365), .B(n12364), .Z(n12370) );
  XOR U14218 ( .A(n12371), .B(n12370), .Z(n12349) );
  NANDN U14219 ( .A(n12326), .B(n12325), .Z(n12330) );
  NANDN U14220 ( .A(n12328), .B(n12327), .Z(n12329) );
  AND U14221 ( .A(n12330), .B(n12329), .Z(n12348) );
  XNOR U14222 ( .A(n12349), .B(n12348), .Z(n12350) );
  NANDN U14223 ( .A(n12332), .B(n12331), .Z(n12336) );
  NAND U14224 ( .A(n12334), .B(n12333), .Z(n12335) );
  NAND U14225 ( .A(n12336), .B(n12335), .Z(n12351) );
  XNOR U14226 ( .A(n12350), .B(n12351), .Z(n12342) );
  XNOR U14227 ( .A(n12343), .B(n12342), .Z(n12344) );
  XNOR U14228 ( .A(n12345), .B(n12344), .Z(n12374) );
  XNOR U14229 ( .A(sreg[1239]), .B(n12374), .Z(n12376) );
  NANDN U14230 ( .A(sreg[1238]), .B(n12337), .Z(n12341) );
  NAND U14231 ( .A(n12339), .B(n12338), .Z(n12340) );
  NAND U14232 ( .A(n12341), .B(n12340), .Z(n12375) );
  XNOR U14233 ( .A(n12376), .B(n12375), .Z(c[1239]) );
  NANDN U14234 ( .A(n12343), .B(n12342), .Z(n12347) );
  NANDN U14235 ( .A(n12345), .B(n12344), .Z(n12346) );
  AND U14236 ( .A(n12347), .B(n12346), .Z(n12382) );
  NANDN U14237 ( .A(n12349), .B(n12348), .Z(n12353) );
  NANDN U14238 ( .A(n12351), .B(n12350), .Z(n12352) );
  AND U14239 ( .A(n12353), .B(n12352), .Z(n12380) );
  NAND U14240 ( .A(n42143), .B(n12354), .Z(n12356) );
  XNOR U14241 ( .A(a[218]), .B(n4103), .Z(n12391) );
  NAND U14242 ( .A(n42144), .B(n12391), .Z(n12355) );
  AND U14243 ( .A(n12356), .B(n12355), .Z(n12406) );
  XOR U14244 ( .A(a[222]), .B(n42012), .Z(n12394) );
  XNOR U14245 ( .A(n12406), .B(n12405), .Z(n12408) );
  AND U14246 ( .A(a[224]), .B(b[0]), .Z(n12358) );
  XNOR U14247 ( .A(n12358), .B(n4071), .Z(n12360) );
  NANDN U14248 ( .A(b[0]), .B(a[223]), .Z(n12359) );
  NAND U14249 ( .A(n12360), .B(n12359), .Z(n12402) );
  XOR U14250 ( .A(a[220]), .B(n42085), .Z(n12395) );
  AND U14251 ( .A(a[216]), .B(b[7]), .Z(n12399) );
  XNOR U14252 ( .A(n12400), .B(n12399), .Z(n12401) );
  XNOR U14253 ( .A(n12402), .B(n12401), .Z(n12407) );
  XOR U14254 ( .A(n12408), .B(n12407), .Z(n12386) );
  NANDN U14255 ( .A(n12363), .B(n12362), .Z(n12367) );
  NANDN U14256 ( .A(n12365), .B(n12364), .Z(n12366) );
  AND U14257 ( .A(n12367), .B(n12366), .Z(n12385) );
  XNOR U14258 ( .A(n12386), .B(n12385), .Z(n12387) );
  NANDN U14259 ( .A(n12369), .B(n12368), .Z(n12373) );
  NAND U14260 ( .A(n12371), .B(n12370), .Z(n12372) );
  NAND U14261 ( .A(n12373), .B(n12372), .Z(n12388) );
  XNOR U14262 ( .A(n12387), .B(n12388), .Z(n12379) );
  XNOR U14263 ( .A(n12380), .B(n12379), .Z(n12381) );
  XNOR U14264 ( .A(n12382), .B(n12381), .Z(n12411) );
  XNOR U14265 ( .A(sreg[1240]), .B(n12411), .Z(n12413) );
  NANDN U14266 ( .A(sreg[1239]), .B(n12374), .Z(n12378) );
  NAND U14267 ( .A(n12376), .B(n12375), .Z(n12377) );
  NAND U14268 ( .A(n12378), .B(n12377), .Z(n12412) );
  XNOR U14269 ( .A(n12413), .B(n12412), .Z(c[1240]) );
  NANDN U14270 ( .A(n12380), .B(n12379), .Z(n12384) );
  NANDN U14271 ( .A(n12382), .B(n12381), .Z(n12383) );
  AND U14272 ( .A(n12384), .B(n12383), .Z(n12419) );
  NANDN U14273 ( .A(n12386), .B(n12385), .Z(n12390) );
  NANDN U14274 ( .A(n12388), .B(n12387), .Z(n12389) );
  AND U14275 ( .A(n12390), .B(n12389), .Z(n12417) );
  NAND U14276 ( .A(n42143), .B(n12391), .Z(n12393) );
  XNOR U14277 ( .A(a[219]), .B(n4103), .Z(n12428) );
  NAND U14278 ( .A(n42144), .B(n12428), .Z(n12392) );
  AND U14279 ( .A(n12393), .B(n12392), .Z(n12443) );
  XOR U14280 ( .A(a[223]), .B(n42012), .Z(n12431) );
  XNOR U14281 ( .A(n12443), .B(n12442), .Z(n12445) );
  XOR U14282 ( .A(a[221]), .B(n42085), .Z(n12435) );
  AND U14283 ( .A(a[217]), .B(b[7]), .Z(n12436) );
  XNOR U14284 ( .A(n12437), .B(n12436), .Z(n12438) );
  AND U14285 ( .A(a[225]), .B(b[0]), .Z(n12396) );
  XNOR U14286 ( .A(n12396), .B(n4071), .Z(n12398) );
  NANDN U14287 ( .A(b[0]), .B(a[224]), .Z(n12397) );
  NAND U14288 ( .A(n12398), .B(n12397), .Z(n12439) );
  XNOR U14289 ( .A(n12438), .B(n12439), .Z(n12444) );
  XOR U14290 ( .A(n12445), .B(n12444), .Z(n12423) );
  NANDN U14291 ( .A(n12400), .B(n12399), .Z(n12404) );
  NANDN U14292 ( .A(n12402), .B(n12401), .Z(n12403) );
  AND U14293 ( .A(n12404), .B(n12403), .Z(n12422) );
  XNOR U14294 ( .A(n12423), .B(n12422), .Z(n12424) );
  NANDN U14295 ( .A(n12406), .B(n12405), .Z(n12410) );
  NAND U14296 ( .A(n12408), .B(n12407), .Z(n12409) );
  NAND U14297 ( .A(n12410), .B(n12409), .Z(n12425) );
  XNOR U14298 ( .A(n12424), .B(n12425), .Z(n12416) );
  XNOR U14299 ( .A(n12417), .B(n12416), .Z(n12418) );
  XNOR U14300 ( .A(n12419), .B(n12418), .Z(n12448) );
  XNOR U14301 ( .A(sreg[1241]), .B(n12448), .Z(n12450) );
  NANDN U14302 ( .A(sreg[1240]), .B(n12411), .Z(n12415) );
  NAND U14303 ( .A(n12413), .B(n12412), .Z(n12414) );
  NAND U14304 ( .A(n12415), .B(n12414), .Z(n12449) );
  XNOR U14305 ( .A(n12450), .B(n12449), .Z(c[1241]) );
  NANDN U14306 ( .A(n12417), .B(n12416), .Z(n12421) );
  NANDN U14307 ( .A(n12419), .B(n12418), .Z(n12420) );
  AND U14308 ( .A(n12421), .B(n12420), .Z(n12456) );
  NANDN U14309 ( .A(n12423), .B(n12422), .Z(n12427) );
  NANDN U14310 ( .A(n12425), .B(n12424), .Z(n12426) );
  AND U14311 ( .A(n12427), .B(n12426), .Z(n12454) );
  NAND U14312 ( .A(n42143), .B(n12428), .Z(n12430) );
  XNOR U14313 ( .A(a[220]), .B(n4103), .Z(n12465) );
  NAND U14314 ( .A(n42144), .B(n12465), .Z(n12429) );
  AND U14315 ( .A(n12430), .B(n12429), .Z(n12480) );
  XOR U14316 ( .A(a[224]), .B(n42012), .Z(n12468) );
  XNOR U14317 ( .A(n12480), .B(n12479), .Z(n12482) );
  AND U14318 ( .A(a[226]), .B(b[0]), .Z(n12432) );
  XNOR U14319 ( .A(n12432), .B(n4071), .Z(n12434) );
  NANDN U14320 ( .A(b[0]), .B(a[225]), .Z(n12433) );
  NAND U14321 ( .A(n12434), .B(n12433), .Z(n12476) );
  XOR U14322 ( .A(a[222]), .B(n42085), .Z(n12472) );
  AND U14323 ( .A(a[218]), .B(b[7]), .Z(n12473) );
  XNOR U14324 ( .A(n12474), .B(n12473), .Z(n12475) );
  XNOR U14325 ( .A(n12476), .B(n12475), .Z(n12481) );
  XOR U14326 ( .A(n12482), .B(n12481), .Z(n12460) );
  NANDN U14327 ( .A(n12437), .B(n12436), .Z(n12441) );
  NANDN U14328 ( .A(n12439), .B(n12438), .Z(n12440) );
  AND U14329 ( .A(n12441), .B(n12440), .Z(n12459) );
  XNOR U14330 ( .A(n12460), .B(n12459), .Z(n12461) );
  NANDN U14331 ( .A(n12443), .B(n12442), .Z(n12447) );
  NAND U14332 ( .A(n12445), .B(n12444), .Z(n12446) );
  NAND U14333 ( .A(n12447), .B(n12446), .Z(n12462) );
  XNOR U14334 ( .A(n12461), .B(n12462), .Z(n12453) );
  XNOR U14335 ( .A(n12454), .B(n12453), .Z(n12455) );
  XNOR U14336 ( .A(n12456), .B(n12455), .Z(n12485) );
  XNOR U14337 ( .A(sreg[1242]), .B(n12485), .Z(n12487) );
  NANDN U14338 ( .A(sreg[1241]), .B(n12448), .Z(n12452) );
  NAND U14339 ( .A(n12450), .B(n12449), .Z(n12451) );
  NAND U14340 ( .A(n12452), .B(n12451), .Z(n12486) );
  XNOR U14341 ( .A(n12487), .B(n12486), .Z(c[1242]) );
  NANDN U14342 ( .A(n12454), .B(n12453), .Z(n12458) );
  NANDN U14343 ( .A(n12456), .B(n12455), .Z(n12457) );
  AND U14344 ( .A(n12458), .B(n12457), .Z(n12493) );
  NANDN U14345 ( .A(n12460), .B(n12459), .Z(n12464) );
  NANDN U14346 ( .A(n12462), .B(n12461), .Z(n12463) );
  AND U14347 ( .A(n12464), .B(n12463), .Z(n12491) );
  NAND U14348 ( .A(n42143), .B(n12465), .Z(n12467) );
  XNOR U14349 ( .A(a[221]), .B(n4103), .Z(n12502) );
  NAND U14350 ( .A(n42144), .B(n12502), .Z(n12466) );
  AND U14351 ( .A(n12467), .B(n12466), .Z(n12517) );
  XOR U14352 ( .A(a[225]), .B(n42012), .Z(n12505) );
  XNOR U14353 ( .A(n12517), .B(n12516), .Z(n12519) );
  AND U14354 ( .A(a[227]), .B(b[0]), .Z(n12469) );
  XNOR U14355 ( .A(n12469), .B(n4071), .Z(n12471) );
  NANDN U14356 ( .A(b[0]), .B(a[226]), .Z(n12470) );
  NAND U14357 ( .A(n12471), .B(n12470), .Z(n12513) );
  XOR U14358 ( .A(a[223]), .B(n42085), .Z(n12506) );
  AND U14359 ( .A(a[219]), .B(b[7]), .Z(n12510) );
  XNOR U14360 ( .A(n12511), .B(n12510), .Z(n12512) );
  XNOR U14361 ( .A(n12513), .B(n12512), .Z(n12518) );
  XOR U14362 ( .A(n12519), .B(n12518), .Z(n12497) );
  NANDN U14363 ( .A(n12474), .B(n12473), .Z(n12478) );
  NANDN U14364 ( .A(n12476), .B(n12475), .Z(n12477) );
  AND U14365 ( .A(n12478), .B(n12477), .Z(n12496) );
  XNOR U14366 ( .A(n12497), .B(n12496), .Z(n12498) );
  NANDN U14367 ( .A(n12480), .B(n12479), .Z(n12484) );
  NAND U14368 ( .A(n12482), .B(n12481), .Z(n12483) );
  NAND U14369 ( .A(n12484), .B(n12483), .Z(n12499) );
  XNOR U14370 ( .A(n12498), .B(n12499), .Z(n12490) );
  XNOR U14371 ( .A(n12491), .B(n12490), .Z(n12492) );
  XNOR U14372 ( .A(n12493), .B(n12492), .Z(n12522) );
  XNOR U14373 ( .A(sreg[1243]), .B(n12522), .Z(n12524) );
  NANDN U14374 ( .A(sreg[1242]), .B(n12485), .Z(n12489) );
  NAND U14375 ( .A(n12487), .B(n12486), .Z(n12488) );
  NAND U14376 ( .A(n12489), .B(n12488), .Z(n12523) );
  XNOR U14377 ( .A(n12524), .B(n12523), .Z(c[1243]) );
  NANDN U14378 ( .A(n12491), .B(n12490), .Z(n12495) );
  NANDN U14379 ( .A(n12493), .B(n12492), .Z(n12494) );
  AND U14380 ( .A(n12495), .B(n12494), .Z(n12530) );
  NANDN U14381 ( .A(n12497), .B(n12496), .Z(n12501) );
  NANDN U14382 ( .A(n12499), .B(n12498), .Z(n12500) );
  AND U14383 ( .A(n12501), .B(n12500), .Z(n12528) );
  NAND U14384 ( .A(n42143), .B(n12502), .Z(n12504) );
  XNOR U14385 ( .A(a[222]), .B(n4103), .Z(n12539) );
  NAND U14386 ( .A(n42144), .B(n12539), .Z(n12503) );
  AND U14387 ( .A(n12504), .B(n12503), .Z(n12554) );
  XOR U14388 ( .A(a[226]), .B(n42012), .Z(n12542) );
  XNOR U14389 ( .A(n12554), .B(n12553), .Z(n12556) );
  XOR U14390 ( .A(a[224]), .B(n42085), .Z(n12546) );
  AND U14391 ( .A(a[220]), .B(b[7]), .Z(n12547) );
  XNOR U14392 ( .A(n12548), .B(n12547), .Z(n12549) );
  AND U14393 ( .A(a[228]), .B(b[0]), .Z(n12507) );
  XNOR U14394 ( .A(n12507), .B(n4071), .Z(n12509) );
  NANDN U14395 ( .A(b[0]), .B(a[227]), .Z(n12508) );
  NAND U14396 ( .A(n12509), .B(n12508), .Z(n12550) );
  XNOR U14397 ( .A(n12549), .B(n12550), .Z(n12555) );
  XOR U14398 ( .A(n12556), .B(n12555), .Z(n12534) );
  NANDN U14399 ( .A(n12511), .B(n12510), .Z(n12515) );
  NANDN U14400 ( .A(n12513), .B(n12512), .Z(n12514) );
  AND U14401 ( .A(n12515), .B(n12514), .Z(n12533) );
  XNOR U14402 ( .A(n12534), .B(n12533), .Z(n12535) );
  NANDN U14403 ( .A(n12517), .B(n12516), .Z(n12521) );
  NAND U14404 ( .A(n12519), .B(n12518), .Z(n12520) );
  NAND U14405 ( .A(n12521), .B(n12520), .Z(n12536) );
  XNOR U14406 ( .A(n12535), .B(n12536), .Z(n12527) );
  XNOR U14407 ( .A(n12528), .B(n12527), .Z(n12529) );
  XNOR U14408 ( .A(n12530), .B(n12529), .Z(n12559) );
  XNOR U14409 ( .A(sreg[1244]), .B(n12559), .Z(n12561) );
  NANDN U14410 ( .A(sreg[1243]), .B(n12522), .Z(n12526) );
  NAND U14411 ( .A(n12524), .B(n12523), .Z(n12525) );
  NAND U14412 ( .A(n12526), .B(n12525), .Z(n12560) );
  XNOR U14413 ( .A(n12561), .B(n12560), .Z(c[1244]) );
  NANDN U14414 ( .A(n12528), .B(n12527), .Z(n12532) );
  NANDN U14415 ( .A(n12530), .B(n12529), .Z(n12531) );
  AND U14416 ( .A(n12532), .B(n12531), .Z(n12567) );
  NANDN U14417 ( .A(n12534), .B(n12533), .Z(n12538) );
  NANDN U14418 ( .A(n12536), .B(n12535), .Z(n12537) );
  AND U14419 ( .A(n12538), .B(n12537), .Z(n12565) );
  NAND U14420 ( .A(n42143), .B(n12539), .Z(n12541) );
  XNOR U14421 ( .A(a[223]), .B(n4103), .Z(n12576) );
  NAND U14422 ( .A(n42144), .B(n12576), .Z(n12540) );
  AND U14423 ( .A(n12541), .B(n12540), .Z(n12591) );
  XOR U14424 ( .A(a[227]), .B(n42012), .Z(n12579) );
  XNOR U14425 ( .A(n12591), .B(n12590), .Z(n12593) );
  AND U14426 ( .A(a[229]), .B(b[0]), .Z(n12543) );
  XNOR U14427 ( .A(n12543), .B(n4071), .Z(n12545) );
  NANDN U14428 ( .A(b[0]), .B(a[228]), .Z(n12544) );
  NAND U14429 ( .A(n12545), .B(n12544), .Z(n12587) );
  XOR U14430 ( .A(a[225]), .B(n42085), .Z(n12580) );
  AND U14431 ( .A(a[221]), .B(b[7]), .Z(n12584) );
  XNOR U14432 ( .A(n12585), .B(n12584), .Z(n12586) );
  XNOR U14433 ( .A(n12587), .B(n12586), .Z(n12592) );
  XOR U14434 ( .A(n12593), .B(n12592), .Z(n12571) );
  NANDN U14435 ( .A(n12548), .B(n12547), .Z(n12552) );
  NANDN U14436 ( .A(n12550), .B(n12549), .Z(n12551) );
  AND U14437 ( .A(n12552), .B(n12551), .Z(n12570) );
  XNOR U14438 ( .A(n12571), .B(n12570), .Z(n12572) );
  NANDN U14439 ( .A(n12554), .B(n12553), .Z(n12558) );
  NAND U14440 ( .A(n12556), .B(n12555), .Z(n12557) );
  NAND U14441 ( .A(n12558), .B(n12557), .Z(n12573) );
  XNOR U14442 ( .A(n12572), .B(n12573), .Z(n12564) );
  XNOR U14443 ( .A(n12565), .B(n12564), .Z(n12566) );
  XNOR U14444 ( .A(n12567), .B(n12566), .Z(n12596) );
  XNOR U14445 ( .A(sreg[1245]), .B(n12596), .Z(n12598) );
  NANDN U14446 ( .A(sreg[1244]), .B(n12559), .Z(n12563) );
  NAND U14447 ( .A(n12561), .B(n12560), .Z(n12562) );
  NAND U14448 ( .A(n12563), .B(n12562), .Z(n12597) );
  XNOR U14449 ( .A(n12598), .B(n12597), .Z(c[1245]) );
  NANDN U14450 ( .A(n12565), .B(n12564), .Z(n12569) );
  NANDN U14451 ( .A(n12567), .B(n12566), .Z(n12568) );
  AND U14452 ( .A(n12569), .B(n12568), .Z(n12604) );
  NANDN U14453 ( .A(n12571), .B(n12570), .Z(n12575) );
  NANDN U14454 ( .A(n12573), .B(n12572), .Z(n12574) );
  AND U14455 ( .A(n12575), .B(n12574), .Z(n12602) );
  NAND U14456 ( .A(n42143), .B(n12576), .Z(n12578) );
  XNOR U14457 ( .A(a[224]), .B(n4103), .Z(n12613) );
  NAND U14458 ( .A(n42144), .B(n12613), .Z(n12577) );
  AND U14459 ( .A(n12578), .B(n12577), .Z(n12628) );
  XOR U14460 ( .A(a[228]), .B(n42012), .Z(n12616) );
  XNOR U14461 ( .A(n12628), .B(n12627), .Z(n12630) );
  XOR U14462 ( .A(a[226]), .B(n42085), .Z(n12620) );
  AND U14463 ( .A(a[222]), .B(b[7]), .Z(n12621) );
  XNOR U14464 ( .A(n12622), .B(n12621), .Z(n12623) );
  AND U14465 ( .A(a[230]), .B(b[0]), .Z(n12581) );
  XNOR U14466 ( .A(n12581), .B(n4071), .Z(n12583) );
  NANDN U14467 ( .A(b[0]), .B(a[229]), .Z(n12582) );
  NAND U14468 ( .A(n12583), .B(n12582), .Z(n12624) );
  XNOR U14469 ( .A(n12623), .B(n12624), .Z(n12629) );
  XOR U14470 ( .A(n12630), .B(n12629), .Z(n12608) );
  NANDN U14471 ( .A(n12585), .B(n12584), .Z(n12589) );
  NANDN U14472 ( .A(n12587), .B(n12586), .Z(n12588) );
  AND U14473 ( .A(n12589), .B(n12588), .Z(n12607) );
  XNOR U14474 ( .A(n12608), .B(n12607), .Z(n12609) );
  NANDN U14475 ( .A(n12591), .B(n12590), .Z(n12595) );
  NAND U14476 ( .A(n12593), .B(n12592), .Z(n12594) );
  NAND U14477 ( .A(n12595), .B(n12594), .Z(n12610) );
  XNOR U14478 ( .A(n12609), .B(n12610), .Z(n12601) );
  XNOR U14479 ( .A(n12602), .B(n12601), .Z(n12603) );
  XNOR U14480 ( .A(n12604), .B(n12603), .Z(n12633) );
  XNOR U14481 ( .A(sreg[1246]), .B(n12633), .Z(n12635) );
  NANDN U14482 ( .A(sreg[1245]), .B(n12596), .Z(n12600) );
  NAND U14483 ( .A(n12598), .B(n12597), .Z(n12599) );
  NAND U14484 ( .A(n12600), .B(n12599), .Z(n12634) );
  XNOR U14485 ( .A(n12635), .B(n12634), .Z(c[1246]) );
  NANDN U14486 ( .A(n12602), .B(n12601), .Z(n12606) );
  NANDN U14487 ( .A(n12604), .B(n12603), .Z(n12605) );
  AND U14488 ( .A(n12606), .B(n12605), .Z(n12641) );
  NANDN U14489 ( .A(n12608), .B(n12607), .Z(n12612) );
  NANDN U14490 ( .A(n12610), .B(n12609), .Z(n12611) );
  AND U14491 ( .A(n12612), .B(n12611), .Z(n12639) );
  NAND U14492 ( .A(n42143), .B(n12613), .Z(n12615) );
  XNOR U14493 ( .A(a[225]), .B(n4104), .Z(n12650) );
  NAND U14494 ( .A(n42144), .B(n12650), .Z(n12614) );
  AND U14495 ( .A(n12615), .B(n12614), .Z(n12665) );
  XOR U14496 ( .A(a[229]), .B(n42012), .Z(n12653) );
  XNOR U14497 ( .A(n12665), .B(n12664), .Z(n12667) );
  AND U14498 ( .A(a[231]), .B(b[0]), .Z(n12617) );
  XNOR U14499 ( .A(n12617), .B(n4071), .Z(n12619) );
  NANDN U14500 ( .A(b[0]), .B(a[230]), .Z(n12618) );
  NAND U14501 ( .A(n12619), .B(n12618), .Z(n12661) );
  XOR U14502 ( .A(a[227]), .B(n42085), .Z(n12657) );
  AND U14503 ( .A(a[223]), .B(b[7]), .Z(n12658) );
  XNOR U14504 ( .A(n12659), .B(n12658), .Z(n12660) );
  XNOR U14505 ( .A(n12661), .B(n12660), .Z(n12666) );
  XOR U14506 ( .A(n12667), .B(n12666), .Z(n12645) );
  NANDN U14507 ( .A(n12622), .B(n12621), .Z(n12626) );
  NANDN U14508 ( .A(n12624), .B(n12623), .Z(n12625) );
  AND U14509 ( .A(n12626), .B(n12625), .Z(n12644) );
  XNOR U14510 ( .A(n12645), .B(n12644), .Z(n12646) );
  NANDN U14511 ( .A(n12628), .B(n12627), .Z(n12632) );
  NAND U14512 ( .A(n12630), .B(n12629), .Z(n12631) );
  NAND U14513 ( .A(n12632), .B(n12631), .Z(n12647) );
  XNOR U14514 ( .A(n12646), .B(n12647), .Z(n12638) );
  XNOR U14515 ( .A(n12639), .B(n12638), .Z(n12640) );
  XNOR U14516 ( .A(n12641), .B(n12640), .Z(n12670) );
  XNOR U14517 ( .A(sreg[1247]), .B(n12670), .Z(n12672) );
  NANDN U14518 ( .A(sreg[1246]), .B(n12633), .Z(n12637) );
  NAND U14519 ( .A(n12635), .B(n12634), .Z(n12636) );
  NAND U14520 ( .A(n12637), .B(n12636), .Z(n12671) );
  XNOR U14521 ( .A(n12672), .B(n12671), .Z(c[1247]) );
  NANDN U14522 ( .A(n12639), .B(n12638), .Z(n12643) );
  NANDN U14523 ( .A(n12641), .B(n12640), .Z(n12642) );
  AND U14524 ( .A(n12643), .B(n12642), .Z(n12678) );
  NANDN U14525 ( .A(n12645), .B(n12644), .Z(n12649) );
  NANDN U14526 ( .A(n12647), .B(n12646), .Z(n12648) );
  AND U14527 ( .A(n12649), .B(n12648), .Z(n12676) );
  NAND U14528 ( .A(n42143), .B(n12650), .Z(n12652) );
  XNOR U14529 ( .A(a[226]), .B(n4104), .Z(n12687) );
  NAND U14530 ( .A(n42144), .B(n12687), .Z(n12651) );
  AND U14531 ( .A(n12652), .B(n12651), .Z(n12702) );
  XOR U14532 ( .A(a[230]), .B(n42012), .Z(n12690) );
  XNOR U14533 ( .A(n12702), .B(n12701), .Z(n12704) );
  AND U14534 ( .A(a[232]), .B(b[0]), .Z(n12654) );
  XNOR U14535 ( .A(n12654), .B(n4071), .Z(n12656) );
  NANDN U14536 ( .A(b[0]), .B(a[231]), .Z(n12655) );
  NAND U14537 ( .A(n12656), .B(n12655), .Z(n12698) );
  XOR U14538 ( .A(a[228]), .B(n42085), .Z(n12694) );
  AND U14539 ( .A(a[224]), .B(b[7]), .Z(n12695) );
  XNOR U14540 ( .A(n12696), .B(n12695), .Z(n12697) );
  XNOR U14541 ( .A(n12698), .B(n12697), .Z(n12703) );
  XOR U14542 ( .A(n12704), .B(n12703), .Z(n12682) );
  NANDN U14543 ( .A(n12659), .B(n12658), .Z(n12663) );
  NANDN U14544 ( .A(n12661), .B(n12660), .Z(n12662) );
  AND U14545 ( .A(n12663), .B(n12662), .Z(n12681) );
  XNOR U14546 ( .A(n12682), .B(n12681), .Z(n12683) );
  NANDN U14547 ( .A(n12665), .B(n12664), .Z(n12669) );
  NAND U14548 ( .A(n12667), .B(n12666), .Z(n12668) );
  NAND U14549 ( .A(n12669), .B(n12668), .Z(n12684) );
  XNOR U14550 ( .A(n12683), .B(n12684), .Z(n12675) );
  XNOR U14551 ( .A(n12676), .B(n12675), .Z(n12677) );
  XNOR U14552 ( .A(n12678), .B(n12677), .Z(n12707) );
  XNOR U14553 ( .A(sreg[1248]), .B(n12707), .Z(n12709) );
  NANDN U14554 ( .A(sreg[1247]), .B(n12670), .Z(n12674) );
  NAND U14555 ( .A(n12672), .B(n12671), .Z(n12673) );
  NAND U14556 ( .A(n12674), .B(n12673), .Z(n12708) );
  XNOR U14557 ( .A(n12709), .B(n12708), .Z(c[1248]) );
  NANDN U14558 ( .A(n12676), .B(n12675), .Z(n12680) );
  NANDN U14559 ( .A(n12678), .B(n12677), .Z(n12679) );
  AND U14560 ( .A(n12680), .B(n12679), .Z(n12715) );
  NANDN U14561 ( .A(n12682), .B(n12681), .Z(n12686) );
  NANDN U14562 ( .A(n12684), .B(n12683), .Z(n12685) );
  AND U14563 ( .A(n12686), .B(n12685), .Z(n12713) );
  NAND U14564 ( .A(n42143), .B(n12687), .Z(n12689) );
  XNOR U14565 ( .A(a[227]), .B(n4104), .Z(n12724) );
  NAND U14566 ( .A(n42144), .B(n12724), .Z(n12688) );
  AND U14567 ( .A(n12689), .B(n12688), .Z(n12739) );
  XOR U14568 ( .A(a[231]), .B(n42012), .Z(n12727) );
  XNOR U14569 ( .A(n12739), .B(n12738), .Z(n12741) );
  AND U14570 ( .A(a[233]), .B(b[0]), .Z(n12691) );
  XNOR U14571 ( .A(n12691), .B(n4071), .Z(n12693) );
  NANDN U14572 ( .A(b[0]), .B(a[232]), .Z(n12692) );
  NAND U14573 ( .A(n12693), .B(n12692), .Z(n12735) );
  XOR U14574 ( .A(a[229]), .B(n42085), .Z(n12731) );
  AND U14575 ( .A(a[225]), .B(b[7]), .Z(n12732) );
  XNOR U14576 ( .A(n12733), .B(n12732), .Z(n12734) );
  XNOR U14577 ( .A(n12735), .B(n12734), .Z(n12740) );
  XOR U14578 ( .A(n12741), .B(n12740), .Z(n12719) );
  NANDN U14579 ( .A(n12696), .B(n12695), .Z(n12700) );
  NANDN U14580 ( .A(n12698), .B(n12697), .Z(n12699) );
  AND U14581 ( .A(n12700), .B(n12699), .Z(n12718) );
  XNOR U14582 ( .A(n12719), .B(n12718), .Z(n12720) );
  NANDN U14583 ( .A(n12702), .B(n12701), .Z(n12706) );
  NAND U14584 ( .A(n12704), .B(n12703), .Z(n12705) );
  NAND U14585 ( .A(n12706), .B(n12705), .Z(n12721) );
  XNOR U14586 ( .A(n12720), .B(n12721), .Z(n12712) );
  XNOR U14587 ( .A(n12713), .B(n12712), .Z(n12714) );
  XNOR U14588 ( .A(n12715), .B(n12714), .Z(n12744) );
  XNOR U14589 ( .A(sreg[1249]), .B(n12744), .Z(n12746) );
  NANDN U14590 ( .A(sreg[1248]), .B(n12707), .Z(n12711) );
  NAND U14591 ( .A(n12709), .B(n12708), .Z(n12710) );
  NAND U14592 ( .A(n12711), .B(n12710), .Z(n12745) );
  XNOR U14593 ( .A(n12746), .B(n12745), .Z(c[1249]) );
  NANDN U14594 ( .A(n12713), .B(n12712), .Z(n12717) );
  NANDN U14595 ( .A(n12715), .B(n12714), .Z(n12716) );
  AND U14596 ( .A(n12717), .B(n12716), .Z(n12752) );
  NANDN U14597 ( .A(n12719), .B(n12718), .Z(n12723) );
  NANDN U14598 ( .A(n12721), .B(n12720), .Z(n12722) );
  AND U14599 ( .A(n12723), .B(n12722), .Z(n12750) );
  NAND U14600 ( .A(n42143), .B(n12724), .Z(n12726) );
  XNOR U14601 ( .A(a[228]), .B(n4104), .Z(n12761) );
  NAND U14602 ( .A(n42144), .B(n12761), .Z(n12725) );
  AND U14603 ( .A(n12726), .B(n12725), .Z(n12776) );
  XOR U14604 ( .A(a[232]), .B(n42012), .Z(n12764) );
  XNOR U14605 ( .A(n12776), .B(n12775), .Z(n12778) );
  AND U14606 ( .A(a[234]), .B(b[0]), .Z(n12728) );
  XNOR U14607 ( .A(n12728), .B(n4071), .Z(n12730) );
  NANDN U14608 ( .A(b[0]), .B(a[233]), .Z(n12729) );
  NAND U14609 ( .A(n12730), .B(n12729), .Z(n12772) );
  XOR U14610 ( .A(a[230]), .B(n42085), .Z(n12768) );
  AND U14611 ( .A(a[226]), .B(b[7]), .Z(n12769) );
  XNOR U14612 ( .A(n12770), .B(n12769), .Z(n12771) );
  XNOR U14613 ( .A(n12772), .B(n12771), .Z(n12777) );
  XOR U14614 ( .A(n12778), .B(n12777), .Z(n12756) );
  NANDN U14615 ( .A(n12733), .B(n12732), .Z(n12737) );
  NANDN U14616 ( .A(n12735), .B(n12734), .Z(n12736) );
  AND U14617 ( .A(n12737), .B(n12736), .Z(n12755) );
  XNOR U14618 ( .A(n12756), .B(n12755), .Z(n12757) );
  NANDN U14619 ( .A(n12739), .B(n12738), .Z(n12743) );
  NAND U14620 ( .A(n12741), .B(n12740), .Z(n12742) );
  NAND U14621 ( .A(n12743), .B(n12742), .Z(n12758) );
  XNOR U14622 ( .A(n12757), .B(n12758), .Z(n12749) );
  XNOR U14623 ( .A(n12750), .B(n12749), .Z(n12751) );
  XNOR U14624 ( .A(n12752), .B(n12751), .Z(n12781) );
  XNOR U14625 ( .A(sreg[1250]), .B(n12781), .Z(n12783) );
  NANDN U14626 ( .A(sreg[1249]), .B(n12744), .Z(n12748) );
  NAND U14627 ( .A(n12746), .B(n12745), .Z(n12747) );
  NAND U14628 ( .A(n12748), .B(n12747), .Z(n12782) );
  XNOR U14629 ( .A(n12783), .B(n12782), .Z(c[1250]) );
  NANDN U14630 ( .A(n12750), .B(n12749), .Z(n12754) );
  NANDN U14631 ( .A(n12752), .B(n12751), .Z(n12753) );
  AND U14632 ( .A(n12754), .B(n12753), .Z(n12789) );
  NANDN U14633 ( .A(n12756), .B(n12755), .Z(n12760) );
  NANDN U14634 ( .A(n12758), .B(n12757), .Z(n12759) );
  AND U14635 ( .A(n12760), .B(n12759), .Z(n12787) );
  NAND U14636 ( .A(n42143), .B(n12761), .Z(n12763) );
  XNOR U14637 ( .A(a[229]), .B(n4104), .Z(n12798) );
  NAND U14638 ( .A(n42144), .B(n12798), .Z(n12762) );
  AND U14639 ( .A(n12763), .B(n12762), .Z(n12813) );
  XOR U14640 ( .A(a[233]), .B(n42012), .Z(n12801) );
  XNOR U14641 ( .A(n12813), .B(n12812), .Z(n12815) );
  AND U14642 ( .A(a[235]), .B(b[0]), .Z(n12765) );
  XNOR U14643 ( .A(n12765), .B(n4071), .Z(n12767) );
  NANDN U14644 ( .A(b[0]), .B(a[234]), .Z(n12766) );
  NAND U14645 ( .A(n12767), .B(n12766), .Z(n12809) );
  XOR U14646 ( .A(a[231]), .B(n42085), .Z(n12805) );
  AND U14647 ( .A(a[227]), .B(b[7]), .Z(n12806) );
  XNOR U14648 ( .A(n12807), .B(n12806), .Z(n12808) );
  XNOR U14649 ( .A(n12809), .B(n12808), .Z(n12814) );
  XOR U14650 ( .A(n12815), .B(n12814), .Z(n12793) );
  NANDN U14651 ( .A(n12770), .B(n12769), .Z(n12774) );
  NANDN U14652 ( .A(n12772), .B(n12771), .Z(n12773) );
  AND U14653 ( .A(n12774), .B(n12773), .Z(n12792) );
  XNOR U14654 ( .A(n12793), .B(n12792), .Z(n12794) );
  NANDN U14655 ( .A(n12776), .B(n12775), .Z(n12780) );
  NAND U14656 ( .A(n12778), .B(n12777), .Z(n12779) );
  NAND U14657 ( .A(n12780), .B(n12779), .Z(n12795) );
  XNOR U14658 ( .A(n12794), .B(n12795), .Z(n12786) );
  XNOR U14659 ( .A(n12787), .B(n12786), .Z(n12788) );
  XNOR U14660 ( .A(n12789), .B(n12788), .Z(n12818) );
  XNOR U14661 ( .A(sreg[1251]), .B(n12818), .Z(n12820) );
  NANDN U14662 ( .A(sreg[1250]), .B(n12781), .Z(n12785) );
  NAND U14663 ( .A(n12783), .B(n12782), .Z(n12784) );
  NAND U14664 ( .A(n12785), .B(n12784), .Z(n12819) );
  XNOR U14665 ( .A(n12820), .B(n12819), .Z(c[1251]) );
  NANDN U14666 ( .A(n12787), .B(n12786), .Z(n12791) );
  NANDN U14667 ( .A(n12789), .B(n12788), .Z(n12790) );
  AND U14668 ( .A(n12791), .B(n12790), .Z(n12826) );
  NANDN U14669 ( .A(n12793), .B(n12792), .Z(n12797) );
  NANDN U14670 ( .A(n12795), .B(n12794), .Z(n12796) );
  AND U14671 ( .A(n12797), .B(n12796), .Z(n12824) );
  NAND U14672 ( .A(n42143), .B(n12798), .Z(n12800) );
  XNOR U14673 ( .A(a[230]), .B(n4104), .Z(n12835) );
  NAND U14674 ( .A(n42144), .B(n12835), .Z(n12799) );
  AND U14675 ( .A(n12800), .B(n12799), .Z(n12850) );
  XOR U14676 ( .A(a[234]), .B(n42012), .Z(n12838) );
  XNOR U14677 ( .A(n12850), .B(n12849), .Z(n12852) );
  AND U14678 ( .A(a[236]), .B(b[0]), .Z(n12802) );
  XNOR U14679 ( .A(n12802), .B(n4071), .Z(n12804) );
  NANDN U14680 ( .A(b[0]), .B(a[235]), .Z(n12803) );
  NAND U14681 ( .A(n12804), .B(n12803), .Z(n12846) );
  XOR U14682 ( .A(a[232]), .B(n42085), .Z(n12842) );
  AND U14683 ( .A(a[228]), .B(b[7]), .Z(n12843) );
  XNOR U14684 ( .A(n12844), .B(n12843), .Z(n12845) );
  XNOR U14685 ( .A(n12846), .B(n12845), .Z(n12851) );
  XOR U14686 ( .A(n12852), .B(n12851), .Z(n12830) );
  NANDN U14687 ( .A(n12807), .B(n12806), .Z(n12811) );
  NANDN U14688 ( .A(n12809), .B(n12808), .Z(n12810) );
  AND U14689 ( .A(n12811), .B(n12810), .Z(n12829) );
  XNOR U14690 ( .A(n12830), .B(n12829), .Z(n12831) );
  NANDN U14691 ( .A(n12813), .B(n12812), .Z(n12817) );
  NAND U14692 ( .A(n12815), .B(n12814), .Z(n12816) );
  NAND U14693 ( .A(n12817), .B(n12816), .Z(n12832) );
  XNOR U14694 ( .A(n12831), .B(n12832), .Z(n12823) );
  XNOR U14695 ( .A(n12824), .B(n12823), .Z(n12825) );
  XNOR U14696 ( .A(n12826), .B(n12825), .Z(n12855) );
  XNOR U14697 ( .A(sreg[1252]), .B(n12855), .Z(n12857) );
  NANDN U14698 ( .A(sreg[1251]), .B(n12818), .Z(n12822) );
  NAND U14699 ( .A(n12820), .B(n12819), .Z(n12821) );
  NAND U14700 ( .A(n12822), .B(n12821), .Z(n12856) );
  XNOR U14701 ( .A(n12857), .B(n12856), .Z(c[1252]) );
  NANDN U14702 ( .A(n12824), .B(n12823), .Z(n12828) );
  NANDN U14703 ( .A(n12826), .B(n12825), .Z(n12827) );
  AND U14704 ( .A(n12828), .B(n12827), .Z(n12863) );
  NANDN U14705 ( .A(n12830), .B(n12829), .Z(n12834) );
  NANDN U14706 ( .A(n12832), .B(n12831), .Z(n12833) );
  AND U14707 ( .A(n12834), .B(n12833), .Z(n12861) );
  NAND U14708 ( .A(n42143), .B(n12835), .Z(n12837) );
  XNOR U14709 ( .A(a[231]), .B(n4104), .Z(n12872) );
  NAND U14710 ( .A(n42144), .B(n12872), .Z(n12836) );
  AND U14711 ( .A(n12837), .B(n12836), .Z(n12887) );
  XOR U14712 ( .A(a[235]), .B(n42012), .Z(n12875) );
  XNOR U14713 ( .A(n12887), .B(n12886), .Z(n12889) );
  AND U14714 ( .A(a[237]), .B(b[0]), .Z(n12839) );
  XNOR U14715 ( .A(n12839), .B(n4071), .Z(n12841) );
  NANDN U14716 ( .A(b[0]), .B(a[236]), .Z(n12840) );
  NAND U14717 ( .A(n12841), .B(n12840), .Z(n12883) );
  XOR U14718 ( .A(a[233]), .B(n42085), .Z(n12879) );
  AND U14719 ( .A(a[229]), .B(b[7]), .Z(n12880) );
  XNOR U14720 ( .A(n12881), .B(n12880), .Z(n12882) );
  XNOR U14721 ( .A(n12883), .B(n12882), .Z(n12888) );
  XOR U14722 ( .A(n12889), .B(n12888), .Z(n12867) );
  NANDN U14723 ( .A(n12844), .B(n12843), .Z(n12848) );
  NANDN U14724 ( .A(n12846), .B(n12845), .Z(n12847) );
  AND U14725 ( .A(n12848), .B(n12847), .Z(n12866) );
  XNOR U14726 ( .A(n12867), .B(n12866), .Z(n12868) );
  NANDN U14727 ( .A(n12850), .B(n12849), .Z(n12854) );
  NAND U14728 ( .A(n12852), .B(n12851), .Z(n12853) );
  NAND U14729 ( .A(n12854), .B(n12853), .Z(n12869) );
  XNOR U14730 ( .A(n12868), .B(n12869), .Z(n12860) );
  XNOR U14731 ( .A(n12861), .B(n12860), .Z(n12862) );
  XNOR U14732 ( .A(n12863), .B(n12862), .Z(n12892) );
  XNOR U14733 ( .A(sreg[1253]), .B(n12892), .Z(n12894) );
  NANDN U14734 ( .A(sreg[1252]), .B(n12855), .Z(n12859) );
  NAND U14735 ( .A(n12857), .B(n12856), .Z(n12858) );
  NAND U14736 ( .A(n12859), .B(n12858), .Z(n12893) );
  XNOR U14737 ( .A(n12894), .B(n12893), .Z(c[1253]) );
  NANDN U14738 ( .A(n12861), .B(n12860), .Z(n12865) );
  NANDN U14739 ( .A(n12863), .B(n12862), .Z(n12864) );
  AND U14740 ( .A(n12865), .B(n12864), .Z(n12900) );
  NANDN U14741 ( .A(n12867), .B(n12866), .Z(n12871) );
  NANDN U14742 ( .A(n12869), .B(n12868), .Z(n12870) );
  AND U14743 ( .A(n12871), .B(n12870), .Z(n12898) );
  NAND U14744 ( .A(n42143), .B(n12872), .Z(n12874) );
  XNOR U14745 ( .A(a[232]), .B(n4105), .Z(n12909) );
  NAND U14746 ( .A(n42144), .B(n12909), .Z(n12873) );
  AND U14747 ( .A(n12874), .B(n12873), .Z(n12924) );
  XOR U14748 ( .A(a[236]), .B(n42012), .Z(n12912) );
  XNOR U14749 ( .A(n12924), .B(n12923), .Z(n12926) );
  AND U14750 ( .A(a[238]), .B(b[0]), .Z(n12876) );
  XNOR U14751 ( .A(n12876), .B(n4071), .Z(n12878) );
  NANDN U14752 ( .A(b[0]), .B(a[237]), .Z(n12877) );
  NAND U14753 ( .A(n12878), .B(n12877), .Z(n12920) );
  XOR U14754 ( .A(a[234]), .B(n42085), .Z(n12916) );
  AND U14755 ( .A(a[230]), .B(b[7]), .Z(n12917) );
  XNOR U14756 ( .A(n12918), .B(n12917), .Z(n12919) );
  XNOR U14757 ( .A(n12920), .B(n12919), .Z(n12925) );
  XOR U14758 ( .A(n12926), .B(n12925), .Z(n12904) );
  NANDN U14759 ( .A(n12881), .B(n12880), .Z(n12885) );
  NANDN U14760 ( .A(n12883), .B(n12882), .Z(n12884) );
  AND U14761 ( .A(n12885), .B(n12884), .Z(n12903) );
  XNOR U14762 ( .A(n12904), .B(n12903), .Z(n12905) );
  NANDN U14763 ( .A(n12887), .B(n12886), .Z(n12891) );
  NAND U14764 ( .A(n12889), .B(n12888), .Z(n12890) );
  NAND U14765 ( .A(n12891), .B(n12890), .Z(n12906) );
  XNOR U14766 ( .A(n12905), .B(n12906), .Z(n12897) );
  XNOR U14767 ( .A(n12898), .B(n12897), .Z(n12899) );
  XNOR U14768 ( .A(n12900), .B(n12899), .Z(n12929) );
  XNOR U14769 ( .A(sreg[1254]), .B(n12929), .Z(n12931) );
  NANDN U14770 ( .A(sreg[1253]), .B(n12892), .Z(n12896) );
  NAND U14771 ( .A(n12894), .B(n12893), .Z(n12895) );
  NAND U14772 ( .A(n12896), .B(n12895), .Z(n12930) );
  XNOR U14773 ( .A(n12931), .B(n12930), .Z(c[1254]) );
  NANDN U14774 ( .A(n12898), .B(n12897), .Z(n12902) );
  NANDN U14775 ( .A(n12900), .B(n12899), .Z(n12901) );
  AND U14776 ( .A(n12902), .B(n12901), .Z(n12937) );
  NANDN U14777 ( .A(n12904), .B(n12903), .Z(n12908) );
  NANDN U14778 ( .A(n12906), .B(n12905), .Z(n12907) );
  AND U14779 ( .A(n12908), .B(n12907), .Z(n12935) );
  NAND U14780 ( .A(n42143), .B(n12909), .Z(n12911) );
  XNOR U14781 ( .A(a[233]), .B(n4105), .Z(n12946) );
  NAND U14782 ( .A(n42144), .B(n12946), .Z(n12910) );
  AND U14783 ( .A(n12911), .B(n12910), .Z(n12961) );
  XOR U14784 ( .A(a[237]), .B(n42012), .Z(n12949) );
  XNOR U14785 ( .A(n12961), .B(n12960), .Z(n12963) );
  AND U14786 ( .A(a[239]), .B(b[0]), .Z(n12913) );
  XNOR U14787 ( .A(n12913), .B(n4071), .Z(n12915) );
  NANDN U14788 ( .A(b[0]), .B(a[238]), .Z(n12914) );
  NAND U14789 ( .A(n12915), .B(n12914), .Z(n12957) );
  XOR U14790 ( .A(a[235]), .B(n42085), .Z(n12950) );
  AND U14791 ( .A(a[231]), .B(b[7]), .Z(n12954) );
  XNOR U14792 ( .A(n12955), .B(n12954), .Z(n12956) );
  XNOR U14793 ( .A(n12957), .B(n12956), .Z(n12962) );
  XOR U14794 ( .A(n12963), .B(n12962), .Z(n12941) );
  NANDN U14795 ( .A(n12918), .B(n12917), .Z(n12922) );
  NANDN U14796 ( .A(n12920), .B(n12919), .Z(n12921) );
  AND U14797 ( .A(n12922), .B(n12921), .Z(n12940) );
  XNOR U14798 ( .A(n12941), .B(n12940), .Z(n12942) );
  NANDN U14799 ( .A(n12924), .B(n12923), .Z(n12928) );
  NAND U14800 ( .A(n12926), .B(n12925), .Z(n12927) );
  NAND U14801 ( .A(n12928), .B(n12927), .Z(n12943) );
  XNOR U14802 ( .A(n12942), .B(n12943), .Z(n12934) );
  XNOR U14803 ( .A(n12935), .B(n12934), .Z(n12936) );
  XNOR U14804 ( .A(n12937), .B(n12936), .Z(n12966) );
  XNOR U14805 ( .A(sreg[1255]), .B(n12966), .Z(n12968) );
  NANDN U14806 ( .A(sreg[1254]), .B(n12929), .Z(n12933) );
  NAND U14807 ( .A(n12931), .B(n12930), .Z(n12932) );
  NAND U14808 ( .A(n12933), .B(n12932), .Z(n12967) );
  XNOR U14809 ( .A(n12968), .B(n12967), .Z(c[1255]) );
  NANDN U14810 ( .A(n12935), .B(n12934), .Z(n12939) );
  NANDN U14811 ( .A(n12937), .B(n12936), .Z(n12938) );
  AND U14812 ( .A(n12939), .B(n12938), .Z(n12974) );
  NANDN U14813 ( .A(n12941), .B(n12940), .Z(n12945) );
  NANDN U14814 ( .A(n12943), .B(n12942), .Z(n12944) );
  AND U14815 ( .A(n12945), .B(n12944), .Z(n12972) );
  NAND U14816 ( .A(n42143), .B(n12946), .Z(n12948) );
  XNOR U14817 ( .A(a[234]), .B(n4105), .Z(n12983) );
  NAND U14818 ( .A(n42144), .B(n12983), .Z(n12947) );
  AND U14819 ( .A(n12948), .B(n12947), .Z(n12998) );
  XOR U14820 ( .A(a[238]), .B(n42012), .Z(n12986) );
  XNOR U14821 ( .A(n12998), .B(n12997), .Z(n13000) );
  XOR U14822 ( .A(a[236]), .B(n42085), .Z(n12990) );
  AND U14823 ( .A(a[232]), .B(b[7]), .Z(n12991) );
  XNOR U14824 ( .A(n12992), .B(n12991), .Z(n12993) );
  AND U14825 ( .A(a[240]), .B(b[0]), .Z(n12951) );
  XNOR U14826 ( .A(n12951), .B(n4071), .Z(n12953) );
  NANDN U14827 ( .A(b[0]), .B(a[239]), .Z(n12952) );
  NAND U14828 ( .A(n12953), .B(n12952), .Z(n12994) );
  XNOR U14829 ( .A(n12993), .B(n12994), .Z(n12999) );
  XOR U14830 ( .A(n13000), .B(n12999), .Z(n12978) );
  NANDN U14831 ( .A(n12955), .B(n12954), .Z(n12959) );
  NANDN U14832 ( .A(n12957), .B(n12956), .Z(n12958) );
  AND U14833 ( .A(n12959), .B(n12958), .Z(n12977) );
  XNOR U14834 ( .A(n12978), .B(n12977), .Z(n12979) );
  NANDN U14835 ( .A(n12961), .B(n12960), .Z(n12965) );
  NAND U14836 ( .A(n12963), .B(n12962), .Z(n12964) );
  NAND U14837 ( .A(n12965), .B(n12964), .Z(n12980) );
  XNOR U14838 ( .A(n12979), .B(n12980), .Z(n12971) );
  XNOR U14839 ( .A(n12972), .B(n12971), .Z(n12973) );
  XNOR U14840 ( .A(n12974), .B(n12973), .Z(n13003) );
  XNOR U14841 ( .A(sreg[1256]), .B(n13003), .Z(n13005) );
  NANDN U14842 ( .A(sreg[1255]), .B(n12966), .Z(n12970) );
  NAND U14843 ( .A(n12968), .B(n12967), .Z(n12969) );
  NAND U14844 ( .A(n12970), .B(n12969), .Z(n13004) );
  XNOR U14845 ( .A(n13005), .B(n13004), .Z(c[1256]) );
  NANDN U14846 ( .A(n12972), .B(n12971), .Z(n12976) );
  NANDN U14847 ( .A(n12974), .B(n12973), .Z(n12975) );
  AND U14848 ( .A(n12976), .B(n12975), .Z(n13011) );
  NANDN U14849 ( .A(n12978), .B(n12977), .Z(n12982) );
  NANDN U14850 ( .A(n12980), .B(n12979), .Z(n12981) );
  AND U14851 ( .A(n12982), .B(n12981), .Z(n13009) );
  NAND U14852 ( .A(n42143), .B(n12983), .Z(n12985) );
  XNOR U14853 ( .A(a[235]), .B(n4105), .Z(n13020) );
  NAND U14854 ( .A(n42144), .B(n13020), .Z(n12984) );
  AND U14855 ( .A(n12985), .B(n12984), .Z(n13035) );
  XOR U14856 ( .A(a[239]), .B(n42012), .Z(n13023) );
  XNOR U14857 ( .A(n13035), .B(n13034), .Z(n13037) );
  AND U14858 ( .A(a[241]), .B(b[0]), .Z(n12987) );
  XNOR U14859 ( .A(n12987), .B(n4071), .Z(n12989) );
  NANDN U14860 ( .A(b[0]), .B(a[240]), .Z(n12988) );
  NAND U14861 ( .A(n12989), .B(n12988), .Z(n13031) );
  XOR U14862 ( .A(a[237]), .B(n42085), .Z(n13024) );
  AND U14863 ( .A(a[233]), .B(b[7]), .Z(n13028) );
  XNOR U14864 ( .A(n13029), .B(n13028), .Z(n13030) );
  XNOR U14865 ( .A(n13031), .B(n13030), .Z(n13036) );
  XOR U14866 ( .A(n13037), .B(n13036), .Z(n13015) );
  NANDN U14867 ( .A(n12992), .B(n12991), .Z(n12996) );
  NANDN U14868 ( .A(n12994), .B(n12993), .Z(n12995) );
  AND U14869 ( .A(n12996), .B(n12995), .Z(n13014) );
  XNOR U14870 ( .A(n13015), .B(n13014), .Z(n13016) );
  NANDN U14871 ( .A(n12998), .B(n12997), .Z(n13002) );
  NAND U14872 ( .A(n13000), .B(n12999), .Z(n13001) );
  NAND U14873 ( .A(n13002), .B(n13001), .Z(n13017) );
  XNOR U14874 ( .A(n13016), .B(n13017), .Z(n13008) );
  XNOR U14875 ( .A(n13009), .B(n13008), .Z(n13010) );
  XNOR U14876 ( .A(n13011), .B(n13010), .Z(n13040) );
  XNOR U14877 ( .A(sreg[1257]), .B(n13040), .Z(n13042) );
  NANDN U14878 ( .A(sreg[1256]), .B(n13003), .Z(n13007) );
  NAND U14879 ( .A(n13005), .B(n13004), .Z(n13006) );
  NAND U14880 ( .A(n13007), .B(n13006), .Z(n13041) );
  XNOR U14881 ( .A(n13042), .B(n13041), .Z(c[1257]) );
  NANDN U14882 ( .A(n13009), .B(n13008), .Z(n13013) );
  NANDN U14883 ( .A(n13011), .B(n13010), .Z(n13012) );
  AND U14884 ( .A(n13013), .B(n13012), .Z(n13048) );
  NANDN U14885 ( .A(n13015), .B(n13014), .Z(n13019) );
  NANDN U14886 ( .A(n13017), .B(n13016), .Z(n13018) );
  AND U14887 ( .A(n13019), .B(n13018), .Z(n13046) );
  NAND U14888 ( .A(n42143), .B(n13020), .Z(n13022) );
  XNOR U14889 ( .A(a[236]), .B(n4105), .Z(n13057) );
  NAND U14890 ( .A(n42144), .B(n13057), .Z(n13021) );
  AND U14891 ( .A(n13022), .B(n13021), .Z(n13072) );
  XOR U14892 ( .A(a[240]), .B(n42012), .Z(n13060) );
  XNOR U14893 ( .A(n13072), .B(n13071), .Z(n13074) );
  XOR U14894 ( .A(a[238]), .B(n42085), .Z(n13064) );
  AND U14895 ( .A(a[234]), .B(b[7]), .Z(n13065) );
  XNOR U14896 ( .A(n13066), .B(n13065), .Z(n13067) );
  AND U14897 ( .A(a[242]), .B(b[0]), .Z(n13025) );
  XNOR U14898 ( .A(n13025), .B(n4071), .Z(n13027) );
  NANDN U14899 ( .A(b[0]), .B(a[241]), .Z(n13026) );
  NAND U14900 ( .A(n13027), .B(n13026), .Z(n13068) );
  XNOR U14901 ( .A(n13067), .B(n13068), .Z(n13073) );
  XOR U14902 ( .A(n13074), .B(n13073), .Z(n13052) );
  NANDN U14903 ( .A(n13029), .B(n13028), .Z(n13033) );
  NANDN U14904 ( .A(n13031), .B(n13030), .Z(n13032) );
  AND U14905 ( .A(n13033), .B(n13032), .Z(n13051) );
  XNOR U14906 ( .A(n13052), .B(n13051), .Z(n13053) );
  NANDN U14907 ( .A(n13035), .B(n13034), .Z(n13039) );
  NAND U14908 ( .A(n13037), .B(n13036), .Z(n13038) );
  NAND U14909 ( .A(n13039), .B(n13038), .Z(n13054) );
  XNOR U14910 ( .A(n13053), .B(n13054), .Z(n13045) );
  XNOR U14911 ( .A(n13046), .B(n13045), .Z(n13047) );
  XNOR U14912 ( .A(n13048), .B(n13047), .Z(n13077) );
  XNOR U14913 ( .A(sreg[1258]), .B(n13077), .Z(n13079) );
  NANDN U14914 ( .A(sreg[1257]), .B(n13040), .Z(n13044) );
  NAND U14915 ( .A(n13042), .B(n13041), .Z(n13043) );
  NAND U14916 ( .A(n13044), .B(n13043), .Z(n13078) );
  XNOR U14917 ( .A(n13079), .B(n13078), .Z(c[1258]) );
  NANDN U14918 ( .A(n13046), .B(n13045), .Z(n13050) );
  NANDN U14919 ( .A(n13048), .B(n13047), .Z(n13049) );
  AND U14920 ( .A(n13050), .B(n13049), .Z(n13085) );
  NANDN U14921 ( .A(n13052), .B(n13051), .Z(n13056) );
  NANDN U14922 ( .A(n13054), .B(n13053), .Z(n13055) );
  AND U14923 ( .A(n13056), .B(n13055), .Z(n13083) );
  NAND U14924 ( .A(n42143), .B(n13057), .Z(n13059) );
  XNOR U14925 ( .A(a[237]), .B(n4105), .Z(n13094) );
  NAND U14926 ( .A(n42144), .B(n13094), .Z(n13058) );
  AND U14927 ( .A(n13059), .B(n13058), .Z(n13109) );
  XOR U14928 ( .A(a[241]), .B(n42012), .Z(n13097) );
  XNOR U14929 ( .A(n13109), .B(n13108), .Z(n13111) );
  AND U14930 ( .A(b[0]), .B(a[243]), .Z(n13061) );
  XOR U14931 ( .A(b[1]), .B(n13061), .Z(n13063) );
  NANDN U14932 ( .A(b[0]), .B(a[242]), .Z(n13062) );
  AND U14933 ( .A(n13063), .B(n13062), .Z(n13104) );
  XOR U14934 ( .A(a[239]), .B(n42085), .Z(n13101) );
  AND U14935 ( .A(a[235]), .B(b[7]), .Z(n13102) );
  XOR U14936 ( .A(n13103), .B(n13102), .Z(n13105) );
  XNOR U14937 ( .A(n13104), .B(n13105), .Z(n13110) );
  XOR U14938 ( .A(n13111), .B(n13110), .Z(n13089) );
  NANDN U14939 ( .A(n13066), .B(n13065), .Z(n13070) );
  NANDN U14940 ( .A(n13068), .B(n13067), .Z(n13069) );
  AND U14941 ( .A(n13070), .B(n13069), .Z(n13088) );
  XNOR U14942 ( .A(n13089), .B(n13088), .Z(n13090) );
  NANDN U14943 ( .A(n13072), .B(n13071), .Z(n13076) );
  NAND U14944 ( .A(n13074), .B(n13073), .Z(n13075) );
  NAND U14945 ( .A(n13076), .B(n13075), .Z(n13091) );
  XNOR U14946 ( .A(n13090), .B(n13091), .Z(n13082) );
  XNOR U14947 ( .A(n13083), .B(n13082), .Z(n13084) );
  XNOR U14948 ( .A(n13085), .B(n13084), .Z(n13114) );
  XNOR U14949 ( .A(sreg[1259]), .B(n13114), .Z(n13116) );
  NANDN U14950 ( .A(sreg[1258]), .B(n13077), .Z(n13081) );
  NAND U14951 ( .A(n13079), .B(n13078), .Z(n13080) );
  NAND U14952 ( .A(n13081), .B(n13080), .Z(n13115) );
  XNOR U14953 ( .A(n13116), .B(n13115), .Z(c[1259]) );
  NANDN U14954 ( .A(n13083), .B(n13082), .Z(n13087) );
  NANDN U14955 ( .A(n13085), .B(n13084), .Z(n13086) );
  AND U14956 ( .A(n13087), .B(n13086), .Z(n13122) );
  NANDN U14957 ( .A(n13089), .B(n13088), .Z(n13093) );
  NANDN U14958 ( .A(n13091), .B(n13090), .Z(n13092) );
  AND U14959 ( .A(n13093), .B(n13092), .Z(n13120) );
  NAND U14960 ( .A(n42143), .B(n13094), .Z(n13096) );
  XNOR U14961 ( .A(a[238]), .B(n4105), .Z(n13131) );
  NAND U14962 ( .A(n42144), .B(n13131), .Z(n13095) );
  AND U14963 ( .A(n13096), .B(n13095), .Z(n13146) );
  XOR U14964 ( .A(a[242]), .B(n42012), .Z(n13134) );
  XNOR U14965 ( .A(n13146), .B(n13145), .Z(n13148) );
  AND U14966 ( .A(a[244]), .B(b[0]), .Z(n13098) );
  XNOR U14967 ( .A(n13098), .B(n4071), .Z(n13100) );
  NANDN U14968 ( .A(b[0]), .B(a[243]), .Z(n13099) );
  NAND U14969 ( .A(n13100), .B(n13099), .Z(n13142) );
  XOR U14970 ( .A(a[240]), .B(n42085), .Z(n13138) );
  AND U14971 ( .A(a[236]), .B(b[7]), .Z(n13139) );
  XNOR U14972 ( .A(n13140), .B(n13139), .Z(n13141) );
  XNOR U14973 ( .A(n13142), .B(n13141), .Z(n13147) );
  XOR U14974 ( .A(n13148), .B(n13147), .Z(n13126) );
  NANDN U14975 ( .A(n13103), .B(n13102), .Z(n13107) );
  NANDN U14976 ( .A(n13105), .B(n13104), .Z(n13106) );
  AND U14977 ( .A(n13107), .B(n13106), .Z(n13125) );
  XNOR U14978 ( .A(n13126), .B(n13125), .Z(n13127) );
  NANDN U14979 ( .A(n13109), .B(n13108), .Z(n13113) );
  NAND U14980 ( .A(n13111), .B(n13110), .Z(n13112) );
  NAND U14981 ( .A(n13113), .B(n13112), .Z(n13128) );
  XNOR U14982 ( .A(n13127), .B(n13128), .Z(n13119) );
  XNOR U14983 ( .A(n13120), .B(n13119), .Z(n13121) );
  XNOR U14984 ( .A(n13122), .B(n13121), .Z(n13151) );
  XNOR U14985 ( .A(sreg[1260]), .B(n13151), .Z(n13153) );
  NANDN U14986 ( .A(sreg[1259]), .B(n13114), .Z(n13118) );
  NAND U14987 ( .A(n13116), .B(n13115), .Z(n13117) );
  NAND U14988 ( .A(n13118), .B(n13117), .Z(n13152) );
  XNOR U14989 ( .A(n13153), .B(n13152), .Z(c[1260]) );
  NANDN U14990 ( .A(n13120), .B(n13119), .Z(n13124) );
  NANDN U14991 ( .A(n13122), .B(n13121), .Z(n13123) );
  AND U14992 ( .A(n13124), .B(n13123), .Z(n13159) );
  NANDN U14993 ( .A(n13126), .B(n13125), .Z(n13130) );
  NANDN U14994 ( .A(n13128), .B(n13127), .Z(n13129) );
  AND U14995 ( .A(n13130), .B(n13129), .Z(n13157) );
  NAND U14996 ( .A(n42143), .B(n13131), .Z(n13133) );
  XNOR U14997 ( .A(a[239]), .B(n4106), .Z(n13168) );
  NAND U14998 ( .A(n42144), .B(n13168), .Z(n13132) );
  AND U14999 ( .A(n13133), .B(n13132), .Z(n13183) );
  XOR U15000 ( .A(a[243]), .B(n42012), .Z(n13171) );
  XNOR U15001 ( .A(n13183), .B(n13182), .Z(n13185) );
  AND U15002 ( .A(a[245]), .B(b[0]), .Z(n13135) );
  XNOR U15003 ( .A(n13135), .B(n4071), .Z(n13137) );
  NANDN U15004 ( .A(b[0]), .B(a[244]), .Z(n13136) );
  NAND U15005 ( .A(n13137), .B(n13136), .Z(n13179) );
  XOR U15006 ( .A(a[241]), .B(n42085), .Z(n13175) );
  AND U15007 ( .A(a[237]), .B(b[7]), .Z(n13176) );
  XNOR U15008 ( .A(n13177), .B(n13176), .Z(n13178) );
  XNOR U15009 ( .A(n13179), .B(n13178), .Z(n13184) );
  XOR U15010 ( .A(n13185), .B(n13184), .Z(n13163) );
  NANDN U15011 ( .A(n13140), .B(n13139), .Z(n13144) );
  NANDN U15012 ( .A(n13142), .B(n13141), .Z(n13143) );
  AND U15013 ( .A(n13144), .B(n13143), .Z(n13162) );
  XNOR U15014 ( .A(n13163), .B(n13162), .Z(n13164) );
  NANDN U15015 ( .A(n13146), .B(n13145), .Z(n13150) );
  NAND U15016 ( .A(n13148), .B(n13147), .Z(n13149) );
  NAND U15017 ( .A(n13150), .B(n13149), .Z(n13165) );
  XNOR U15018 ( .A(n13164), .B(n13165), .Z(n13156) );
  XNOR U15019 ( .A(n13157), .B(n13156), .Z(n13158) );
  XNOR U15020 ( .A(n13159), .B(n13158), .Z(n13188) );
  XNOR U15021 ( .A(sreg[1261]), .B(n13188), .Z(n13190) );
  NANDN U15022 ( .A(sreg[1260]), .B(n13151), .Z(n13155) );
  NAND U15023 ( .A(n13153), .B(n13152), .Z(n13154) );
  NAND U15024 ( .A(n13155), .B(n13154), .Z(n13189) );
  XNOR U15025 ( .A(n13190), .B(n13189), .Z(c[1261]) );
  NANDN U15026 ( .A(n13157), .B(n13156), .Z(n13161) );
  NANDN U15027 ( .A(n13159), .B(n13158), .Z(n13160) );
  AND U15028 ( .A(n13161), .B(n13160), .Z(n13196) );
  NANDN U15029 ( .A(n13163), .B(n13162), .Z(n13167) );
  NANDN U15030 ( .A(n13165), .B(n13164), .Z(n13166) );
  AND U15031 ( .A(n13167), .B(n13166), .Z(n13194) );
  NAND U15032 ( .A(n42143), .B(n13168), .Z(n13170) );
  XNOR U15033 ( .A(a[240]), .B(n4106), .Z(n13205) );
  NAND U15034 ( .A(n42144), .B(n13205), .Z(n13169) );
  AND U15035 ( .A(n13170), .B(n13169), .Z(n13220) );
  XOR U15036 ( .A(a[244]), .B(n42012), .Z(n13208) );
  XNOR U15037 ( .A(n13220), .B(n13219), .Z(n13222) );
  AND U15038 ( .A(a[246]), .B(b[0]), .Z(n13172) );
  XNOR U15039 ( .A(n13172), .B(n4071), .Z(n13174) );
  NANDN U15040 ( .A(b[0]), .B(a[245]), .Z(n13173) );
  NAND U15041 ( .A(n13174), .B(n13173), .Z(n13216) );
  XOR U15042 ( .A(a[242]), .B(n42085), .Z(n13212) );
  AND U15043 ( .A(a[238]), .B(b[7]), .Z(n13213) );
  XNOR U15044 ( .A(n13214), .B(n13213), .Z(n13215) );
  XNOR U15045 ( .A(n13216), .B(n13215), .Z(n13221) );
  XOR U15046 ( .A(n13222), .B(n13221), .Z(n13200) );
  NANDN U15047 ( .A(n13177), .B(n13176), .Z(n13181) );
  NANDN U15048 ( .A(n13179), .B(n13178), .Z(n13180) );
  AND U15049 ( .A(n13181), .B(n13180), .Z(n13199) );
  XNOR U15050 ( .A(n13200), .B(n13199), .Z(n13201) );
  NANDN U15051 ( .A(n13183), .B(n13182), .Z(n13187) );
  NAND U15052 ( .A(n13185), .B(n13184), .Z(n13186) );
  NAND U15053 ( .A(n13187), .B(n13186), .Z(n13202) );
  XNOR U15054 ( .A(n13201), .B(n13202), .Z(n13193) );
  XNOR U15055 ( .A(n13194), .B(n13193), .Z(n13195) );
  XNOR U15056 ( .A(n13196), .B(n13195), .Z(n13225) );
  XNOR U15057 ( .A(sreg[1262]), .B(n13225), .Z(n13227) );
  NANDN U15058 ( .A(sreg[1261]), .B(n13188), .Z(n13192) );
  NAND U15059 ( .A(n13190), .B(n13189), .Z(n13191) );
  NAND U15060 ( .A(n13192), .B(n13191), .Z(n13226) );
  XNOR U15061 ( .A(n13227), .B(n13226), .Z(c[1262]) );
  NANDN U15062 ( .A(n13194), .B(n13193), .Z(n13198) );
  NANDN U15063 ( .A(n13196), .B(n13195), .Z(n13197) );
  AND U15064 ( .A(n13198), .B(n13197), .Z(n13233) );
  NANDN U15065 ( .A(n13200), .B(n13199), .Z(n13204) );
  NANDN U15066 ( .A(n13202), .B(n13201), .Z(n13203) );
  AND U15067 ( .A(n13204), .B(n13203), .Z(n13231) );
  NAND U15068 ( .A(n42143), .B(n13205), .Z(n13207) );
  XNOR U15069 ( .A(a[241]), .B(n4106), .Z(n13242) );
  NAND U15070 ( .A(n42144), .B(n13242), .Z(n13206) );
  AND U15071 ( .A(n13207), .B(n13206), .Z(n13257) );
  XOR U15072 ( .A(a[245]), .B(n42012), .Z(n13245) );
  XNOR U15073 ( .A(n13257), .B(n13256), .Z(n13259) );
  AND U15074 ( .A(a[247]), .B(b[0]), .Z(n13209) );
  XNOR U15075 ( .A(n13209), .B(n4071), .Z(n13211) );
  NANDN U15076 ( .A(b[0]), .B(a[246]), .Z(n13210) );
  NAND U15077 ( .A(n13211), .B(n13210), .Z(n13253) );
  XOR U15078 ( .A(a[243]), .B(n42085), .Z(n13249) );
  AND U15079 ( .A(a[239]), .B(b[7]), .Z(n13250) );
  XNOR U15080 ( .A(n13251), .B(n13250), .Z(n13252) );
  XNOR U15081 ( .A(n13253), .B(n13252), .Z(n13258) );
  XOR U15082 ( .A(n13259), .B(n13258), .Z(n13237) );
  NANDN U15083 ( .A(n13214), .B(n13213), .Z(n13218) );
  NANDN U15084 ( .A(n13216), .B(n13215), .Z(n13217) );
  AND U15085 ( .A(n13218), .B(n13217), .Z(n13236) );
  XNOR U15086 ( .A(n13237), .B(n13236), .Z(n13238) );
  NANDN U15087 ( .A(n13220), .B(n13219), .Z(n13224) );
  NAND U15088 ( .A(n13222), .B(n13221), .Z(n13223) );
  NAND U15089 ( .A(n13224), .B(n13223), .Z(n13239) );
  XNOR U15090 ( .A(n13238), .B(n13239), .Z(n13230) );
  XNOR U15091 ( .A(n13231), .B(n13230), .Z(n13232) );
  XNOR U15092 ( .A(n13233), .B(n13232), .Z(n13262) );
  XNOR U15093 ( .A(sreg[1263]), .B(n13262), .Z(n13264) );
  NANDN U15094 ( .A(sreg[1262]), .B(n13225), .Z(n13229) );
  NAND U15095 ( .A(n13227), .B(n13226), .Z(n13228) );
  NAND U15096 ( .A(n13229), .B(n13228), .Z(n13263) );
  XNOR U15097 ( .A(n13264), .B(n13263), .Z(c[1263]) );
  NANDN U15098 ( .A(n13231), .B(n13230), .Z(n13235) );
  NANDN U15099 ( .A(n13233), .B(n13232), .Z(n13234) );
  AND U15100 ( .A(n13235), .B(n13234), .Z(n13270) );
  NANDN U15101 ( .A(n13237), .B(n13236), .Z(n13241) );
  NANDN U15102 ( .A(n13239), .B(n13238), .Z(n13240) );
  AND U15103 ( .A(n13241), .B(n13240), .Z(n13268) );
  NAND U15104 ( .A(n42143), .B(n13242), .Z(n13244) );
  XNOR U15105 ( .A(a[242]), .B(n4106), .Z(n13279) );
  NAND U15106 ( .A(n42144), .B(n13279), .Z(n13243) );
  AND U15107 ( .A(n13244), .B(n13243), .Z(n13294) );
  XOR U15108 ( .A(a[246]), .B(n42012), .Z(n13282) );
  XNOR U15109 ( .A(n13294), .B(n13293), .Z(n13296) );
  AND U15110 ( .A(a[248]), .B(b[0]), .Z(n13246) );
  XNOR U15111 ( .A(n13246), .B(n4071), .Z(n13248) );
  NANDN U15112 ( .A(b[0]), .B(a[247]), .Z(n13247) );
  NAND U15113 ( .A(n13248), .B(n13247), .Z(n13290) );
  XOR U15114 ( .A(a[244]), .B(n42085), .Z(n13286) );
  AND U15115 ( .A(a[240]), .B(b[7]), .Z(n13287) );
  XNOR U15116 ( .A(n13288), .B(n13287), .Z(n13289) );
  XNOR U15117 ( .A(n13290), .B(n13289), .Z(n13295) );
  XOR U15118 ( .A(n13296), .B(n13295), .Z(n13274) );
  NANDN U15119 ( .A(n13251), .B(n13250), .Z(n13255) );
  NANDN U15120 ( .A(n13253), .B(n13252), .Z(n13254) );
  AND U15121 ( .A(n13255), .B(n13254), .Z(n13273) );
  XNOR U15122 ( .A(n13274), .B(n13273), .Z(n13275) );
  NANDN U15123 ( .A(n13257), .B(n13256), .Z(n13261) );
  NAND U15124 ( .A(n13259), .B(n13258), .Z(n13260) );
  NAND U15125 ( .A(n13261), .B(n13260), .Z(n13276) );
  XNOR U15126 ( .A(n13275), .B(n13276), .Z(n13267) );
  XNOR U15127 ( .A(n13268), .B(n13267), .Z(n13269) );
  XNOR U15128 ( .A(n13270), .B(n13269), .Z(n13299) );
  XNOR U15129 ( .A(sreg[1264]), .B(n13299), .Z(n13301) );
  NANDN U15130 ( .A(sreg[1263]), .B(n13262), .Z(n13266) );
  NAND U15131 ( .A(n13264), .B(n13263), .Z(n13265) );
  NAND U15132 ( .A(n13266), .B(n13265), .Z(n13300) );
  XNOR U15133 ( .A(n13301), .B(n13300), .Z(c[1264]) );
  NANDN U15134 ( .A(n13268), .B(n13267), .Z(n13272) );
  NANDN U15135 ( .A(n13270), .B(n13269), .Z(n13271) );
  AND U15136 ( .A(n13272), .B(n13271), .Z(n13307) );
  NANDN U15137 ( .A(n13274), .B(n13273), .Z(n13278) );
  NANDN U15138 ( .A(n13276), .B(n13275), .Z(n13277) );
  AND U15139 ( .A(n13278), .B(n13277), .Z(n13305) );
  NAND U15140 ( .A(n42143), .B(n13279), .Z(n13281) );
  XNOR U15141 ( .A(a[243]), .B(n4106), .Z(n13316) );
  NAND U15142 ( .A(n42144), .B(n13316), .Z(n13280) );
  AND U15143 ( .A(n13281), .B(n13280), .Z(n13331) );
  XOR U15144 ( .A(a[247]), .B(n42012), .Z(n13319) );
  XNOR U15145 ( .A(n13331), .B(n13330), .Z(n13333) );
  AND U15146 ( .A(a[249]), .B(b[0]), .Z(n13283) );
  XNOR U15147 ( .A(n13283), .B(n4071), .Z(n13285) );
  NANDN U15148 ( .A(b[0]), .B(a[248]), .Z(n13284) );
  NAND U15149 ( .A(n13285), .B(n13284), .Z(n13327) );
  XOR U15150 ( .A(a[245]), .B(n42085), .Z(n13320) );
  AND U15151 ( .A(a[241]), .B(b[7]), .Z(n13324) );
  XNOR U15152 ( .A(n13325), .B(n13324), .Z(n13326) );
  XNOR U15153 ( .A(n13327), .B(n13326), .Z(n13332) );
  XOR U15154 ( .A(n13333), .B(n13332), .Z(n13311) );
  NANDN U15155 ( .A(n13288), .B(n13287), .Z(n13292) );
  NANDN U15156 ( .A(n13290), .B(n13289), .Z(n13291) );
  AND U15157 ( .A(n13292), .B(n13291), .Z(n13310) );
  XNOR U15158 ( .A(n13311), .B(n13310), .Z(n13312) );
  NANDN U15159 ( .A(n13294), .B(n13293), .Z(n13298) );
  NAND U15160 ( .A(n13296), .B(n13295), .Z(n13297) );
  NAND U15161 ( .A(n13298), .B(n13297), .Z(n13313) );
  XNOR U15162 ( .A(n13312), .B(n13313), .Z(n13304) );
  XNOR U15163 ( .A(n13305), .B(n13304), .Z(n13306) );
  XNOR U15164 ( .A(n13307), .B(n13306), .Z(n13336) );
  XNOR U15165 ( .A(sreg[1265]), .B(n13336), .Z(n13338) );
  NANDN U15166 ( .A(sreg[1264]), .B(n13299), .Z(n13303) );
  NAND U15167 ( .A(n13301), .B(n13300), .Z(n13302) );
  NAND U15168 ( .A(n13303), .B(n13302), .Z(n13337) );
  XNOR U15169 ( .A(n13338), .B(n13337), .Z(c[1265]) );
  NANDN U15170 ( .A(n13305), .B(n13304), .Z(n13309) );
  NANDN U15171 ( .A(n13307), .B(n13306), .Z(n13308) );
  AND U15172 ( .A(n13309), .B(n13308), .Z(n13344) );
  NANDN U15173 ( .A(n13311), .B(n13310), .Z(n13315) );
  NANDN U15174 ( .A(n13313), .B(n13312), .Z(n13314) );
  AND U15175 ( .A(n13315), .B(n13314), .Z(n13342) );
  NAND U15176 ( .A(n42143), .B(n13316), .Z(n13318) );
  XNOR U15177 ( .A(a[244]), .B(n4106), .Z(n13353) );
  NAND U15178 ( .A(n42144), .B(n13353), .Z(n13317) );
  AND U15179 ( .A(n13318), .B(n13317), .Z(n13368) );
  XOR U15180 ( .A(a[248]), .B(n42012), .Z(n13356) );
  XNOR U15181 ( .A(n13368), .B(n13367), .Z(n13370) );
  XOR U15182 ( .A(a[246]), .B(n42085), .Z(n13360) );
  AND U15183 ( .A(a[242]), .B(b[7]), .Z(n13361) );
  XNOR U15184 ( .A(n13362), .B(n13361), .Z(n13363) );
  AND U15185 ( .A(a[250]), .B(b[0]), .Z(n13321) );
  XNOR U15186 ( .A(n13321), .B(n4071), .Z(n13323) );
  NANDN U15187 ( .A(b[0]), .B(a[249]), .Z(n13322) );
  NAND U15188 ( .A(n13323), .B(n13322), .Z(n13364) );
  XNOR U15189 ( .A(n13363), .B(n13364), .Z(n13369) );
  XOR U15190 ( .A(n13370), .B(n13369), .Z(n13348) );
  NANDN U15191 ( .A(n13325), .B(n13324), .Z(n13329) );
  NANDN U15192 ( .A(n13327), .B(n13326), .Z(n13328) );
  AND U15193 ( .A(n13329), .B(n13328), .Z(n13347) );
  XNOR U15194 ( .A(n13348), .B(n13347), .Z(n13349) );
  NANDN U15195 ( .A(n13331), .B(n13330), .Z(n13335) );
  NAND U15196 ( .A(n13333), .B(n13332), .Z(n13334) );
  NAND U15197 ( .A(n13335), .B(n13334), .Z(n13350) );
  XNOR U15198 ( .A(n13349), .B(n13350), .Z(n13341) );
  XNOR U15199 ( .A(n13342), .B(n13341), .Z(n13343) );
  XNOR U15200 ( .A(n13344), .B(n13343), .Z(n13373) );
  XNOR U15201 ( .A(sreg[1266]), .B(n13373), .Z(n13375) );
  NANDN U15202 ( .A(sreg[1265]), .B(n13336), .Z(n13340) );
  NAND U15203 ( .A(n13338), .B(n13337), .Z(n13339) );
  NAND U15204 ( .A(n13340), .B(n13339), .Z(n13374) );
  XNOR U15205 ( .A(n13375), .B(n13374), .Z(c[1266]) );
  NANDN U15206 ( .A(n13342), .B(n13341), .Z(n13346) );
  NANDN U15207 ( .A(n13344), .B(n13343), .Z(n13345) );
  AND U15208 ( .A(n13346), .B(n13345), .Z(n13381) );
  NANDN U15209 ( .A(n13348), .B(n13347), .Z(n13352) );
  NANDN U15210 ( .A(n13350), .B(n13349), .Z(n13351) );
  AND U15211 ( .A(n13352), .B(n13351), .Z(n13379) );
  NAND U15212 ( .A(n42143), .B(n13353), .Z(n13355) );
  XNOR U15213 ( .A(a[245]), .B(n4106), .Z(n13390) );
  NAND U15214 ( .A(n42144), .B(n13390), .Z(n13354) );
  AND U15215 ( .A(n13355), .B(n13354), .Z(n13405) );
  XOR U15216 ( .A(a[249]), .B(n42012), .Z(n13393) );
  XNOR U15217 ( .A(n13405), .B(n13404), .Z(n13407) );
  AND U15218 ( .A(a[251]), .B(b[0]), .Z(n13357) );
  XNOR U15219 ( .A(n13357), .B(n4071), .Z(n13359) );
  NANDN U15220 ( .A(b[0]), .B(a[250]), .Z(n13358) );
  NAND U15221 ( .A(n13359), .B(n13358), .Z(n13401) );
  XOR U15222 ( .A(a[247]), .B(n42085), .Z(n13397) );
  AND U15223 ( .A(a[243]), .B(b[7]), .Z(n13398) );
  XNOR U15224 ( .A(n13399), .B(n13398), .Z(n13400) );
  XNOR U15225 ( .A(n13401), .B(n13400), .Z(n13406) );
  XOR U15226 ( .A(n13407), .B(n13406), .Z(n13385) );
  NANDN U15227 ( .A(n13362), .B(n13361), .Z(n13366) );
  NANDN U15228 ( .A(n13364), .B(n13363), .Z(n13365) );
  AND U15229 ( .A(n13366), .B(n13365), .Z(n13384) );
  XNOR U15230 ( .A(n13385), .B(n13384), .Z(n13386) );
  NANDN U15231 ( .A(n13368), .B(n13367), .Z(n13372) );
  NAND U15232 ( .A(n13370), .B(n13369), .Z(n13371) );
  NAND U15233 ( .A(n13372), .B(n13371), .Z(n13387) );
  XNOR U15234 ( .A(n13386), .B(n13387), .Z(n13378) );
  XNOR U15235 ( .A(n13379), .B(n13378), .Z(n13380) );
  XNOR U15236 ( .A(n13381), .B(n13380), .Z(n13410) );
  XNOR U15237 ( .A(sreg[1267]), .B(n13410), .Z(n13412) );
  NANDN U15238 ( .A(sreg[1266]), .B(n13373), .Z(n13377) );
  NAND U15239 ( .A(n13375), .B(n13374), .Z(n13376) );
  NAND U15240 ( .A(n13377), .B(n13376), .Z(n13411) );
  XNOR U15241 ( .A(n13412), .B(n13411), .Z(c[1267]) );
  NANDN U15242 ( .A(n13379), .B(n13378), .Z(n13383) );
  NANDN U15243 ( .A(n13381), .B(n13380), .Z(n13382) );
  AND U15244 ( .A(n13383), .B(n13382), .Z(n13418) );
  NANDN U15245 ( .A(n13385), .B(n13384), .Z(n13389) );
  NANDN U15246 ( .A(n13387), .B(n13386), .Z(n13388) );
  AND U15247 ( .A(n13389), .B(n13388), .Z(n13416) );
  NAND U15248 ( .A(n42143), .B(n13390), .Z(n13392) );
  XNOR U15249 ( .A(a[246]), .B(n4107), .Z(n13427) );
  NAND U15250 ( .A(n42144), .B(n13427), .Z(n13391) );
  AND U15251 ( .A(n13392), .B(n13391), .Z(n13442) );
  XOR U15252 ( .A(a[250]), .B(n42012), .Z(n13430) );
  XNOR U15253 ( .A(n13442), .B(n13441), .Z(n13444) );
  AND U15254 ( .A(a[252]), .B(b[0]), .Z(n13394) );
  XNOR U15255 ( .A(n13394), .B(n4071), .Z(n13396) );
  NANDN U15256 ( .A(b[0]), .B(a[251]), .Z(n13395) );
  NAND U15257 ( .A(n13396), .B(n13395), .Z(n13438) );
  XOR U15258 ( .A(a[248]), .B(n42085), .Z(n13431) );
  AND U15259 ( .A(a[244]), .B(b[7]), .Z(n13435) );
  XNOR U15260 ( .A(n13436), .B(n13435), .Z(n13437) );
  XNOR U15261 ( .A(n13438), .B(n13437), .Z(n13443) );
  XOR U15262 ( .A(n13444), .B(n13443), .Z(n13422) );
  NANDN U15263 ( .A(n13399), .B(n13398), .Z(n13403) );
  NANDN U15264 ( .A(n13401), .B(n13400), .Z(n13402) );
  AND U15265 ( .A(n13403), .B(n13402), .Z(n13421) );
  XNOR U15266 ( .A(n13422), .B(n13421), .Z(n13423) );
  NANDN U15267 ( .A(n13405), .B(n13404), .Z(n13409) );
  NAND U15268 ( .A(n13407), .B(n13406), .Z(n13408) );
  NAND U15269 ( .A(n13409), .B(n13408), .Z(n13424) );
  XNOR U15270 ( .A(n13423), .B(n13424), .Z(n13415) );
  XNOR U15271 ( .A(n13416), .B(n13415), .Z(n13417) );
  XNOR U15272 ( .A(n13418), .B(n13417), .Z(n13447) );
  XNOR U15273 ( .A(sreg[1268]), .B(n13447), .Z(n13449) );
  NANDN U15274 ( .A(sreg[1267]), .B(n13410), .Z(n13414) );
  NAND U15275 ( .A(n13412), .B(n13411), .Z(n13413) );
  NAND U15276 ( .A(n13414), .B(n13413), .Z(n13448) );
  XNOR U15277 ( .A(n13449), .B(n13448), .Z(c[1268]) );
  NANDN U15278 ( .A(n13416), .B(n13415), .Z(n13420) );
  NANDN U15279 ( .A(n13418), .B(n13417), .Z(n13419) );
  AND U15280 ( .A(n13420), .B(n13419), .Z(n13455) );
  NANDN U15281 ( .A(n13422), .B(n13421), .Z(n13426) );
  NANDN U15282 ( .A(n13424), .B(n13423), .Z(n13425) );
  AND U15283 ( .A(n13426), .B(n13425), .Z(n13453) );
  NAND U15284 ( .A(n42143), .B(n13427), .Z(n13429) );
  XNOR U15285 ( .A(a[247]), .B(n4107), .Z(n13464) );
  NAND U15286 ( .A(n42144), .B(n13464), .Z(n13428) );
  AND U15287 ( .A(n13429), .B(n13428), .Z(n13479) );
  XOR U15288 ( .A(a[251]), .B(n42012), .Z(n13467) );
  XNOR U15289 ( .A(n13479), .B(n13478), .Z(n13481) );
  XOR U15290 ( .A(a[249]), .B(n42085), .Z(n13471) );
  AND U15291 ( .A(a[245]), .B(b[7]), .Z(n13472) );
  XNOR U15292 ( .A(n13473), .B(n13472), .Z(n13474) );
  AND U15293 ( .A(a[253]), .B(b[0]), .Z(n13432) );
  XNOR U15294 ( .A(n13432), .B(n4071), .Z(n13434) );
  NANDN U15295 ( .A(b[0]), .B(a[252]), .Z(n13433) );
  NAND U15296 ( .A(n13434), .B(n13433), .Z(n13475) );
  XNOR U15297 ( .A(n13474), .B(n13475), .Z(n13480) );
  XOR U15298 ( .A(n13481), .B(n13480), .Z(n13459) );
  NANDN U15299 ( .A(n13436), .B(n13435), .Z(n13440) );
  NANDN U15300 ( .A(n13438), .B(n13437), .Z(n13439) );
  AND U15301 ( .A(n13440), .B(n13439), .Z(n13458) );
  XNOR U15302 ( .A(n13459), .B(n13458), .Z(n13460) );
  NANDN U15303 ( .A(n13442), .B(n13441), .Z(n13446) );
  NAND U15304 ( .A(n13444), .B(n13443), .Z(n13445) );
  NAND U15305 ( .A(n13446), .B(n13445), .Z(n13461) );
  XNOR U15306 ( .A(n13460), .B(n13461), .Z(n13452) );
  XNOR U15307 ( .A(n13453), .B(n13452), .Z(n13454) );
  XNOR U15308 ( .A(n13455), .B(n13454), .Z(n13484) );
  XNOR U15309 ( .A(sreg[1269]), .B(n13484), .Z(n13486) );
  NANDN U15310 ( .A(sreg[1268]), .B(n13447), .Z(n13451) );
  NAND U15311 ( .A(n13449), .B(n13448), .Z(n13450) );
  NAND U15312 ( .A(n13451), .B(n13450), .Z(n13485) );
  XNOR U15313 ( .A(n13486), .B(n13485), .Z(c[1269]) );
  NANDN U15314 ( .A(n13453), .B(n13452), .Z(n13457) );
  NANDN U15315 ( .A(n13455), .B(n13454), .Z(n13456) );
  AND U15316 ( .A(n13457), .B(n13456), .Z(n13492) );
  NANDN U15317 ( .A(n13459), .B(n13458), .Z(n13463) );
  NANDN U15318 ( .A(n13461), .B(n13460), .Z(n13462) );
  AND U15319 ( .A(n13463), .B(n13462), .Z(n13490) );
  NAND U15320 ( .A(n42143), .B(n13464), .Z(n13466) );
  XNOR U15321 ( .A(a[248]), .B(n4107), .Z(n13501) );
  NAND U15322 ( .A(n42144), .B(n13501), .Z(n13465) );
  AND U15323 ( .A(n13466), .B(n13465), .Z(n13516) );
  XOR U15324 ( .A(a[252]), .B(n42012), .Z(n13504) );
  XNOR U15325 ( .A(n13516), .B(n13515), .Z(n13518) );
  AND U15326 ( .A(a[254]), .B(b[0]), .Z(n13468) );
  XNOR U15327 ( .A(n13468), .B(n4071), .Z(n13470) );
  NANDN U15328 ( .A(b[0]), .B(a[253]), .Z(n13469) );
  NAND U15329 ( .A(n13470), .B(n13469), .Z(n13512) );
  XOR U15330 ( .A(a[250]), .B(n42085), .Z(n13505) );
  AND U15331 ( .A(a[246]), .B(b[7]), .Z(n13509) );
  XNOR U15332 ( .A(n13510), .B(n13509), .Z(n13511) );
  XNOR U15333 ( .A(n13512), .B(n13511), .Z(n13517) );
  XOR U15334 ( .A(n13518), .B(n13517), .Z(n13496) );
  NANDN U15335 ( .A(n13473), .B(n13472), .Z(n13477) );
  NANDN U15336 ( .A(n13475), .B(n13474), .Z(n13476) );
  AND U15337 ( .A(n13477), .B(n13476), .Z(n13495) );
  XNOR U15338 ( .A(n13496), .B(n13495), .Z(n13497) );
  NANDN U15339 ( .A(n13479), .B(n13478), .Z(n13483) );
  NAND U15340 ( .A(n13481), .B(n13480), .Z(n13482) );
  NAND U15341 ( .A(n13483), .B(n13482), .Z(n13498) );
  XNOR U15342 ( .A(n13497), .B(n13498), .Z(n13489) );
  XNOR U15343 ( .A(n13490), .B(n13489), .Z(n13491) );
  XNOR U15344 ( .A(n13492), .B(n13491), .Z(n13521) );
  XNOR U15345 ( .A(sreg[1270]), .B(n13521), .Z(n13523) );
  NANDN U15346 ( .A(sreg[1269]), .B(n13484), .Z(n13488) );
  NAND U15347 ( .A(n13486), .B(n13485), .Z(n13487) );
  NAND U15348 ( .A(n13488), .B(n13487), .Z(n13522) );
  XNOR U15349 ( .A(n13523), .B(n13522), .Z(c[1270]) );
  NANDN U15350 ( .A(n13490), .B(n13489), .Z(n13494) );
  NANDN U15351 ( .A(n13492), .B(n13491), .Z(n13493) );
  AND U15352 ( .A(n13494), .B(n13493), .Z(n13529) );
  NANDN U15353 ( .A(n13496), .B(n13495), .Z(n13500) );
  NANDN U15354 ( .A(n13498), .B(n13497), .Z(n13499) );
  AND U15355 ( .A(n13500), .B(n13499), .Z(n13527) );
  NAND U15356 ( .A(n42143), .B(n13501), .Z(n13503) );
  XNOR U15357 ( .A(a[249]), .B(n4107), .Z(n13538) );
  NAND U15358 ( .A(n42144), .B(n13538), .Z(n13502) );
  AND U15359 ( .A(n13503), .B(n13502), .Z(n13553) );
  XOR U15360 ( .A(a[253]), .B(n42012), .Z(n13541) );
  XNOR U15361 ( .A(n13553), .B(n13552), .Z(n13555) );
  XOR U15362 ( .A(a[251]), .B(n42085), .Z(n13545) );
  AND U15363 ( .A(a[247]), .B(b[7]), .Z(n13546) );
  XNOR U15364 ( .A(n13547), .B(n13546), .Z(n13548) );
  AND U15365 ( .A(a[255]), .B(b[0]), .Z(n13506) );
  XNOR U15366 ( .A(n13506), .B(n4071), .Z(n13508) );
  NANDN U15367 ( .A(b[0]), .B(a[254]), .Z(n13507) );
  NAND U15368 ( .A(n13508), .B(n13507), .Z(n13549) );
  XNOR U15369 ( .A(n13548), .B(n13549), .Z(n13554) );
  XOR U15370 ( .A(n13555), .B(n13554), .Z(n13533) );
  NANDN U15371 ( .A(n13510), .B(n13509), .Z(n13514) );
  NANDN U15372 ( .A(n13512), .B(n13511), .Z(n13513) );
  AND U15373 ( .A(n13514), .B(n13513), .Z(n13532) );
  XNOR U15374 ( .A(n13533), .B(n13532), .Z(n13534) );
  NANDN U15375 ( .A(n13516), .B(n13515), .Z(n13520) );
  NAND U15376 ( .A(n13518), .B(n13517), .Z(n13519) );
  NAND U15377 ( .A(n13520), .B(n13519), .Z(n13535) );
  XNOR U15378 ( .A(n13534), .B(n13535), .Z(n13526) );
  XNOR U15379 ( .A(n13527), .B(n13526), .Z(n13528) );
  XNOR U15380 ( .A(n13529), .B(n13528), .Z(n13558) );
  XNOR U15381 ( .A(sreg[1271]), .B(n13558), .Z(n13560) );
  NANDN U15382 ( .A(sreg[1270]), .B(n13521), .Z(n13525) );
  NAND U15383 ( .A(n13523), .B(n13522), .Z(n13524) );
  NAND U15384 ( .A(n13525), .B(n13524), .Z(n13559) );
  XNOR U15385 ( .A(n13560), .B(n13559), .Z(c[1271]) );
  NANDN U15386 ( .A(n13527), .B(n13526), .Z(n13531) );
  NANDN U15387 ( .A(n13529), .B(n13528), .Z(n13530) );
  AND U15388 ( .A(n13531), .B(n13530), .Z(n13566) );
  NANDN U15389 ( .A(n13533), .B(n13532), .Z(n13537) );
  NANDN U15390 ( .A(n13535), .B(n13534), .Z(n13536) );
  AND U15391 ( .A(n13537), .B(n13536), .Z(n13564) );
  NAND U15392 ( .A(n42143), .B(n13538), .Z(n13540) );
  XNOR U15393 ( .A(a[250]), .B(n4107), .Z(n13575) );
  NAND U15394 ( .A(n42144), .B(n13575), .Z(n13539) );
  AND U15395 ( .A(n13540), .B(n13539), .Z(n13590) );
  XOR U15396 ( .A(a[254]), .B(n42012), .Z(n13578) );
  XNOR U15397 ( .A(n13590), .B(n13589), .Z(n13592) );
  AND U15398 ( .A(a[256]), .B(b[0]), .Z(n13542) );
  XNOR U15399 ( .A(n13542), .B(n4071), .Z(n13544) );
  NANDN U15400 ( .A(b[0]), .B(a[255]), .Z(n13543) );
  NAND U15401 ( .A(n13544), .B(n13543), .Z(n13586) );
  XOR U15402 ( .A(a[252]), .B(n42085), .Z(n13582) );
  AND U15403 ( .A(a[248]), .B(b[7]), .Z(n13583) );
  XNOR U15404 ( .A(n13584), .B(n13583), .Z(n13585) );
  XNOR U15405 ( .A(n13586), .B(n13585), .Z(n13591) );
  XOR U15406 ( .A(n13592), .B(n13591), .Z(n13570) );
  NANDN U15407 ( .A(n13547), .B(n13546), .Z(n13551) );
  NANDN U15408 ( .A(n13549), .B(n13548), .Z(n13550) );
  AND U15409 ( .A(n13551), .B(n13550), .Z(n13569) );
  XNOR U15410 ( .A(n13570), .B(n13569), .Z(n13571) );
  NANDN U15411 ( .A(n13553), .B(n13552), .Z(n13557) );
  NAND U15412 ( .A(n13555), .B(n13554), .Z(n13556) );
  NAND U15413 ( .A(n13557), .B(n13556), .Z(n13572) );
  XNOR U15414 ( .A(n13571), .B(n13572), .Z(n13563) );
  XNOR U15415 ( .A(n13564), .B(n13563), .Z(n13565) );
  XNOR U15416 ( .A(n13566), .B(n13565), .Z(n13595) );
  XNOR U15417 ( .A(sreg[1272]), .B(n13595), .Z(n13597) );
  NANDN U15418 ( .A(sreg[1271]), .B(n13558), .Z(n13562) );
  NAND U15419 ( .A(n13560), .B(n13559), .Z(n13561) );
  NAND U15420 ( .A(n13562), .B(n13561), .Z(n13596) );
  XNOR U15421 ( .A(n13597), .B(n13596), .Z(c[1272]) );
  NANDN U15422 ( .A(n13564), .B(n13563), .Z(n13568) );
  NANDN U15423 ( .A(n13566), .B(n13565), .Z(n13567) );
  AND U15424 ( .A(n13568), .B(n13567), .Z(n13603) );
  NANDN U15425 ( .A(n13570), .B(n13569), .Z(n13574) );
  NANDN U15426 ( .A(n13572), .B(n13571), .Z(n13573) );
  AND U15427 ( .A(n13574), .B(n13573), .Z(n13601) );
  NAND U15428 ( .A(n42143), .B(n13575), .Z(n13577) );
  XNOR U15429 ( .A(a[251]), .B(n4107), .Z(n13612) );
  NAND U15430 ( .A(n42144), .B(n13612), .Z(n13576) );
  AND U15431 ( .A(n13577), .B(n13576), .Z(n13627) );
  XOR U15432 ( .A(a[255]), .B(n42012), .Z(n13615) );
  XNOR U15433 ( .A(n13627), .B(n13626), .Z(n13629) );
  AND U15434 ( .A(a[257]), .B(b[0]), .Z(n13579) );
  XNOR U15435 ( .A(n13579), .B(n4071), .Z(n13581) );
  NANDN U15436 ( .A(b[0]), .B(a[256]), .Z(n13580) );
  NAND U15437 ( .A(n13581), .B(n13580), .Z(n13623) );
  XOR U15438 ( .A(a[253]), .B(n42085), .Z(n13619) );
  AND U15439 ( .A(a[249]), .B(b[7]), .Z(n13620) );
  XNOR U15440 ( .A(n13621), .B(n13620), .Z(n13622) );
  XNOR U15441 ( .A(n13623), .B(n13622), .Z(n13628) );
  XOR U15442 ( .A(n13629), .B(n13628), .Z(n13607) );
  NANDN U15443 ( .A(n13584), .B(n13583), .Z(n13588) );
  NANDN U15444 ( .A(n13586), .B(n13585), .Z(n13587) );
  AND U15445 ( .A(n13588), .B(n13587), .Z(n13606) );
  XNOR U15446 ( .A(n13607), .B(n13606), .Z(n13608) );
  NANDN U15447 ( .A(n13590), .B(n13589), .Z(n13594) );
  NAND U15448 ( .A(n13592), .B(n13591), .Z(n13593) );
  NAND U15449 ( .A(n13594), .B(n13593), .Z(n13609) );
  XNOR U15450 ( .A(n13608), .B(n13609), .Z(n13600) );
  XNOR U15451 ( .A(n13601), .B(n13600), .Z(n13602) );
  XNOR U15452 ( .A(n13603), .B(n13602), .Z(n13632) );
  XNOR U15453 ( .A(sreg[1273]), .B(n13632), .Z(n13634) );
  NANDN U15454 ( .A(sreg[1272]), .B(n13595), .Z(n13599) );
  NAND U15455 ( .A(n13597), .B(n13596), .Z(n13598) );
  NAND U15456 ( .A(n13599), .B(n13598), .Z(n13633) );
  XNOR U15457 ( .A(n13634), .B(n13633), .Z(c[1273]) );
  NANDN U15458 ( .A(n13601), .B(n13600), .Z(n13605) );
  NANDN U15459 ( .A(n13603), .B(n13602), .Z(n13604) );
  AND U15460 ( .A(n13605), .B(n13604), .Z(n13640) );
  NANDN U15461 ( .A(n13607), .B(n13606), .Z(n13611) );
  NANDN U15462 ( .A(n13609), .B(n13608), .Z(n13610) );
  AND U15463 ( .A(n13611), .B(n13610), .Z(n13638) );
  NAND U15464 ( .A(n42143), .B(n13612), .Z(n13614) );
  XNOR U15465 ( .A(a[252]), .B(n4107), .Z(n13649) );
  NAND U15466 ( .A(n42144), .B(n13649), .Z(n13613) );
  AND U15467 ( .A(n13614), .B(n13613), .Z(n13664) );
  XOR U15468 ( .A(a[256]), .B(n42012), .Z(n13652) );
  XNOR U15469 ( .A(n13664), .B(n13663), .Z(n13666) );
  AND U15470 ( .A(a[258]), .B(b[0]), .Z(n13616) );
  XNOR U15471 ( .A(n13616), .B(n4071), .Z(n13618) );
  NANDN U15472 ( .A(b[0]), .B(a[257]), .Z(n13617) );
  NAND U15473 ( .A(n13618), .B(n13617), .Z(n13660) );
  XOR U15474 ( .A(a[254]), .B(n42085), .Z(n13656) );
  AND U15475 ( .A(a[250]), .B(b[7]), .Z(n13657) );
  XNOR U15476 ( .A(n13658), .B(n13657), .Z(n13659) );
  XNOR U15477 ( .A(n13660), .B(n13659), .Z(n13665) );
  XOR U15478 ( .A(n13666), .B(n13665), .Z(n13644) );
  NANDN U15479 ( .A(n13621), .B(n13620), .Z(n13625) );
  NANDN U15480 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U15481 ( .A(n13625), .B(n13624), .Z(n13643) );
  XNOR U15482 ( .A(n13644), .B(n13643), .Z(n13645) );
  NANDN U15483 ( .A(n13627), .B(n13626), .Z(n13631) );
  NAND U15484 ( .A(n13629), .B(n13628), .Z(n13630) );
  NAND U15485 ( .A(n13631), .B(n13630), .Z(n13646) );
  XNOR U15486 ( .A(n13645), .B(n13646), .Z(n13637) );
  XNOR U15487 ( .A(n13638), .B(n13637), .Z(n13639) );
  XNOR U15488 ( .A(n13640), .B(n13639), .Z(n13669) );
  XNOR U15489 ( .A(sreg[1274]), .B(n13669), .Z(n13671) );
  NANDN U15490 ( .A(sreg[1273]), .B(n13632), .Z(n13636) );
  NAND U15491 ( .A(n13634), .B(n13633), .Z(n13635) );
  NAND U15492 ( .A(n13636), .B(n13635), .Z(n13670) );
  XNOR U15493 ( .A(n13671), .B(n13670), .Z(c[1274]) );
  NANDN U15494 ( .A(n13638), .B(n13637), .Z(n13642) );
  NANDN U15495 ( .A(n13640), .B(n13639), .Z(n13641) );
  AND U15496 ( .A(n13642), .B(n13641), .Z(n13677) );
  NANDN U15497 ( .A(n13644), .B(n13643), .Z(n13648) );
  NANDN U15498 ( .A(n13646), .B(n13645), .Z(n13647) );
  AND U15499 ( .A(n13648), .B(n13647), .Z(n13675) );
  NAND U15500 ( .A(n42143), .B(n13649), .Z(n13651) );
  XNOR U15501 ( .A(a[253]), .B(n4108), .Z(n13686) );
  NAND U15502 ( .A(n42144), .B(n13686), .Z(n13650) );
  AND U15503 ( .A(n13651), .B(n13650), .Z(n13701) );
  XOR U15504 ( .A(a[257]), .B(n42012), .Z(n13689) );
  XNOR U15505 ( .A(n13701), .B(n13700), .Z(n13703) );
  AND U15506 ( .A(a[259]), .B(b[0]), .Z(n13653) );
  XNOR U15507 ( .A(n13653), .B(n4071), .Z(n13655) );
  NANDN U15508 ( .A(b[0]), .B(a[258]), .Z(n13654) );
  NAND U15509 ( .A(n13655), .B(n13654), .Z(n13697) );
  XOR U15510 ( .A(a[255]), .B(n42085), .Z(n13693) );
  AND U15511 ( .A(a[251]), .B(b[7]), .Z(n13694) );
  XNOR U15512 ( .A(n13695), .B(n13694), .Z(n13696) );
  XNOR U15513 ( .A(n13697), .B(n13696), .Z(n13702) );
  XOR U15514 ( .A(n13703), .B(n13702), .Z(n13681) );
  NANDN U15515 ( .A(n13658), .B(n13657), .Z(n13662) );
  NANDN U15516 ( .A(n13660), .B(n13659), .Z(n13661) );
  AND U15517 ( .A(n13662), .B(n13661), .Z(n13680) );
  XNOR U15518 ( .A(n13681), .B(n13680), .Z(n13682) );
  NANDN U15519 ( .A(n13664), .B(n13663), .Z(n13668) );
  NAND U15520 ( .A(n13666), .B(n13665), .Z(n13667) );
  NAND U15521 ( .A(n13668), .B(n13667), .Z(n13683) );
  XNOR U15522 ( .A(n13682), .B(n13683), .Z(n13674) );
  XNOR U15523 ( .A(n13675), .B(n13674), .Z(n13676) );
  XNOR U15524 ( .A(n13677), .B(n13676), .Z(n13706) );
  XNOR U15525 ( .A(sreg[1275]), .B(n13706), .Z(n13708) );
  NANDN U15526 ( .A(sreg[1274]), .B(n13669), .Z(n13673) );
  NAND U15527 ( .A(n13671), .B(n13670), .Z(n13672) );
  NAND U15528 ( .A(n13673), .B(n13672), .Z(n13707) );
  XNOR U15529 ( .A(n13708), .B(n13707), .Z(c[1275]) );
  NANDN U15530 ( .A(n13675), .B(n13674), .Z(n13679) );
  NANDN U15531 ( .A(n13677), .B(n13676), .Z(n13678) );
  AND U15532 ( .A(n13679), .B(n13678), .Z(n13714) );
  NANDN U15533 ( .A(n13681), .B(n13680), .Z(n13685) );
  NANDN U15534 ( .A(n13683), .B(n13682), .Z(n13684) );
  AND U15535 ( .A(n13685), .B(n13684), .Z(n13712) );
  NAND U15536 ( .A(n42143), .B(n13686), .Z(n13688) );
  XNOR U15537 ( .A(a[254]), .B(n4108), .Z(n13723) );
  NAND U15538 ( .A(n42144), .B(n13723), .Z(n13687) );
  AND U15539 ( .A(n13688), .B(n13687), .Z(n13738) );
  XOR U15540 ( .A(a[258]), .B(n42012), .Z(n13726) );
  XNOR U15541 ( .A(n13738), .B(n13737), .Z(n13740) );
  AND U15542 ( .A(a[260]), .B(b[0]), .Z(n13690) );
  XNOR U15543 ( .A(n13690), .B(n4071), .Z(n13692) );
  NANDN U15544 ( .A(b[0]), .B(a[259]), .Z(n13691) );
  NAND U15545 ( .A(n13692), .B(n13691), .Z(n13734) );
  XOR U15546 ( .A(a[256]), .B(n42085), .Z(n13727) );
  AND U15547 ( .A(a[252]), .B(b[7]), .Z(n13731) );
  XNOR U15548 ( .A(n13732), .B(n13731), .Z(n13733) );
  XNOR U15549 ( .A(n13734), .B(n13733), .Z(n13739) );
  XOR U15550 ( .A(n13740), .B(n13739), .Z(n13718) );
  NANDN U15551 ( .A(n13695), .B(n13694), .Z(n13699) );
  NANDN U15552 ( .A(n13697), .B(n13696), .Z(n13698) );
  AND U15553 ( .A(n13699), .B(n13698), .Z(n13717) );
  XNOR U15554 ( .A(n13718), .B(n13717), .Z(n13719) );
  NANDN U15555 ( .A(n13701), .B(n13700), .Z(n13705) );
  NAND U15556 ( .A(n13703), .B(n13702), .Z(n13704) );
  NAND U15557 ( .A(n13705), .B(n13704), .Z(n13720) );
  XNOR U15558 ( .A(n13719), .B(n13720), .Z(n13711) );
  XNOR U15559 ( .A(n13712), .B(n13711), .Z(n13713) );
  XNOR U15560 ( .A(n13714), .B(n13713), .Z(n13743) );
  XNOR U15561 ( .A(sreg[1276]), .B(n13743), .Z(n13745) );
  NANDN U15562 ( .A(sreg[1275]), .B(n13706), .Z(n13710) );
  NAND U15563 ( .A(n13708), .B(n13707), .Z(n13709) );
  NAND U15564 ( .A(n13710), .B(n13709), .Z(n13744) );
  XNOR U15565 ( .A(n13745), .B(n13744), .Z(c[1276]) );
  NANDN U15566 ( .A(n13712), .B(n13711), .Z(n13716) );
  NANDN U15567 ( .A(n13714), .B(n13713), .Z(n13715) );
  AND U15568 ( .A(n13716), .B(n13715), .Z(n13751) );
  NANDN U15569 ( .A(n13718), .B(n13717), .Z(n13722) );
  NANDN U15570 ( .A(n13720), .B(n13719), .Z(n13721) );
  AND U15571 ( .A(n13722), .B(n13721), .Z(n13749) );
  NAND U15572 ( .A(n42143), .B(n13723), .Z(n13725) );
  XNOR U15573 ( .A(a[255]), .B(n4108), .Z(n13760) );
  NAND U15574 ( .A(n42144), .B(n13760), .Z(n13724) );
  AND U15575 ( .A(n13725), .B(n13724), .Z(n13775) );
  XOR U15576 ( .A(a[259]), .B(n42012), .Z(n13763) );
  XNOR U15577 ( .A(n13775), .B(n13774), .Z(n13777) );
  XOR U15578 ( .A(a[257]), .B(n42085), .Z(n13767) );
  AND U15579 ( .A(a[253]), .B(b[7]), .Z(n13768) );
  XNOR U15580 ( .A(n13769), .B(n13768), .Z(n13770) );
  AND U15581 ( .A(a[261]), .B(b[0]), .Z(n13728) );
  XNOR U15582 ( .A(n13728), .B(n4071), .Z(n13730) );
  NANDN U15583 ( .A(b[0]), .B(a[260]), .Z(n13729) );
  NAND U15584 ( .A(n13730), .B(n13729), .Z(n13771) );
  XNOR U15585 ( .A(n13770), .B(n13771), .Z(n13776) );
  XOR U15586 ( .A(n13777), .B(n13776), .Z(n13755) );
  NANDN U15587 ( .A(n13732), .B(n13731), .Z(n13736) );
  NANDN U15588 ( .A(n13734), .B(n13733), .Z(n13735) );
  AND U15589 ( .A(n13736), .B(n13735), .Z(n13754) );
  XNOR U15590 ( .A(n13755), .B(n13754), .Z(n13756) );
  NANDN U15591 ( .A(n13738), .B(n13737), .Z(n13742) );
  NAND U15592 ( .A(n13740), .B(n13739), .Z(n13741) );
  NAND U15593 ( .A(n13742), .B(n13741), .Z(n13757) );
  XNOR U15594 ( .A(n13756), .B(n13757), .Z(n13748) );
  XNOR U15595 ( .A(n13749), .B(n13748), .Z(n13750) );
  XNOR U15596 ( .A(n13751), .B(n13750), .Z(n13780) );
  XNOR U15597 ( .A(sreg[1277]), .B(n13780), .Z(n13782) );
  NANDN U15598 ( .A(sreg[1276]), .B(n13743), .Z(n13747) );
  NAND U15599 ( .A(n13745), .B(n13744), .Z(n13746) );
  NAND U15600 ( .A(n13747), .B(n13746), .Z(n13781) );
  XNOR U15601 ( .A(n13782), .B(n13781), .Z(c[1277]) );
  NANDN U15602 ( .A(n13749), .B(n13748), .Z(n13753) );
  NANDN U15603 ( .A(n13751), .B(n13750), .Z(n13752) );
  AND U15604 ( .A(n13753), .B(n13752), .Z(n13788) );
  NANDN U15605 ( .A(n13755), .B(n13754), .Z(n13759) );
  NANDN U15606 ( .A(n13757), .B(n13756), .Z(n13758) );
  AND U15607 ( .A(n13759), .B(n13758), .Z(n13786) );
  NAND U15608 ( .A(n42143), .B(n13760), .Z(n13762) );
  XNOR U15609 ( .A(a[256]), .B(n4108), .Z(n13797) );
  NAND U15610 ( .A(n42144), .B(n13797), .Z(n13761) );
  AND U15611 ( .A(n13762), .B(n13761), .Z(n13812) );
  XOR U15612 ( .A(a[260]), .B(n42012), .Z(n13800) );
  XNOR U15613 ( .A(n13812), .B(n13811), .Z(n13814) );
  AND U15614 ( .A(a[262]), .B(b[0]), .Z(n13764) );
  XNOR U15615 ( .A(n13764), .B(n4071), .Z(n13766) );
  NANDN U15616 ( .A(b[0]), .B(a[261]), .Z(n13765) );
  NAND U15617 ( .A(n13766), .B(n13765), .Z(n13808) );
  XOR U15618 ( .A(a[258]), .B(n42085), .Z(n13804) );
  AND U15619 ( .A(a[254]), .B(b[7]), .Z(n13805) );
  XNOR U15620 ( .A(n13806), .B(n13805), .Z(n13807) );
  XNOR U15621 ( .A(n13808), .B(n13807), .Z(n13813) );
  XOR U15622 ( .A(n13814), .B(n13813), .Z(n13792) );
  NANDN U15623 ( .A(n13769), .B(n13768), .Z(n13773) );
  NANDN U15624 ( .A(n13771), .B(n13770), .Z(n13772) );
  AND U15625 ( .A(n13773), .B(n13772), .Z(n13791) );
  XNOR U15626 ( .A(n13792), .B(n13791), .Z(n13793) );
  NANDN U15627 ( .A(n13775), .B(n13774), .Z(n13779) );
  NAND U15628 ( .A(n13777), .B(n13776), .Z(n13778) );
  NAND U15629 ( .A(n13779), .B(n13778), .Z(n13794) );
  XNOR U15630 ( .A(n13793), .B(n13794), .Z(n13785) );
  XNOR U15631 ( .A(n13786), .B(n13785), .Z(n13787) );
  XNOR U15632 ( .A(n13788), .B(n13787), .Z(n13817) );
  XNOR U15633 ( .A(sreg[1278]), .B(n13817), .Z(n13819) );
  NANDN U15634 ( .A(sreg[1277]), .B(n13780), .Z(n13784) );
  NAND U15635 ( .A(n13782), .B(n13781), .Z(n13783) );
  NAND U15636 ( .A(n13784), .B(n13783), .Z(n13818) );
  XNOR U15637 ( .A(n13819), .B(n13818), .Z(c[1278]) );
  NANDN U15638 ( .A(n13786), .B(n13785), .Z(n13790) );
  NANDN U15639 ( .A(n13788), .B(n13787), .Z(n13789) );
  AND U15640 ( .A(n13790), .B(n13789), .Z(n13825) );
  NANDN U15641 ( .A(n13792), .B(n13791), .Z(n13796) );
  NANDN U15642 ( .A(n13794), .B(n13793), .Z(n13795) );
  AND U15643 ( .A(n13796), .B(n13795), .Z(n13823) );
  NAND U15644 ( .A(n42143), .B(n13797), .Z(n13799) );
  XNOR U15645 ( .A(a[257]), .B(n4108), .Z(n13834) );
  NAND U15646 ( .A(n42144), .B(n13834), .Z(n13798) );
  AND U15647 ( .A(n13799), .B(n13798), .Z(n13849) );
  XOR U15648 ( .A(a[261]), .B(n42012), .Z(n13837) );
  XNOR U15649 ( .A(n13849), .B(n13848), .Z(n13851) );
  AND U15650 ( .A(a[263]), .B(b[0]), .Z(n13801) );
  XNOR U15651 ( .A(n13801), .B(n4071), .Z(n13803) );
  NANDN U15652 ( .A(b[0]), .B(a[262]), .Z(n13802) );
  NAND U15653 ( .A(n13803), .B(n13802), .Z(n13845) );
  XOR U15654 ( .A(a[259]), .B(n42085), .Z(n13841) );
  AND U15655 ( .A(a[255]), .B(b[7]), .Z(n13842) );
  XNOR U15656 ( .A(n13843), .B(n13842), .Z(n13844) );
  XNOR U15657 ( .A(n13845), .B(n13844), .Z(n13850) );
  XOR U15658 ( .A(n13851), .B(n13850), .Z(n13829) );
  NANDN U15659 ( .A(n13806), .B(n13805), .Z(n13810) );
  NANDN U15660 ( .A(n13808), .B(n13807), .Z(n13809) );
  AND U15661 ( .A(n13810), .B(n13809), .Z(n13828) );
  XNOR U15662 ( .A(n13829), .B(n13828), .Z(n13830) );
  NANDN U15663 ( .A(n13812), .B(n13811), .Z(n13816) );
  NAND U15664 ( .A(n13814), .B(n13813), .Z(n13815) );
  NAND U15665 ( .A(n13816), .B(n13815), .Z(n13831) );
  XNOR U15666 ( .A(n13830), .B(n13831), .Z(n13822) );
  XNOR U15667 ( .A(n13823), .B(n13822), .Z(n13824) );
  XNOR U15668 ( .A(n13825), .B(n13824), .Z(n13854) );
  XNOR U15669 ( .A(sreg[1279]), .B(n13854), .Z(n13856) );
  NANDN U15670 ( .A(sreg[1278]), .B(n13817), .Z(n13821) );
  NAND U15671 ( .A(n13819), .B(n13818), .Z(n13820) );
  NAND U15672 ( .A(n13821), .B(n13820), .Z(n13855) );
  XNOR U15673 ( .A(n13856), .B(n13855), .Z(c[1279]) );
  NANDN U15674 ( .A(n13823), .B(n13822), .Z(n13827) );
  NANDN U15675 ( .A(n13825), .B(n13824), .Z(n13826) );
  AND U15676 ( .A(n13827), .B(n13826), .Z(n13862) );
  NANDN U15677 ( .A(n13829), .B(n13828), .Z(n13833) );
  NANDN U15678 ( .A(n13831), .B(n13830), .Z(n13832) );
  AND U15679 ( .A(n13833), .B(n13832), .Z(n13860) );
  NAND U15680 ( .A(n42143), .B(n13834), .Z(n13836) );
  XNOR U15681 ( .A(a[258]), .B(n4108), .Z(n13871) );
  NAND U15682 ( .A(n42144), .B(n13871), .Z(n13835) );
  AND U15683 ( .A(n13836), .B(n13835), .Z(n13886) );
  XOR U15684 ( .A(a[262]), .B(n42012), .Z(n13874) );
  XNOR U15685 ( .A(n13886), .B(n13885), .Z(n13888) );
  AND U15686 ( .A(a[264]), .B(b[0]), .Z(n13838) );
  XNOR U15687 ( .A(n13838), .B(n4071), .Z(n13840) );
  NANDN U15688 ( .A(b[0]), .B(a[263]), .Z(n13839) );
  NAND U15689 ( .A(n13840), .B(n13839), .Z(n13882) );
  XOR U15690 ( .A(a[260]), .B(n42085), .Z(n13878) );
  AND U15691 ( .A(a[256]), .B(b[7]), .Z(n13879) );
  XNOR U15692 ( .A(n13880), .B(n13879), .Z(n13881) );
  XNOR U15693 ( .A(n13882), .B(n13881), .Z(n13887) );
  XOR U15694 ( .A(n13888), .B(n13887), .Z(n13866) );
  NANDN U15695 ( .A(n13843), .B(n13842), .Z(n13847) );
  NANDN U15696 ( .A(n13845), .B(n13844), .Z(n13846) );
  AND U15697 ( .A(n13847), .B(n13846), .Z(n13865) );
  XNOR U15698 ( .A(n13866), .B(n13865), .Z(n13867) );
  NANDN U15699 ( .A(n13849), .B(n13848), .Z(n13853) );
  NAND U15700 ( .A(n13851), .B(n13850), .Z(n13852) );
  NAND U15701 ( .A(n13853), .B(n13852), .Z(n13868) );
  XNOR U15702 ( .A(n13867), .B(n13868), .Z(n13859) );
  XNOR U15703 ( .A(n13860), .B(n13859), .Z(n13861) );
  XNOR U15704 ( .A(n13862), .B(n13861), .Z(n13891) );
  XNOR U15705 ( .A(sreg[1280]), .B(n13891), .Z(n13893) );
  NANDN U15706 ( .A(sreg[1279]), .B(n13854), .Z(n13858) );
  NAND U15707 ( .A(n13856), .B(n13855), .Z(n13857) );
  NAND U15708 ( .A(n13858), .B(n13857), .Z(n13892) );
  XNOR U15709 ( .A(n13893), .B(n13892), .Z(c[1280]) );
  NANDN U15710 ( .A(n13860), .B(n13859), .Z(n13864) );
  NANDN U15711 ( .A(n13862), .B(n13861), .Z(n13863) );
  AND U15712 ( .A(n13864), .B(n13863), .Z(n13899) );
  NANDN U15713 ( .A(n13866), .B(n13865), .Z(n13870) );
  NANDN U15714 ( .A(n13868), .B(n13867), .Z(n13869) );
  AND U15715 ( .A(n13870), .B(n13869), .Z(n13897) );
  NAND U15716 ( .A(n42143), .B(n13871), .Z(n13873) );
  XNOR U15717 ( .A(a[259]), .B(n4108), .Z(n13908) );
  NAND U15718 ( .A(n42144), .B(n13908), .Z(n13872) );
  AND U15719 ( .A(n13873), .B(n13872), .Z(n13923) );
  XOR U15720 ( .A(a[263]), .B(n42012), .Z(n13911) );
  XNOR U15721 ( .A(n13923), .B(n13922), .Z(n13925) );
  AND U15722 ( .A(a[265]), .B(b[0]), .Z(n13875) );
  XNOR U15723 ( .A(n13875), .B(n4071), .Z(n13877) );
  NANDN U15724 ( .A(b[0]), .B(a[264]), .Z(n13876) );
  NAND U15725 ( .A(n13877), .B(n13876), .Z(n13919) );
  XOR U15726 ( .A(a[261]), .B(n42085), .Z(n13915) );
  AND U15727 ( .A(a[257]), .B(b[7]), .Z(n13916) );
  XNOR U15728 ( .A(n13917), .B(n13916), .Z(n13918) );
  XNOR U15729 ( .A(n13919), .B(n13918), .Z(n13924) );
  XOR U15730 ( .A(n13925), .B(n13924), .Z(n13903) );
  NANDN U15731 ( .A(n13880), .B(n13879), .Z(n13884) );
  NANDN U15732 ( .A(n13882), .B(n13881), .Z(n13883) );
  AND U15733 ( .A(n13884), .B(n13883), .Z(n13902) );
  XNOR U15734 ( .A(n13903), .B(n13902), .Z(n13904) );
  NANDN U15735 ( .A(n13886), .B(n13885), .Z(n13890) );
  NAND U15736 ( .A(n13888), .B(n13887), .Z(n13889) );
  NAND U15737 ( .A(n13890), .B(n13889), .Z(n13905) );
  XNOR U15738 ( .A(n13904), .B(n13905), .Z(n13896) );
  XNOR U15739 ( .A(n13897), .B(n13896), .Z(n13898) );
  XNOR U15740 ( .A(n13899), .B(n13898), .Z(n13928) );
  XNOR U15741 ( .A(sreg[1281]), .B(n13928), .Z(n13930) );
  NANDN U15742 ( .A(sreg[1280]), .B(n13891), .Z(n13895) );
  NAND U15743 ( .A(n13893), .B(n13892), .Z(n13894) );
  NAND U15744 ( .A(n13895), .B(n13894), .Z(n13929) );
  XNOR U15745 ( .A(n13930), .B(n13929), .Z(c[1281]) );
  NANDN U15746 ( .A(n13897), .B(n13896), .Z(n13901) );
  NANDN U15747 ( .A(n13899), .B(n13898), .Z(n13900) );
  AND U15748 ( .A(n13901), .B(n13900), .Z(n13936) );
  NANDN U15749 ( .A(n13903), .B(n13902), .Z(n13907) );
  NANDN U15750 ( .A(n13905), .B(n13904), .Z(n13906) );
  AND U15751 ( .A(n13907), .B(n13906), .Z(n13934) );
  NAND U15752 ( .A(n42143), .B(n13908), .Z(n13910) );
  XNOR U15753 ( .A(a[260]), .B(n4109), .Z(n13945) );
  NAND U15754 ( .A(n42144), .B(n13945), .Z(n13909) );
  AND U15755 ( .A(n13910), .B(n13909), .Z(n13960) );
  XOR U15756 ( .A(a[264]), .B(n42012), .Z(n13948) );
  XNOR U15757 ( .A(n13960), .B(n13959), .Z(n13962) );
  AND U15758 ( .A(a[266]), .B(b[0]), .Z(n13912) );
  XNOR U15759 ( .A(n13912), .B(n4071), .Z(n13914) );
  NANDN U15760 ( .A(b[0]), .B(a[265]), .Z(n13913) );
  NAND U15761 ( .A(n13914), .B(n13913), .Z(n13956) );
  XOR U15762 ( .A(a[262]), .B(n42085), .Z(n13952) );
  AND U15763 ( .A(a[258]), .B(b[7]), .Z(n13953) );
  XNOR U15764 ( .A(n13954), .B(n13953), .Z(n13955) );
  XNOR U15765 ( .A(n13956), .B(n13955), .Z(n13961) );
  XOR U15766 ( .A(n13962), .B(n13961), .Z(n13940) );
  NANDN U15767 ( .A(n13917), .B(n13916), .Z(n13921) );
  NANDN U15768 ( .A(n13919), .B(n13918), .Z(n13920) );
  AND U15769 ( .A(n13921), .B(n13920), .Z(n13939) );
  XNOR U15770 ( .A(n13940), .B(n13939), .Z(n13941) );
  NANDN U15771 ( .A(n13923), .B(n13922), .Z(n13927) );
  NAND U15772 ( .A(n13925), .B(n13924), .Z(n13926) );
  NAND U15773 ( .A(n13927), .B(n13926), .Z(n13942) );
  XNOR U15774 ( .A(n13941), .B(n13942), .Z(n13933) );
  XNOR U15775 ( .A(n13934), .B(n13933), .Z(n13935) );
  XNOR U15776 ( .A(n13936), .B(n13935), .Z(n13965) );
  XNOR U15777 ( .A(sreg[1282]), .B(n13965), .Z(n13967) );
  NANDN U15778 ( .A(sreg[1281]), .B(n13928), .Z(n13932) );
  NAND U15779 ( .A(n13930), .B(n13929), .Z(n13931) );
  NAND U15780 ( .A(n13932), .B(n13931), .Z(n13966) );
  XNOR U15781 ( .A(n13967), .B(n13966), .Z(c[1282]) );
  NANDN U15782 ( .A(n13934), .B(n13933), .Z(n13938) );
  NANDN U15783 ( .A(n13936), .B(n13935), .Z(n13937) );
  AND U15784 ( .A(n13938), .B(n13937), .Z(n13973) );
  NANDN U15785 ( .A(n13940), .B(n13939), .Z(n13944) );
  NANDN U15786 ( .A(n13942), .B(n13941), .Z(n13943) );
  AND U15787 ( .A(n13944), .B(n13943), .Z(n13971) );
  NAND U15788 ( .A(n42143), .B(n13945), .Z(n13947) );
  XNOR U15789 ( .A(a[261]), .B(n4109), .Z(n13982) );
  NAND U15790 ( .A(n42144), .B(n13982), .Z(n13946) );
  AND U15791 ( .A(n13947), .B(n13946), .Z(n13997) );
  XOR U15792 ( .A(a[265]), .B(n42012), .Z(n13985) );
  XNOR U15793 ( .A(n13997), .B(n13996), .Z(n13999) );
  AND U15794 ( .A(a[267]), .B(b[0]), .Z(n13949) );
  XNOR U15795 ( .A(n13949), .B(n4071), .Z(n13951) );
  NANDN U15796 ( .A(b[0]), .B(a[266]), .Z(n13950) );
  NAND U15797 ( .A(n13951), .B(n13950), .Z(n13993) );
  XOR U15798 ( .A(a[263]), .B(n42085), .Z(n13986) );
  AND U15799 ( .A(a[259]), .B(b[7]), .Z(n13990) );
  XNOR U15800 ( .A(n13991), .B(n13990), .Z(n13992) );
  XNOR U15801 ( .A(n13993), .B(n13992), .Z(n13998) );
  XOR U15802 ( .A(n13999), .B(n13998), .Z(n13977) );
  NANDN U15803 ( .A(n13954), .B(n13953), .Z(n13958) );
  NANDN U15804 ( .A(n13956), .B(n13955), .Z(n13957) );
  AND U15805 ( .A(n13958), .B(n13957), .Z(n13976) );
  XNOR U15806 ( .A(n13977), .B(n13976), .Z(n13978) );
  NANDN U15807 ( .A(n13960), .B(n13959), .Z(n13964) );
  NAND U15808 ( .A(n13962), .B(n13961), .Z(n13963) );
  NAND U15809 ( .A(n13964), .B(n13963), .Z(n13979) );
  XNOR U15810 ( .A(n13978), .B(n13979), .Z(n13970) );
  XNOR U15811 ( .A(n13971), .B(n13970), .Z(n13972) );
  XNOR U15812 ( .A(n13973), .B(n13972), .Z(n14002) );
  XNOR U15813 ( .A(sreg[1283]), .B(n14002), .Z(n14004) );
  NANDN U15814 ( .A(sreg[1282]), .B(n13965), .Z(n13969) );
  NAND U15815 ( .A(n13967), .B(n13966), .Z(n13968) );
  NAND U15816 ( .A(n13969), .B(n13968), .Z(n14003) );
  XNOR U15817 ( .A(n14004), .B(n14003), .Z(c[1283]) );
  NANDN U15818 ( .A(n13971), .B(n13970), .Z(n13975) );
  NANDN U15819 ( .A(n13973), .B(n13972), .Z(n13974) );
  AND U15820 ( .A(n13975), .B(n13974), .Z(n14010) );
  NANDN U15821 ( .A(n13977), .B(n13976), .Z(n13981) );
  NANDN U15822 ( .A(n13979), .B(n13978), .Z(n13980) );
  AND U15823 ( .A(n13981), .B(n13980), .Z(n14008) );
  NAND U15824 ( .A(n42143), .B(n13982), .Z(n13984) );
  XNOR U15825 ( .A(a[262]), .B(n4109), .Z(n14019) );
  NAND U15826 ( .A(n42144), .B(n14019), .Z(n13983) );
  AND U15827 ( .A(n13984), .B(n13983), .Z(n14034) );
  XOR U15828 ( .A(a[266]), .B(n42012), .Z(n14022) );
  XNOR U15829 ( .A(n14034), .B(n14033), .Z(n14036) );
  XOR U15830 ( .A(a[264]), .B(n42085), .Z(n14026) );
  AND U15831 ( .A(a[260]), .B(b[7]), .Z(n14027) );
  XNOR U15832 ( .A(n14028), .B(n14027), .Z(n14029) );
  AND U15833 ( .A(a[268]), .B(b[0]), .Z(n13987) );
  XNOR U15834 ( .A(n13987), .B(n4071), .Z(n13989) );
  NANDN U15835 ( .A(b[0]), .B(a[267]), .Z(n13988) );
  NAND U15836 ( .A(n13989), .B(n13988), .Z(n14030) );
  XNOR U15837 ( .A(n14029), .B(n14030), .Z(n14035) );
  XOR U15838 ( .A(n14036), .B(n14035), .Z(n14014) );
  NANDN U15839 ( .A(n13991), .B(n13990), .Z(n13995) );
  NANDN U15840 ( .A(n13993), .B(n13992), .Z(n13994) );
  AND U15841 ( .A(n13995), .B(n13994), .Z(n14013) );
  XNOR U15842 ( .A(n14014), .B(n14013), .Z(n14015) );
  NANDN U15843 ( .A(n13997), .B(n13996), .Z(n14001) );
  NAND U15844 ( .A(n13999), .B(n13998), .Z(n14000) );
  NAND U15845 ( .A(n14001), .B(n14000), .Z(n14016) );
  XNOR U15846 ( .A(n14015), .B(n14016), .Z(n14007) );
  XNOR U15847 ( .A(n14008), .B(n14007), .Z(n14009) );
  XNOR U15848 ( .A(n14010), .B(n14009), .Z(n14039) );
  XNOR U15849 ( .A(sreg[1284]), .B(n14039), .Z(n14041) );
  NANDN U15850 ( .A(sreg[1283]), .B(n14002), .Z(n14006) );
  NAND U15851 ( .A(n14004), .B(n14003), .Z(n14005) );
  NAND U15852 ( .A(n14006), .B(n14005), .Z(n14040) );
  XNOR U15853 ( .A(n14041), .B(n14040), .Z(c[1284]) );
  NANDN U15854 ( .A(n14008), .B(n14007), .Z(n14012) );
  NANDN U15855 ( .A(n14010), .B(n14009), .Z(n14011) );
  AND U15856 ( .A(n14012), .B(n14011), .Z(n14047) );
  NANDN U15857 ( .A(n14014), .B(n14013), .Z(n14018) );
  NANDN U15858 ( .A(n14016), .B(n14015), .Z(n14017) );
  AND U15859 ( .A(n14018), .B(n14017), .Z(n14045) );
  NAND U15860 ( .A(n42143), .B(n14019), .Z(n14021) );
  XNOR U15861 ( .A(a[263]), .B(n4109), .Z(n14056) );
  NAND U15862 ( .A(n42144), .B(n14056), .Z(n14020) );
  AND U15863 ( .A(n14021), .B(n14020), .Z(n14071) );
  XOR U15864 ( .A(a[267]), .B(n42012), .Z(n14059) );
  XNOR U15865 ( .A(n14071), .B(n14070), .Z(n14073) );
  AND U15866 ( .A(a[269]), .B(b[0]), .Z(n14023) );
  XNOR U15867 ( .A(n14023), .B(n4071), .Z(n14025) );
  NANDN U15868 ( .A(b[0]), .B(a[268]), .Z(n14024) );
  NAND U15869 ( .A(n14025), .B(n14024), .Z(n14067) );
  XOR U15870 ( .A(a[265]), .B(n42085), .Z(n14063) );
  AND U15871 ( .A(a[261]), .B(b[7]), .Z(n14064) );
  XNOR U15872 ( .A(n14065), .B(n14064), .Z(n14066) );
  XNOR U15873 ( .A(n14067), .B(n14066), .Z(n14072) );
  XOR U15874 ( .A(n14073), .B(n14072), .Z(n14051) );
  NANDN U15875 ( .A(n14028), .B(n14027), .Z(n14032) );
  NANDN U15876 ( .A(n14030), .B(n14029), .Z(n14031) );
  AND U15877 ( .A(n14032), .B(n14031), .Z(n14050) );
  XNOR U15878 ( .A(n14051), .B(n14050), .Z(n14052) );
  NANDN U15879 ( .A(n14034), .B(n14033), .Z(n14038) );
  NAND U15880 ( .A(n14036), .B(n14035), .Z(n14037) );
  NAND U15881 ( .A(n14038), .B(n14037), .Z(n14053) );
  XNOR U15882 ( .A(n14052), .B(n14053), .Z(n14044) );
  XNOR U15883 ( .A(n14045), .B(n14044), .Z(n14046) );
  XNOR U15884 ( .A(n14047), .B(n14046), .Z(n14076) );
  XNOR U15885 ( .A(sreg[1285]), .B(n14076), .Z(n14078) );
  NANDN U15886 ( .A(sreg[1284]), .B(n14039), .Z(n14043) );
  NAND U15887 ( .A(n14041), .B(n14040), .Z(n14042) );
  NAND U15888 ( .A(n14043), .B(n14042), .Z(n14077) );
  XNOR U15889 ( .A(n14078), .B(n14077), .Z(c[1285]) );
  NANDN U15890 ( .A(n14045), .B(n14044), .Z(n14049) );
  NANDN U15891 ( .A(n14047), .B(n14046), .Z(n14048) );
  AND U15892 ( .A(n14049), .B(n14048), .Z(n14089) );
  NANDN U15893 ( .A(n14051), .B(n14050), .Z(n14055) );
  NANDN U15894 ( .A(n14053), .B(n14052), .Z(n14054) );
  AND U15895 ( .A(n14055), .B(n14054), .Z(n14087) );
  NAND U15896 ( .A(n42143), .B(n14056), .Z(n14058) );
  XNOR U15897 ( .A(a[264]), .B(n4109), .Z(n14098) );
  NAND U15898 ( .A(n42144), .B(n14098), .Z(n14057) );
  AND U15899 ( .A(n14058), .B(n14057), .Z(n14113) );
  XOR U15900 ( .A(a[268]), .B(n42012), .Z(n14101) );
  XNOR U15901 ( .A(n14113), .B(n14112), .Z(n14115) );
  AND U15902 ( .A(a[270]), .B(b[0]), .Z(n14060) );
  XNOR U15903 ( .A(n14060), .B(n4071), .Z(n14062) );
  NANDN U15904 ( .A(b[0]), .B(a[269]), .Z(n14061) );
  NAND U15905 ( .A(n14062), .B(n14061), .Z(n14109) );
  XOR U15906 ( .A(a[266]), .B(n42085), .Z(n14105) );
  AND U15907 ( .A(a[262]), .B(b[7]), .Z(n14106) );
  XNOR U15908 ( .A(n14107), .B(n14106), .Z(n14108) );
  XNOR U15909 ( .A(n14109), .B(n14108), .Z(n14114) );
  XOR U15910 ( .A(n14115), .B(n14114), .Z(n14093) );
  NANDN U15911 ( .A(n14065), .B(n14064), .Z(n14069) );
  NANDN U15912 ( .A(n14067), .B(n14066), .Z(n14068) );
  AND U15913 ( .A(n14069), .B(n14068), .Z(n14092) );
  XNOR U15914 ( .A(n14093), .B(n14092), .Z(n14094) );
  NANDN U15915 ( .A(n14071), .B(n14070), .Z(n14075) );
  NAND U15916 ( .A(n14073), .B(n14072), .Z(n14074) );
  NAND U15917 ( .A(n14075), .B(n14074), .Z(n14095) );
  XNOR U15918 ( .A(n14094), .B(n14095), .Z(n14086) );
  XNOR U15919 ( .A(n14087), .B(n14086), .Z(n14088) );
  XNOR U15920 ( .A(n14089), .B(n14088), .Z(n14081) );
  XNOR U15921 ( .A(sreg[1286]), .B(n14081), .Z(n14083) );
  NANDN U15922 ( .A(sreg[1285]), .B(n14076), .Z(n14080) );
  NAND U15923 ( .A(n14078), .B(n14077), .Z(n14079) );
  NAND U15924 ( .A(n14080), .B(n14079), .Z(n14082) );
  XNOR U15925 ( .A(n14083), .B(n14082), .Z(c[1286]) );
  NANDN U15926 ( .A(sreg[1286]), .B(n14081), .Z(n14085) );
  NAND U15927 ( .A(n14083), .B(n14082), .Z(n14084) );
  AND U15928 ( .A(n14085), .B(n14084), .Z(n14120) );
  NANDN U15929 ( .A(n14087), .B(n14086), .Z(n14091) );
  NANDN U15930 ( .A(n14089), .B(n14088), .Z(n14090) );
  AND U15931 ( .A(n14091), .B(n14090), .Z(n14125) );
  NANDN U15932 ( .A(n14093), .B(n14092), .Z(n14097) );
  NANDN U15933 ( .A(n14095), .B(n14094), .Z(n14096) );
  AND U15934 ( .A(n14097), .B(n14096), .Z(n14124) );
  NAND U15935 ( .A(n42143), .B(n14098), .Z(n14100) );
  XNOR U15936 ( .A(a[265]), .B(n4109), .Z(n14135) );
  NAND U15937 ( .A(n42144), .B(n14135), .Z(n14099) );
  AND U15938 ( .A(n14100), .B(n14099), .Z(n14150) );
  XOR U15939 ( .A(a[269]), .B(n42012), .Z(n14138) );
  XNOR U15940 ( .A(n14150), .B(n14149), .Z(n14152) );
  AND U15941 ( .A(a[271]), .B(b[0]), .Z(n14102) );
  XNOR U15942 ( .A(n14102), .B(n4071), .Z(n14104) );
  NANDN U15943 ( .A(b[0]), .B(a[270]), .Z(n14103) );
  NAND U15944 ( .A(n14104), .B(n14103), .Z(n14146) );
  XOR U15945 ( .A(a[267]), .B(n42085), .Z(n14139) );
  AND U15946 ( .A(a[263]), .B(b[7]), .Z(n14143) );
  XNOR U15947 ( .A(n14144), .B(n14143), .Z(n14145) );
  XNOR U15948 ( .A(n14146), .B(n14145), .Z(n14151) );
  XOR U15949 ( .A(n14152), .B(n14151), .Z(n14130) );
  NANDN U15950 ( .A(n14107), .B(n14106), .Z(n14111) );
  NANDN U15951 ( .A(n14109), .B(n14108), .Z(n14110) );
  AND U15952 ( .A(n14111), .B(n14110), .Z(n14129) );
  XNOR U15953 ( .A(n14130), .B(n14129), .Z(n14131) );
  NANDN U15954 ( .A(n14113), .B(n14112), .Z(n14117) );
  NAND U15955 ( .A(n14115), .B(n14114), .Z(n14116) );
  NAND U15956 ( .A(n14117), .B(n14116), .Z(n14132) );
  XNOR U15957 ( .A(n14131), .B(n14132), .Z(n14123) );
  XOR U15958 ( .A(n14124), .B(n14123), .Z(n14126) );
  XOR U15959 ( .A(n14125), .B(n14126), .Z(n14118) );
  XNOR U15960 ( .A(n14118), .B(sreg[1287]), .Z(n14119) );
  XOR U15961 ( .A(n14120), .B(n14119), .Z(c[1287]) );
  NANDN U15962 ( .A(n14118), .B(sreg[1287]), .Z(n14122) );
  NAND U15963 ( .A(n14120), .B(n14119), .Z(n14121) );
  AND U15964 ( .A(n14122), .B(n14121), .Z(n14189) );
  NANDN U15965 ( .A(n14124), .B(n14123), .Z(n14128) );
  OR U15966 ( .A(n14126), .B(n14125), .Z(n14127) );
  AND U15967 ( .A(n14128), .B(n14127), .Z(n14158) );
  NANDN U15968 ( .A(n14130), .B(n14129), .Z(n14134) );
  NANDN U15969 ( .A(n14132), .B(n14131), .Z(n14133) );
  AND U15970 ( .A(n14134), .B(n14133), .Z(n14156) );
  NAND U15971 ( .A(n42143), .B(n14135), .Z(n14137) );
  XNOR U15972 ( .A(a[266]), .B(n4109), .Z(n14167) );
  NAND U15973 ( .A(n42144), .B(n14167), .Z(n14136) );
  AND U15974 ( .A(n14137), .B(n14136), .Z(n14182) );
  XOR U15975 ( .A(a[270]), .B(n42012), .Z(n14170) );
  XNOR U15976 ( .A(n14182), .B(n14181), .Z(n14184) );
  XOR U15977 ( .A(a[268]), .B(n42085), .Z(n14174) );
  AND U15978 ( .A(a[264]), .B(b[7]), .Z(n14175) );
  XNOR U15979 ( .A(n14176), .B(n14175), .Z(n14177) );
  AND U15980 ( .A(a[272]), .B(b[0]), .Z(n14140) );
  XNOR U15981 ( .A(n14140), .B(n4071), .Z(n14142) );
  NANDN U15982 ( .A(b[0]), .B(a[271]), .Z(n14141) );
  NAND U15983 ( .A(n14142), .B(n14141), .Z(n14178) );
  XNOR U15984 ( .A(n14177), .B(n14178), .Z(n14183) );
  XOR U15985 ( .A(n14184), .B(n14183), .Z(n14162) );
  NANDN U15986 ( .A(n14144), .B(n14143), .Z(n14148) );
  NANDN U15987 ( .A(n14146), .B(n14145), .Z(n14147) );
  AND U15988 ( .A(n14148), .B(n14147), .Z(n14161) );
  XNOR U15989 ( .A(n14162), .B(n14161), .Z(n14163) );
  NANDN U15990 ( .A(n14150), .B(n14149), .Z(n14154) );
  NAND U15991 ( .A(n14152), .B(n14151), .Z(n14153) );
  NAND U15992 ( .A(n14154), .B(n14153), .Z(n14164) );
  XNOR U15993 ( .A(n14163), .B(n14164), .Z(n14155) );
  XNOR U15994 ( .A(n14156), .B(n14155), .Z(n14157) );
  XNOR U15995 ( .A(n14158), .B(n14157), .Z(n14187) );
  XNOR U15996 ( .A(sreg[1288]), .B(n14187), .Z(n14188) );
  XNOR U15997 ( .A(n14189), .B(n14188), .Z(c[1288]) );
  NANDN U15998 ( .A(n14156), .B(n14155), .Z(n14160) );
  NANDN U15999 ( .A(n14158), .B(n14157), .Z(n14159) );
  AND U16000 ( .A(n14160), .B(n14159), .Z(n14195) );
  NANDN U16001 ( .A(n14162), .B(n14161), .Z(n14166) );
  NANDN U16002 ( .A(n14164), .B(n14163), .Z(n14165) );
  AND U16003 ( .A(n14166), .B(n14165), .Z(n14193) );
  NAND U16004 ( .A(n42143), .B(n14167), .Z(n14169) );
  XNOR U16005 ( .A(a[267]), .B(n4110), .Z(n14204) );
  NAND U16006 ( .A(n42144), .B(n14204), .Z(n14168) );
  AND U16007 ( .A(n14169), .B(n14168), .Z(n14219) );
  XOR U16008 ( .A(a[271]), .B(n42012), .Z(n14207) );
  XNOR U16009 ( .A(n14219), .B(n14218), .Z(n14221) );
  AND U16010 ( .A(a[273]), .B(b[0]), .Z(n14171) );
  XNOR U16011 ( .A(n14171), .B(n4071), .Z(n14173) );
  NANDN U16012 ( .A(b[0]), .B(a[272]), .Z(n14172) );
  NAND U16013 ( .A(n14173), .B(n14172), .Z(n14215) );
  XOR U16014 ( .A(a[269]), .B(n42085), .Z(n14211) );
  AND U16015 ( .A(a[265]), .B(b[7]), .Z(n14212) );
  XNOR U16016 ( .A(n14213), .B(n14212), .Z(n14214) );
  XNOR U16017 ( .A(n14215), .B(n14214), .Z(n14220) );
  XOR U16018 ( .A(n14221), .B(n14220), .Z(n14199) );
  NANDN U16019 ( .A(n14176), .B(n14175), .Z(n14180) );
  NANDN U16020 ( .A(n14178), .B(n14177), .Z(n14179) );
  AND U16021 ( .A(n14180), .B(n14179), .Z(n14198) );
  XNOR U16022 ( .A(n14199), .B(n14198), .Z(n14200) );
  NANDN U16023 ( .A(n14182), .B(n14181), .Z(n14186) );
  NAND U16024 ( .A(n14184), .B(n14183), .Z(n14185) );
  NAND U16025 ( .A(n14186), .B(n14185), .Z(n14201) );
  XNOR U16026 ( .A(n14200), .B(n14201), .Z(n14192) );
  XNOR U16027 ( .A(n14193), .B(n14192), .Z(n14194) );
  XNOR U16028 ( .A(n14195), .B(n14194), .Z(n14224) );
  XNOR U16029 ( .A(sreg[1289]), .B(n14224), .Z(n14226) );
  NANDN U16030 ( .A(sreg[1288]), .B(n14187), .Z(n14191) );
  NAND U16031 ( .A(n14189), .B(n14188), .Z(n14190) );
  NAND U16032 ( .A(n14191), .B(n14190), .Z(n14225) );
  XNOR U16033 ( .A(n14226), .B(n14225), .Z(c[1289]) );
  NANDN U16034 ( .A(n14193), .B(n14192), .Z(n14197) );
  NANDN U16035 ( .A(n14195), .B(n14194), .Z(n14196) );
  AND U16036 ( .A(n14197), .B(n14196), .Z(n14236) );
  NANDN U16037 ( .A(n14199), .B(n14198), .Z(n14203) );
  NANDN U16038 ( .A(n14201), .B(n14200), .Z(n14202) );
  AND U16039 ( .A(n14203), .B(n14202), .Z(n14235) );
  NAND U16040 ( .A(n42143), .B(n14204), .Z(n14206) );
  XNOR U16041 ( .A(a[268]), .B(n4110), .Z(n14246) );
  NAND U16042 ( .A(n42144), .B(n14246), .Z(n14205) );
  AND U16043 ( .A(n14206), .B(n14205), .Z(n14261) );
  XOR U16044 ( .A(a[272]), .B(n42012), .Z(n14249) );
  XNOR U16045 ( .A(n14261), .B(n14260), .Z(n14263) );
  AND U16046 ( .A(a[274]), .B(b[0]), .Z(n14208) );
  XNOR U16047 ( .A(n14208), .B(n4071), .Z(n14210) );
  NANDN U16048 ( .A(b[0]), .B(a[273]), .Z(n14209) );
  NAND U16049 ( .A(n14210), .B(n14209), .Z(n14257) );
  XOR U16050 ( .A(a[270]), .B(n42085), .Z(n14253) );
  AND U16051 ( .A(a[266]), .B(b[7]), .Z(n14254) );
  XNOR U16052 ( .A(n14255), .B(n14254), .Z(n14256) );
  XNOR U16053 ( .A(n14257), .B(n14256), .Z(n14262) );
  XOR U16054 ( .A(n14263), .B(n14262), .Z(n14241) );
  NANDN U16055 ( .A(n14213), .B(n14212), .Z(n14217) );
  NANDN U16056 ( .A(n14215), .B(n14214), .Z(n14216) );
  AND U16057 ( .A(n14217), .B(n14216), .Z(n14240) );
  XNOR U16058 ( .A(n14241), .B(n14240), .Z(n14242) );
  NANDN U16059 ( .A(n14219), .B(n14218), .Z(n14223) );
  NAND U16060 ( .A(n14221), .B(n14220), .Z(n14222) );
  NAND U16061 ( .A(n14223), .B(n14222), .Z(n14243) );
  XNOR U16062 ( .A(n14242), .B(n14243), .Z(n14234) );
  XOR U16063 ( .A(n14235), .B(n14234), .Z(n14237) );
  XOR U16064 ( .A(n14236), .B(n14237), .Z(n14229) );
  XNOR U16065 ( .A(n14229), .B(sreg[1290]), .Z(n14231) );
  NANDN U16066 ( .A(sreg[1289]), .B(n14224), .Z(n14228) );
  NAND U16067 ( .A(n14226), .B(n14225), .Z(n14227) );
  AND U16068 ( .A(n14228), .B(n14227), .Z(n14230) );
  XOR U16069 ( .A(n14231), .B(n14230), .Z(c[1290]) );
  NANDN U16070 ( .A(n14229), .B(sreg[1290]), .Z(n14233) );
  NAND U16071 ( .A(n14231), .B(n14230), .Z(n14232) );
  AND U16072 ( .A(n14233), .B(n14232), .Z(n14300) );
  NANDN U16073 ( .A(n14235), .B(n14234), .Z(n14239) );
  OR U16074 ( .A(n14237), .B(n14236), .Z(n14238) );
  AND U16075 ( .A(n14239), .B(n14238), .Z(n14269) );
  NANDN U16076 ( .A(n14241), .B(n14240), .Z(n14245) );
  NANDN U16077 ( .A(n14243), .B(n14242), .Z(n14244) );
  AND U16078 ( .A(n14245), .B(n14244), .Z(n14267) );
  NAND U16079 ( .A(n42143), .B(n14246), .Z(n14248) );
  XNOR U16080 ( .A(a[269]), .B(n4110), .Z(n14278) );
  NAND U16081 ( .A(n42144), .B(n14278), .Z(n14247) );
  AND U16082 ( .A(n14248), .B(n14247), .Z(n14293) );
  XOR U16083 ( .A(a[273]), .B(n42012), .Z(n14281) );
  XNOR U16084 ( .A(n14293), .B(n14292), .Z(n14295) );
  AND U16085 ( .A(a[275]), .B(b[0]), .Z(n14250) );
  XNOR U16086 ( .A(n14250), .B(n4071), .Z(n14252) );
  NANDN U16087 ( .A(b[0]), .B(a[274]), .Z(n14251) );
  NAND U16088 ( .A(n14252), .B(n14251), .Z(n14289) );
  XOR U16089 ( .A(a[271]), .B(n42085), .Z(n14285) );
  AND U16090 ( .A(a[267]), .B(b[7]), .Z(n14286) );
  XNOR U16091 ( .A(n14287), .B(n14286), .Z(n14288) );
  XNOR U16092 ( .A(n14289), .B(n14288), .Z(n14294) );
  XOR U16093 ( .A(n14295), .B(n14294), .Z(n14273) );
  NANDN U16094 ( .A(n14255), .B(n14254), .Z(n14259) );
  NANDN U16095 ( .A(n14257), .B(n14256), .Z(n14258) );
  AND U16096 ( .A(n14259), .B(n14258), .Z(n14272) );
  XNOR U16097 ( .A(n14273), .B(n14272), .Z(n14274) );
  NANDN U16098 ( .A(n14261), .B(n14260), .Z(n14265) );
  NAND U16099 ( .A(n14263), .B(n14262), .Z(n14264) );
  NAND U16100 ( .A(n14265), .B(n14264), .Z(n14275) );
  XNOR U16101 ( .A(n14274), .B(n14275), .Z(n14266) );
  XNOR U16102 ( .A(n14267), .B(n14266), .Z(n14268) );
  XNOR U16103 ( .A(n14269), .B(n14268), .Z(n14298) );
  XNOR U16104 ( .A(sreg[1291]), .B(n14298), .Z(n14299) );
  XNOR U16105 ( .A(n14300), .B(n14299), .Z(c[1291]) );
  NANDN U16106 ( .A(n14267), .B(n14266), .Z(n14271) );
  NANDN U16107 ( .A(n14269), .B(n14268), .Z(n14270) );
  AND U16108 ( .A(n14271), .B(n14270), .Z(n14306) );
  NANDN U16109 ( .A(n14273), .B(n14272), .Z(n14277) );
  NANDN U16110 ( .A(n14275), .B(n14274), .Z(n14276) );
  AND U16111 ( .A(n14277), .B(n14276), .Z(n14304) );
  NAND U16112 ( .A(n42143), .B(n14278), .Z(n14280) );
  XNOR U16113 ( .A(a[270]), .B(n4110), .Z(n14315) );
  NAND U16114 ( .A(n42144), .B(n14315), .Z(n14279) );
  AND U16115 ( .A(n14280), .B(n14279), .Z(n14330) );
  XOR U16116 ( .A(a[274]), .B(n42012), .Z(n14318) );
  XNOR U16117 ( .A(n14330), .B(n14329), .Z(n14332) );
  AND U16118 ( .A(a[276]), .B(b[0]), .Z(n14282) );
  XNOR U16119 ( .A(n14282), .B(n4071), .Z(n14284) );
  NANDN U16120 ( .A(b[0]), .B(a[275]), .Z(n14283) );
  NAND U16121 ( .A(n14284), .B(n14283), .Z(n14326) );
  XOR U16122 ( .A(a[272]), .B(n42085), .Z(n14319) );
  AND U16123 ( .A(a[268]), .B(b[7]), .Z(n14323) );
  XNOR U16124 ( .A(n14324), .B(n14323), .Z(n14325) );
  XNOR U16125 ( .A(n14326), .B(n14325), .Z(n14331) );
  XOR U16126 ( .A(n14332), .B(n14331), .Z(n14310) );
  NANDN U16127 ( .A(n14287), .B(n14286), .Z(n14291) );
  NANDN U16128 ( .A(n14289), .B(n14288), .Z(n14290) );
  AND U16129 ( .A(n14291), .B(n14290), .Z(n14309) );
  XNOR U16130 ( .A(n14310), .B(n14309), .Z(n14311) );
  NANDN U16131 ( .A(n14293), .B(n14292), .Z(n14297) );
  NAND U16132 ( .A(n14295), .B(n14294), .Z(n14296) );
  NAND U16133 ( .A(n14297), .B(n14296), .Z(n14312) );
  XNOR U16134 ( .A(n14311), .B(n14312), .Z(n14303) );
  XNOR U16135 ( .A(n14304), .B(n14303), .Z(n14305) );
  XNOR U16136 ( .A(n14306), .B(n14305), .Z(n14335) );
  XNOR U16137 ( .A(sreg[1292]), .B(n14335), .Z(n14337) );
  NANDN U16138 ( .A(sreg[1291]), .B(n14298), .Z(n14302) );
  NAND U16139 ( .A(n14300), .B(n14299), .Z(n14301) );
  NAND U16140 ( .A(n14302), .B(n14301), .Z(n14336) );
  XNOR U16141 ( .A(n14337), .B(n14336), .Z(c[1292]) );
  NANDN U16142 ( .A(n14304), .B(n14303), .Z(n14308) );
  NANDN U16143 ( .A(n14306), .B(n14305), .Z(n14307) );
  AND U16144 ( .A(n14308), .B(n14307), .Z(n14343) );
  NANDN U16145 ( .A(n14310), .B(n14309), .Z(n14314) );
  NANDN U16146 ( .A(n14312), .B(n14311), .Z(n14313) );
  AND U16147 ( .A(n14314), .B(n14313), .Z(n14341) );
  NAND U16148 ( .A(n42143), .B(n14315), .Z(n14317) );
  XNOR U16149 ( .A(a[271]), .B(n4110), .Z(n14352) );
  NAND U16150 ( .A(n42144), .B(n14352), .Z(n14316) );
  AND U16151 ( .A(n14317), .B(n14316), .Z(n14367) );
  XOR U16152 ( .A(a[275]), .B(n42012), .Z(n14355) );
  XNOR U16153 ( .A(n14367), .B(n14366), .Z(n14369) );
  XOR U16154 ( .A(a[273]), .B(n42085), .Z(n14359) );
  AND U16155 ( .A(a[269]), .B(b[7]), .Z(n14360) );
  XNOR U16156 ( .A(n14361), .B(n14360), .Z(n14362) );
  AND U16157 ( .A(a[277]), .B(b[0]), .Z(n14320) );
  XNOR U16158 ( .A(n14320), .B(n4071), .Z(n14322) );
  NANDN U16159 ( .A(b[0]), .B(a[276]), .Z(n14321) );
  NAND U16160 ( .A(n14322), .B(n14321), .Z(n14363) );
  XNOR U16161 ( .A(n14362), .B(n14363), .Z(n14368) );
  XOR U16162 ( .A(n14369), .B(n14368), .Z(n14347) );
  NANDN U16163 ( .A(n14324), .B(n14323), .Z(n14328) );
  NANDN U16164 ( .A(n14326), .B(n14325), .Z(n14327) );
  AND U16165 ( .A(n14328), .B(n14327), .Z(n14346) );
  XNOR U16166 ( .A(n14347), .B(n14346), .Z(n14348) );
  NANDN U16167 ( .A(n14330), .B(n14329), .Z(n14334) );
  NAND U16168 ( .A(n14332), .B(n14331), .Z(n14333) );
  NAND U16169 ( .A(n14334), .B(n14333), .Z(n14349) );
  XNOR U16170 ( .A(n14348), .B(n14349), .Z(n14340) );
  XNOR U16171 ( .A(n14341), .B(n14340), .Z(n14342) );
  XNOR U16172 ( .A(n14343), .B(n14342), .Z(n14372) );
  XNOR U16173 ( .A(sreg[1293]), .B(n14372), .Z(n14374) );
  NANDN U16174 ( .A(sreg[1292]), .B(n14335), .Z(n14339) );
  NAND U16175 ( .A(n14337), .B(n14336), .Z(n14338) );
  NAND U16176 ( .A(n14339), .B(n14338), .Z(n14373) );
  XNOR U16177 ( .A(n14374), .B(n14373), .Z(c[1293]) );
  NANDN U16178 ( .A(n14341), .B(n14340), .Z(n14345) );
  NANDN U16179 ( .A(n14343), .B(n14342), .Z(n14344) );
  AND U16180 ( .A(n14345), .B(n14344), .Z(n14380) );
  NANDN U16181 ( .A(n14347), .B(n14346), .Z(n14351) );
  NANDN U16182 ( .A(n14349), .B(n14348), .Z(n14350) );
  AND U16183 ( .A(n14351), .B(n14350), .Z(n14378) );
  NAND U16184 ( .A(n42143), .B(n14352), .Z(n14354) );
  XNOR U16185 ( .A(a[272]), .B(n4110), .Z(n14389) );
  NAND U16186 ( .A(n42144), .B(n14389), .Z(n14353) );
  AND U16187 ( .A(n14354), .B(n14353), .Z(n14404) );
  XOR U16188 ( .A(a[276]), .B(n42012), .Z(n14392) );
  XNOR U16189 ( .A(n14404), .B(n14403), .Z(n14406) );
  AND U16190 ( .A(a[278]), .B(b[0]), .Z(n14356) );
  XNOR U16191 ( .A(n14356), .B(n4071), .Z(n14358) );
  NANDN U16192 ( .A(b[0]), .B(a[277]), .Z(n14357) );
  NAND U16193 ( .A(n14358), .B(n14357), .Z(n14400) );
  XOR U16194 ( .A(a[274]), .B(n42085), .Z(n14396) );
  AND U16195 ( .A(a[270]), .B(b[7]), .Z(n14397) );
  XNOR U16196 ( .A(n14398), .B(n14397), .Z(n14399) );
  XNOR U16197 ( .A(n14400), .B(n14399), .Z(n14405) );
  XOR U16198 ( .A(n14406), .B(n14405), .Z(n14384) );
  NANDN U16199 ( .A(n14361), .B(n14360), .Z(n14365) );
  NANDN U16200 ( .A(n14363), .B(n14362), .Z(n14364) );
  AND U16201 ( .A(n14365), .B(n14364), .Z(n14383) );
  XNOR U16202 ( .A(n14384), .B(n14383), .Z(n14385) );
  NANDN U16203 ( .A(n14367), .B(n14366), .Z(n14371) );
  NAND U16204 ( .A(n14369), .B(n14368), .Z(n14370) );
  NAND U16205 ( .A(n14371), .B(n14370), .Z(n14386) );
  XNOR U16206 ( .A(n14385), .B(n14386), .Z(n14377) );
  XNOR U16207 ( .A(n14378), .B(n14377), .Z(n14379) );
  XNOR U16208 ( .A(n14380), .B(n14379), .Z(n14409) );
  XNOR U16209 ( .A(sreg[1294]), .B(n14409), .Z(n14411) );
  NANDN U16210 ( .A(sreg[1293]), .B(n14372), .Z(n14376) );
  NAND U16211 ( .A(n14374), .B(n14373), .Z(n14375) );
  NAND U16212 ( .A(n14376), .B(n14375), .Z(n14410) );
  XNOR U16213 ( .A(n14411), .B(n14410), .Z(c[1294]) );
  NANDN U16214 ( .A(n14378), .B(n14377), .Z(n14382) );
  NANDN U16215 ( .A(n14380), .B(n14379), .Z(n14381) );
  AND U16216 ( .A(n14382), .B(n14381), .Z(n14417) );
  NANDN U16217 ( .A(n14384), .B(n14383), .Z(n14388) );
  NANDN U16218 ( .A(n14386), .B(n14385), .Z(n14387) );
  AND U16219 ( .A(n14388), .B(n14387), .Z(n14415) );
  NAND U16220 ( .A(n42143), .B(n14389), .Z(n14391) );
  XNOR U16221 ( .A(a[273]), .B(n4110), .Z(n14426) );
  NAND U16222 ( .A(n42144), .B(n14426), .Z(n14390) );
  AND U16223 ( .A(n14391), .B(n14390), .Z(n14441) );
  XOR U16224 ( .A(a[277]), .B(n42012), .Z(n14429) );
  XNOR U16225 ( .A(n14441), .B(n14440), .Z(n14443) );
  AND U16226 ( .A(b[0]), .B(a[279]), .Z(n14393) );
  XOR U16227 ( .A(b[1]), .B(n14393), .Z(n14395) );
  NANDN U16228 ( .A(b[0]), .B(b[1]), .Z(n29564) );
  NANDN U16229 ( .A(n29564), .B(a[278]), .Z(n14394) );
  AND U16230 ( .A(n14395), .B(n14394), .Z(n14436) );
  XOR U16231 ( .A(a[275]), .B(n42085), .Z(n14433) );
  AND U16232 ( .A(a[271]), .B(b[7]), .Z(n14434) );
  XOR U16233 ( .A(n14435), .B(n14434), .Z(n14437) );
  XNOR U16234 ( .A(n14436), .B(n14437), .Z(n14442) );
  XOR U16235 ( .A(n14443), .B(n14442), .Z(n14421) );
  NANDN U16236 ( .A(n14398), .B(n14397), .Z(n14402) );
  NANDN U16237 ( .A(n14400), .B(n14399), .Z(n14401) );
  AND U16238 ( .A(n14402), .B(n14401), .Z(n14420) );
  XNOR U16239 ( .A(n14421), .B(n14420), .Z(n14422) );
  NANDN U16240 ( .A(n14404), .B(n14403), .Z(n14408) );
  NAND U16241 ( .A(n14406), .B(n14405), .Z(n14407) );
  NAND U16242 ( .A(n14408), .B(n14407), .Z(n14423) );
  XNOR U16243 ( .A(n14422), .B(n14423), .Z(n14414) );
  XNOR U16244 ( .A(n14415), .B(n14414), .Z(n14416) );
  XNOR U16245 ( .A(n14417), .B(n14416), .Z(n14446) );
  XNOR U16246 ( .A(sreg[1295]), .B(n14446), .Z(n14448) );
  NANDN U16247 ( .A(sreg[1294]), .B(n14409), .Z(n14413) );
  NAND U16248 ( .A(n14411), .B(n14410), .Z(n14412) );
  NAND U16249 ( .A(n14413), .B(n14412), .Z(n14447) );
  XNOR U16250 ( .A(n14448), .B(n14447), .Z(c[1295]) );
  NANDN U16251 ( .A(n14415), .B(n14414), .Z(n14419) );
  NANDN U16252 ( .A(n14417), .B(n14416), .Z(n14418) );
  AND U16253 ( .A(n14419), .B(n14418), .Z(n14454) );
  NANDN U16254 ( .A(n14421), .B(n14420), .Z(n14425) );
  NANDN U16255 ( .A(n14423), .B(n14422), .Z(n14424) );
  AND U16256 ( .A(n14425), .B(n14424), .Z(n14452) );
  NAND U16257 ( .A(n42143), .B(n14426), .Z(n14428) );
  XNOR U16258 ( .A(a[274]), .B(n4111), .Z(n14463) );
  NAND U16259 ( .A(n42144), .B(n14463), .Z(n14427) );
  AND U16260 ( .A(n14428), .B(n14427), .Z(n14478) );
  XOR U16261 ( .A(a[278]), .B(n42012), .Z(n14466) );
  XNOR U16262 ( .A(n14478), .B(n14477), .Z(n14480) );
  AND U16263 ( .A(a[280]), .B(b[0]), .Z(n14430) );
  XNOR U16264 ( .A(n14430), .B(n4071), .Z(n14432) );
  NANDN U16265 ( .A(b[0]), .B(a[279]), .Z(n14431) );
  NAND U16266 ( .A(n14432), .B(n14431), .Z(n14474) );
  XOR U16267 ( .A(a[276]), .B(n42085), .Z(n14470) );
  AND U16268 ( .A(a[272]), .B(b[7]), .Z(n14471) );
  XNOR U16269 ( .A(n14472), .B(n14471), .Z(n14473) );
  XNOR U16270 ( .A(n14474), .B(n14473), .Z(n14479) );
  XOR U16271 ( .A(n14480), .B(n14479), .Z(n14458) );
  NANDN U16272 ( .A(n14435), .B(n14434), .Z(n14439) );
  NANDN U16273 ( .A(n14437), .B(n14436), .Z(n14438) );
  AND U16274 ( .A(n14439), .B(n14438), .Z(n14457) );
  XNOR U16275 ( .A(n14458), .B(n14457), .Z(n14459) );
  NANDN U16276 ( .A(n14441), .B(n14440), .Z(n14445) );
  NAND U16277 ( .A(n14443), .B(n14442), .Z(n14444) );
  NAND U16278 ( .A(n14445), .B(n14444), .Z(n14460) );
  XNOR U16279 ( .A(n14459), .B(n14460), .Z(n14451) );
  XNOR U16280 ( .A(n14452), .B(n14451), .Z(n14453) );
  XNOR U16281 ( .A(n14454), .B(n14453), .Z(n14483) );
  XNOR U16282 ( .A(sreg[1296]), .B(n14483), .Z(n14485) );
  NANDN U16283 ( .A(sreg[1295]), .B(n14446), .Z(n14450) );
  NAND U16284 ( .A(n14448), .B(n14447), .Z(n14449) );
  NAND U16285 ( .A(n14450), .B(n14449), .Z(n14484) );
  XNOR U16286 ( .A(n14485), .B(n14484), .Z(c[1296]) );
  NANDN U16287 ( .A(n14452), .B(n14451), .Z(n14456) );
  NANDN U16288 ( .A(n14454), .B(n14453), .Z(n14455) );
  AND U16289 ( .A(n14456), .B(n14455), .Z(n14491) );
  NANDN U16290 ( .A(n14458), .B(n14457), .Z(n14462) );
  NANDN U16291 ( .A(n14460), .B(n14459), .Z(n14461) );
  AND U16292 ( .A(n14462), .B(n14461), .Z(n14489) );
  NAND U16293 ( .A(n42143), .B(n14463), .Z(n14465) );
  XNOR U16294 ( .A(a[275]), .B(n4111), .Z(n14500) );
  NAND U16295 ( .A(n42144), .B(n14500), .Z(n14464) );
  AND U16296 ( .A(n14465), .B(n14464), .Z(n14515) );
  XOR U16297 ( .A(a[279]), .B(n42012), .Z(n14503) );
  XNOR U16298 ( .A(n14515), .B(n14514), .Z(n14517) );
  AND U16299 ( .A(a[281]), .B(b[0]), .Z(n14467) );
  XNOR U16300 ( .A(n14467), .B(n4071), .Z(n14469) );
  NANDN U16301 ( .A(b[0]), .B(a[280]), .Z(n14468) );
  NAND U16302 ( .A(n14469), .B(n14468), .Z(n14511) );
  XOR U16303 ( .A(a[277]), .B(n42085), .Z(n14504) );
  AND U16304 ( .A(a[273]), .B(b[7]), .Z(n14508) );
  XNOR U16305 ( .A(n14509), .B(n14508), .Z(n14510) );
  XNOR U16306 ( .A(n14511), .B(n14510), .Z(n14516) );
  XOR U16307 ( .A(n14517), .B(n14516), .Z(n14495) );
  NANDN U16308 ( .A(n14472), .B(n14471), .Z(n14476) );
  NANDN U16309 ( .A(n14474), .B(n14473), .Z(n14475) );
  AND U16310 ( .A(n14476), .B(n14475), .Z(n14494) );
  XNOR U16311 ( .A(n14495), .B(n14494), .Z(n14496) );
  NANDN U16312 ( .A(n14478), .B(n14477), .Z(n14482) );
  NAND U16313 ( .A(n14480), .B(n14479), .Z(n14481) );
  NAND U16314 ( .A(n14482), .B(n14481), .Z(n14497) );
  XNOR U16315 ( .A(n14496), .B(n14497), .Z(n14488) );
  XNOR U16316 ( .A(n14489), .B(n14488), .Z(n14490) );
  XNOR U16317 ( .A(n14491), .B(n14490), .Z(n14520) );
  XNOR U16318 ( .A(sreg[1297]), .B(n14520), .Z(n14522) );
  NANDN U16319 ( .A(sreg[1296]), .B(n14483), .Z(n14487) );
  NAND U16320 ( .A(n14485), .B(n14484), .Z(n14486) );
  NAND U16321 ( .A(n14487), .B(n14486), .Z(n14521) );
  XNOR U16322 ( .A(n14522), .B(n14521), .Z(c[1297]) );
  NANDN U16323 ( .A(n14489), .B(n14488), .Z(n14493) );
  NANDN U16324 ( .A(n14491), .B(n14490), .Z(n14492) );
  AND U16325 ( .A(n14493), .B(n14492), .Z(n14528) );
  NANDN U16326 ( .A(n14495), .B(n14494), .Z(n14499) );
  NANDN U16327 ( .A(n14497), .B(n14496), .Z(n14498) );
  AND U16328 ( .A(n14499), .B(n14498), .Z(n14526) );
  NAND U16329 ( .A(n42143), .B(n14500), .Z(n14502) );
  XNOR U16330 ( .A(a[276]), .B(n4111), .Z(n14537) );
  NAND U16331 ( .A(n42144), .B(n14537), .Z(n14501) );
  AND U16332 ( .A(n14502), .B(n14501), .Z(n14552) );
  XOR U16333 ( .A(a[280]), .B(n42012), .Z(n14540) );
  XNOR U16334 ( .A(n14552), .B(n14551), .Z(n14554) );
  XOR U16335 ( .A(a[278]), .B(n42085), .Z(n14541) );
  AND U16336 ( .A(a[274]), .B(b[7]), .Z(n14545) );
  XNOR U16337 ( .A(n14546), .B(n14545), .Z(n14547) );
  AND U16338 ( .A(a[282]), .B(b[0]), .Z(n14505) );
  XNOR U16339 ( .A(n14505), .B(n4071), .Z(n14507) );
  NANDN U16340 ( .A(b[0]), .B(a[281]), .Z(n14506) );
  NAND U16341 ( .A(n14507), .B(n14506), .Z(n14548) );
  XNOR U16342 ( .A(n14547), .B(n14548), .Z(n14553) );
  XOR U16343 ( .A(n14554), .B(n14553), .Z(n14532) );
  NANDN U16344 ( .A(n14509), .B(n14508), .Z(n14513) );
  NANDN U16345 ( .A(n14511), .B(n14510), .Z(n14512) );
  AND U16346 ( .A(n14513), .B(n14512), .Z(n14531) );
  XNOR U16347 ( .A(n14532), .B(n14531), .Z(n14533) );
  NANDN U16348 ( .A(n14515), .B(n14514), .Z(n14519) );
  NAND U16349 ( .A(n14517), .B(n14516), .Z(n14518) );
  NAND U16350 ( .A(n14519), .B(n14518), .Z(n14534) );
  XNOR U16351 ( .A(n14533), .B(n14534), .Z(n14525) );
  XNOR U16352 ( .A(n14526), .B(n14525), .Z(n14527) );
  XNOR U16353 ( .A(n14528), .B(n14527), .Z(n14557) );
  XNOR U16354 ( .A(sreg[1298]), .B(n14557), .Z(n14559) );
  NANDN U16355 ( .A(sreg[1297]), .B(n14520), .Z(n14524) );
  NAND U16356 ( .A(n14522), .B(n14521), .Z(n14523) );
  NAND U16357 ( .A(n14524), .B(n14523), .Z(n14558) );
  XNOR U16358 ( .A(n14559), .B(n14558), .Z(c[1298]) );
  NANDN U16359 ( .A(n14526), .B(n14525), .Z(n14530) );
  NANDN U16360 ( .A(n14528), .B(n14527), .Z(n14529) );
  AND U16361 ( .A(n14530), .B(n14529), .Z(n14565) );
  NANDN U16362 ( .A(n14532), .B(n14531), .Z(n14536) );
  NANDN U16363 ( .A(n14534), .B(n14533), .Z(n14535) );
  AND U16364 ( .A(n14536), .B(n14535), .Z(n14563) );
  NAND U16365 ( .A(n42143), .B(n14537), .Z(n14539) );
  XNOR U16366 ( .A(a[277]), .B(n4111), .Z(n14574) );
  NAND U16367 ( .A(n42144), .B(n14574), .Z(n14538) );
  AND U16368 ( .A(n14539), .B(n14538), .Z(n14589) );
  XOR U16369 ( .A(a[281]), .B(n42012), .Z(n14577) );
  XNOR U16370 ( .A(n14589), .B(n14588), .Z(n14591) );
  XOR U16371 ( .A(a[279]), .B(n42085), .Z(n14581) );
  AND U16372 ( .A(a[275]), .B(b[7]), .Z(n14582) );
  XNOR U16373 ( .A(n14583), .B(n14582), .Z(n14584) );
  AND U16374 ( .A(a[283]), .B(b[0]), .Z(n14542) );
  XNOR U16375 ( .A(n14542), .B(n4071), .Z(n14544) );
  NANDN U16376 ( .A(b[0]), .B(a[282]), .Z(n14543) );
  NAND U16377 ( .A(n14544), .B(n14543), .Z(n14585) );
  XNOR U16378 ( .A(n14584), .B(n14585), .Z(n14590) );
  XOR U16379 ( .A(n14591), .B(n14590), .Z(n14569) );
  NANDN U16380 ( .A(n14546), .B(n14545), .Z(n14550) );
  NANDN U16381 ( .A(n14548), .B(n14547), .Z(n14549) );
  AND U16382 ( .A(n14550), .B(n14549), .Z(n14568) );
  XNOR U16383 ( .A(n14569), .B(n14568), .Z(n14570) );
  NANDN U16384 ( .A(n14552), .B(n14551), .Z(n14556) );
  NAND U16385 ( .A(n14554), .B(n14553), .Z(n14555) );
  NAND U16386 ( .A(n14556), .B(n14555), .Z(n14571) );
  XNOR U16387 ( .A(n14570), .B(n14571), .Z(n14562) );
  XNOR U16388 ( .A(n14563), .B(n14562), .Z(n14564) );
  XNOR U16389 ( .A(n14565), .B(n14564), .Z(n14594) );
  XNOR U16390 ( .A(sreg[1299]), .B(n14594), .Z(n14596) );
  NANDN U16391 ( .A(sreg[1298]), .B(n14557), .Z(n14561) );
  NAND U16392 ( .A(n14559), .B(n14558), .Z(n14560) );
  NAND U16393 ( .A(n14561), .B(n14560), .Z(n14595) );
  XNOR U16394 ( .A(n14596), .B(n14595), .Z(c[1299]) );
  NANDN U16395 ( .A(n14563), .B(n14562), .Z(n14567) );
  NANDN U16396 ( .A(n14565), .B(n14564), .Z(n14566) );
  AND U16397 ( .A(n14567), .B(n14566), .Z(n14602) );
  NANDN U16398 ( .A(n14569), .B(n14568), .Z(n14573) );
  NANDN U16399 ( .A(n14571), .B(n14570), .Z(n14572) );
  AND U16400 ( .A(n14573), .B(n14572), .Z(n14600) );
  NAND U16401 ( .A(n42143), .B(n14574), .Z(n14576) );
  XNOR U16402 ( .A(a[278]), .B(n4111), .Z(n14611) );
  NAND U16403 ( .A(n42144), .B(n14611), .Z(n14575) );
  AND U16404 ( .A(n14576), .B(n14575), .Z(n14626) );
  XOR U16405 ( .A(a[282]), .B(n42012), .Z(n14614) );
  XNOR U16406 ( .A(n14626), .B(n14625), .Z(n14628) );
  AND U16407 ( .A(a[284]), .B(b[0]), .Z(n14578) );
  XNOR U16408 ( .A(n14578), .B(n4071), .Z(n14580) );
  NANDN U16409 ( .A(b[0]), .B(a[283]), .Z(n14579) );
  NAND U16410 ( .A(n14580), .B(n14579), .Z(n14622) );
  XOR U16411 ( .A(a[280]), .B(n42085), .Z(n14618) );
  AND U16412 ( .A(a[276]), .B(b[7]), .Z(n14619) );
  XNOR U16413 ( .A(n14620), .B(n14619), .Z(n14621) );
  XNOR U16414 ( .A(n14622), .B(n14621), .Z(n14627) );
  XOR U16415 ( .A(n14628), .B(n14627), .Z(n14606) );
  NANDN U16416 ( .A(n14583), .B(n14582), .Z(n14587) );
  NANDN U16417 ( .A(n14585), .B(n14584), .Z(n14586) );
  AND U16418 ( .A(n14587), .B(n14586), .Z(n14605) );
  XNOR U16419 ( .A(n14606), .B(n14605), .Z(n14607) );
  NANDN U16420 ( .A(n14589), .B(n14588), .Z(n14593) );
  NAND U16421 ( .A(n14591), .B(n14590), .Z(n14592) );
  NAND U16422 ( .A(n14593), .B(n14592), .Z(n14608) );
  XNOR U16423 ( .A(n14607), .B(n14608), .Z(n14599) );
  XNOR U16424 ( .A(n14600), .B(n14599), .Z(n14601) );
  XNOR U16425 ( .A(n14602), .B(n14601), .Z(n14631) );
  XNOR U16426 ( .A(sreg[1300]), .B(n14631), .Z(n14633) );
  NANDN U16427 ( .A(sreg[1299]), .B(n14594), .Z(n14598) );
  NAND U16428 ( .A(n14596), .B(n14595), .Z(n14597) );
  NAND U16429 ( .A(n14598), .B(n14597), .Z(n14632) );
  XNOR U16430 ( .A(n14633), .B(n14632), .Z(c[1300]) );
  NANDN U16431 ( .A(n14600), .B(n14599), .Z(n14604) );
  NANDN U16432 ( .A(n14602), .B(n14601), .Z(n14603) );
  AND U16433 ( .A(n14604), .B(n14603), .Z(n14639) );
  NANDN U16434 ( .A(n14606), .B(n14605), .Z(n14610) );
  NANDN U16435 ( .A(n14608), .B(n14607), .Z(n14609) );
  AND U16436 ( .A(n14610), .B(n14609), .Z(n14637) );
  NAND U16437 ( .A(n42143), .B(n14611), .Z(n14613) );
  XNOR U16438 ( .A(a[279]), .B(n4111), .Z(n14648) );
  NAND U16439 ( .A(n42144), .B(n14648), .Z(n14612) );
  AND U16440 ( .A(n14613), .B(n14612), .Z(n14663) );
  XOR U16441 ( .A(a[283]), .B(n42012), .Z(n14651) );
  XNOR U16442 ( .A(n14663), .B(n14662), .Z(n14665) );
  AND U16443 ( .A(a[285]), .B(b[0]), .Z(n14615) );
  XNOR U16444 ( .A(n14615), .B(n4071), .Z(n14617) );
  NANDN U16445 ( .A(b[0]), .B(a[284]), .Z(n14616) );
  NAND U16446 ( .A(n14617), .B(n14616), .Z(n14659) );
  XOR U16447 ( .A(a[281]), .B(n42085), .Z(n14655) );
  AND U16448 ( .A(a[277]), .B(b[7]), .Z(n14656) );
  XNOR U16449 ( .A(n14657), .B(n14656), .Z(n14658) );
  XNOR U16450 ( .A(n14659), .B(n14658), .Z(n14664) );
  XOR U16451 ( .A(n14665), .B(n14664), .Z(n14643) );
  NANDN U16452 ( .A(n14620), .B(n14619), .Z(n14624) );
  NANDN U16453 ( .A(n14622), .B(n14621), .Z(n14623) );
  AND U16454 ( .A(n14624), .B(n14623), .Z(n14642) );
  XNOR U16455 ( .A(n14643), .B(n14642), .Z(n14644) );
  NANDN U16456 ( .A(n14626), .B(n14625), .Z(n14630) );
  NAND U16457 ( .A(n14628), .B(n14627), .Z(n14629) );
  NAND U16458 ( .A(n14630), .B(n14629), .Z(n14645) );
  XNOR U16459 ( .A(n14644), .B(n14645), .Z(n14636) );
  XNOR U16460 ( .A(n14637), .B(n14636), .Z(n14638) );
  XNOR U16461 ( .A(n14639), .B(n14638), .Z(n14668) );
  XNOR U16462 ( .A(sreg[1301]), .B(n14668), .Z(n14670) );
  NANDN U16463 ( .A(sreg[1300]), .B(n14631), .Z(n14635) );
  NAND U16464 ( .A(n14633), .B(n14632), .Z(n14634) );
  NAND U16465 ( .A(n14635), .B(n14634), .Z(n14669) );
  XNOR U16466 ( .A(n14670), .B(n14669), .Z(c[1301]) );
  NANDN U16467 ( .A(n14637), .B(n14636), .Z(n14641) );
  NANDN U16468 ( .A(n14639), .B(n14638), .Z(n14640) );
  AND U16469 ( .A(n14641), .B(n14640), .Z(n14676) );
  NANDN U16470 ( .A(n14643), .B(n14642), .Z(n14647) );
  NANDN U16471 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U16472 ( .A(n14647), .B(n14646), .Z(n14674) );
  NAND U16473 ( .A(n42143), .B(n14648), .Z(n14650) );
  XNOR U16474 ( .A(a[280]), .B(n4111), .Z(n14685) );
  NAND U16475 ( .A(n42144), .B(n14685), .Z(n14649) );
  AND U16476 ( .A(n14650), .B(n14649), .Z(n14700) );
  XOR U16477 ( .A(a[284]), .B(n42012), .Z(n14688) );
  XNOR U16478 ( .A(n14700), .B(n14699), .Z(n14702) );
  AND U16479 ( .A(a[286]), .B(b[0]), .Z(n14652) );
  XNOR U16480 ( .A(n14652), .B(n4071), .Z(n14654) );
  NANDN U16481 ( .A(b[0]), .B(a[285]), .Z(n14653) );
  NAND U16482 ( .A(n14654), .B(n14653), .Z(n14696) );
  XOR U16483 ( .A(a[282]), .B(n42085), .Z(n14692) );
  AND U16484 ( .A(a[278]), .B(b[7]), .Z(n14693) );
  XNOR U16485 ( .A(n14694), .B(n14693), .Z(n14695) );
  XNOR U16486 ( .A(n14696), .B(n14695), .Z(n14701) );
  XOR U16487 ( .A(n14702), .B(n14701), .Z(n14680) );
  NANDN U16488 ( .A(n14657), .B(n14656), .Z(n14661) );
  NANDN U16489 ( .A(n14659), .B(n14658), .Z(n14660) );
  AND U16490 ( .A(n14661), .B(n14660), .Z(n14679) );
  XNOR U16491 ( .A(n14680), .B(n14679), .Z(n14681) );
  NANDN U16492 ( .A(n14663), .B(n14662), .Z(n14667) );
  NAND U16493 ( .A(n14665), .B(n14664), .Z(n14666) );
  NAND U16494 ( .A(n14667), .B(n14666), .Z(n14682) );
  XNOR U16495 ( .A(n14681), .B(n14682), .Z(n14673) );
  XNOR U16496 ( .A(n14674), .B(n14673), .Z(n14675) );
  XNOR U16497 ( .A(n14676), .B(n14675), .Z(n14705) );
  XNOR U16498 ( .A(sreg[1302]), .B(n14705), .Z(n14707) );
  NANDN U16499 ( .A(sreg[1301]), .B(n14668), .Z(n14672) );
  NAND U16500 ( .A(n14670), .B(n14669), .Z(n14671) );
  NAND U16501 ( .A(n14672), .B(n14671), .Z(n14706) );
  XNOR U16502 ( .A(n14707), .B(n14706), .Z(c[1302]) );
  NANDN U16503 ( .A(n14674), .B(n14673), .Z(n14678) );
  NANDN U16504 ( .A(n14676), .B(n14675), .Z(n14677) );
  AND U16505 ( .A(n14678), .B(n14677), .Z(n14713) );
  NANDN U16506 ( .A(n14680), .B(n14679), .Z(n14684) );
  NANDN U16507 ( .A(n14682), .B(n14681), .Z(n14683) );
  AND U16508 ( .A(n14684), .B(n14683), .Z(n14711) );
  NAND U16509 ( .A(n42143), .B(n14685), .Z(n14687) );
  XNOR U16510 ( .A(a[281]), .B(n4112), .Z(n14722) );
  NAND U16511 ( .A(n42144), .B(n14722), .Z(n14686) );
  AND U16512 ( .A(n14687), .B(n14686), .Z(n14737) );
  XOR U16513 ( .A(a[285]), .B(n42012), .Z(n14725) );
  XNOR U16514 ( .A(n14737), .B(n14736), .Z(n14739) );
  AND U16515 ( .A(a[287]), .B(b[0]), .Z(n14689) );
  XNOR U16516 ( .A(n14689), .B(n4071), .Z(n14691) );
  NANDN U16517 ( .A(b[0]), .B(a[286]), .Z(n14690) );
  NAND U16518 ( .A(n14691), .B(n14690), .Z(n14733) );
  XOR U16519 ( .A(a[283]), .B(n42085), .Z(n14729) );
  AND U16520 ( .A(a[279]), .B(b[7]), .Z(n14730) );
  XNOR U16521 ( .A(n14731), .B(n14730), .Z(n14732) );
  XNOR U16522 ( .A(n14733), .B(n14732), .Z(n14738) );
  XOR U16523 ( .A(n14739), .B(n14738), .Z(n14717) );
  NANDN U16524 ( .A(n14694), .B(n14693), .Z(n14698) );
  NANDN U16525 ( .A(n14696), .B(n14695), .Z(n14697) );
  AND U16526 ( .A(n14698), .B(n14697), .Z(n14716) );
  XNOR U16527 ( .A(n14717), .B(n14716), .Z(n14718) );
  NANDN U16528 ( .A(n14700), .B(n14699), .Z(n14704) );
  NAND U16529 ( .A(n14702), .B(n14701), .Z(n14703) );
  NAND U16530 ( .A(n14704), .B(n14703), .Z(n14719) );
  XNOR U16531 ( .A(n14718), .B(n14719), .Z(n14710) );
  XNOR U16532 ( .A(n14711), .B(n14710), .Z(n14712) );
  XNOR U16533 ( .A(n14713), .B(n14712), .Z(n14742) );
  XNOR U16534 ( .A(sreg[1303]), .B(n14742), .Z(n14744) );
  NANDN U16535 ( .A(sreg[1302]), .B(n14705), .Z(n14709) );
  NAND U16536 ( .A(n14707), .B(n14706), .Z(n14708) );
  NAND U16537 ( .A(n14709), .B(n14708), .Z(n14743) );
  XNOR U16538 ( .A(n14744), .B(n14743), .Z(c[1303]) );
  NANDN U16539 ( .A(n14711), .B(n14710), .Z(n14715) );
  NANDN U16540 ( .A(n14713), .B(n14712), .Z(n14714) );
  AND U16541 ( .A(n14715), .B(n14714), .Z(n14750) );
  NANDN U16542 ( .A(n14717), .B(n14716), .Z(n14721) );
  NANDN U16543 ( .A(n14719), .B(n14718), .Z(n14720) );
  AND U16544 ( .A(n14721), .B(n14720), .Z(n14748) );
  NAND U16545 ( .A(n42143), .B(n14722), .Z(n14724) );
  XNOR U16546 ( .A(a[282]), .B(n4112), .Z(n14759) );
  NAND U16547 ( .A(n42144), .B(n14759), .Z(n14723) );
  AND U16548 ( .A(n14724), .B(n14723), .Z(n14774) );
  XOR U16549 ( .A(a[286]), .B(n42012), .Z(n14762) );
  XNOR U16550 ( .A(n14774), .B(n14773), .Z(n14776) );
  AND U16551 ( .A(a[288]), .B(b[0]), .Z(n14726) );
  XNOR U16552 ( .A(n14726), .B(n4071), .Z(n14728) );
  NANDN U16553 ( .A(b[0]), .B(a[287]), .Z(n14727) );
  NAND U16554 ( .A(n14728), .B(n14727), .Z(n14770) );
  XOR U16555 ( .A(a[284]), .B(n42085), .Z(n14766) );
  AND U16556 ( .A(a[280]), .B(b[7]), .Z(n14767) );
  XNOR U16557 ( .A(n14768), .B(n14767), .Z(n14769) );
  XNOR U16558 ( .A(n14770), .B(n14769), .Z(n14775) );
  XOR U16559 ( .A(n14776), .B(n14775), .Z(n14754) );
  NANDN U16560 ( .A(n14731), .B(n14730), .Z(n14735) );
  NANDN U16561 ( .A(n14733), .B(n14732), .Z(n14734) );
  AND U16562 ( .A(n14735), .B(n14734), .Z(n14753) );
  XNOR U16563 ( .A(n14754), .B(n14753), .Z(n14755) );
  NANDN U16564 ( .A(n14737), .B(n14736), .Z(n14741) );
  NAND U16565 ( .A(n14739), .B(n14738), .Z(n14740) );
  NAND U16566 ( .A(n14741), .B(n14740), .Z(n14756) );
  XNOR U16567 ( .A(n14755), .B(n14756), .Z(n14747) );
  XNOR U16568 ( .A(n14748), .B(n14747), .Z(n14749) );
  XNOR U16569 ( .A(n14750), .B(n14749), .Z(n14779) );
  XNOR U16570 ( .A(sreg[1304]), .B(n14779), .Z(n14781) );
  NANDN U16571 ( .A(sreg[1303]), .B(n14742), .Z(n14746) );
  NAND U16572 ( .A(n14744), .B(n14743), .Z(n14745) );
  NAND U16573 ( .A(n14746), .B(n14745), .Z(n14780) );
  XNOR U16574 ( .A(n14781), .B(n14780), .Z(c[1304]) );
  NANDN U16575 ( .A(n14748), .B(n14747), .Z(n14752) );
  NANDN U16576 ( .A(n14750), .B(n14749), .Z(n14751) );
  AND U16577 ( .A(n14752), .B(n14751), .Z(n14787) );
  NANDN U16578 ( .A(n14754), .B(n14753), .Z(n14758) );
  NANDN U16579 ( .A(n14756), .B(n14755), .Z(n14757) );
  AND U16580 ( .A(n14758), .B(n14757), .Z(n14785) );
  NAND U16581 ( .A(n42143), .B(n14759), .Z(n14761) );
  XNOR U16582 ( .A(a[283]), .B(n4112), .Z(n14796) );
  NAND U16583 ( .A(n42144), .B(n14796), .Z(n14760) );
  AND U16584 ( .A(n14761), .B(n14760), .Z(n14811) );
  XOR U16585 ( .A(a[287]), .B(n42012), .Z(n14799) );
  XNOR U16586 ( .A(n14811), .B(n14810), .Z(n14813) );
  AND U16587 ( .A(a[289]), .B(b[0]), .Z(n14763) );
  XNOR U16588 ( .A(n14763), .B(n4071), .Z(n14765) );
  NANDN U16589 ( .A(b[0]), .B(a[288]), .Z(n14764) );
  NAND U16590 ( .A(n14765), .B(n14764), .Z(n14807) );
  XOR U16591 ( .A(a[285]), .B(n42085), .Z(n14800) );
  AND U16592 ( .A(a[281]), .B(b[7]), .Z(n14804) );
  XNOR U16593 ( .A(n14805), .B(n14804), .Z(n14806) );
  XNOR U16594 ( .A(n14807), .B(n14806), .Z(n14812) );
  XOR U16595 ( .A(n14813), .B(n14812), .Z(n14791) );
  NANDN U16596 ( .A(n14768), .B(n14767), .Z(n14772) );
  NANDN U16597 ( .A(n14770), .B(n14769), .Z(n14771) );
  AND U16598 ( .A(n14772), .B(n14771), .Z(n14790) );
  XNOR U16599 ( .A(n14791), .B(n14790), .Z(n14792) );
  NANDN U16600 ( .A(n14774), .B(n14773), .Z(n14778) );
  NAND U16601 ( .A(n14776), .B(n14775), .Z(n14777) );
  NAND U16602 ( .A(n14778), .B(n14777), .Z(n14793) );
  XNOR U16603 ( .A(n14792), .B(n14793), .Z(n14784) );
  XNOR U16604 ( .A(n14785), .B(n14784), .Z(n14786) );
  XNOR U16605 ( .A(n14787), .B(n14786), .Z(n14816) );
  XNOR U16606 ( .A(sreg[1305]), .B(n14816), .Z(n14818) );
  NANDN U16607 ( .A(sreg[1304]), .B(n14779), .Z(n14783) );
  NAND U16608 ( .A(n14781), .B(n14780), .Z(n14782) );
  NAND U16609 ( .A(n14783), .B(n14782), .Z(n14817) );
  XNOR U16610 ( .A(n14818), .B(n14817), .Z(c[1305]) );
  NANDN U16611 ( .A(n14785), .B(n14784), .Z(n14789) );
  NANDN U16612 ( .A(n14787), .B(n14786), .Z(n14788) );
  AND U16613 ( .A(n14789), .B(n14788), .Z(n14824) );
  NANDN U16614 ( .A(n14791), .B(n14790), .Z(n14795) );
  NANDN U16615 ( .A(n14793), .B(n14792), .Z(n14794) );
  AND U16616 ( .A(n14795), .B(n14794), .Z(n14822) );
  NAND U16617 ( .A(n42143), .B(n14796), .Z(n14798) );
  XNOR U16618 ( .A(a[284]), .B(n4112), .Z(n14833) );
  NAND U16619 ( .A(n42144), .B(n14833), .Z(n14797) );
  AND U16620 ( .A(n14798), .B(n14797), .Z(n14848) );
  XOR U16621 ( .A(a[288]), .B(n42012), .Z(n14836) );
  XNOR U16622 ( .A(n14848), .B(n14847), .Z(n14850) );
  XOR U16623 ( .A(a[286]), .B(n42085), .Z(n14837) );
  AND U16624 ( .A(a[282]), .B(b[7]), .Z(n14841) );
  XNOR U16625 ( .A(n14842), .B(n14841), .Z(n14843) );
  AND U16626 ( .A(a[290]), .B(b[0]), .Z(n14801) );
  XNOR U16627 ( .A(n14801), .B(n4071), .Z(n14803) );
  NANDN U16628 ( .A(b[0]), .B(a[289]), .Z(n14802) );
  NAND U16629 ( .A(n14803), .B(n14802), .Z(n14844) );
  XNOR U16630 ( .A(n14843), .B(n14844), .Z(n14849) );
  XOR U16631 ( .A(n14850), .B(n14849), .Z(n14828) );
  NANDN U16632 ( .A(n14805), .B(n14804), .Z(n14809) );
  NANDN U16633 ( .A(n14807), .B(n14806), .Z(n14808) );
  AND U16634 ( .A(n14809), .B(n14808), .Z(n14827) );
  XNOR U16635 ( .A(n14828), .B(n14827), .Z(n14829) );
  NANDN U16636 ( .A(n14811), .B(n14810), .Z(n14815) );
  NAND U16637 ( .A(n14813), .B(n14812), .Z(n14814) );
  NAND U16638 ( .A(n14815), .B(n14814), .Z(n14830) );
  XNOR U16639 ( .A(n14829), .B(n14830), .Z(n14821) );
  XNOR U16640 ( .A(n14822), .B(n14821), .Z(n14823) );
  XNOR U16641 ( .A(n14824), .B(n14823), .Z(n14853) );
  XNOR U16642 ( .A(sreg[1306]), .B(n14853), .Z(n14855) );
  NANDN U16643 ( .A(sreg[1305]), .B(n14816), .Z(n14820) );
  NAND U16644 ( .A(n14818), .B(n14817), .Z(n14819) );
  NAND U16645 ( .A(n14820), .B(n14819), .Z(n14854) );
  XNOR U16646 ( .A(n14855), .B(n14854), .Z(c[1306]) );
  NANDN U16647 ( .A(n14822), .B(n14821), .Z(n14826) );
  NANDN U16648 ( .A(n14824), .B(n14823), .Z(n14825) );
  AND U16649 ( .A(n14826), .B(n14825), .Z(n14861) );
  NANDN U16650 ( .A(n14828), .B(n14827), .Z(n14832) );
  NANDN U16651 ( .A(n14830), .B(n14829), .Z(n14831) );
  AND U16652 ( .A(n14832), .B(n14831), .Z(n14859) );
  NAND U16653 ( .A(n42143), .B(n14833), .Z(n14835) );
  XNOR U16654 ( .A(a[285]), .B(n4112), .Z(n14870) );
  NAND U16655 ( .A(n42144), .B(n14870), .Z(n14834) );
  AND U16656 ( .A(n14835), .B(n14834), .Z(n14885) );
  XOR U16657 ( .A(a[289]), .B(n42012), .Z(n14873) );
  XNOR U16658 ( .A(n14885), .B(n14884), .Z(n14887) );
  XOR U16659 ( .A(a[287]), .B(n42085), .Z(n14877) );
  AND U16660 ( .A(a[283]), .B(b[7]), .Z(n14878) );
  XNOR U16661 ( .A(n14879), .B(n14878), .Z(n14880) );
  AND U16662 ( .A(a[291]), .B(b[0]), .Z(n14838) );
  XNOR U16663 ( .A(n14838), .B(n4071), .Z(n14840) );
  NANDN U16664 ( .A(b[0]), .B(a[290]), .Z(n14839) );
  NAND U16665 ( .A(n14840), .B(n14839), .Z(n14881) );
  XNOR U16666 ( .A(n14880), .B(n14881), .Z(n14886) );
  XOR U16667 ( .A(n14887), .B(n14886), .Z(n14865) );
  NANDN U16668 ( .A(n14842), .B(n14841), .Z(n14846) );
  NANDN U16669 ( .A(n14844), .B(n14843), .Z(n14845) );
  AND U16670 ( .A(n14846), .B(n14845), .Z(n14864) );
  XNOR U16671 ( .A(n14865), .B(n14864), .Z(n14866) );
  NANDN U16672 ( .A(n14848), .B(n14847), .Z(n14852) );
  NAND U16673 ( .A(n14850), .B(n14849), .Z(n14851) );
  NAND U16674 ( .A(n14852), .B(n14851), .Z(n14867) );
  XNOR U16675 ( .A(n14866), .B(n14867), .Z(n14858) );
  XNOR U16676 ( .A(n14859), .B(n14858), .Z(n14860) );
  XNOR U16677 ( .A(n14861), .B(n14860), .Z(n14890) );
  XNOR U16678 ( .A(sreg[1307]), .B(n14890), .Z(n14892) );
  NANDN U16679 ( .A(sreg[1306]), .B(n14853), .Z(n14857) );
  NAND U16680 ( .A(n14855), .B(n14854), .Z(n14856) );
  NAND U16681 ( .A(n14857), .B(n14856), .Z(n14891) );
  XNOR U16682 ( .A(n14892), .B(n14891), .Z(c[1307]) );
  NANDN U16683 ( .A(n14859), .B(n14858), .Z(n14863) );
  NANDN U16684 ( .A(n14861), .B(n14860), .Z(n14862) );
  AND U16685 ( .A(n14863), .B(n14862), .Z(n14898) );
  NANDN U16686 ( .A(n14865), .B(n14864), .Z(n14869) );
  NANDN U16687 ( .A(n14867), .B(n14866), .Z(n14868) );
  AND U16688 ( .A(n14869), .B(n14868), .Z(n14896) );
  NAND U16689 ( .A(n42143), .B(n14870), .Z(n14872) );
  XNOR U16690 ( .A(a[286]), .B(n4112), .Z(n14907) );
  NAND U16691 ( .A(n42144), .B(n14907), .Z(n14871) );
  AND U16692 ( .A(n14872), .B(n14871), .Z(n14922) );
  XOR U16693 ( .A(a[290]), .B(n42012), .Z(n14910) );
  XNOR U16694 ( .A(n14922), .B(n14921), .Z(n14924) );
  AND U16695 ( .A(a[292]), .B(b[0]), .Z(n14874) );
  XNOR U16696 ( .A(n14874), .B(n4071), .Z(n14876) );
  NANDN U16697 ( .A(b[0]), .B(a[291]), .Z(n14875) );
  NAND U16698 ( .A(n14876), .B(n14875), .Z(n14918) );
  XOR U16699 ( .A(a[288]), .B(n42085), .Z(n14914) );
  AND U16700 ( .A(a[284]), .B(b[7]), .Z(n14915) );
  XNOR U16701 ( .A(n14916), .B(n14915), .Z(n14917) );
  XNOR U16702 ( .A(n14918), .B(n14917), .Z(n14923) );
  XOR U16703 ( .A(n14924), .B(n14923), .Z(n14902) );
  NANDN U16704 ( .A(n14879), .B(n14878), .Z(n14883) );
  NANDN U16705 ( .A(n14881), .B(n14880), .Z(n14882) );
  AND U16706 ( .A(n14883), .B(n14882), .Z(n14901) );
  XNOR U16707 ( .A(n14902), .B(n14901), .Z(n14903) );
  NANDN U16708 ( .A(n14885), .B(n14884), .Z(n14889) );
  NAND U16709 ( .A(n14887), .B(n14886), .Z(n14888) );
  NAND U16710 ( .A(n14889), .B(n14888), .Z(n14904) );
  XNOR U16711 ( .A(n14903), .B(n14904), .Z(n14895) );
  XNOR U16712 ( .A(n14896), .B(n14895), .Z(n14897) );
  XNOR U16713 ( .A(n14898), .B(n14897), .Z(n14927) );
  XNOR U16714 ( .A(sreg[1308]), .B(n14927), .Z(n14929) );
  NANDN U16715 ( .A(sreg[1307]), .B(n14890), .Z(n14894) );
  NAND U16716 ( .A(n14892), .B(n14891), .Z(n14893) );
  NAND U16717 ( .A(n14894), .B(n14893), .Z(n14928) );
  XNOR U16718 ( .A(n14929), .B(n14928), .Z(c[1308]) );
  NANDN U16719 ( .A(n14896), .B(n14895), .Z(n14900) );
  NANDN U16720 ( .A(n14898), .B(n14897), .Z(n14899) );
  AND U16721 ( .A(n14900), .B(n14899), .Z(n14935) );
  NANDN U16722 ( .A(n14902), .B(n14901), .Z(n14906) );
  NANDN U16723 ( .A(n14904), .B(n14903), .Z(n14905) );
  AND U16724 ( .A(n14906), .B(n14905), .Z(n14933) );
  NAND U16725 ( .A(n42143), .B(n14907), .Z(n14909) );
  XNOR U16726 ( .A(a[287]), .B(n4112), .Z(n14944) );
  NAND U16727 ( .A(n42144), .B(n14944), .Z(n14908) );
  AND U16728 ( .A(n14909), .B(n14908), .Z(n14959) );
  XOR U16729 ( .A(a[291]), .B(n42012), .Z(n14947) );
  XNOR U16730 ( .A(n14959), .B(n14958), .Z(n14961) );
  AND U16731 ( .A(a[293]), .B(b[0]), .Z(n14911) );
  XNOR U16732 ( .A(n14911), .B(n4071), .Z(n14913) );
  NANDN U16733 ( .A(b[0]), .B(a[292]), .Z(n14912) );
  NAND U16734 ( .A(n14913), .B(n14912), .Z(n14955) );
  XOR U16735 ( .A(a[289]), .B(n42085), .Z(n14951) );
  AND U16736 ( .A(a[285]), .B(b[7]), .Z(n14952) );
  XNOR U16737 ( .A(n14953), .B(n14952), .Z(n14954) );
  XNOR U16738 ( .A(n14955), .B(n14954), .Z(n14960) );
  XOR U16739 ( .A(n14961), .B(n14960), .Z(n14939) );
  NANDN U16740 ( .A(n14916), .B(n14915), .Z(n14920) );
  NANDN U16741 ( .A(n14918), .B(n14917), .Z(n14919) );
  AND U16742 ( .A(n14920), .B(n14919), .Z(n14938) );
  XNOR U16743 ( .A(n14939), .B(n14938), .Z(n14940) );
  NANDN U16744 ( .A(n14922), .B(n14921), .Z(n14926) );
  NAND U16745 ( .A(n14924), .B(n14923), .Z(n14925) );
  NAND U16746 ( .A(n14926), .B(n14925), .Z(n14941) );
  XNOR U16747 ( .A(n14940), .B(n14941), .Z(n14932) );
  XNOR U16748 ( .A(n14933), .B(n14932), .Z(n14934) );
  XNOR U16749 ( .A(n14935), .B(n14934), .Z(n14964) );
  XNOR U16750 ( .A(sreg[1309]), .B(n14964), .Z(n14966) );
  NANDN U16751 ( .A(sreg[1308]), .B(n14927), .Z(n14931) );
  NAND U16752 ( .A(n14929), .B(n14928), .Z(n14930) );
  NAND U16753 ( .A(n14931), .B(n14930), .Z(n14965) );
  XNOR U16754 ( .A(n14966), .B(n14965), .Z(c[1309]) );
  NANDN U16755 ( .A(n14933), .B(n14932), .Z(n14937) );
  NANDN U16756 ( .A(n14935), .B(n14934), .Z(n14936) );
  AND U16757 ( .A(n14937), .B(n14936), .Z(n14972) );
  NANDN U16758 ( .A(n14939), .B(n14938), .Z(n14943) );
  NANDN U16759 ( .A(n14941), .B(n14940), .Z(n14942) );
  AND U16760 ( .A(n14943), .B(n14942), .Z(n14970) );
  NAND U16761 ( .A(n42143), .B(n14944), .Z(n14946) );
  XNOR U16762 ( .A(a[288]), .B(n4113), .Z(n14981) );
  NAND U16763 ( .A(n42144), .B(n14981), .Z(n14945) );
  AND U16764 ( .A(n14946), .B(n14945), .Z(n14996) );
  XOR U16765 ( .A(a[292]), .B(n42012), .Z(n14984) );
  XNOR U16766 ( .A(n14996), .B(n14995), .Z(n14998) );
  AND U16767 ( .A(a[294]), .B(b[0]), .Z(n14948) );
  XNOR U16768 ( .A(n14948), .B(n4071), .Z(n14950) );
  NANDN U16769 ( .A(b[0]), .B(a[293]), .Z(n14949) );
  NAND U16770 ( .A(n14950), .B(n14949), .Z(n14992) );
  XOR U16771 ( .A(a[290]), .B(n42085), .Z(n14985) );
  AND U16772 ( .A(a[286]), .B(b[7]), .Z(n14989) );
  XNOR U16773 ( .A(n14990), .B(n14989), .Z(n14991) );
  XNOR U16774 ( .A(n14992), .B(n14991), .Z(n14997) );
  XOR U16775 ( .A(n14998), .B(n14997), .Z(n14976) );
  NANDN U16776 ( .A(n14953), .B(n14952), .Z(n14957) );
  NANDN U16777 ( .A(n14955), .B(n14954), .Z(n14956) );
  AND U16778 ( .A(n14957), .B(n14956), .Z(n14975) );
  XNOR U16779 ( .A(n14976), .B(n14975), .Z(n14977) );
  NANDN U16780 ( .A(n14959), .B(n14958), .Z(n14963) );
  NAND U16781 ( .A(n14961), .B(n14960), .Z(n14962) );
  NAND U16782 ( .A(n14963), .B(n14962), .Z(n14978) );
  XNOR U16783 ( .A(n14977), .B(n14978), .Z(n14969) );
  XNOR U16784 ( .A(n14970), .B(n14969), .Z(n14971) );
  XNOR U16785 ( .A(n14972), .B(n14971), .Z(n15001) );
  XNOR U16786 ( .A(sreg[1310]), .B(n15001), .Z(n15003) );
  NANDN U16787 ( .A(sreg[1309]), .B(n14964), .Z(n14968) );
  NAND U16788 ( .A(n14966), .B(n14965), .Z(n14967) );
  NAND U16789 ( .A(n14968), .B(n14967), .Z(n15002) );
  XNOR U16790 ( .A(n15003), .B(n15002), .Z(c[1310]) );
  NANDN U16791 ( .A(n14970), .B(n14969), .Z(n14974) );
  NANDN U16792 ( .A(n14972), .B(n14971), .Z(n14973) );
  AND U16793 ( .A(n14974), .B(n14973), .Z(n15009) );
  NANDN U16794 ( .A(n14976), .B(n14975), .Z(n14980) );
  NANDN U16795 ( .A(n14978), .B(n14977), .Z(n14979) );
  AND U16796 ( .A(n14980), .B(n14979), .Z(n15007) );
  NAND U16797 ( .A(n42143), .B(n14981), .Z(n14983) );
  XNOR U16798 ( .A(a[289]), .B(n4113), .Z(n15018) );
  NAND U16799 ( .A(n42144), .B(n15018), .Z(n14982) );
  AND U16800 ( .A(n14983), .B(n14982), .Z(n15033) );
  XOR U16801 ( .A(a[293]), .B(n42012), .Z(n15021) );
  XNOR U16802 ( .A(n15033), .B(n15032), .Z(n15035) );
  XOR U16803 ( .A(a[291]), .B(n42085), .Z(n15025) );
  AND U16804 ( .A(a[287]), .B(b[7]), .Z(n15026) );
  XNOR U16805 ( .A(n15027), .B(n15026), .Z(n15028) );
  AND U16806 ( .A(a[295]), .B(b[0]), .Z(n14986) );
  XNOR U16807 ( .A(n14986), .B(n4071), .Z(n14988) );
  NANDN U16808 ( .A(b[0]), .B(a[294]), .Z(n14987) );
  NAND U16809 ( .A(n14988), .B(n14987), .Z(n15029) );
  XNOR U16810 ( .A(n15028), .B(n15029), .Z(n15034) );
  XOR U16811 ( .A(n15035), .B(n15034), .Z(n15013) );
  NANDN U16812 ( .A(n14990), .B(n14989), .Z(n14994) );
  NANDN U16813 ( .A(n14992), .B(n14991), .Z(n14993) );
  AND U16814 ( .A(n14994), .B(n14993), .Z(n15012) );
  XNOR U16815 ( .A(n15013), .B(n15012), .Z(n15014) );
  NANDN U16816 ( .A(n14996), .B(n14995), .Z(n15000) );
  NAND U16817 ( .A(n14998), .B(n14997), .Z(n14999) );
  NAND U16818 ( .A(n15000), .B(n14999), .Z(n15015) );
  XNOR U16819 ( .A(n15014), .B(n15015), .Z(n15006) );
  XNOR U16820 ( .A(n15007), .B(n15006), .Z(n15008) );
  XNOR U16821 ( .A(n15009), .B(n15008), .Z(n15038) );
  XNOR U16822 ( .A(sreg[1311]), .B(n15038), .Z(n15040) );
  NANDN U16823 ( .A(sreg[1310]), .B(n15001), .Z(n15005) );
  NAND U16824 ( .A(n15003), .B(n15002), .Z(n15004) );
  NAND U16825 ( .A(n15005), .B(n15004), .Z(n15039) );
  XNOR U16826 ( .A(n15040), .B(n15039), .Z(c[1311]) );
  NANDN U16827 ( .A(n15007), .B(n15006), .Z(n15011) );
  NANDN U16828 ( .A(n15009), .B(n15008), .Z(n15010) );
  AND U16829 ( .A(n15011), .B(n15010), .Z(n15046) );
  NANDN U16830 ( .A(n15013), .B(n15012), .Z(n15017) );
  NANDN U16831 ( .A(n15015), .B(n15014), .Z(n15016) );
  AND U16832 ( .A(n15017), .B(n15016), .Z(n15044) );
  NAND U16833 ( .A(n42143), .B(n15018), .Z(n15020) );
  XNOR U16834 ( .A(a[290]), .B(n4113), .Z(n15055) );
  NAND U16835 ( .A(n42144), .B(n15055), .Z(n15019) );
  AND U16836 ( .A(n15020), .B(n15019), .Z(n15070) );
  XOR U16837 ( .A(a[294]), .B(n42012), .Z(n15058) );
  XNOR U16838 ( .A(n15070), .B(n15069), .Z(n15072) );
  AND U16839 ( .A(a[296]), .B(b[0]), .Z(n15022) );
  XNOR U16840 ( .A(n15022), .B(n4071), .Z(n15024) );
  NANDN U16841 ( .A(b[0]), .B(a[295]), .Z(n15023) );
  NAND U16842 ( .A(n15024), .B(n15023), .Z(n15066) );
  XOR U16843 ( .A(a[292]), .B(n42085), .Z(n15062) );
  AND U16844 ( .A(a[288]), .B(b[7]), .Z(n15063) );
  XNOR U16845 ( .A(n15064), .B(n15063), .Z(n15065) );
  XNOR U16846 ( .A(n15066), .B(n15065), .Z(n15071) );
  XOR U16847 ( .A(n15072), .B(n15071), .Z(n15050) );
  NANDN U16848 ( .A(n15027), .B(n15026), .Z(n15031) );
  NANDN U16849 ( .A(n15029), .B(n15028), .Z(n15030) );
  AND U16850 ( .A(n15031), .B(n15030), .Z(n15049) );
  XNOR U16851 ( .A(n15050), .B(n15049), .Z(n15051) );
  NANDN U16852 ( .A(n15033), .B(n15032), .Z(n15037) );
  NAND U16853 ( .A(n15035), .B(n15034), .Z(n15036) );
  NAND U16854 ( .A(n15037), .B(n15036), .Z(n15052) );
  XNOR U16855 ( .A(n15051), .B(n15052), .Z(n15043) );
  XNOR U16856 ( .A(n15044), .B(n15043), .Z(n15045) );
  XNOR U16857 ( .A(n15046), .B(n15045), .Z(n15075) );
  XNOR U16858 ( .A(sreg[1312]), .B(n15075), .Z(n15077) );
  NANDN U16859 ( .A(sreg[1311]), .B(n15038), .Z(n15042) );
  NAND U16860 ( .A(n15040), .B(n15039), .Z(n15041) );
  NAND U16861 ( .A(n15042), .B(n15041), .Z(n15076) );
  XNOR U16862 ( .A(n15077), .B(n15076), .Z(c[1312]) );
  NANDN U16863 ( .A(n15044), .B(n15043), .Z(n15048) );
  NANDN U16864 ( .A(n15046), .B(n15045), .Z(n15047) );
  AND U16865 ( .A(n15048), .B(n15047), .Z(n15083) );
  NANDN U16866 ( .A(n15050), .B(n15049), .Z(n15054) );
  NANDN U16867 ( .A(n15052), .B(n15051), .Z(n15053) );
  AND U16868 ( .A(n15054), .B(n15053), .Z(n15081) );
  NAND U16869 ( .A(n42143), .B(n15055), .Z(n15057) );
  XNOR U16870 ( .A(a[291]), .B(n4113), .Z(n15092) );
  NAND U16871 ( .A(n42144), .B(n15092), .Z(n15056) );
  AND U16872 ( .A(n15057), .B(n15056), .Z(n15107) );
  XOR U16873 ( .A(a[295]), .B(n42012), .Z(n15095) );
  XNOR U16874 ( .A(n15107), .B(n15106), .Z(n15109) );
  AND U16875 ( .A(a[297]), .B(b[0]), .Z(n15059) );
  XNOR U16876 ( .A(n15059), .B(n4071), .Z(n15061) );
  NANDN U16877 ( .A(b[0]), .B(a[296]), .Z(n15060) );
  NAND U16878 ( .A(n15061), .B(n15060), .Z(n15103) );
  XOR U16879 ( .A(a[293]), .B(n42085), .Z(n15099) );
  AND U16880 ( .A(a[289]), .B(b[7]), .Z(n15100) );
  XNOR U16881 ( .A(n15101), .B(n15100), .Z(n15102) );
  XNOR U16882 ( .A(n15103), .B(n15102), .Z(n15108) );
  XOR U16883 ( .A(n15109), .B(n15108), .Z(n15087) );
  NANDN U16884 ( .A(n15064), .B(n15063), .Z(n15068) );
  NANDN U16885 ( .A(n15066), .B(n15065), .Z(n15067) );
  AND U16886 ( .A(n15068), .B(n15067), .Z(n15086) );
  XNOR U16887 ( .A(n15087), .B(n15086), .Z(n15088) );
  NANDN U16888 ( .A(n15070), .B(n15069), .Z(n15074) );
  NAND U16889 ( .A(n15072), .B(n15071), .Z(n15073) );
  NAND U16890 ( .A(n15074), .B(n15073), .Z(n15089) );
  XNOR U16891 ( .A(n15088), .B(n15089), .Z(n15080) );
  XNOR U16892 ( .A(n15081), .B(n15080), .Z(n15082) );
  XNOR U16893 ( .A(n15083), .B(n15082), .Z(n15112) );
  XNOR U16894 ( .A(sreg[1313]), .B(n15112), .Z(n15114) );
  NANDN U16895 ( .A(sreg[1312]), .B(n15075), .Z(n15079) );
  NAND U16896 ( .A(n15077), .B(n15076), .Z(n15078) );
  NAND U16897 ( .A(n15079), .B(n15078), .Z(n15113) );
  XNOR U16898 ( .A(n15114), .B(n15113), .Z(c[1313]) );
  NANDN U16899 ( .A(n15081), .B(n15080), .Z(n15085) );
  NANDN U16900 ( .A(n15083), .B(n15082), .Z(n15084) );
  AND U16901 ( .A(n15085), .B(n15084), .Z(n15120) );
  NANDN U16902 ( .A(n15087), .B(n15086), .Z(n15091) );
  NANDN U16903 ( .A(n15089), .B(n15088), .Z(n15090) );
  AND U16904 ( .A(n15091), .B(n15090), .Z(n15118) );
  NAND U16905 ( .A(n42143), .B(n15092), .Z(n15094) );
  XNOR U16906 ( .A(a[292]), .B(n4113), .Z(n15129) );
  NAND U16907 ( .A(n42144), .B(n15129), .Z(n15093) );
  AND U16908 ( .A(n15094), .B(n15093), .Z(n15144) );
  XOR U16909 ( .A(a[296]), .B(n42012), .Z(n15132) );
  XNOR U16910 ( .A(n15144), .B(n15143), .Z(n15146) );
  AND U16911 ( .A(a[298]), .B(b[0]), .Z(n15096) );
  XNOR U16912 ( .A(n15096), .B(n4071), .Z(n15098) );
  NANDN U16913 ( .A(b[0]), .B(a[297]), .Z(n15097) );
  NAND U16914 ( .A(n15098), .B(n15097), .Z(n15140) );
  XOR U16915 ( .A(a[294]), .B(n42085), .Z(n15136) );
  AND U16916 ( .A(a[290]), .B(b[7]), .Z(n15137) );
  XNOR U16917 ( .A(n15138), .B(n15137), .Z(n15139) );
  XNOR U16918 ( .A(n15140), .B(n15139), .Z(n15145) );
  XOR U16919 ( .A(n15146), .B(n15145), .Z(n15124) );
  NANDN U16920 ( .A(n15101), .B(n15100), .Z(n15105) );
  NANDN U16921 ( .A(n15103), .B(n15102), .Z(n15104) );
  AND U16922 ( .A(n15105), .B(n15104), .Z(n15123) );
  XNOR U16923 ( .A(n15124), .B(n15123), .Z(n15125) );
  NANDN U16924 ( .A(n15107), .B(n15106), .Z(n15111) );
  NAND U16925 ( .A(n15109), .B(n15108), .Z(n15110) );
  NAND U16926 ( .A(n15111), .B(n15110), .Z(n15126) );
  XNOR U16927 ( .A(n15125), .B(n15126), .Z(n15117) );
  XNOR U16928 ( .A(n15118), .B(n15117), .Z(n15119) );
  XNOR U16929 ( .A(n15120), .B(n15119), .Z(n15149) );
  XNOR U16930 ( .A(sreg[1314]), .B(n15149), .Z(n15151) );
  NANDN U16931 ( .A(sreg[1313]), .B(n15112), .Z(n15116) );
  NAND U16932 ( .A(n15114), .B(n15113), .Z(n15115) );
  NAND U16933 ( .A(n15116), .B(n15115), .Z(n15150) );
  XNOR U16934 ( .A(n15151), .B(n15150), .Z(c[1314]) );
  NANDN U16935 ( .A(n15118), .B(n15117), .Z(n15122) );
  NANDN U16936 ( .A(n15120), .B(n15119), .Z(n15121) );
  AND U16937 ( .A(n15122), .B(n15121), .Z(n15157) );
  NANDN U16938 ( .A(n15124), .B(n15123), .Z(n15128) );
  NANDN U16939 ( .A(n15126), .B(n15125), .Z(n15127) );
  AND U16940 ( .A(n15128), .B(n15127), .Z(n15155) );
  NAND U16941 ( .A(n42143), .B(n15129), .Z(n15131) );
  XNOR U16942 ( .A(a[293]), .B(n4113), .Z(n15166) );
  NAND U16943 ( .A(n42144), .B(n15166), .Z(n15130) );
  AND U16944 ( .A(n15131), .B(n15130), .Z(n15181) );
  XOR U16945 ( .A(a[297]), .B(n42012), .Z(n15169) );
  XNOR U16946 ( .A(n15181), .B(n15180), .Z(n15183) );
  AND U16947 ( .A(a[299]), .B(b[0]), .Z(n15133) );
  XNOR U16948 ( .A(n15133), .B(n4071), .Z(n15135) );
  NANDN U16949 ( .A(b[0]), .B(a[298]), .Z(n15134) );
  NAND U16950 ( .A(n15135), .B(n15134), .Z(n15177) );
  XOR U16951 ( .A(a[295]), .B(n42085), .Z(n15170) );
  AND U16952 ( .A(a[291]), .B(b[7]), .Z(n15174) );
  XNOR U16953 ( .A(n15175), .B(n15174), .Z(n15176) );
  XNOR U16954 ( .A(n15177), .B(n15176), .Z(n15182) );
  XOR U16955 ( .A(n15183), .B(n15182), .Z(n15161) );
  NANDN U16956 ( .A(n15138), .B(n15137), .Z(n15142) );
  NANDN U16957 ( .A(n15140), .B(n15139), .Z(n15141) );
  AND U16958 ( .A(n15142), .B(n15141), .Z(n15160) );
  XNOR U16959 ( .A(n15161), .B(n15160), .Z(n15162) );
  NANDN U16960 ( .A(n15144), .B(n15143), .Z(n15148) );
  NAND U16961 ( .A(n15146), .B(n15145), .Z(n15147) );
  NAND U16962 ( .A(n15148), .B(n15147), .Z(n15163) );
  XNOR U16963 ( .A(n15162), .B(n15163), .Z(n15154) );
  XNOR U16964 ( .A(n15155), .B(n15154), .Z(n15156) );
  XNOR U16965 ( .A(n15157), .B(n15156), .Z(n15186) );
  XNOR U16966 ( .A(sreg[1315]), .B(n15186), .Z(n15188) );
  NANDN U16967 ( .A(sreg[1314]), .B(n15149), .Z(n15153) );
  NAND U16968 ( .A(n15151), .B(n15150), .Z(n15152) );
  NAND U16969 ( .A(n15153), .B(n15152), .Z(n15187) );
  XNOR U16970 ( .A(n15188), .B(n15187), .Z(c[1315]) );
  NANDN U16971 ( .A(n15155), .B(n15154), .Z(n15159) );
  NANDN U16972 ( .A(n15157), .B(n15156), .Z(n15158) );
  AND U16973 ( .A(n15159), .B(n15158), .Z(n15194) );
  NANDN U16974 ( .A(n15161), .B(n15160), .Z(n15165) );
  NANDN U16975 ( .A(n15163), .B(n15162), .Z(n15164) );
  AND U16976 ( .A(n15165), .B(n15164), .Z(n15192) );
  NAND U16977 ( .A(n42143), .B(n15166), .Z(n15168) );
  XNOR U16978 ( .A(a[294]), .B(n4113), .Z(n15203) );
  NAND U16979 ( .A(n42144), .B(n15203), .Z(n15167) );
  AND U16980 ( .A(n15168), .B(n15167), .Z(n15218) );
  XOR U16981 ( .A(a[298]), .B(n42012), .Z(n15206) );
  XNOR U16982 ( .A(n15218), .B(n15217), .Z(n15220) );
  XOR U16983 ( .A(a[296]), .B(n42085), .Z(n15210) );
  AND U16984 ( .A(a[292]), .B(b[7]), .Z(n15211) );
  XNOR U16985 ( .A(n15212), .B(n15211), .Z(n15213) );
  AND U16986 ( .A(a[300]), .B(b[0]), .Z(n15171) );
  XNOR U16987 ( .A(n15171), .B(n4071), .Z(n15173) );
  NANDN U16988 ( .A(b[0]), .B(a[299]), .Z(n15172) );
  NAND U16989 ( .A(n15173), .B(n15172), .Z(n15214) );
  XNOR U16990 ( .A(n15213), .B(n15214), .Z(n15219) );
  XOR U16991 ( .A(n15220), .B(n15219), .Z(n15198) );
  NANDN U16992 ( .A(n15175), .B(n15174), .Z(n15179) );
  NANDN U16993 ( .A(n15177), .B(n15176), .Z(n15178) );
  AND U16994 ( .A(n15179), .B(n15178), .Z(n15197) );
  XNOR U16995 ( .A(n15198), .B(n15197), .Z(n15199) );
  NANDN U16996 ( .A(n15181), .B(n15180), .Z(n15185) );
  NAND U16997 ( .A(n15183), .B(n15182), .Z(n15184) );
  NAND U16998 ( .A(n15185), .B(n15184), .Z(n15200) );
  XNOR U16999 ( .A(n15199), .B(n15200), .Z(n15191) );
  XNOR U17000 ( .A(n15192), .B(n15191), .Z(n15193) );
  XNOR U17001 ( .A(n15194), .B(n15193), .Z(n15223) );
  XNOR U17002 ( .A(sreg[1316]), .B(n15223), .Z(n15225) );
  NANDN U17003 ( .A(sreg[1315]), .B(n15186), .Z(n15190) );
  NAND U17004 ( .A(n15188), .B(n15187), .Z(n15189) );
  NAND U17005 ( .A(n15190), .B(n15189), .Z(n15224) );
  XNOR U17006 ( .A(n15225), .B(n15224), .Z(c[1316]) );
  NANDN U17007 ( .A(n15192), .B(n15191), .Z(n15196) );
  NANDN U17008 ( .A(n15194), .B(n15193), .Z(n15195) );
  AND U17009 ( .A(n15196), .B(n15195), .Z(n15231) );
  NANDN U17010 ( .A(n15198), .B(n15197), .Z(n15202) );
  NANDN U17011 ( .A(n15200), .B(n15199), .Z(n15201) );
  AND U17012 ( .A(n15202), .B(n15201), .Z(n15229) );
  NAND U17013 ( .A(n42143), .B(n15203), .Z(n15205) );
  XNOR U17014 ( .A(a[295]), .B(n4114), .Z(n15240) );
  NAND U17015 ( .A(n42144), .B(n15240), .Z(n15204) );
  AND U17016 ( .A(n15205), .B(n15204), .Z(n15255) );
  XOR U17017 ( .A(a[299]), .B(n42012), .Z(n15243) );
  XNOR U17018 ( .A(n15255), .B(n15254), .Z(n15257) );
  AND U17019 ( .A(a[301]), .B(b[0]), .Z(n15207) );
  XNOR U17020 ( .A(n15207), .B(n4071), .Z(n15209) );
  NANDN U17021 ( .A(b[0]), .B(a[300]), .Z(n15208) );
  NAND U17022 ( .A(n15209), .B(n15208), .Z(n15251) );
  XOR U17023 ( .A(a[297]), .B(n42085), .Z(n15244) );
  AND U17024 ( .A(a[293]), .B(b[7]), .Z(n15248) );
  XNOR U17025 ( .A(n15249), .B(n15248), .Z(n15250) );
  XNOR U17026 ( .A(n15251), .B(n15250), .Z(n15256) );
  XOR U17027 ( .A(n15257), .B(n15256), .Z(n15235) );
  NANDN U17028 ( .A(n15212), .B(n15211), .Z(n15216) );
  NANDN U17029 ( .A(n15214), .B(n15213), .Z(n15215) );
  AND U17030 ( .A(n15216), .B(n15215), .Z(n15234) );
  XNOR U17031 ( .A(n15235), .B(n15234), .Z(n15236) );
  NANDN U17032 ( .A(n15218), .B(n15217), .Z(n15222) );
  NAND U17033 ( .A(n15220), .B(n15219), .Z(n15221) );
  NAND U17034 ( .A(n15222), .B(n15221), .Z(n15237) );
  XNOR U17035 ( .A(n15236), .B(n15237), .Z(n15228) );
  XNOR U17036 ( .A(n15229), .B(n15228), .Z(n15230) );
  XNOR U17037 ( .A(n15231), .B(n15230), .Z(n15260) );
  XNOR U17038 ( .A(sreg[1317]), .B(n15260), .Z(n15262) );
  NANDN U17039 ( .A(sreg[1316]), .B(n15223), .Z(n15227) );
  NAND U17040 ( .A(n15225), .B(n15224), .Z(n15226) );
  NAND U17041 ( .A(n15227), .B(n15226), .Z(n15261) );
  XNOR U17042 ( .A(n15262), .B(n15261), .Z(c[1317]) );
  NANDN U17043 ( .A(n15229), .B(n15228), .Z(n15233) );
  NANDN U17044 ( .A(n15231), .B(n15230), .Z(n15232) );
  AND U17045 ( .A(n15233), .B(n15232), .Z(n15268) );
  NANDN U17046 ( .A(n15235), .B(n15234), .Z(n15239) );
  NANDN U17047 ( .A(n15237), .B(n15236), .Z(n15238) );
  AND U17048 ( .A(n15239), .B(n15238), .Z(n15266) );
  NAND U17049 ( .A(n42143), .B(n15240), .Z(n15242) );
  XNOR U17050 ( .A(a[296]), .B(n4114), .Z(n15277) );
  NAND U17051 ( .A(n42144), .B(n15277), .Z(n15241) );
  AND U17052 ( .A(n15242), .B(n15241), .Z(n15292) );
  XOR U17053 ( .A(a[300]), .B(n42012), .Z(n15280) );
  XNOR U17054 ( .A(n15292), .B(n15291), .Z(n15294) );
  XOR U17055 ( .A(a[298]), .B(n42085), .Z(n15284) );
  AND U17056 ( .A(a[294]), .B(b[7]), .Z(n15285) );
  XNOR U17057 ( .A(n15286), .B(n15285), .Z(n15287) );
  AND U17058 ( .A(a[302]), .B(b[0]), .Z(n15245) );
  XNOR U17059 ( .A(n15245), .B(n4071), .Z(n15247) );
  NANDN U17060 ( .A(b[0]), .B(a[301]), .Z(n15246) );
  NAND U17061 ( .A(n15247), .B(n15246), .Z(n15288) );
  XNOR U17062 ( .A(n15287), .B(n15288), .Z(n15293) );
  XOR U17063 ( .A(n15294), .B(n15293), .Z(n15272) );
  NANDN U17064 ( .A(n15249), .B(n15248), .Z(n15253) );
  NANDN U17065 ( .A(n15251), .B(n15250), .Z(n15252) );
  AND U17066 ( .A(n15253), .B(n15252), .Z(n15271) );
  XNOR U17067 ( .A(n15272), .B(n15271), .Z(n15273) );
  NANDN U17068 ( .A(n15255), .B(n15254), .Z(n15259) );
  NAND U17069 ( .A(n15257), .B(n15256), .Z(n15258) );
  NAND U17070 ( .A(n15259), .B(n15258), .Z(n15274) );
  XNOR U17071 ( .A(n15273), .B(n15274), .Z(n15265) );
  XNOR U17072 ( .A(n15266), .B(n15265), .Z(n15267) );
  XNOR U17073 ( .A(n15268), .B(n15267), .Z(n15297) );
  XNOR U17074 ( .A(sreg[1318]), .B(n15297), .Z(n15299) );
  NANDN U17075 ( .A(sreg[1317]), .B(n15260), .Z(n15264) );
  NAND U17076 ( .A(n15262), .B(n15261), .Z(n15263) );
  NAND U17077 ( .A(n15264), .B(n15263), .Z(n15298) );
  XNOR U17078 ( .A(n15299), .B(n15298), .Z(c[1318]) );
  NANDN U17079 ( .A(n15266), .B(n15265), .Z(n15270) );
  NANDN U17080 ( .A(n15268), .B(n15267), .Z(n15269) );
  AND U17081 ( .A(n15270), .B(n15269), .Z(n15305) );
  NANDN U17082 ( .A(n15272), .B(n15271), .Z(n15276) );
  NANDN U17083 ( .A(n15274), .B(n15273), .Z(n15275) );
  AND U17084 ( .A(n15276), .B(n15275), .Z(n15303) );
  NAND U17085 ( .A(n42143), .B(n15277), .Z(n15279) );
  XNOR U17086 ( .A(a[297]), .B(n4114), .Z(n15314) );
  NAND U17087 ( .A(n42144), .B(n15314), .Z(n15278) );
  AND U17088 ( .A(n15279), .B(n15278), .Z(n15329) );
  XOR U17089 ( .A(a[301]), .B(n42012), .Z(n15317) );
  XNOR U17090 ( .A(n15329), .B(n15328), .Z(n15331) );
  AND U17091 ( .A(a[303]), .B(b[0]), .Z(n15281) );
  XNOR U17092 ( .A(n15281), .B(n4071), .Z(n15283) );
  NANDN U17093 ( .A(b[0]), .B(a[302]), .Z(n15282) );
  NAND U17094 ( .A(n15283), .B(n15282), .Z(n15325) );
  XOR U17095 ( .A(a[299]), .B(n42085), .Z(n15318) );
  AND U17096 ( .A(a[295]), .B(b[7]), .Z(n15322) );
  XNOR U17097 ( .A(n15323), .B(n15322), .Z(n15324) );
  XNOR U17098 ( .A(n15325), .B(n15324), .Z(n15330) );
  XOR U17099 ( .A(n15331), .B(n15330), .Z(n15309) );
  NANDN U17100 ( .A(n15286), .B(n15285), .Z(n15290) );
  NANDN U17101 ( .A(n15288), .B(n15287), .Z(n15289) );
  AND U17102 ( .A(n15290), .B(n15289), .Z(n15308) );
  XNOR U17103 ( .A(n15309), .B(n15308), .Z(n15310) );
  NANDN U17104 ( .A(n15292), .B(n15291), .Z(n15296) );
  NAND U17105 ( .A(n15294), .B(n15293), .Z(n15295) );
  NAND U17106 ( .A(n15296), .B(n15295), .Z(n15311) );
  XNOR U17107 ( .A(n15310), .B(n15311), .Z(n15302) );
  XNOR U17108 ( .A(n15303), .B(n15302), .Z(n15304) );
  XNOR U17109 ( .A(n15305), .B(n15304), .Z(n15334) );
  XNOR U17110 ( .A(sreg[1319]), .B(n15334), .Z(n15336) );
  NANDN U17111 ( .A(sreg[1318]), .B(n15297), .Z(n15301) );
  NAND U17112 ( .A(n15299), .B(n15298), .Z(n15300) );
  NAND U17113 ( .A(n15301), .B(n15300), .Z(n15335) );
  XNOR U17114 ( .A(n15336), .B(n15335), .Z(c[1319]) );
  NANDN U17115 ( .A(n15303), .B(n15302), .Z(n15307) );
  NANDN U17116 ( .A(n15305), .B(n15304), .Z(n15306) );
  AND U17117 ( .A(n15307), .B(n15306), .Z(n15342) );
  NANDN U17118 ( .A(n15309), .B(n15308), .Z(n15313) );
  NANDN U17119 ( .A(n15311), .B(n15310), .Z(n15312) );
  AND U17120 ( .A(n15313), .B(n15312), .Z(n15340) );
  NAND U17121 ( .A(n42143), .B(n15314), .Z(n15316) );
  XNOR U17122 ( .A(a[298]), .B(n4114), .Z(n15351) );
  NAND U17123 ( .A(n42144), .B(n15351), .Z(n15315) );
  AND U17124 ( .A(n15316), .B(n15315), .Z(n15366) );
  XOR U17125 ( .A(a[302]), .B(n42012), .Z(n15354) );
  XNOR U17126 ( .A(n15366), .B(n15365), .Z(n15368) );
  XOR U17127 ( .A(a[300]), .B(n42085), .Z(n15355) );
  AND U17128 ( .A(a[296]), .B(b[7]), .Z(n15359) );
  XNOR U17129 ( .A(n15360), .B(n15359), .Z(n15361) );
  AND U17130 ( .A(a[304]), .B(b[0]), .Z(n15319) );
  XNOR U17131 ( .A(n15319), .B(n4071), .Z(n15321) );
  NANDN U17132 ( .A(b[0]), .B(a[303]), .Z(n15320) );
  NAND U17133 ( .A(n15321), .B(n15320), .Z(n15362) );
  XNOR U17134 ( .A(n15361), .B(n15362), .Z(n15367) );
  XOR U17135 ( .A(n15368), .B(n15367), .Z(n15346) );
  NANDN U17136 ( .A(n15323), .B(n15322), .Z(n15327) );
  NANDN U17137 ( .A(n15325), .B(n15324), .Z(n15326) );
  AND U17138 ( .A(n15327), .B(n15326), .Z(n15345) );
  XNOR U17139 ( .A(n15346), .B(n15345), .Z(n15347) );
  NANDN U17140 ( .A(n15329), .B(n15328), .Z(n15333) );
  NAND U17141 ( .A(n15331), .B(n15330), .Z(n15332) );
  NAND U17142 ( .A(n15333), .B(n15332), .Z(n15348) );
  XNOR U17143 ( .A(n15347), .B(n15348), .Z(n15339) );
  XNOR U17144 ( .A(n15340), .B(n15339), .Z(n15341) );
  XNOR U17145 ( .A(n15342), .B(n15341), .Z(n15371) );
  XNOR U17146 ( .A(sreg[1320]), .B(n15371), .Z(n15373) );
  NANDN U17147 ( .A(sreg[1319]), .B(n15334), .Z(n15338) );
  NAND U17148 ( .A(n15336), .B(n15335), .Z(n15337) );
  NAND U17149 ( .A(n15338), .B(n15337), .Z(n15372) );
  XNOR U17150 ( .A(n15373), .B(n15372), .Z(c[1320]) );
  NANDN U17151 ( .A(n15340), .B(n15339), .Z(n15344) );
  NANDN U17152 ( .A(n15342), .B(n15341), .Z(n15343) );
  AND U17153 ( .A(n15344), .B(n15343), .Z(n15379) );
  NANDN U17154 ( .A(n15346), .B(n15345), .Z(n15350) );
  NANDN U17155 ( .A(n15348), .B(n15347), .Z(n15349) );
  AND U17156 ( .A(n15350), .B(n15349), .Z(n15377) );
  NAND U17157 ( .A(n42143), .B(n15351), .Z(n15353) );
  XNOR U17158 ( .A(a[299]), .B(n4114), .Z(n15388) );
  NAND U17159 ( .A(n42144), .B(n15388), .Z(n15352) );
  AND U17160 ( .A(n15353), .B(n15352), .Z(n15403) );
  XOR U17161 ( .A(a[303]), .B(n42012), .Z(n15391) );
  XNOR U17162 ( .A(n15403), .B(n15402), .Z(n15405) );
  XOR U17163 ( .A(a[301]), .B(n42085), .Z(n15395) );
  AND U17164 ( .A(a[297]), .B(b[7]), .Z(n15396) );
  XNOR U17165 ( .A(n15397), .B(n15396), .Z(n15398) );
  AND U17166 ( .A(a[305]), .B(b[0]), .Z(n15356) );
  XNOR U17167 ( .A(n15356), .B(n4071), .Z(n15358) );
  NANDN U17168 ( .A(b[0]), .B(a[304]), .Z(n15357) );
  NAND U17169 ( .A(n15358), .B(n15357), .Z(n15399) );
  XNOR U17170 ( .A(n15398), .B(n15399), .Z(n15404) );
  XOR U17171 ( .A(n15405), .B(n15404), .Z(n15383) );
  NANDN U17172 ( .A(n15360), .B(n15359), .Z(n15364) );
  NANDN U17173 ( .A(n15362), .B(n15361), .Z(n15363) );
  AND U17174 ( .A(n15364), .B(n15363), .Z(n15382) );
  XNOR U17175 ( .A(n15383), .B(n15382), .Z(n15384) );
  NANDN U17176 ( .A(n15366), .B(n15365), .Z(n15370) );
  NAND U17177 ( .A(n15368), .B(n15367), .Z(n15369) );
  NAND U17178 ( .A(n15370), .B(n15369), .Z(n15385) );
  XNOR U17179 ( .A(n15384), .B(n15385), .Z(n15376) );
  XNOR U17180 ( .A(n15377), .B(n15376), .Z(n15378) );
  XNOR U17181 ( .A(n15379), .B(n15378), .Z(n15408) );
  XNOR U17182 ( .A(sreg[1321]), .B(n15408), .Z(n15410) );
  NANDN U17183 ( .A(sreg[1320]), .B(n15371), .Z(n15375) );
  NAND U17184 ( .A(n15373), .B(n15372), .Z(n15374) );
  NAND U17185 ( .A(n15375), .B(n15374), .Z(n15409) );
  XNOR U17186 ( .A(n15410), .B(n15409), .Z(c[1321]) );
  NANDN U17187 ( .A(n15377), .B(n15376), .Z(n15381) );
  NANDN U17188 ( .A(n15379), .B(n15378), .Z(n15380) );
  AND U17189 ( .A(n15381), .B(n15380), .Z(n15416) );
  NANDN U17190 ( .A(n15383), .B(n15382), .Z(n15387) );
  NANDN U17191 ( .A(n15385), .B(n15384), .Z(n15386) );
  AND U17192 ( .A(n15387), .B(n15386), .Z(n15414) );
  NAND U17193 ( .A(n42143), .B(n15388), .Z(n15390) );
  XNOR U17194 ( .A(a[300]), .B(n4114), .Z(n15425) );
  NAND U17195 ( .A(n42144), .B(n15425), .Z(n15389) );
  AND U17196 ( .A(n15390), .B(n15389), .Z(n15440) );
  XOR U17197 ( .A(a[304]), .B(n42012), .Z(n15428) );
  XNOR U17198 ( .A(n15440), .B(n15439), .Z(n15442) );
  AND U17199 ( .A(a[306]), .B(b[0]), .Z(n15392) );
  XNOR U17200 ( .A(n15392), .B(n4071), .Z(n15394) );
  NANDN U17201 ( .A(b[0]), .B(a[305]), .Z(n15393) );
  NAND U17202 ( .A(n15394), .B(n15393), .Z(n15436) );
  XOR U17203 ( .A(a[302]), .B(n42085), .Z(n15429) );
  AND U17204 ( .A(a[298]), .B(b[7]), .Z(n15433) );
  XNOR U17205 ( .A(n15434), .B(n15433), .Z(n15435) );
  XNOR U17206 ( .A(n15436), .B(n15435), .Z(n15441) );
  XOR U17207 ( .A(n15442), .B(n15441), .Z(n15420) );
  NANDN U17208 ( .A(n15397), .B(n15396), .Z(n15401) );
  NANDN U17209 ( .A(n15399), .B(n15398), .Z(n15400) );
  AND U17210 ( .A(n15401), .B(n15400), .Z(n15419) );
  XNOR U17211 ( .A(n15420), .B(n15419), .Z(n15421) );
  NANDN U17212 ( .A(n15403), .B(n15402), .Z(n15407) );
  NAND U17213 ( .A(n15405), .B(n15404), .Z(n15406) );
  NAND U17214 ( .A(n15407), .B(n15406), .Z(n15422) );
  XNOR U17215 ( .A(n15421), .B(n15422), .Z(n15413) );
  XNOR U17216 ( .A(n15414), .B(n15413), .Z(n15415) );
  XNOR U17217 ( .A(n15416), .B(n15415), .Z(n15445) );
  XNOR U17218 ( .A(sreg[1322]), .B(n15445), .Z(n15447) );
  NANDN U17219 ( .A(sreg[1321]), .B(n15408), .Z(n15412) );
  NAND U17220 ( .A(n15410), .B(n15409), .Z(n15411) );
  NAND U17221 ( .A(n15412), .B(n15411), .Z(n15446) );
  XNOR U17222 ( .A(n15447), .B(n15446), .Z(c[1322]) );
  NANDN U17223 ( .A(n15414), .B(n15413), .Z(n15418) );
  NANDN U17224 ( .A(n15416), .B(n15415), .Z(n15417) );
  AND U17225 ( .A(n15418), .B(n15417), .Z(n15453) );
  NANDN U17226 ( .A(n15420), .B(n15419), .Z(n15424) );
  NANDN U17227 ( .A(n15422), .B(n15421), .Z(n15423) );
  AND U17228 ( .A(n15424), .B(n15423), .Z(n15451) );
  NAND U17229 ( .A(n42143), .B(n15425), .Z(n15427) );
  XNOR U17230 ( .A(a[301]), .B(n4114), .Z(n15462) );
  NAND U17231 ( .A(n42144), .B(n15462), .Z(n15426) );
  AND U17232 ( .A(n15427), .B(n15426), .Z(n15477) );
  XOR U17233 ( .A(a[305]), .B(n42012), .Z(n15465) );
  XNOR U17234 ( .A(n15477), .B(n15476), .Z(n15479) );
  XOR U17235 ( .A(a[303]), .B(n42085), .Z(n15469) );
  AND U17236 ( .A(a[299]), .B(b[7]), .Z(n15470) );
  XNOR U17237 ( .A(n15471), .B(n15470), .Z(n15472) );
  AND U17238 ( .A(a[307]), .B(b[0]), .Z(n15430) );
  XNOR U17239 ( .A(n15430), .B(n4071), .Z(n15432) );
  NANDN U17240 ( .A(b[0]), .B(a[306]), .Z(n15431) );
  NAND U17241 ( .A(n15432), .B(n15431), .Z(n15473) );
  XNOR U17242 ( .A(n15472), .B(n15473), .Z(n15478) );
  XOR U17243 ( .A(n15479), .B(n15478), .Z(n15457) );
  NANDN U17244 ( .A(n15434), .B(n15433), .Z(n15438) );
  NANDN U17245 ( .A(n15436), .B(n15435), .Z(n15437) );
  AND U17246 ( .A(n15438), .B(n15437), .Z(n15456) );
  XNOR U17247 ( .A(n15457), .B(n15456), .Z(n15458) );
  NANDN U17248 ( .A(n15440), .B(n15439), .Z(n15444) );
  NAND U17249 ( .A(n15442), .B(n15441), .Z(n15443) );
  NAND U17250 ( .A(n15444), .B(n15443), .Z(n15459) );
  XNOR U17251 ( .A(n15458), .B(n15459), .Z(n15450) );
  XNOR U17252 ( .A(n15451), .B(n15450), .Z(n15452) );
  XNOR U17253 ( .A(n15453), .B(n15452), .Z(n15482) );
  XNOR U17254 ( .A(sreg[1323]), .B(n15482), .Z(n15484) );
  NANDN U17255 ( .A(sreg[1322]), .B(n15445), .Z(n15449) );
  NAND U17256 ( .A(n15447), .B(n15446), .Z(n15448) );
  NAND U17257 ( .A(n15449), .B(n15448), .Z(n15483) );
  XNOR U17258 ( .A(n15484), .B(n15483), .Z(c[1323]) );
  NANDN U17259 ( .A(n15451), .B(n15450), .Z(n15455) );
  NANDN U17260 ( .A(n15453), .B(n15452), .Z(n15454) );
  AND U17261 ( .A(n15455), .B(n15454), .Z(n15490) );
  NANDN U17262 ( .A(n15457), .B(n15456), .Z(n15461) );
  NANDN U17263 ( .A(n15459), .B(n15458), .Z(n15460) );
  AND U17264 ( .A(n15461), .B(n15460), .Z(n15488) );
  NAND U17265 ( .A(n42143), .B(n15462), .Z(n15464) );
  XNOR U17266 ( .A(a[302]), .B(n4115), .Z(n15499) );
  NAND U17267 ( .A(n42144), .B(n15499), .Z(n15463) );
  AND U17268 ( .A(n15464), .B(n15463), .Z(n15514) );
  XOR U17269 ( .A(a[306]), .B(n42012), .Z(n15502) );
  XNOR U17270 ( .A(n15514), .B(n15513), .Z(n15516) );
  AND U17271 ( .A(a[308]), .B(b[0]), .Z(n15466) );
  XNOR U17272 ( .A(n15466), .B(n4071), .Z(n15468) );
  NANDN U17273 ( .A(b[0]), .B(a[307]), .Z(n15467) );
  NAND U17274 ( .A(n15468), .B(n15467), .Z(n15510) );
  XOR U17275 ( .A(a[304]), .B(n42085), .Z(n15503) );
  AND U17276 ( .A(a[300]), .B(b[7]), .Z(n15507) );
  XNOR U17277 ( .A(n15508), .B(n15507), .Z(n15509) );
  XNOR U17278 ( .A(n15510), .B(n15509), .Z(n15515) );
  XOR U17279 ( .A(n15516), .B(n15515), .Z(n15494) );
  NANDN U17280 ( .A(n15471), .B(n15470), .Z(n15475) );
  NANDN U17281 ( .A(n15473), .B(n15472), .Z(n15474) );
  AND U17282 ( .A(n15475), .B(n15474), .Z(n15493) );
  XNOR U17283 ( .A(n15494), .B(n15493), .Z(n15495) );
  NANDN U17284 ( .A(n15477), .B(n15476), .Z(n15481) );
  NAND U17285 ( .A(n15479), .B(n15478), .Z(n15480) );
  NAND U17286 ( .A(n15481), .B(n15480), .Z(n15496) );
  XNOR U17287 ( .A(n15495), .B(n15496), .Z(n15487) );
  XNOR U17288 ( .A(n15488), .B(n15487), .Z(n15489) );
  XNOR U17289 ( .A(n15490), .B(n15489), .Z(n15519) );
  XNOR U17290 ( .A(sreg[1324]), .B(n15519), .Z(n15521) );
  NANDN U17291 ( .A(sreg[1323]), .B(n15482), .Z(n15486) );
  NAND U17292 ( .A(n15484), .B(n15483), .Z(n15485) );
  NAND U17293 ( .A(n15486), .B(n15485), .Z(n15520) );
  XNOR U17294 ( .A(n15521), .B(n15520), .Z(c[1324]) );
  NANDN U17295 ( .A(n15488), .B(n15487), .Z(n15492) );
  NANDN U17296 ( .A(n15490), .B(n15489), .Z(n15491) );
  AND U17297 ( .A(n15492), .B(n15491), .Z(n15527) );
  NANDN U17298 ( .A(n15494), .B(n15493), .Z(n15498) );
  NANDN U17299 ( .A(n15496), .B(n15495), .Z(n15497) );
  AND U17300 ( .A(n15498), .B(n15497), .Z(n15525) );
  NAND U17301 ( .A(n42143), .B(n15499), .Z(n15501) );
  XNOR U17302 ( .A(a[303]), .B(n4115), .Z(n15536) );
  NAND U17303 ( .A(n42144), .B(n15536), .Z(n15500) );
  AND U17304 ( .A(n15501), .B(n15500), .Z(n15551) );
  XOR U17305 ( .A(a[307]), .B(n42012), .Z(n15539) );
  XNOR U17306 ( .A(n15551), .B(n15550), .Z(n15553) );
  XOR U17307 ( .A(a[305]), .B(n42085), .Z(n15543) );
  AND U17308 ( .A(a[301]), .B(b[7]), .Z(n15544) );
  XNOR U17309 ( .A(n15545), .B(n15544), .Z(n15546) );
  AND U17310 ( .A(a[309]), .B(b[0]), .Z(n15504) );
  XNOR U17311 ( .A(n15504), .B(n4071), .Z(n15506) );
  NANDN U17312 ( .A(b[0]), .B(a[308]), .Z(n15505) );
  NAND U17313 ( .A(n15506), .B(n15505), .Z(n15547) );
  XNOR U17314 ( .A(n15546), .B(n15547), .Z(n15552) );
  XOR U17315 ( .A(n15553), .B(n15552), .Z(n15531) );
  NANDN U17316 ( .A(n15508), .B(n15507), .Z(n15512) );
  NANDN U17317 ( .A(n15510), .B(n15509), .Z(n15511) );
  AND U17318 ( .A(n15512), .B(n15511), .Z(n15530) );
  XNOR U17319 ( .A(n15531), .B(n15530), .Z(n15532) );
  NANDN U17320 ( .A(n15514), .B(n15513), .Z(n15518) );
  NAND U17321 ( .A(n15516), .B(n15515), .Z(n15517) );
  NAND U17322 ( .A(n15518), .B(n15517), .Z(n15533) );
  XNOR U17323 ( .A(n15532), .B(n15533), .Z(n15524) );
  XNOR U17324 ( .A(n15525), .B(n15524), .Z(n15526) );
  XNOR U17325 ( .A(n15527), .B(n15526), .Z(n15556) );
  XNOR U17326 ( .A(sreg[1325]), .B(n15556), .Z(n15558) );
  NANDN U17327 ( .A(sreg[1324]), .B(n15519), .Z(n15523) );
  NAND U17328 ( .A(n15521), .B(n15520), .Z(n15522) );
  NAND U17329 ( .A(n15523), .B(n15522), .Z(n15557) );
  XNOR U17330 ( .A(n15558), .B(n15557), .Z(c[1325]) );
  NANDN U17331 ( .A(n15525), .B(n15524), .Z(n15529) );
  NANDN U17332 ( .A(n15527), .B(n15526), .Z(n15528) );
  AND U17333 ( .A(n15529), .B(n15528), .Z(n15564) );
  NANDN U17334 ( .A(n15531), .B(n15530), .Z(n15535) );
  NANDN U17335 ( .A(n15533), .B(n15532), .Z(n15534) );
  AND U17336 ( .A(n15535), .B(n15534), .Z(n15562) );
  NAND U17337 ( .A(n42143), .B(n15536), .Z(n15538) );
  XNOR U17338 ( .A(a[304]), .B(n4115), .Z(n15573) );
  NAND U17339 ( .A(n42144), .B(n15573), .Z(n15537) );
  AND U17340 ( .A(n15538), .B(n15537), .Z(n15588) );
  XOR U17341 ( .A(a[308]), .B(n42012), .Z(n15576) );
  XNOR U17342 ( .A(n15588), .B(n15587), .Z(n15590) );
  AND U17343 ( .A(a[310]), .B(b[0]), .Z(n15540) );
  XNOR U17344 ( .A(n15540), .B(n4071), .Z(n15542) );
  NANDN U17345 ( .A(b[0]), .B(a[309]), .Z(n15541) );
  NAND U17346 ( .A(n15542), .B(n15541), .Z(n15584) );
  XOR U17347 ( .A(a[306]), .B(n42085), .Z(n15580) );
  AND U17348 ( .A(a[302]), .B(b[7]), .Z(n15581) );
  XNOR U17349 ( .A(n15582), .B(n15581), .Z(n15583) );
  XNOR U17350 ( .A(n15584), .B(n15583), .Z(n15589) );
  XOR U17351 ( .A(n15590), .B(n15589), .Z(n15568) );
  NANDN U17352 ( .A(n15545), .B(n15544), .Z(n15549) );
  NANDN U17353 ( .A(n15547), .B(n15546), .Z(n15548) );
  AND U17354 ( .A(n15549), .B(n15548), .Z(n15567) );
  XNOR U17355 ( .A(n15568), .B(n15567), .Z(n15569) );
  NANDN U17356 ( .A(n15551), .B(n15550), .Z(n15555) );
  NAND U17357 ( .A(n15553), .B(n15552), .Z(n15554) );
  NAND U17358 ( .A(n15555), .B(n15554), .Z(n15570) );
  XNOR U17359 ( .A(n15569), .B(n15570), .Z(n15561) );
  XNOR U17360 ( .A(n15562), .B(n15561), .Z(n15563) );
  XNOR U17361 ( .A(n15564), .B(n15563), .Z(n15593) );
  XNOR U17362 ( .A(sreg[1326]), .B(n15593), .Z(n15595) );
  NANDN U17363 ( .A(sreg[1325]), .B(n15556), .Z(n15560) );
  NAND U17364 ( .A(n15558), .B(n15557), .Z(n15559) );
  NAND U17365 ( .A(n15560), .B(n15559), .Z(n15594) );
  XNOR U17366 ( .A(n15595), .B(n15594), .Z(c[1326]) );
  NANDN U17367 ( .A(n15562), .B(n15561), .Z(n15566) );
  NANDN U17368 ( .A(n15564), .B(n15563), .Z(n15565) );
  AND U17369 ( .A(n15566), .B(n15565), .Z(n15601) );
  NANDN U17370 ( .A(n15568), .B(n15567), .Z(n15572) );
  NANDN U17371 ( .A(n15570), .B(n15569), .Z(n15571) );
  AND U17372 ( .A(n15572), .B(n15571), .Z(n15599) );
  NAND U17373 ( .A(n42143), .B(n15573), .Z(n15575) );
  XNOR U17374 ( .A(a[305]), .B(n4115), .Z(n15610) );
  NAND U17375 ( .A(n42144), .B(n15610), .Z(n15574) );
  AND U17376 ( .A(n15575), .B(n15574), .Z(n15625) );
  XOR U17377 ( .A(a[309]), .B(n42012), .Z(n15613) );
  XNOR U17378 ( .A(n15625), .B(n15624), .Z(n15627) );
  AND U17379 ( .A(a[311]), .B(b[0]), .Z(n15577) );
  XNOR U17380 ( .A(n15577), .B(n4071), .Z(n15579) );
  NANDN U17381 ( .A(b[0]), .B(a[310]), .Z(n15578) );
  NAND U17382 ( .A(n15579), .B(n15578), .Z(n15621) );
  XOR U17383 ( .A(a[307]), .B(n42085), .Z(n15617) );
  AND U17384 ( .A(a[303]), .B(b[7]), .Z(n15618) );
  XNOR U17385 ( .A(n15619), .B(n15618), .Z(n15620) );
  XNOR U17386 ( .A(n15621), .B(n15620), .Z(n15626) );
  XOR U17387 ( .A(n15627), .B(n15626), .Z(n15605) );
  NANDN U17388 ( .A(n15582), .B(n15581), .Z(n15586) );
  NANDN U17389 ( .A(n15584), .B(n15583), .Z(n15585) );
  AND U17390 ( .A(n15586), .B(n15585), .Z(n15604) );
  XNOR U17391 ( .A(n15605), .B(n15604), .Z(n15606) );
  NANDN U17392 ( .A(n15588), .B(n15587), .Z(n15592) );
  NAND U17393 ( .A(n15590), .B(n15589), .Z(n15591) );
  NAND U17394 ( .A(n15592), .B(n15591), .Z(n15607) );
  XNOR U17395 ( .A(n15606), .B(n15607), .Z(n15598) );
  XNOR U17396 ( .A(n15599), .B(n15598), .Z(n15600) );
  XNOR U17397 ( .A(n15601), .B(n15600), .Z(n15630) );
  XNOR U17398 ( .A(sreg[1327]), .B(n15630), .Z(n15632) );
  NANDN U17399 ( .A(sreg[1326]), .B(n15593), .Z(n15597) );
  NAND U17400 ( .A(n15595), .B(n15594), .Z(n15596) );
  NAND U17401 ( .A(n15597), .B(n15596), .Z(n15631) );
  XNOR U17402 ( .A(n15632), .B(n15631), .Z(c[1327]) );
  NANDN U17403 ( .A(n15599), .B(n15598), .Z(n15603) );
  NANDN U17404 ( .A(n15601), .B(n15600), .Z(n15602) );
  AND U17405 ( .A(n15603), .B(n15602), .Z(n15638) );
  NANDN U17406 ( .A(n15605), .B(n15604), .Z(n15609) );
  NANDN U17407 ( .A(n15607), .B(n15606), .Z(n15608) );
  AND U17408 ( .A(n15609), .B(n15608), .Z(n15636) );
  NAND U17409 ( .A(n42143), .B(n15610), .Z(n15612) );
  XNOR U17410 ( .A(a[306]), .B(n4115), .Z(n15647) );
  NAND U17411 ( .A(n42144), .B(n15647), .Z(n15611) );
  AND U17412 ( .A(n15612), .B(n15611), .Z(n15662) );
  XOR U17413 ( .A(a[310]), .B(n42012), .Z(n15650) );
  XNOR U17414 ( .A(n15662), .B(n15661), .Z(n15664) );
  AND U17415 ( .A(a[312]), .B(b[0]), .Z(n15614) );
  XNOR U17416 ( .A(n15614), .B(n4071), .Z(n15616) );
  NANDN U17417 ( .A(b[0]), .B(a[311]), .Z(n15615) );
  NAND U17418 ( .A(n15616), .B(n15615), .Z(n15658) );
  XOR U17419 ( .A(a[308]), .B(n42085), .Z(n15651) );
  AND U17420 ( .A(a[304]), .B(b[7]), .Z(n15655) );
  XNOR U17421 ( .A(n15656), .B(n15655), .Z(n15657) );
  XNOR U17422 ( .A(n15658), .B(n15657), .Z(n15663) );
  XOR U17423 ( .A(n15664), .B(n15663), .Z(n15642) );
  NANDN U17424 ( .A(n15619), .B(n15618), .Z(n15623) );
  NANDN U17425 ( .A(n15621), .B(n15620), .Z(n15622) );
  AND U17426 ( .A(n15623), .B(n15622), .Z(n15641) );
  XNOR U17427 ( .A(n15642), .B(n15641), .Z(n15643) );
  NANDN U17428 ( .A(n15625), .B(n15624), .Z(n15629) );
  NAND U17429 ( .A(n15627), .B(n15626), .Z(n15628) );
  NAND U17430 ( .A(n15629), .B(n15628), .Z(n15644) );
  XNOR U17431 ( .A(n15643), .B(n15644), .Z(n15635) );
  XNOR U17432 ( .A(n15636), .B(n15635), .Z(n15637) );
  XNOR U17433 ( .A(n15638), .B(n15637), .Z(n15667) );
  XNOR U17434 ( .A(sreg[1328]), .B(n15667), .Z(n15669) );
  NANDN U17435 ( .A(sreg[1327]), .B(n15630), .Z(n15634) );
  NAND U17436 ( .A(n15632), .B(n15631), .Z(n15633) );
  NAND U17437 ( .A(n15634), .B(n15633), .Z(n15668) );
  XNOR U17438 ( .A(n15669), .B(n15668), .Z(c[1328]) );
  NANDN U17439 ( .A(n15636), .B(n15635), .Z(n15640) );
  NANDN U17440 ( .A(n15638), .B(n15637), .Z(n15639) );
  AND U17441 ( .A(n15640), .B(n15639), .Z(n15675) );
  NANDN U17442 ( .A(n15642), .B(n15641), .Z(n15646) );
  NANDN U17443 ( .A(n15644), .B(n15643), .Z(n15645) );
  AND U17444 ( .A(n15646), .B(n15645), .Z(n15673) );
  NAND U17445 ( .A(n42143), .B(n15647), .Z(n15649) );
  XNOR U17446 ( .A(a[307]), .B(n4115), .Z(n15684) );
  NAND U17447 ( .A(n42144), .B(n15684), .Z(n15648) );
  AND U17448 ( .A(n15649), .B(n15648), .Z(n15699) );
  XOR U17449 ( .A(a[311]), .B(n42012), .Z(n15687) );
  XNOR U17450 ( .A(n15699), .B(n15698), .Z(n15701) );
  XOR U17451 ( .A(a[309]), .B(n42085), .Z(n15691) );
  AND U17452 ( .A(a[305]), .B(b[7]), .Z(n15692) );
  XNOR U17453 ( .A(n15693), .B(n15692), .Z(n15694) );
  AND U17454 ( .A(a[313]), .B(b[0]), .Z(n15652) );
  XNOR U17455 ( .A(n15652), .B(n4071), .Z(n15654) );
  NANDN U17456 ( .A(b[0]), .B(a[312]), .Z(n15653) );
  NAND U17457 ( .A(n15654), .B(n15653), .Z(n15695) );
  XNOR U17458 ( .A(n15694), .B(n15695), .Z(n15700) );
  XOR U17459 ( .A(n15701), .B(n15700), .Z(n15679) );
  NANDN U17460 ( .A(n15656), .B(n15655), .Z(n15660) );
  NANDN U17461 ( .A(n15658), .B(n15657), .Z(n15659) );
  AND U17462 ( .A(n15660), .B(n15659), .Z(n15678) );
  XNOR U17463 ( .A(n15679), .B(n15678), .Z(n15680) );
  NANDN U17464 ( .A(n15662), .B(n15661), .Z(n15666) );
  NAND U17465 ( .A(n15664), .B(n15663), .Z(n15665) );
  NAND U17466 ( .A(n15666), .B(n15665), .Z(n15681) );
  XNOR U17467 ( .A(n15680), .B(n15681), .Z(n15672) );
  XNOR U17468 ( .A(n15673), .B(n15672), .Z(n15674) );
  XNOR U17469 ( .A(n15675), .B(n15674), .Z(n15704) );
  XNOR U17470 ( .A(sreg[1329]), .B(n15704), .Z(n15706) );
  NANDN U17471 ( .A(sreg[1328]), .B(n15667), .Z(n15671) );
  NAND U17472 ( .A(n15669), .B(n15668), .Z(n15670) );
  NAND U17473 ( .A(n15671), .B(n15670), .Z(n15705) );
  XNOR U17474 ( .A(n15706), .B(n15705), .Z(c[1329]) );
  NANDN U17475 ( .A(n15673), .B(n15672), .Z(n15677) );
  NANDN U17476 ( .A(n15675), .B(n15674), .Z(n15676) );
  AND U17477 ( .A(n15677), .B(n15676), .Z(n15712) );
  NANDN U17478 ( .A(n15679), .B(n15678), .Z(n15683) );
  NANDN U17479 ( .A(n15681), .B(n15680), .Z(n15682) );
  AND U17480 ( .A(n15683), .B(n15682), .Z(n15710) );
  NAND U17481 ( .A(n42143), .B(n15684), .Z(n15686) );
  XNOR U17482 ( .A(a[308]), .B(n4115), .Z(n15721) );
  NAND U17483 ( .A(n42144), .B(n15721), .Z(n15685) );
  AND U17484 ( .A(n15686), .B(n15685), .Z(n15736) );
  XOR U17485 ( .A(a[312]), .B(n42012), .Z(n15724) );
  XNOR U17486 ( .A(n15736), .B(n15735), .Z(n15738) );
  AND U17487 ( .A(a[314]), .B(b[0]), .Z(n15688) );
  XNOR U17488 ( .A(n15688), .B(n4071), .Z(n15690) );
  NANDN U17489 ( .A(b[0]), .B(a[313]), .Z(n15689) );
  NAND U17490 ( .A(n15690), .B(n15689), .Z(n15732) );
  XOR U17491 ( .A(a[310]), .B(n42085), .Z(n15728) );
  AND U17492 ( .A(a[306]), .B(b[7]), .Z(n15729) );
  XNOR U17493 ( .A(n15730), .B(n15729), .Z(n15731) );
  XNOR U17494 ( .A(n15732), .B(n15731), .Z(n15737) );
  XOR U17495 ( .A(n15738), .B(n15737), .Z(n15716) );
  NANDN U17496 ( .A(n15693), .B(n15692), .Z(n15697) );
  NANDN U17497 ( .A(n15695), .B(n15694), .Z(n15696) );
  AND U17498 ( .A(n15697), .B(n15696), .Z(n15715) );
  XNOR U17499 ( .A(n15716), .B(n15715), .Z(n15717) );
  NANDN U17500 ( .A(n15699), .B(n15698), .Z(n15703) );
  NAND U17501 ( .A(n15701), .B(n15700), .Z(n15702) );
  NAND U17502 ( .A(n15703), .B(n15702), .Z(n15718) );
  XNOR U17503 ( .A(n15717), .B(n15718), .Z(n15709) );
  XNOR U17504 ( .A(n15710), .B(n15709), .Z(n15711) );
  XNOR U17505 ( .A(n15712), .B(n15711), .Z(n15741) );
  XNOR U17506 ( .A(sreg[1330]), .B(n15741), .Z(n15743) );
  NANDN U17507 ( .A(sreg[1329]), .B(n15704), .Z(n15708) );
  NAND U17508 ( .A(n15706), .B(n15705), .Z(n15707) );
  NAND U17509 ( .A(n15708), .B(n15707), .Z(n15742) );
  XNOR U17510 ( .A(n15743), .B(n15742), .Z(c[1330]) );
  NANDN U17511 ( .A(n15710), .B(n15709), .Z(n15714) );
  NANDN U17512 ( .A(n15712), .B(n15711), .Z(n15713) );
  AND U17513 ( .A(n15714), .B(n15713), .Z(n15749) );
  NANDN U17514 ( .A(n15716), .B(n15715), .Z(n15720) );
  NANDN U17515 ( .A(n15718), .B(n15717), .Z(n15719) );
  AND U17516 ( .A(n15720), .B(n15719), .Z(n15747) );
  NAND U17517 ( .A(n42143), .B(n15721), .Z(n15723) );
  XNOR U17518 ( .A(a[309]), .B(n4116), .Z(n15758) );
  NAND U17519 ( .A(n42144), .B(n15758), .Z(n15722) );
  AND U17520 ( .A(n15723), .B(n15722), .Z(n15773) );
  XOR U17521 ( .A(a[313]), .B(n42012), .Z(n15761) );
  XNOR U17522 ( .A(n15773), .B(n15772), .Z(n15775) );
  AND U17523 ( .A(a[315]), .B(b[0]), .Z(n15725) );
  XNOR U17524 ( .A(n15725), .B(n4071), .Z(n15727) );
  NANDN U17525 ( .A(b[0]), .B(a[314]), .Z(n15726) );
  NAND U17526 ( .A(n15727), .B(n15726), .Z(n15769) );
  XOR U17527 ( .A(a[311]), .B(n42085), .Z(n15762) );
  AND U17528 ( .A(a[307]), .B(b[7]), .Z(n15766) );
  XNOR U17529 ( .A(n15767), .B(n15766), .Z(n15768) );
  XNOR U17530 ( .A(n15769), .B(n15768), .Z(n15774) );
  XOR U17531 ( .A(n15775), .B(n15774), .Z(n15753) );
  NANDN U17532 ( .A(n15730), .B(n15729), .Z(n15734) );
  NANDN U17533 ( .A(n15732), .B(n15731), .Z(n15733) );
  AND U17534 ( .A(n15734), .B(n15733), .Z(n15752) );
  XNOR U17535 ( .A(n15753), .B(n15752), .Z(n15754) );
  NANDN U17536 ( .A(n15736), .B(n15735), .Z(n15740) );
  NAND U17537 ( .A(n15738), .B(n15737), .Z(n15739) );
  NAND U17538 ( .A(n15740), .B(n15739), .Z(n15755) );
  XNOR U17539 ( .A(n15754), .B(n15755), .Z(n15746) );
  XNOR U17540 ( .A(n15747), .B(n15746), .Z(n15748) );
  XNOR U17541 ( .A(n15749), .B(n15748), .Z(n15778) );
  XNOR U17542 ( .A(sreg[1331]), .B(n15778), .Z(n15780) );
  NANDN U17543 ( .A(sreg[1330]), .B(n15741), .Z(n15745) );
  NAND U17544 ( .A(n15743), .B(n15742), .Z(n15744) );
  NAND U17545 ( .A(n15745), .B(n15744), .Z(n15779) );
  XNOR U17546 ( .A(n15780), .B(n15779), .Z(c[1331]) );
  NANDN U17547 ( .A(n15747), .B(n15746), .Z(n15751) );
  NANDN U17548 ( .A(n15749), .B(n15748), .Z(n15750) );
  AND U17549 ( .A(n15751), .B(n15750), .Z(n15786) );
  NANDN U17550 ( .A(n15753), .B(n15752), .Z(n15757) );
  NANDN U17551 ( .A(n15755), .B(n15754), .Z(n15756) );
  AND U17552 ( .A(n15757), .B(n15756), .Z(n15784) );
  NAND U17553 ( .A(n42143), .B(n15758), .Z(n15760) );
  XNOR U17554 ( .A(a[310]), .B(n4116), .Z(n15795) );
  NAND U17555 ( .A(n42144), .B(n15795), .Z(n15759) );
  AND U17556 ( .A(n15760), .B(n15759), .Z(n15810) );
  XOR U17557 ( .A(a[314]), .B(n42012), .Z(n15798) );
  XNOR U17558 ( .A(n15810), .B(n15809), .Z(n15812) );
  XOR U17559 ( .A(a[312]), .B(n42085), .Z(n15802) );
  AND U17560 ( .A(a[308]), .B(b[7]), .Z(n15803) );
  XNOR U17561 ( .A(n15804), .B(n15803), .Z(n15805) );
  AND U17562 ( .A(a[316]), .B(b[0]), .Z(n15763) );
  XNOR U17563 ( .A(n15763), .B(n4071), .Z(n15765) );
  NANDN U17564 ( .A(b[0]), .B(a[315]), .Z(n15764) );
  NAND U17565 ( .A(n15765), .B(n15764), .Z(n15806) );
  XNOR U17566 ( .A(n15805), .B(n15806), .Z(n15811) );
  XOR U17567 ( .A(n15812), .B(n15811), .Z(n15790) );
  NANDN U17568 ( .A(n15767), .B(n15766), .Z(n15771) );
  NANDN U17569 ( .A(n15769), .B(n15768), .Z(n15770) );
  AND U17570 ( .A(n15771), .B(n15770), .Z(n15789) );
  XNOR U17571 ( .A(n15790), .B(n15789), .Z(n15791) );
  NANDN U17572 ( .A(n15773), .B(n15772), .Z(n15777) );
  NAND U17573 ( .A(n15775), .B(n15774), .Z(n15776) );
  NAND U17574 ( .A(n15777), .B(n15776), .Z(n15792) );
  XNOR U17575 ( .A(n15791), .B(n15792), .Z(n15783) );
  XNOR U17576 ( .A(n15784), .B(n15783), .Z(n15785) );
  XNOR U17577 ( .A(n15786), .B(n15785), .Z(n15815) );
  XNOR U17578 ( .A(sreg[1332]), .B(n15815), .Z(n15817) );
  NANDN U17579 ( .A(sreg[1331]), .B(n15778), .Z(n15782) );
  NAND U17580 ( .A(n15780), .B(n15779), .Z(n15781) );
  NAND U17581 ( .A(n15782), .B(n15781), .Z(n15816) );
  XNOR U17582 ( .A(n15817), .B(n15816), .Z(c[1332]) );
  NANDN U17583 ( .A(n15784), .B(n15783), .Z(n15788) );
  NANDN U17584 ( .A(n15786), .B(n15785), .Z(n15787) );
  AND U17585 ( .A(n15788), .B(n15787), .Z(n15823) );
  NANDN U17586 ( .A(n15790), .B(n15789), .Z(n15794) );
  NANDN U17587 ( .A(n15792), .B(n15791), .Z(n15793) );
  AND U17588 ( .A(n15794), .B(n15793), .Z(n15821) );
  NAND U17589 ( .A(n42143), .B(n15795), .Z(n15797) );
  XNOR U17590 ( .A(a[311]), .B(n4116), .Z(n15832) );
  NAND U17591 ( .A(n42144), .B(n15832), .Z(n15796) );
  AND U17592 ( .A(n15797), .B(n15796), .Z(n15847) );
  XOR U17593 ( .A(a[315]), .B(n42012), .Z(n15835) );
  XNOR U17594 ( .A(n15847), .B(n15846), .Z(n15849) );
  AND U17595 ( .A(a[317]), .B(b[0]), .Z(n15799) );
  XNOR U17596 ( .A(n15799), .B(n4071), .Z(n15801) );
  NANDN U17597 ( .A(b[0]), .B(a[316]), .Z(n15800) );
  NAND U17598 ( .A(n15801), .B(n15800), .Z(n15843) );
  XOR U17599 ( .A(a[313]), .B(n42085), .Z(n15836) );
  AND U17600 ( .A(a[309]), .B(b[7]), .Z(n15840) );
  XNOR U17601 ( .A(n15841), .B(n15840), .Z(n15842) );
  XNOR U17602 ( .A(n15843), .B(n15842), .Z(n15848) );
  XOR U17603 ( .A(n15849), .B(n15848), .Z(n15827) );
  NANDN U17604 ( .A(n15804), .B(n15803), .Z(n15808) );
  NANDN U17605 ( .A(n15806), .B(n15805), .Z(n15807) );
  AND U17606 ( .A(n15808), .B(n15807), .Z(n15826) );
  XNOR U17607 ( .A(n15827), .B(n15826), .Z(n15828) );
  NANDN U17608 ( .A(n15810), .B(n15809), .Z(n15814) );
  NAND U17609 ( .A(n15812), .B(n15811), .Z(n15813) );
  NAND U17610 ( .A(n15814), .B(n15813), .Z(n15829) );
  XNOR U17611 ( .A(n15828), .B(n15829), .Z(n15820) );
  XNOR U17612 ( .A(n15821), .B(n15820), .Z(n15822) );
  XNOR U17613 ( .A(n15823), .B(n15822), .Z(n15852) );
  XNOR U17614 ( .A(sreg[1333]), .B(n15852), .Z(n15854) );
  NANDN U17615 ( .A(sreg[1332]), .B(n15815), .Z(n15819) );
  NAND U17616 ( .A(n15817), .B(n15816), .Z(n15818) );
  NAND U17617 ( .A(n15819), .B(n15818), .Z(n15853) );
  XNOR U17618 ( .A(n15854), .B(n15853), .Z(c[1333]) );
  NANDN U17619 ( .A(n15821), .B(n15820), .Z(n15825) );
  NANDN U17620 ( .A(n15823), .B(n15822), .Z(n15824) );
  AND U17621 ( .A(n15825), .B(n15824), .Z(n15860) );
  NANDN U17622 ( .A(n15827), .B(n15826), .Z(n15831) );
  NANDN U17623 ( .A(n15829), .B(n15828), .Z(n15830) );
  AND U17624 ( .A(n15831), .B(n15830), .Z(n15858) );
  NAND U17625 ( .A(n42143), .B(n15832), .Z(n15834) );
  XNOR U17626 ( .A(a[312]), .B(n4116), .Z(n15869) );
  NAND U17627 ( .A(n42144), .B(n15869), .Z(n15833) );
  AND U17628 ( .A(n15834), .B(n15833), .Z(n15884) );
  XOR U17629 ( .A(a[316]), .B(n42012), .Z(n15872) );
  XNOR U17630 ( .A(n15884), .B(n15883), .Z(n15886) );
  XOR U17631 ( .A(a[314]), .B(n42085), .Z(n15876) );
  AND U17632 ( .A(a[310]), .B(b[7]), .Z(n15877) );
  XNOR U17633 ( .A(n15878), .B(n15877), .Z(n15879) );
  AND U17634 ( .A(a[318]), .B(b[0]), .Z(n15837) );
  XNOR U17635 ( .A(n15837), .B(n4071), .Z(n15839) );
  NANDN U17636 ( .A(b[0]), .B(a[317]), .Z(n15838) );
  NAND U17637 ( .A(n15839), .B(n15838), .Z(n15880) );
  XNOR U17638 ( .A(n15879), .B(n15880), .Z(n15885) );
  XOR U17639 ( .A(n15886), .B(n15885), .Z(n15864) );
  NANDN U17640 ( .A(n15841), .B(n15840), .Z(n15845) );
  NANDN U17641 ( .A(n15843), .B(n15842), .Z(n15844) );
  AND U17642 ( .A(n15845), .B(n15844), .Z(n15863) );
  XNOR U17643 ( .A(n15864), .B(n15863), .Z(n15865) );
  NANDN U17644 ( .A(n15847), .B(n15846), .Z(n15851) );
  NAND U17645 ( .A(n15849), .B(n15848), .Z(n15850) );
  NAND U17646 ( .A(n15851), .B(n15850), .Z(n15866) );
  XNOR U17647 ( .A(n15865), .B(n15866), .Z(n15857) );
  XNOR U17648 ( .A(n15858), .B(n15857), .Z(n15859) );
  XNOR U17649 ( .A(n15860), .B(n15859), .Z(n15889) );
  XNOR U17650 ( .A(sreg[1334]), .B(n15889), .Z(n15891) );
  NANDN U17651 ( .A(sreg[1333]), .B(n15852), .Z(n15856) );
  NAND U17652 ( .A(n15854), .B(n15853), .Z(n15855) );
  NAND U17653 ( .A(n15856), .B(n15855), .Z(n15890) );
  XNOR U17654 ( .A(n15891), .B(n15890), .Z(c[1334]) );
  NANDN U17655 ( .A(n15858), .B(n15857), .Z(n15862) );
  NANDN U17656 ( .A(n15860), .B(n15859), .Z(n15861) );
  AND U17657 ( .A(n15862), .B(n15861), .Z(n15897) );
  NANDN U17658 ( .A(n15864), .B(n15863), .Z(n15868) );
  NANDN U17659 ( .A(n15866), .B(n15865), .Z(n15867) );
  AND U17660 ( .A(n15868), .B(n15867), .Z(n15895) );
  NAND U17661 ( .A(n42143), .B(n15869), .Z(n15871) );
  XNOR U17662 ( .A(a[313]), .B(n4116), .Z(n15906) );
  NAND U17663 ( .A(n42144), .B(n15906), .Z(n15870) );
  AND U17664 ( .A(n15871), .B(n15870), .Z(n15921) );
  XOR U17665 ( .A(a[317]), .B(n42012), .Z(n15909) );
  XNOR U17666 ( .A(n15921), .B(n15920), .Z(n15923) );
  AND U17667 ( .A(a[319]), .B(b[0]), .Z(n15873) );
  XNOR U17668 ( .A(n15873), .B(n4071), .Z(n15875) );
  NANDN U17669 ( .A(b[0]), .B(a[318]), .Z(n15874) );
  NAND U17670 ( .A(n15875), .B(n15874), .Z(n15917) );
  XOR U17671 ( .A(a[315]), .B(n42085), .Z(n15913) );
  AND U17672 ( .A(a[311]), .B(b[7]), .Z(n15914) );
  XNOR U17673 ( .A(n15915), .B(n15914), .Z(n15916) );
  XNOR U17674 ( .A(n15917), .B(n15916), .Z(n15922) );
  XOR U17675 ( .A(n15923), .B(n15922), .Z(n15901) );
  NANDN U17676 ( .A(n15878), .B(n15877), .Z(n15882) );
  NANDN U17677 ( .A(n15880), .B(n15879), .Z(n15881) );
  AND U17678 ( .A(n15882), .B(n15881), .Z(n15900) );
  XNOR U17679 ( .A(n15901), .B(n15900), .Z(n15902) );
  NANDN U17680 ( .A(n15884), .B(n15883), .Z(n15888) );
  NAND U17681 ( .A(n15886), .B(n15885), .Z(n15887) );
  NAND U17682 ( .A(n15888), .B(n15887), .Z(n15903) );
  XNOR U17683 ( .A(n15902), .B(n15903), .Z(n15894) );
  XNOR U17684 ( .A(n15895), .B(n15894), .Z(n15896) );
  XNOR U17685 ( .A(n15897), .B(n15896), .Z(n15926) );
  XNOR U17686 ( .A(sreg[1335]), .B(n15926), .Z(n15928) );
  NANDN U17687 ( .A(sreg[1334]), .B(n15889), .Z(n15893) );
  NAND U17688 ( .A(n15891), .B(n15890), .Z(n15892) );
  NAND U17689 ( .A(n15893), .B(n15892), .Z(n15927) );
  XNOR U17690 ( .A(n15928), .B(n15927), .Z(c[1335]) );
  NANDN U17691 ( .A(n15895), .B(n15894), .Z(n15899) );
  NANDN U17692 ( .A(n15897), .B(n15896), .Z(n15898) );
  AND U17693 ( .A(n15899), .B(n15898), .Z(n15934) );
  NANDN U17694 ( .A(n15901), .B(n15900), .Z(n15905) );
  NANDN U17695 ( .A(n15903), .B(n15902), .Z(n15904) );
  AND U17696 ( .A(n15905), .B(n15904), .Z(n15932) );
  NAND U17697 ( .A(n42143), .B(n15906), .Z(n15908) );
  XNOR U17698 ( .A(a[314]), .B(n4116), .Z(n15943) );
  NAND U17699 ( .A(n42144), .B(n15943), .Z(n15907) );
  AND U17700 ( .A(n15908), .B(n15907), .Z(n15958) );
  XOR U17701 ( .A(a[318]), .B(n42012), .Z(n15946) );
  XNOR U17702 ( .A(n15958), .B(n15957), .Z(n15960) );
  AND U17703 ( .A(b[0]), .B(a[320]), .Z(n15910) );
  XOR U17704 ( .A(b[1]), .B(n15910), .Z(n15912) );
  NANDN U17705 ( .A(b[0]), .B(a[319]), .Z(n15911) );
  AND U17706 ( .A(n15912), .B(n15911), .Z(n15953) );
  XOR U17707 ( .A(a[316]), .B(n42085), .Z(n15950) );
  AND U17708 ( .A(a[312]), .B(b[7]), .Z(n15951) );
  XOR U17709 ( .A(n15952), .B(n15951), .Z(n15954) );
  XNOR U17710 ( .A(n15953), .B(n15954), .Z(n15959) );
  XOR U17711 ( .A(n15960), .B(n15959), .Z(n15938) );
  NANDN U17712 ( .A(n15915), .B(n15914), .Z(n15919) );
  NANDN U17713 ( .A(n15917), .B(n15916), .Z(n15918) );
  AND U17714 ( .A(n15919), .B(n15918), .Z(n15937) );
  XNOR U17715 ( .A(n15938), .B(n15937), .Z(n15939) );
  NANDN U17716 ( .A(n15921), .B(n15920), .Z(n15925) );
  NAND U17717 ( .A(n15923), .B(n15922), .Z(n15924) );
  NAND U17718 ( .A(n15925), .B(n15924), .Z(n15940) );
  XNOR U17719 ( .A(n15939), .B(n15940), .Z(n15931) );
  XNOR U17720 ( .A(n15932), .B(n15931), .Z(n15933) );
  XNOR U17721 ( .A(n15934), .B(n15933), .Z(n15963) );
  XNOR U17722 ( .A(sreg[1336]), .B(n15963), .Z(n15965) );
  NANDN U17723 ( .A(sreg[1335]), .B(n15926), .Z(n15930) );
  NAND U17724 ( .A(n15928), .B(n15927), .Z(n15929) );
  NAND U17725 ( .A(n15930), .B(n15929), .Z(n15964) );
  XNOR U17726 ( .A(n15965), .B(n15964), .Z(c[1336]) );
  NANDN U17727 ( .A(n15932), .B(n15931), .Z(n15936) );
  NANDN U17728 ( .A(n15934), .B(n15933), .Z(n15935) );
  AND U17729 ( .A(n15936), .B(n15935), .Z(n15971) );
  NANDN U17730 ( .A(n15938), .B(n15937), .Z(n15942) );
  NANDN U17731 ( .A(n15940), .B(n15939), .Z(n15941) );
  AND U17732 ( .A(n15942), .B(n15941), .Z(n15969) );
  NAND U17733 ( .A(n42143), .B(n15943), .Z(n15945) );
  XNOR U17734 ( .A(a[315]), .B(n4116), .Z(n15980) );
  NAND U17735 ( .A(n42144), .B(n15980), .Z(n15944) );
  AND U17736 ( .A(n15945), .B(n15944), .Z(n15995) );
  XOR U17737 ( .A(a[319]), .B(n42012), .Z(n15983) );
  XNOR U17738 ( .A(n15995), .B(n15994), .Z(n15997) );
  AND U17739 ( .A(a[321]), .B(b[0]), .Z(n15947) );
  XNOR U17740 ( .A(n15947), .B(n4071), .Z(n15949) );
  NANDN U17741 ( .A(b[0]), .B(a[320]), .Z(n15948) );
  NAND U17742 ( .A(n15949), .B(n15948), .Z(n15991) );
  XOR U17743 ( .A(a[317]), .B(n42085), .Z(n15984) );
  AND U17744 ( .A(a[313]), .B(b[7]), .Z(n15988) );
  XNOR U17745 ( .A(n15989), .B(n15988), .Z(n15990) );
  XNOR U17746 ( .A(n15991), .B(n15990), .Z(n15996) );
  XOR U17747 ( .A(n15997), .B(n15996), .Z(n15975) );
  NANDN U17748 ( .A(n15952), .B(n15951), .Z(n15956) );
  NANDN U17749 ( .A(n15954), .B(n15953), .Z(n15955) );
  AND U17750 ( .A(n15956), .B(n15955), .Z(n15974) );
  XNOR U17751 ( .A(n15975), .B(n15974), .Z(n15976) );
  NANDN U17752 ( .A(n15958), .B(n15957), .Z(n15962) );
  NAND U17753 ( .A(n15960), .B(n15959), .Z(n15961) );
  NAND U17754 ( .A(n15962), .B(n15961), .Z(n15977) );
  XNOR U17755 ( .A(n15976), .B(n15977), .Z(n15968) );
  XNOR U17756 ( .A(n15969), .B(n15968), .Z(n15970) );
  XNOR U17757 ( .A(n15971), .B(n15970), .Z(n16000) );
  XNOR U17758 ( .A(sreg[1337]), .B(n16000), .Z(n16002) );
  NANDN U17759 ( .A(sreg[1336]), .B(n15963), .Z(n15967) );
  NAND U17760 ( .A(n15965), .B(n15964), .Z(n15966) );
  NAND U17761 ( .A(n15967), .B(n15966), .Z(n16001) );
  XNOR U17762 ( .A(n16002), .B(n16001), .Z(c[1337]) );
  NANDN U17763 ( .A(n15969), .B(n15968), .Z(n15973) );
  NANDN U17764 ( .A(n15971), .B(n15970), .Z(n15972) );
  AND U17765 ( .A(n15973), .B(n15972), .Z(n16008) );
  NANDN U17766 ( .A(n15975), .B(n15974), .Z(n15979) );
  NANDN U17767 ( .A(n15977), .B(n15976), .Z(n15978) );
  AND U17768 ( .A(n15979), .B(n15978), .Z(n16006) );
  NAND U17769 ( .A(n42143), .B(n15980), .Z(n15982) );
  XNOR U17770 ( .A(a[316]), .B(n4117), .Z(n16017) );
  NAND U17771 ( .A(n42144), .B(n16017), .Z(n15981) );
  AND U17772 ( .A(n15982), .B(n15981), .Z(n16032) );
  XOR U17773 ( .A(a[320]), .B(n42012), .Z(n16020) );
  XNOR U17774 ( .A(n16032), .B(n16031), .Z(n16034) );
  XOR U17775 ( .A(a[318]), .B(n42085), .Z(n16024) );
  AND U17776 ( .A(a[314]), .B(b[7]), .Z(n16025) );
  XNOR U17777 ( .A(n16026), .B(n16025), .Z(n16027) );
  AND U17778 ( .A(a[322]), .B(b[0]), .Z(n15985) );
  XNOR U17779 ( .A(n15985), .B(n4071), .Z(n15987) );
  NANDN U17780 ( .A(b[0]), .B(a[321]), .Z(n15986) );
  NAND U17781 ( .A(n15987), .B(n15986), .Z(n16028) );
  XNOR U17782 ( .A(n16027), .B(n16028), .Z(n16033) );
  XOR U17783 ( .A(n16034), .B(n16033), .Z(n16012) );
  NANDN U17784 ( .A(n15989), .B(n15988), .Z(n15993) );
  NANDN U17785 ( .A(n15991), .B(n15990), .Z(n15992) );
  AND U17786 ( .A(n15993), .B(n15992), .Z(n16011) );
  XNOR U17787 ( .A(n16012), .B(n16011), .Z(n16013) );
  NANDN U17788 ( .A(n15995), .B(n15994), .Z(n15999) );
  NAND U17789 ( .A(n15997), .B(n15996), .Z(n15998) );
  NAND U17790 ( .A(n15999), .B(n15998), .Z(n16014) );
  XNOR U17791 ( .A(n16013), .B(n16014), .Z(n16005) );
  XNOR U17792 ( .A(n16006), .B(n16005), .Z(n16007) );
  XNOR U17793 ( .A(n16008), .B(n16007), .Z(n16037) );
  XNOR U17794 ( .A(sreg[1338]), .B(n16037), .Z(n16039) );
  NANDN U17795 ( .A(sreg[1337]), .B(n16000), .Z(n16004) );
  NAND U17796 ( .A(n16002), .B(n16001), .Z(n16003) );
  NAND U17797 ( .A(n16004), .B(n16003), .Z(n16038) );
  XNOR U17798 ( .A(n16039), .B(n16038), .Z(c[1338]) );
  NANDN U17799 ( .A(n16006), .B(n16005), .Z(n16010) );
  NANDN U17800 ( .A(n16008), .B(n16007), .Z(n16009) );
  AND U17801 ( .A(n16010), .B(n16009), .Z(n16045) );
  NANDN U17802 ( .A(n16012), .B(n16011), .Z(n16016) );
  NANDN U17803 ( .A(n16014), .B(n16013), .Z(n16015) );
  AND U17804 ( .A(n16016), .B(n16015), .Z(n16043) );
  NAND U17805 ( .A(n42143), .B(n16017), .Z(n16019) );
  XNOR U17806 ( .A(a[317]), .B(n4117), .Z(n16054) );
  NAND U17807 ( .A(n42144), .B(n16054), .Z(n16018) );
  AND U17808 ( .A(n16019), .B(n16018), .Z(n16069) );
  XOR U17809 ( .A(a[321]), .B(n42012), .Z(n16057) );
  XNOR U17810 ( .A(n16069), .B(n16068), .Z(n16071) );
  AND U17811 ( .A(a[323]), .B(b[0]), .Z(n16021) );
  XNOR U17812 ( .A(n16021), .B(n4071), .Z(n16023) );
  NANDN U17813 ( .A(b[0]), .B(a[322]), .Z(n16022) );
  NAND U17814 ( .A(n16023), .B(n16022), .Z(n16065) );
  XOR U17815 ( .A(a[319]), .B(n42085), .Z(n16058) );
  AND U17816 ( .A(a[315]), .B(b[7]), .Z(n16062) );
  XNOR U17817 ( .A(n16063), .B(n16062), .Z(n16064) );
  XNOR U17818 ( .A(n16065), .B(n16064), .Z(n16070) );
  XOR U17819 ( .A(n16071), .B(n16070), .Z(n16049) );
  NANDN U17820 ( .A(n16026), .B(n16025), .Z(n16030) );
  NANDN U17821 ( .A(n16028), .B(n16027), .Z(n16029) );
  AND U17822 ( .A(n16030), .B(n16029), .Z(n16048) );
  XNOR U17823 ( .A(n16049), .B(n16048), .Z(n16050) );
  NANDN U17824 ( .A(n16032), .B(n16031), .Z(n16036) );
  NAND U17825 ( .A(n16034), .B(n16033), .Z(n16035) );
  NAND U17826 ( .A(n16036), .B(n16035), .Z(n16051) );
  XNOR U17827 ( .A(n16050), .B(n16051), .Z(n16042) );
  XNOR U17828 ( .A(n16043), .B(n16042), .Z(n16044) );
  XNOR U17829 ( .A(n16045), .B(n16044), .Z(n16074) );
  XNOR U17830 ( .A(sreg[1339]), .B(n16074), .Z(n16076) );
  NANDN U17831 ( .A(sreg[1338]), .B(n16037), .Z(n16041) );
  NAND U17832 ( .A(n16039), .B(n16038), .Z(n16040) );
  NAND U17833 ( .A(n16041), .B(n16040), .Z(n16075) );
  XNOR U17834 ( .A(n16076), .B(n16075), .Z(c[1339]) );
  NANDN U17835 ( .A(n16043), .B(n16042), .Z(n16047) );
  NANDN U17836 ( .A(n16045), .B(n16044), .Z(n16046) );
  AND U17837 ( .A(n16047), .B(n16046), .Z(n16082) );
  NANDN U17838 ( .A(n16049), .B(n16048), .Z(n16053) );
  NANDN U17839 ( .A(n16051), .B(n16050), .Z(n16052) );
  AND U17840 ( .A(n16053), .B(n16052), .Z(n16080) );
  NAND U17841 ( .A(n42143), .B(n16054), .Z(n16056) );
  XNOR U17842 ( .A(a[318]), .B(n4117), .Z(n16091) );
  NAND U17843 ( .A(n42144), .B(n16091), .Z(n16055) );
  AND U17844 ( .A(n16056), .B(n16055), .Z(n16106) );
  XOR U17845 ( .A(a[322]), .B(n42012), .Z(n16094) );
  XNOR U17846 ( .A(n16106), .B(n16105), .Z(n16108) );
  XOR U17847 ( .A(a[320]), .B(n42085), .Z(n16098) );
  AND U17848 ( .A(a[316]), .B(b[7]), .Z(n16099) );
  XNOR U17849 ( .A(n16100), .B(n16099), .Z(n16101) );
  AND U17850 ( .A(a[324]), .B(b[0]), .Z(n16059) );
  XNOR U17851 ( .A(n16059), .B(n4071), .Z(n16061) );
  NANDN U17852 ( .A(b[0]), .B(a[323]), .Z(n16060) );
  NAND U17853 ( .A(n16061), .B(n16060), .Z(n16102) );
  XNOR U17854 ( .A(n16101), .B(n16102), .Z(n16107) );
  XOR U17855 ( .A(n16108), .B(n16107), .Z(n16086) );
  NANDN U17856 ( .A(n16063), .B(n16062), .Z(n16067) );
  NANDN U17857 ( .A(n16065), .B(n16064), .Z(n16066) );
  AND U17858 ( .A(n16067), .B(n16066), .Z(n16085) );
  XNOR U17859 ( .A(n16086), .B(n16085), .Z(n16087) );
  NANDN U17860 ( .A(n16069), .B(n16068), .Z(n16073) );
  NAND U17861 ( .A(n16071), .B(n16070), .Z(n16072) );
  NAND U17862 ( .A(n16073), .B(n16072), .Z(n16088) );
  XNOR U17863 ( .A(n16087), .B(n16088), .Z(n16079) );
  XNOR U17864 ( .A(n16080), .B(n16079), .Z(n16081) );
  XNOR U17865 ( .A(n16082), .B(n16081), .Z(n16111) );
  XNOR U17866 ( .A(sreg[1340]), .B(n16111), .Z(n16113) );
  NANDN U17867 ( .A(sreg[1339]), .B(n16074), .Z(n16078) );
  NAND U17868 ( .A(n16076), .B(n16075), .Z(n16077) );
  NAND U17869 ( .A(n16078), .B(n16077), .Z(n16112) );
  XNOR U17870 ( .A(n16113), .B(n16112), .Z(c[1340]) );
  NANDN U17871 ( .A(n16080), .B(n16079), .Z(n16084) );
  NANDN U17872 ( .A(n16082), .B(n16081), .Z(n16083) );
  AND U17873 ( .A(n16084), .B(n16083), .Z(n16119) );
  NANDN U17874 ( .A(n16086), .B(n16085), .Z(n16090) );
  NANDN U17875 ( .A(n16088), .B(n16087), .Z(n16089) );
  AND U17876 ( .A(n16090), .B(n16089), .Z(n16117) );
  NAND U17877 ( .A(n42143), .B(n16091), .Z(n16093) );
  XNOR U17878 ( .A(a[319]), .B(n4117), .Z(n16128) );
  NAND U17879 ( .A(n42144), .B(n16128), .Z(n16092) );
  AND U17880 ( .A(n16093), .B(n16092), .Z(n16143) );
  XOR U17881 ( .A(a[323]), .B(n42012), .Z(n16131) );
  XNOR U17882 ( .A(n16143), .B(n16142), .Z(n16145) );
  NAND U17883 ( .A(a[325]), .B(b[0]), .Z(n16095) );
  XNOR U17884 ( .A(b[1]), .B(n16095), .Z(n16097) );
  NANDN U17885 ( .A(b[0]), .B(a[324]), .Z(n16096) );
  AND U17886 ( .A(n16097), .B(n16096), .Z(n16138) );
  XOR U17887 ( .A(a[321]), .B(n42085), .Z(n16135) );
  AND U17888 ( .A(a[317]), .B(b[7]), .Z(n16136) );
  XOR U17889 ( .A(n16137), .B(n16136), .Z(n16139) );
  XNOR U17890 ( .A(n16138), .B(n16139), .Z(n16144) );
  XOR U17891 ( .A(n16145), .B(n16144), .Z(n16123) );
  NANDN U17892 ( .A(n16100), .B(n16099), .Z(n16104) );
  NANDN U17893 ( .A(n16102), .B(n16101), .Z(n16103) );
  AND U17894 ( .A(n16104), .B(n16103), .Z(n16122) );
  XNOR U17895 ( .A(n16123), .B(n16122), .Z(n16124) );
  NANDN U17896 ( .A(n16106), .B(n16105), .Z(n16110) );
  NAND U17897 ( .A(n16108), .B(n16107), .Z(n16109) );
  NAND U17898 ( .A(n16110), .B(n16109), .Z(n16125) );
  XNOR U17899 ( .A(n16124), .B(n16125), .Z(n16116) );
  XNOR U17900 ( .A(n16117), .B(n16116), .Z(n16118) );
  XNOR U17901 ( .A(n16119), .B(n16118), .Z(n16148) );
  XNOR U17902 ( .A(sreg[1341]), .B(n16148), .Z(n16150) );
  NANDN U17903 ( .A(sreg[1340]), .B(n16111), .Z(n16115) );
  NAND U17904 ( .A(n16113), .B(n16112), .Z(n16114) );
  NAND U17905 ( .A(n16115), .B(n16114), .Z(n16149) );
  XNOR U17906 ( .A(n16150), .B(n16149), .Z(c[1341]) );
  NANDN U17907 ( .A(n16117), .B(n16116), .Z(n16121) );
  NANDN U17908 ( .A(n16119), .B(n16118), .Z(n16120) );
  AND U17909 ( .A(n16121), .B(n16120), .Z(n16156) );
  NANDN U17910 ( .A(n16123), .B(n16122), .Z(n16127) );
  NANDN U17911 ( .A(n16125), .B(n16124), .Z(n16126) );
  AND U17912 ( .A(n16127), .B(n16126), .Z(n16154) );
  NAND U17913 ( .A(n42143), .B(n16128), .Z(n16130) );
  XNOR U17914 ( .A(a[320]), .B(n4117), .Z(n16165) );
  NAND U17915 ( .A(n42144), .B(n16165), .Z(n16129) );
  AND U17916 ( .A(n16130), .B(n16129), .Z(n16180) );
  XOR U17917 ( .A(a[324]), .B(n42012), .Z(n16168) );
  XNOR U17918 ( .A(n16180), .B(n16179), .Z(n16182) );
  AND U17919 ( .A(a[326]), .B(b[0]), .Z(n16132) );
  XNOR U17920 ( .A(n16132), .B(n4071), .Z(n16134) );
  NANDN U17921 ( .A(b[0]), .B(a[325]), .Z(n16133) );
  NAND U17922 ( .A(n16134), .B(n16133), .Z(n16176) );
  XOR U17923 ( .A(a[322]), .B(n42085), .Z(n16172) );
  AND U17924 ( .A(a[318]), .B(b[7]), .Z(n16173) );
  XNOR U17925 ( .A(n16174), .B(n16173), .Z(n16175) );
  XNOR U17926 ( .A(n16176), .B(n16175), .Z(n16181) );
  XOR U17927 ( .A(n16182), .B(n16181), .Z(n16160) );
  NANDN U17928 ( .A(n16137), .B(n16136), .Z(n16141) );
  NANDN U17929 ( .A(n16139), .B(n16138), .Z(n16140) );
  AND U17930 ( .A(n16141), .B(n16140), .Z(n16159) );
  XNOR U17931 ( .A(n16160), .B(n16159), .Z(n16161) );
  NANDN U17932 ( .A(n16143), .B(n16142), .Z(n16147) );
  NAND U17933 ( .A(n16145), .B(n16144), .Z(n16146) );
  NAND U17934 ( .A(n16147), .B(n16146), .Z(n16162) );
  XNOR U17935 ( .A(n16161), .B(n16162), .Z(n16153) );
  XNOR U17936 ( .A(n16154), .B(n16153), .Z(n16155) );
  XNOR U17937 ( .A(n16156), .B(n16155), .Z(n16185) );
  XNOR U17938 ( .A(sreg[1342]), .B(n16185), .Z(n16187) );
  NANDN U17939 ( .A(sreg[1341]), .B(n16148), .Z(n16152) );
  NAND U17940 ( .A(n16150), .B(n16149), .Z(n16151) );
  NAND U17941 ( .A(n16152), .B(n16151), .Z(n16186) );
  XNOR U17942 ( .A(n16187), .B(n16186), .Z(c[1342]) );
  NANDN U17943 ( .A(n16154), .B(n16153), .Z(n16158) );
  NANDN U17944 ( .A(n16156), .B(n16155), .Z(n16157) );
  AND U17945 ( .A(n16158), .B(n16157), .Z(n16193) );
  NANDN U17946 ( .A(n16160), .B(n16159), .Z(n16164) );
  NANDN U17947 ( .A(n16162), .B(n16161), .Z(n16163) );
  AND U17948 ( .A(n16164), .B(n16163), .Z(n16191) );
  NAND U17949 ( .A(n42143), .B(n16165), .Z(n16167) );
  XNOR U17950 ( .A(a[321]), .B(n4117), .Z(n16202) );
  NAND U17951 ( .A(n42144), .B(n16202), .Z(n16166) );
  AND U17952 ( .A(n16167), .B(n16166), .Z(n16217) );
  XOR U17953 ( .A(a[325]), .B(n42012), .Z(n16205) );
  XNOR U17954 ( .A(n16217), .B(n16216), .Z(n16219) );
  AND U17955 ( .A(a[327]), .B(b[0]), .Z(n16169) );
  XNOR U17956 ( .A(n16169), .B(n4071), .Z(n16171) );
  NANDN U17957 ( .A(b[0]), .B(a[326]), .Z(n16170) );
  NAND U17958 ( .A(n16171), .B(n16170), .Z(n16213) );
  XOR U17959 ( .A(a[323]), .B(n42085), .Z(n16209) );
  AND U17960 ( .A(a[319]), .B(b[7]), .Z(n16210) );
  XNOR U17961 ( .A(n16211), .B(n16210), .Z(n16212) );
  XNOR U17962 ( .A(n16213), .B(n16212), .Z(n16218) );
  XOR U17963 ( .A(n16219), .B(n16218), .Z(n16197) );
  NANDN U17964 ( .A(n16174), .B(n16173), .Z(n16178) );
  NANDN U17965 ( .A(n16176), .B(n16175), .Z(n16177) );
  AND U17966 ( .A(n16178), .B(n16177), .Z(n16196) );
  XNOR U17967 ( .A(n16197), .B(n16196), .Z(n16198) );
  NANDN U17968 ( .A(n16180), .B(n16179), .Z(n16184) );
  NAND U17969 ( .A(n16182), .B(n16181), .Z(n16183) );
  NAND U17970 ( .A(n16184), .B(n16183), .Z(n16199) );
  XNOR U17971 ( .A(n16198), .B(n16199), .Z(n16190) );
  XNOR U17972 ( .A(n16191), .B(n16190), .Z(n16192) );
  XNOR U17973 ( .A(n16193), .B(n16192), .Z(n16222) );
  XNOR U17974 ( .A(sreg[1343]), .B(n16222), .Z(n16224) );
  NANDN U17975 ( .A(sreg[1342]), .B(n16185), .Z(n16189) );
  NAND U17976 ( .A(n16187), .B(n16186), .Z(n16188) );
  NAND U17977 ( .A(n16189), .B(n16188), .Z(n16223) );
  XNOR U17978 ( .A(n16224), .B(n16223), .Z(c[1343]) );
  NANDN U17979 ( .A(n16191), .B(n16190), .Z(n16195) );
  NANDN U17980 ( .A(n16193), .B(n16192), .Z(n16194) );
  AND U17981 ( .A(n16195), .B(n16194), .Z(n16230) );
  NANDN U17982 ( .A(n16197), .B(n16196), .Z(n16201) );
  NANDN U17983 ( .A(n16199), .B(n16198), .Z(n16200) );
  AND U17984 ( .A(n16201), .B(n16200), .Z(n16228) );
  NAND U17985 ( .A(n42143), .B(n16202), .Z(n16204) );
  XNOR U17986 ( .A(a[322]), .B(n4117), .Z(n16239) );
  NAND U17987 ( .A(n42144), .B(n16239), .Z(n16203) );
  AND U17988 ( .A(n16204), .B(n16203), .Z(n16254) );
  XOR U17989 ( .A(a[326]), .B(n42012), .Z(n16242) );
  XNOR U17990 ( .A(n16254), .B(n16253), .Z(n16256) );
  AND U17991 ( .A(a[328]), .B(b[0]), .Z(n16206) );
  XNOR U17992 ( .A(n16206), .B(n4071), .Z(n16208) );
  NANDN U17993 ( .A(b[0]), .B(a[327]), .Z(n16207) );
  NAND U17994 ( .A(n16208), .B(n16207), .Z(n16250) );
  XOR U17995 ( .A(a[324]), .B(n42085), .Z(n16243) );
  AND U17996 ( .A(a[320]), .B(b[7]), .Z(n16247) );
  XNOR U17997 ( .A(n16248), .B(n16247), .Z(n16249) );
  XNOR U17998 ( .A(n16250), .B(n16249), .Z(n16255) );
  XOR U17999 ( .A(n16256), .B(n16255), .Z(n16234) );
  NANDN U18000 ( .A(n16211), .B(n16210), .Z(n16215) );
  NANDN U18001 ( .A(n16213), .B(n16212), .Z(n16214) );
  AND U18002 ( .A(n16215), .B(n16214), .Z(n16233) );
  XNOR U18003 ( .A(n16234), .B(n16233), .Z(n16235) );
  NANDN U18004 ( .A(n16217), .B(n16216), .Z(n16221) );
  NAND U18005 ( .A(n16219), .B(n16218), .Z(n16220) );
  NAND U18006 ( .A(n16221), .B(n16220), .Z(n16236) );
  XNOR U18007 ( .A(n16235), .B(n16236), .Z(n16227) );
  XNOR U18008 ( .A(n16228), .B(n16227), .Z(n16229) );
  XNOR U18009 ( .A(n16230), .B(n16229), .Z(n16259) );
  XNOR U18010 ( .A(sreg[1344]), .B(n16259), .Z(n16261) );
  NANDN U18011 ( .A(sreg[1343]), .B(n16222), .Z(n16226) );
  NAND U18012 ( .A(n16224), .B(n16223), .Z(n16225) );
  NAND U18013 ( .A(n16226), .B(n16225), .Z(n16260) );
  XNOR U18014 ( .A(n16261), .B(n16260), .Z(c[1344]) );
  NANDN U18015 ( .A(n16228), .B(n16227), .Z(n16232) );
  NANDN U18016 ( .A(n16230), .B(n16229), .Z(n16231) );
  AND U18017 ( .A(n16232), .B(n16231), .Z(n16267) );
  NANDN U18018 ( .A(n16234), .B(n16233), .Z(n16238) );
  NANDN U18019 ( .A(n16236), .B(n16235), .Z(n16237) );
  AND U18020 ( .A(n16238), .B(n16237), .Z(n16265) );
  NAND U18021 ( .A(n42143), .B(n16239), .Z(n16241) );
  XNOR U18022 ( .A(a[323]), .B(n4118), .Z(n16276) );
  NAND U18023 ( .A(n42144), .B(n16276), .Z(n16240) );
  AND U18024 ( .A(n16241), .B(n16240), .Z(n16291) );
  XOR U18025 ( .A(a[327]), .B(n42012), .Z(n16279) );
  XNOR U18026 ( .A(n16291), .B(n16290), .Z(n16293) );
  XOR U18027 ( .A(a[325]), .B(n42085), .Z(n16283) );
  AND U18028 ( .A(a[321]), .B(b[7]), .Z(n16284) );
  XNOR U18029 ( .A(n16285), .B(n16284), .Z(n16286) );
  AND U18030 ( .A(a[329]), .B(b[0]), .Z(n16244) );
  XNOR U18031 ( .A(n16244), .B(n4071), .Z(n16246) );
  NANDN U18032 ( .A(b[0]), .B(a[328]), .Z(n16245) );
  NAND U18033 ( .A(n16246), .B(n16245), .Z(n16287) );
  XNOR U18034 ( .A(n16286), .B(n16287), .Z(n16292) );
  XOR U18035 ( .A(n16293), .B(n16292), .Z(n16271) );
  NANDN U18036 ( .A(n16248), .B(n16247), .Z(n16252) );
  NANDN U18037 ( .A(n16250), .B(n16249), .Z(n16251) );
  AND U18038 ( .A(n16252), .B(n16251), .Z(n16270) );
  XNOR U18039 ( .A(n16271), .B(n16270), .Z(n16272) );
  NANDN U18040 ( .A(n16254), .B(n16253), .Z(n16258) );
  NAND U18041 ( .A(n16256), .B(n16255), .Z(n16257) );
  NAND U18042 ( .A(n16258), .B(n16257), .Z(n16273) );
  XNOR U18043 ( .A(n16272), .B(n16273), .Z(n16264) );
  XNOR U18044 ( .A(n16265), .B(n16264), .Z(n16266) );
  XNOR U18045 ( .A(n16267), .B(n16266), .Z(n16296) );
  XNOR U18046 ( .A(sreg[1345]), .B(n16296), .Z(n16298) );
  NANDN U18047 ( .A(sreg[1344]), .B(n16259), .Z(n16263) );
  NAND U18048 ( .A(n16261), .B(n16260), .Z(n16262) );
  NAND U18049 ( .A(n16263), .B(n16262), .Z(n16297) );
  XNOR U18050 ( .A(n16298), .B(n16297), .Z(c[1345]) );
  NANDN U18051 ( .A(n16265), .B(n16264), .Z(n16269) );
  NANDN U18052 ( .A(n16267), .B(n16266), .Z(n16268) );
  AND U18053 ( .A(n16269), .B(n16268), .Z(n16304) );
  NANDN U18054 ( .A(n16271), .B(n16270), .Z(n16275) );
  NANDN U18055 ( .A(n16273), .B(n16272), .Z(n16274) );
  AND U18056 ( .A(n16275), .B(n16274), .Z(n16302) );
  NAND U18057 ( .A(n42143), .B(n16276), .Z(n16278) );
  XNOR U18058 ( .A(a[324]), .B(n4118), .Z(n16313) );
  NAND U18059 ( .A(n42144), .B(n16313), .Z(n16277) );
  AND U18060 ( .A(n16278), .B(n16277), .Z(n16328) );
  XOR U18061 ( .A(a[328]), .B(n42012), .Z(n16316) );
  XNOR U18062 ( .A(n16328), .B(n16327), .Z(n16330) );
  AND U18063 ( .A(a[330]), .B(b[0]), .Z(n16280) );
  XNOR U18064 ( .A(n16280), .B(n4071), .Z(n16282) );
  NANDN U18065 ( .A(b[0]), .B(a[329]), .Z(n16281) );
  NAND U18066 ( .A(n16282), .B(n16281), .Z(n16324) );
  XOR U18067 ( .A(a[326]), .B(n42085), .Z(n16320) );
  AND U18068 ( .A(a[322]), .B(b[7]), .Z(n16321) );
  XNOR U18069 ( .A(n16322), .B(n16321), .Z(n16323) );
  XNOR U18070 ( .A(n16324), .B(n16323), .Z(n16329) );
  XOR U18071 ( .A(n16330), .B(n16329), .Z(n16308) );
  NANDN U18072 ( .A(n16285), .B(n16284), .Z(n16289) );
  NANDN U18073 ( .A(n16287), .B(n16286), .Z(n16288) );
  AND U18074 ( .A(n16289), .B(n16288), .Z(n16307) );
  XNOR U18075 ( .A(n16308), .B(n16307), .Z(n16309) );
  NANDN U18076 ( .A(n16291), .B(n16290), .Z(n16295) );
  NAND U18077 ( .A(n16293), .B(n16292), .Z(n16294) );
  NAND U18078 ( .A(n16295), .B(n16294), .Z(n16310) );
  XNOR U18079 ( .A(n16309), .B(n16310), .Z(n16301) );
  XNOR U18080 ( .A(n16302), .B(n16301), .Z(n16303) );
  XNOR U18081 ( .A(n16304), .B(n16303), .Z(n16333) );
  XNOR U18082 ( .A(sreg[1346]), .B(n16333), .Z(n16335) );
  NANDN U18083 ( .A(sreg[1345]), .B(n16296), .Z(n16300) );
  NAND U18084 ( .A(n16298), .B(n16297), .Z(n16299) );
  NAND U18085 ( .A(n16300), .B(n16299), .Z(n16334) );
  XNOR U18086 ( .A(n16335), .B(n16334), .Z(c[1346]) );
  NANDN U18087 ( .A(n16302), .B(n16301), .Z(n16306) );
  NANDN U18088 ( .A(n16304), .B(n16303), .Z(n16305) );
  AND U18089 ( .A(n16306), .B(n16305), .Z(n16341) );
  NANDN U18090 ( .A(n16308), .B(n16307), .Z(n16312) );
  NANDN U18091 ( .A(n16310), .B(n16309), .Z(n16311) );
  AND U18092 ( .A(n16312), .B(n16311), .Z(n16339) );
  NAND U18093 ( .A(n42143), .B(n16313), .Z(n16315) );
  XNOR U18094 ( .A(a[325]), .B(n4118), .Z(n16350) );
  NAND U18095 ( .A(n42144), .B(n16350), .Z(n16314) );
  AND U18096 ( .A(n16315), .B(n16314), .Z(n16365) );
  XOR U18097 ( .A(a[329]), .B(n42012), .Z(n16353) );
  XNOR U18098 ( .A(n16365), .B(n16364), .Z(n16367) );
  AND U18099 ( .A(a[331]), .B(b[0]), .Z(n16317) );
  XNOR U18100 ( .A(n16317), .B(n4071), .Z(n16319) );
  NANDN U18101 ( .A(b[0]), .B(a[330]), .Z(n16318) );
  NAND U18102 ( .A(n16319), .B(n16318), .Z(n16361) );
  XOR U18103 ( .A(a[327]), .B(n42085), .Z(n16357) );
  AND U18104 ( .A(a[323]), .B(b[7]), .Z(n16358) );
  XNOR U18105 ( .A(n16359), .B(n16358), .Z(n16360) );
  XNOR U18106 ( .A(n16361), .B(n16360), .Z(n16366) );
  XOR U18107 ( .A(n16367), .B(n16366), .Z(n16345) );
  NANDN U18108 ( .A(n16322), .B(n16321), .Z(n16326) );
  NANDN U18109 ( .A(n16324), .B(n16323), .Z(n16325) );
  AND U18110 ( .A(n16326), .B(n16325), .Z(n16344) );
  XNOR U18111 ( .A(n16345), .B(n16344), .Z(n16346) );
  NANDN U18112 ( .A(n16328), .B(n16327), .Z(n16332) );
  NAND U18113 ( .A(n16330), .B(n16329), .Z(n16331) );
  NAND U18114 ( .A(n16332), .B(n16331), .Z(n16347) );
  XNOR U18115 ( .A(n16346), .B(n16347), .Z(n16338) );
  XNOR U18116 ( .A(n16339), .B(n16338), .Z(n16340) );
  XNOR U18117 ( .A(n16341), .B(n16340), .Z(n16370) );
  XNOR U18118 ( .A(sreg[1347]), .B(n16370), .Z(n16372) );
  NANDN U18119 ( .A(sreg[1346]), .B(n16333), .Z(n16337) );
  NAND U18120 ( .A(n16335), .B(n16334), .Z(n16336) );
  NAND U18121 ( .A(n16337), .B(n16336), .Z(n16371) );
  XNOR U18122 ( .A(n16372), .B(n16371), .Z(c[1347]) );
  NANDN U18123 ( .A(n16339), .B(n16338), .Z(n16343) );
  NANDN U18124 ( .A(n16341), .B(n16340), .Z(n16342) );
  AND U18125 ( .A(n16343), .B(n16342), .Z(n16378) );
  NANDN U18126 ( .A(n16345), .B(n16344), .Z(n16349) );
  NANDN U18127 ( .A(n16347), .B(n16346), .Z(n16348) );
  AND U18128 ( .A(n16349), .B(n16348), .Z(n16376) );
  NAND U18129 ( .A(n42143), .B(n16350), .Z(n16352) );
  XNOR U18130 ( .A(a[326]), .B(n4118), .Z(n16387) );
  NAND U18131 ( .A(n42144), .B(n16387), .Z(n16351) );
  AND U18132 ( .A(n16352), .B(n16351), .Z(n16402) );
  XOR U18133 ( .A(a[330]), .B(n42012), .Z(n16390) );
  XNOR U18134 ( .A(n16402), .B(n16401), .Z(n16404) );
  AND U18135 ( .A(a[332]), .B(b[0]), .Z(n16354) );
  XNOR U18136 ( .A(n16354), .B(n4071), .Z(n16356) );
  NANDN U18137 ( .A(b[0]), .B(a[331]), .Z(n16355) );
  NAND U18138 ( .A(n16356), .B(n16355), .Z(n16398) );
  XOR U18139 ( .A(a[328]), .B(n42085), .Z(n16391) );
  AND U18140 ( .A(a[324]), .B(b[7]), .Z(n16395) );
  XNOR U18141 ( .A(n16396), .B(n16395), .Z(n16397) );
  XNOR U18142 ( .A(n16398), .B(n16397), .Z(n16403) );
  XOR U18143 ( .A(n16404), .B(n16403), .Z(n16382) );
  NANDN U18144 ( .A(n16359), .B(n16358), .Z(n16363) );
  NANDN U18145 ( .A(n16361), .B(n16360), .Z(n16362) );
  AND U18146 ( .A(n16363), .B(n16362), .Z(n16381) );
  XNOR U18147 ( .A(n16382), .B(n16381), .Z(n16383) );
  NANDN U18148 ( .A(n16365), .B(n16364), .Z(n16369) );
  NAND U18149 ( .A(n16367), .B(n16366), .Z(n16368) );
  NAND U18150 ( .A(n16369), .B(n16368), .Z(n16384) );
  XNOR U18151 ( .A(n16383), .B(n16384), .Z(n16375) );
  XNOR U18152 ( .A(n16376), .B(n16375), .Z(n16377) );
  XNOR U18153 ( .A(n16378), .B(n16377), .Z(n16407) );
  XNOR U18154 ( .A(sreg[1348]), .B(n16407), .Z(n16409) );
  NANDN U18155 ( .A(sreg[1347]), .B(n16370), .Z(n16374) );
  NAND U18156 ( .A(n16372), .B(n16371), .Z(n16373) );
  NAND U18157 ( .A(n16374), .B(n16373), .Z(n16408) );
  XNOR U18158 ( .A(n16409), .B(n16408), .Z(c[1348]) );
  NANDN U18159 ( .A(n16376), .B(n16375), .Z(n16380) );
  NANDN U18160 ( .A(n16378), .B(n16377), .Z(n16379) );
  AND U18161 ( .A(n16380), .B(n16379), .Z(n16415) );
  NANDN U18162 ( .A(n16382), .B(n16381), .Z(n16386) );
  NANDN U18163 ( .A(n16384), .B(n16383), .Z(n16385) );
  AND U18164 ( .A(n16386), .B(n16385), .Z(n16413) );
  NAND U18165 ( .A(n42143), .B(n16387), .Z(n16389) );
  XNOR U18166 ( .A(a[327]), .B(n4118), .Z(n16424) );
  NAND U18167 ( .A(n42144), .B(n16424), .Z(n16388) );
  AND U18168 ( .A(n16389), .B(n16388), .Z(n16439) );
  XOR U18169 ( .A(a[331]), .B(n42012), .Z(n16427) );
  XNOR U18170 ( .A(n16439), .B(n16438), .Z(n16441) );
  XOR U18171 ( .A(a[329]), .B(n42085), .Z(n16431) );
  AND U18172 ( .A(a[325]), .B(b[7]), .Z(n16432) );
  XNOR U18173 ( .A(n16433), .B(n16432), .Z(n16434) );
  AND U18174 ( .A(a[333]), .B(b[0]), .Z(n16392) );
  XNOR U18175 ( .A(n16392), .B(n4071), .Z(n16394) );
  NANDN U18176 ( .A(b[0]), .B(a[332]), .Z(n16393) );
  NAND U18177 ( .A(n16394), .B(n16393), .Z(n16435) );
  XNOR U18178 ( .A(n16434), .B(n16435), .Z(n16440) );
  XOR U18179 ( .A(n16441), .B(n16440), .Z(n16419) );
  NANDN U18180 ( .A(n16396), .B(n16395), .Z(n16400) );
  NANDN U18181 ( .A(n16398), .B(n16397), .Z(n16399) );
  AND U18182 ( .A(n16400), .B(n16399), .Z(n16418) );
  XNOR U18183 ( .A(n16419), .B(n16418), .Z(n16420) );
  NANDN U18184 ( .A(n16402), .B(n16401), .Z(n16406) );
  NAND U18185 ( .A(n16404), .B(n16403), .Z(n16405) );
  NAND U18186 ( .A(n16406), .B(n16405), .Z(n16421) );
  XNOR U18187 ( .A(n16420), .B(n16421), .Z(n16412) );
  XNOR U18188 ( .A(n16413), .B(n16412), .Z(n16414) );
  XNOR U18189 ( .A(n16415), .B(n16414), .Z(n16444) );
  XNOR U18190 ( .A(sreg[1349]), .B(n16444), .Z(n16446) );
  NANDN U18191 ( .A(sreg[1348]), .B(n16407), .Z(n16411) );
  NAND U18192 ( .A(n16409), .B(n16408), .Z(n16410) );
  NAND U18193 ( .A(n16411), .B(n16410), .Z(n16445) );
  XNOR U18194 ( .A(n16446), .B(n16445), .Z(c[1349]) );
  NANDN U18195 ( .A(n16413), .B(n16412), .Z(n16417) );
  NANDN U18196 ( .A(n16415), .B(n16414), .Z(n16416) );
  AND U18197 ( .A(n16417), .B(n16416), .Z(n16452) );
  NANDN U18198 ( .A(n16419), .B(n16418), .Z(n16423) );
  NANDN U18199 ( .A(n16421), .B(n16420), .Z(n16422) );
  AND U18200 ( .A(n16423), .B(n16422), .Z(n16450) );
  NAND U18201 ( .A(n42143), .B(n16424), .Z(n16426) );
  XNOR U18202 ( .A(a[328]), .B(n4118), .Z(n16461) );
  NAND U18203 ( .A(n42144), .B(n16461), .Z(n16425) );
  AND U18204 ( .A(n16426), .B(n16425), .Z(n16476) );
  XOR U18205 ( .A(a[332]), .B(n42012), .Z(n16464) );
  XNOR U18206 ( .A(n16476), .B(n16475), .Z(n16478) );
  AND U18207 ( .A(a[334]), .B(b[0]), .Z(n16428) );
  XNOR U18208 ( .A(n16428), .B(n4071), .Z(n16430) );
  NANDN U18209 ( .A(b[0]), .B(a[333]), .Z(n16429) );
  NAND U18210 ( .A(n16430), .B(n16429), .Z(n16472) );
  XOR U18211 ( .A(a[330]), .B(n42085), .Z(n16465) );
  AND U18212 ( .A(a[326]), .B(b[7]), .Z(n16469) );
  XNOR U18213 ( .A(n16470), .B(n16469), .Z(n16471) );
  XNOR U18214 ( .A(n16472), .B(n16471), .Z(n16477) );
  XOR U18215 ( .A(n16478), .B(n16477), .Z(n16456) );
  NANDN U18216 ( .A(n16433), .B(n16432), .Z(n16437) );
  NANDN U18217 ( .A(n16435), .B(n16434), .Z(n16436) );
  AND U18218 ( .A(n16437), .B(n16436), .Z(n16455) );
  XNOR U18219 ( .A(n16456), .B(n16455), .Z(n16457) );
  NANDN U18220 ( .A(n16439), .B(n16438), .Z(n16443) );
  NAND U18221 ( .A(n16441), .B(n16440), .Z(n16442) );
  NAND U18222 ( .A(n16443), .B(n16442), .Z(n16458) );
  XNOR U18223 ( .A(n16457), .B(n16458), .Z(n16449) );
  XNOR U18224 ( .A(n16450), .B(n16449), .Z(n16451) );
  XNOR U18225 ( .A(n16452), .B(n16451), .Z(n16481) );
  XNOR U18226 ( .A(sreg[1350]), .B(n16481), .Z(n16483) );
  NANDN U18227 ( .A(sreg[1349]), .B(n16444), .Z(n16448) );
  NAND U18228 ( .A(n16446), .B(n16445), .Z(n16447) );
  NAND U18229 ( .A(n16448), .B(n16447), .Z(n16482) );
  XNOR U18230 ( .A(n16483), .B(n16482), .Z(c[1350]) );
  NANDN U18231 ( .A(n16450), .B(n16449), .Z(n16454) );
  NANDN U18232 ( .A(n16452), .B(n16451), .Z(n16453) );
  AND U18233 ( .A(n16454), .B(n16453), .Z(n16489) );
  NANDN U18234 ( .A(n16456), .B(n16455), .Z(n16460) );
  NANDN U18235 ( .A(n16458), .B(n16457), .Z(n16459) );
  AND U18236 ( .A(n16460), .B(n16459), .Z(n16487) );
  NAND U18237 ( .A(n42143), .B(n16461), .Z(n16463) );
  XNOR U18238 ( .A(a[329]), .B(n4118), .Z(n16498) );
  NAND U18239 ( .A(n42144), .B(n16498), .Z(n16462) );
  AND U18240 ( .A(n16463), .B(n16462), .Z(n16513) );
  XOR U18241 ( .A(a[333]), .B(n42012), .Z(n16501) );
  XNOR U18242 ( .A(n16513), .B(n16512), .Z(n16515) );
  XOR U18243 ( .A(a[331]), .B(n42085), .Z(n16505) );
  AND U18244 ( .A(a[327]), .B(b[7]), .Z(n16506) );
  XNOR U18245 ( .A(n16507), .B(n16506), .Z(n16508) );
  AND U18246 ( .A(a[335]), .B(b[0]), .Z(n16466) );
  XNOR U18247 ( .A(n16466), .B(n4071), .Z(n16468) );
  NANDN U18248 ( .A(b[0]), .B(a[334]), .Z(n16467) );
  NAND U18249 ( .A(n16468), .B(n16467), .Z(n16509) );
  XNOR U18250 ( .A(n16508), .B(n16509), .Z(n16514) );
  XOR U18251 ( .A(n16515), .B(n16514), .Z(n16493) );
  NANDN U18252 ( .A(n16470), .B(n16469), .Z(n16474) );
  NANDN U18253 ( .A(n16472), .B(n16471), .Z(n16473) );
  AND U18254 ( .A(n16474), .B(n16473), .Z(n16492) );
  XNOR U18255 ( .A(n16493), .B(n16492), .Z(n16494) );
  NANDN U18256 ( .A(n16476), .B(n16475), .Z(n16480) );
  NAND U18257 ( .A(n16478), .B(n16477), .Z(n16479) );
  NAND U18258 ( .A(n16480), .B(n16479), .Z(n16495) );
  XNOR U18259 ( .A(n16494), .B(n16495), .Z(n16486) );
  XNOR U18260 ( .A(n16487), .B(n16486), .Z(n16488) );
  XNOR U18261 ( .A(n16489), .B(n16488), .Z(n16518) );
  XNOR U18262 ( .A(sreg[1351]), .B(n16518), .Z(n16520) );
  NANDN U18263 ( .A(sreg[1350]), .B(n16481), .Z(n16485) );
  NAND U18264 ( .A(n16483), .B(n16482), .Z(n16484) );
  NAND U18265 ( .A(n16485), .B(n16484), .Z(n16519) );
  XNOR U18266 ( .A(n16520), .B(n16519), .Z(c[1351]) );
  NANDN U18267 ( .A(n16487), .B(n16486), .Z(n16491) );
  NANDN U18268 ( .A(n16489), .B(n16488), .Z(n16490) );
  AND U18269 ( .A(n16491), .B(n16490), .Z(n16526) );
  NANDN U18270 ( .A(n16493), .B(n16492), .Z(n16497) );
  NANDN U18271 ( .A(n16495), .B(n16494), .Z(n16496) );
  AND U18272 ( .A(n16497), .B(n16496), .Z(n16524) );
  NAND U18273 ( .A(n42143), .B(n16498), .Z(n16500) );
  XNOR U18274 ( .A(a[330]), .B(n4119), .Z(n16535) );
  NAND U18275 ( .A(n42144), .B(n16535), .Z(n16499) );
  AND U18276 ( .A(n16500), .B(n16499), .Z(n16550) );
  XOR U18277 ( .A(a[334]), .B(n42012), .Z(n16538) );
  XNOR U18278 ( .A(n16550), .B(n16549), .Z(n16552) );
  AND U18279 ( .A(a[336]), .B(b[0]), .Z(n16502) );
  XNOR U18280 ( .A(n16502), .B(n4071), .Z(n16504) );
  NANDN U18281 ( .A(b[0]), .B(a[335]), .Z(n16503) );
  NAND U18282 ( .A(n16504), .B(n16503), .Z(n16546) );
  XOR U18283 ( .A(a[332]), .B(n42085), .Z(n16539) );
  AND U18284 ( .A(a[328]), .B(b[7]), .Z(n16543) );
  XNOR U18285 ( .A(n16544), .B(n16543), .Z(n16545) );
  XNOR U18286 ( .A(n16546), .B(n16545), .Z(n16551) );
  XOR U18287 ( .A(n16552), .B(n16551), .Z(n16530) );
  NANDN U18288 ( .A(n16507), .B(n16506), .Z(n16511) );
  NANDN U18289 ( .A(n16509), .B(n16508), .Z(n16510) );
  AND U18290 ( .A(n16511), .B(n16510), .Z(n16529) );
  XNOR U18291 ( .A(n16530), .B(n16529), .Z(n16531) );
  NANDN U18292 ( .A(n16513), .B(n16512), .Z(n16517) );
  NAND U18293 ( .A(n16515), .B(n16514), .Z(n16516) );
  NAND U18294 ( .A(n16517), .B(n16516), .Z(n16532) );
  XNOR U18295 ( .A(n16531), .B(n16532), .Z(n16523) );
  XNOR U18296 ( .A(n16524), .B(n16523), .Z(n16525) );
  XNOR U18297 ( .A(n16526), .B(n16525), .Z(n16555) );
  XNOR U18298 ( .A(sreg[1352]), .B(n16555), .Z(n16557) );
  NANDN U18299 ( .A(sreg[1351]), .B(n16518), .Z(n16522) );
  NAND U18300 ( .A(n16520), .B(n16519), .Z(n16521) );
  NAND U18301 ( .A(n16522), .B(n16521), .Z(n16556) );
  XNOR U18302 ( .A(n16557), .B(n16556), .Z(c[1352]) );
  NANDN U18303 ( .A(n16524), .B(n16523), .Z(n16528) );
  NANDN U18304 ( .A(n16526), .B(n16525), .Z(n16527) );
  AND U18305 ( .A(n16528), .B(n16527), .Z(n16563) );
  NANDN U18306 ( .A(n16530), .B(n16529), .Z(n16534) );
  NANDN U18307 ( .A(n16532), .B(n16531), .Z(n16533) );
  AND U18308 ( .A(n16534), .B(n16533), .Z(n16561) );
  NAND U18309 ( .A(n42143), .B(n16535), .Z(n16537) );
  XNOR U18310 ( .A(a[331]), .B(n4119), .Z(n16572) );
  NAND U18311 ( .A(n42144), .B(n16572), .Z(n16536) );
  AND U18312 ( .A(n16537), .B(n16536), .Z(n16587) );
  XOR U18313 ( .A(a[335]), .B(n42012), .Z(n16575) );
  XNOR U18314 ( .A(n16587), .B(n16586), .Z(n16589) );
  XOR U18315 ( .A(a[333]), .B(n42085), .Z(n16579) );
  AND U18316 ( .A(a[329]), .B(b[7]), .Z(n16580) );
  XNOR U18317 ( .A(n16581), .B(n16580), .Z(n16582) );
  AND U18318 ( .A(a[337]), .B(b[0]), .Z(n16540) );
  XNOR U18319 ( .A(n16540), .B(n4071), .Z(n16542) );
  NANDN U18320 ( .A(b[0]), .B(a[336]), .Z(n16541) );
  NAND U18321 ( .A(n16542), .B(n16541), .Z(n16583) );
  XNOR U18322 ( .A(n16582), .B(n16583), .Z(n16588) );
  XOR U18323 ( .A(n16589), .B(n16588), .Z(n16567) );
  NANDN U18324 ( .A(n16544), .B(n16543), .Z(n16548) );
  NANDN U18325 ( .A(n16546), .B(n16545), .Z(n16547) );
  AND U18326 ( .A(n16548), .B(n16547), .Z(n16566) );
  XNOR U18327 ( .A(n16567), .B(n16566), .Z(n16568) );
  NANDN U18328 ( .A(n16550), .B(n16549), .Z(n16554) );
  NAND U18329 ( .A(n16552), .B(n16551), .Z(n16553) );
  NAND U18330 ( .A(n16554), .B(n16553), .Z(n16569) );
  XNOR U18331 ( .A(n16568), .B(n16569), .Z(n16560) );
  XNOR U18332 ( .A(n16561), .B(n16560), .Z(n16562) );
  XNOR U18333 ( .A(n16563), .B(n16562), .Z(n16592) );
  XNOR U18334 ( .A(sreg[1353]), .B(n16592), .Z(n16594) );
  NANDN U18335 ( .A(sreg[1352]), .B(n16555), .Z(n16559) );
  NAND U18336 ( .A(n16557), .B(n16556), .Z(n16558) );
  NAND U18337 ( .A(n16559), .B(n16558), .Z(n16593) );
  XNOR U18338 ( .A(n16594), .B(n16593), .Z(c[1353]) );
  NANDN U18339 ( .A(n16561), .B(n16560), .Z(n16565) );
  NANDN U18340 ( .A(n16563), .B(n16562), .Z(n16564) );
  AND U18341 ( .A(n16565), .B(n16564), .Z(n16600) );
  NANDN U18342 ( .A(n16567), .B(n16566), .Z(n16571) );
  NANDN U18343 ( .A(n16569), .B(n16568), .Z(n16570) );
  AND U18344 ( .A(n16571), .B(n16570), .Z(n16598) );
  NAND U18345 ( .A(n42143), .B(n16572), .Z(n16574) );
  XNOR U18346 ( .A(a[332]), .B(n4119), .Z(n16609) );
  NAND U18347 ( .A(n42144), .B(n16609), .Z(n16573) );
  AND U18348 ( .A(n16574), .B(n16573), .Z(n16624) );
  XOR U18349 ( .A(a[336]), .B(n42012), .Z(n16612) );
  XNOR U18350 ( .A(n16624), .B(n16623), .Z(n16626) );
  AND U18351 ( .A(a[338]), .B(b[0]), .Z(n16576) );
  XNOR U18352 ( .A(n16576), .B(n4071), .Z(n16578) );
  NANDN U18353 ( .A(b[0]), .B(a[337]), .Z(n16577) );
  NAND U18354 ( .A(n16578), .B(n16577), .Z(n16620) );
  XOR U18355 ( .A(a[334]), .B(n42085), .Z(n16616) );
  AND U18356 ( .A(a[330]), .B(b[7]), .Z(n16617) );
  XNOR U18357 ( .A(n16618), .B(n16617), .Z(n16619) );
  XNOR U18358 ( .A(n16620), .B(n16619), .Z(n16625) );
  XOR U18359 ( .A(n16626), .B(n16625), .Z(n16604) );
  NANDN U18360 ( .A(n16581), .B(n16580), .Z(n16585) );
  NANDN U18361 ( .A(n16583), .B(n16582), .Z(n16584) );
  AND U18362 ( .A(n16585), .B(n16584), .Z(n16603) );
  XNOR U18363 ( .A(n16604), .B(n16603), .Z(n16605) );
  NANDN U18364 ( .A(n16587), .B(n16586), .Z(n16591) );
  NAND U18365 ( .A(n16589), .B(n16588), .Z(n16590) );
  NAND U18366 ( .A(n16591), .B(n16590), .Z(n16606) );
  XNOR U18367 ( .A(n16605), .B(n16606), .Z(n16597) );
  XNOR U18368 ( .A(n16598), .B(n16597), .Z(n16599) );
  XNOR U18369 ( .A(n16600), .B(n16599), .Z(n16629) );
  XNOR U18370 ( .A(sreg[1354]), .B(n16629), .Z(n16631) );
  NANDN U18371 ( .A(sreg[1353]), .B(n16592), .Z(n16596) );
  NAND U18372 ( .A(n16594), .B(n16593), .Z(n16595) );
  NAND U18373 ( .A(n16596), .B(n16595), .Z(n16630) );
  XNOR U18374 ( .A(n16631), .B(n16630), .Z(c[1354]) );
  NANDN U18375 ( .A(n16598), .B(n16597), .Z(n16602) );
  NANDN U18376 ( .A(n16600), .B(n16599), .Z(n16601) );
  AND U18377 ( .A(n16602), .B(n16601), .Z(n16637) );
  NANDN U18378 ( .A(n16604), .B(n16603), .Z(n16608) );
  NANDN U18379 ( .A(n16606), .B(n16605), .Z(n16607) );
  AND U18380 ( .A(n16608), .B(n16607), .Z(n16635) );
  NAND U18381 ( .A(n42143), .B(n16609), .Z(n16611) );
  XNOR U18382 ( .A(a[333]), .B(n4119), .Z(n16646) );
  NAND U18383 ( .A(n42144), .B(n16646), .Z(n16610) );
  AND U18384 ( .A(n16611), .B(n16610), .Z(n16661) );
  XOR U18385 ( .A(a[337]), .B(n42012), .Z(n16649) );
  XNOR U18386 ( .A(n16661), .B(n16660), .Z(n16663) );
  AND U18387 ( .A(a[339]), .B(b[0]), .Z(n16613) );
  XNOR U18388 ( .A(n16613), .B(n4071), .Z(n16615) );
  NANDN U18389 ( .A(b[0]), .B(a[338]), .Z(n16614) );
  NAND U18390 ( .A(n16615), .B(n16614), .Z(n16657) );
  XOR U18391 ( .A(a[335]), .B(n42085), .Z(n16653) );
  AND U18392 ( .A(a[331]), .B(b[7]), .Z(n16654) );
  XNOR U18393 ( .A(n16655), .B(n16654), .Z(n16656) );
  XNOR U18394 ( .A(n16657), .B(n16656), .Z(n16662) );
  XOR U18395 ( .A(n16663), .B(n16662), .Z(n16641) );
  NANDN U18396 ( .A(n16618), .B(n16617), .Z(n16622) );
  NANDN U18397 ( .A(n16620), .B(n16619), .Z(n16621) );
  AND U18398 ( .A(n16622), .B(n16621), .Z(n16640) );
  XNOR U18399 ( .A(n16641), .B(n16640), .Z(n16642) );
  NANDN U18400 ( .A(n16624), .B(n16623), .Z(n16628) );
  NAND U18401 ( .A(n16626), .B(n16625), .Z(n16627) );
  NAND U18402 ( .A(n16628), .B(n16627), .Z(n16643) );
  XNOR U18403 ( .A(n16642), .B(n16643), .Z(n16634) );
  XNOR U18404 ( .A(n16635), .B(n16634), .Z(n16636) );
  XNOR U18405 ( .A(n16637), .B(n16636), .Z(n16666) );
  XNOR U18406 ( .A(sreg[1355]), .B(n16666), .Z(n16668) );
  NANDN U18407 ( .A(sreg[1354]), .B(n16629), .Z(n16633) );
  NAND U18408 ( .A(n16631), .B(n16630), .Z(n16632) );
  NAND U18409 ( .A(n16633), .B(n16632), .Z(n16667) );
  XNOR U18410 ( .A(n16668), .B(n16667), .Z(c[1355]) );
  NANDN U18411 ( .A(n16635), .B(n16634), .Z(n16639) );
  NANDN U18412 ( .A(n16637), .B(n16636), .Z(n16638) );
  AND U18413 ( .A(n16639), .B(n16638), .Z(n16674) );
  NANDN U18414 ( .A(n16641), .B(n16640), .Z(n16645) );
  NANDN U18415 ( .A(n16643), .B(n16642), .Z(n16644) );
  AND U18416 ( .A(n16645), .B(n16644), .Z(n16672) );
  NAND U18417 ( .A(n42143), .B(n16646), .Z(n16648) );
  XNOR U18418 ( .A(a[334]), .B(n4119), .Z(n16683) );
  NAND U18419 ( .A(n42144), .B(n16683), .Z(n16647) );
  AND U18420 ( .A(n16648), .B(n16647), .Z(n16698) );
  XOR U18421 ( .A(a[338]), .B(n42012), .Z(n16686) );
  XNOR U18422 ( .A(n16698), .B(n16697), .Z(n16700) );
  AND U18423 ( .A(a[340]), .B(b[0]), .Z(n16650) );
  XNOR U18424 ( .A(n16650), .B(n4071), .Z(n16652) );
  NANDN U18425 ( .A(b[0]), .B(a[339]), .Z(n16651) );
  NAND U18426 ( .A(n16652), .B(n16651), .Z(n16694) );
  XOR U18427 ( .A(a[336]), .B(n42085), .Z(n16690) );
  AND U18428 ( .A(a[332]), .B(b[7]), .Z(n16691) );
  XNOR U18429 ( .A(n16692), .B(n16691), .Z(n16693) );
  XNOR U18430 ( .A(n16694), .B(n16693), .Z(n16699) );
  XOR U18431 ( .A(n16700), .B(n16699), .Z(n16678) );
  NANDN U18432 ( .A(n16655), .B(n16654), .Z(n16659) );
  NANDN U18433 ( .A(n16657), .B(n16656), .Z(n16658) );
  AND U18434 ( .A(n16659), .B(n16658), .Z(n16677) );
  XNOR U18435 ( .A(n16678), .B(n16677), .Z(n16679) );
  NANDN U18436 ( .A(n16661), .B(n16660), .Z(n16665) );
  NAND U18437 ( .A(n16663), .B(n16662), .Z(n16664) );
  NAND U18438 ( .A(n16665), .B(n16664), .Z(n16680) );
  XNOR U18439 ( .A(n16679), .B(n16680), .Z(n16671) );
  XNOR U18440 ( .A(n16672), .B(n16671), .Z(n16673) );
  XNOR U18441 ( .A(n16674), .B(n16673), .Z(n16703) );
  XNOR U18442 ( .A(sreg[1356]), .B(n16703), .Z(n16705) );
  NANDN U18443 ( .A(sreg[1355]), .B(n16666), .Z(n16670) );
  NAND U18444 ( .A(n16668), .B(n16667), .Z(n16669) );
  NAND U18445 ( .A(n16670), .B(n16669), .Z(n16704) );
  XNOR U18446 ( .A(n16705), .B(n16704), .Z(c[1356]) );
  NANDN U18447 ( .A(n16672), .B(n16671), .Z(n16676) );
  NANDN U18448 ( .A(n16674), .B(n16673), .Z(n16675) );
  AND U18449 ( .A(n16676), .B(n16675), .Z(n16711) );
  NANDN U18450 ( .A(n16678), .B(n16677), .Z(n16682) );
  NANDN U18451 ( .A(n16680), .B(n16679), .Z(n16681) );
  AND U18452 ( .A(n16682), .B(n16681), .Z(n16709) );
  NAND U18453 ( .A(n42143), .B(n16683), .Z(n16685) );
  XNOR U18454 ( .A(a[335]), .B(n4119), .Z(n16720) );
  NAND U18455 ( .A(n42144), .B(n16720), .Z(n16684) );
  AND U18456 ( .A(n16685), .B(n16684), .Z(n16735) );
  XOR U18457 ( .A(a[339]), .B(n42012), .Z(n16723) );
  XNOR U18458 ( .A(n16735), .B(n16734), .Z(n16737) );
  AND U18459 ( .A(a[341]), .B(b[0]), .Z(n16687) );
  XNOR U18460 ( .A(n16687), .B(n4071), .Z(n16689) );
  NANDN U18461 ( .A(b[0]), .B(a[340]), .Z(n16688) );
  NAND U18462 ( .A(n16689), .B(n16688), .Z(n16731) );
  XOR U18463 ( .A(a[337]), .B(n42085), .Z(n16727) );
  AND U18464 ( .A(a[333]), .B(b[7]), .Z(n16728) );
  XNOR U18465 ( .A(n16729), .B(n16728), .Z(n16730) );
  XNOR U18466 ( .A(n16731), .B(n16730), .Z(n16736) );
  XOR U18467 ( .A(n16737), .B(n16736), .Z(n16715) );
  NANDN U18468 ( .A(n16692), .B(n16691), .Z(n16696) );
  NANDN U18469 ( .A(n16694), .B(n16693), .Z(n16695) );
  AND U18470 ( .A(n16696), .B(n16695), .Z(n16714) );
  XNOR U18471 ( .A(n16715), .B(n16714), .Z(n16716) );
  NANDN U18472 ( .A(n16698), .B(n16697), .Z(n16702) );
  NAND U18473 ( .A(n16700), .B(n16699), .Z(n16701) );
  NAND U18474 ( .A(n16702), .B(n16701), .Z(n16717) );
  XNOR U18475 ( .A(n16716), .B(n16717), .Z(n16708) );
  XNOR U18476 ( .A(n16709), .B(n16708), .Z(n16710) );
  XNOR U18477 ( .A(n16711), .B(n16710), .Z(n16740) );
  XNOR U18478 ( .A(sreg[1357]), .B(n16740), .Z(n16742) );
  NANDN U18479 ( .A(sreg[1356]), .B(n16703), .Z(n16707) );
  NAND U18480 ( .A(n16705), .B(n16704), .Z(n16706) );
  NAND U18481 ( .A(n16707), .B(n16706), .Z(n16741) );
  XNOR U18482 ( .A(n16742), .B(n16741), .Z(c[1357]) );
  NANDN U18483 ( .A(n16709), .B(n16708), .Z(n16713) );
  NANDN U18484 ( .A(n16711), .B(n16710), .Z(n16712) );
  AND U18485 ( .A(n16713), .B(n16712), .Z(n16748) );
  NANDN U18486 ( .A(n16715), .B(n16714), .Z(n16719) );
  NANDN U18487 ( .A(n16717), .B(n16716), .Z(n16718) );
  AND U18488 ( .A(n16719), .B(n16718), .Z(n16746) );
  NAND U18489 ( .A(n42143), .B(n16720), .Z(n16722) );
  XNOR U18490 ( .A(a[336]), .B(n4119), .Z(n16757) );
  NAND U18491 ( .A(n42144), .B(n16757), .Z(n16721) );
  AND U18492 ( .A(n16722), .B(n16721), .Z(n16772) );
  XOR U18493 ( .A(a[340]), .B(n42012), .Z(n16760) );
  XNOR U18494 ( .A(n16772), .B(n16771), .Z(n16774) );
  AND U18495 ( .A(a[342]), .B(b[0]), .Z(n16724) );
  XNOR U18496 ( .A(n16724), .B(n4071), .Z(n16726) );
  NANDN U18497 ( .A(b[0]), .B(a[341]), .Z(n16725) );
  NAND U18498 ( .A(n16726), .B(n16725), .Z(n16768) );
  XOR U18499 ( .A(a[338]), .B(n42085), .Z(n16764) );
  AND U18500 ( .A(a[334]), .B(b[7]), .Z(n16765) );
  XNOR U18501 ( .A(n16766), .B(n16765), .Z(n16767) );
  XNOR U18502 ( .A(n16768), .B(n16767), .Z(n16773) );
  XOR U18503 ( .A(n16774), .B(n16773), .Z(n16752) );
  NANDN U18504 ( .A(n16729), .B(n16728), .Z(n16733) );
  NANDN U18505 ( .A(n16731), .B(n16730), .Z(n16732) );
  AND U18506 ( .A(n16733), .B(n16732), .Z(n16751) );
  XNOR U18507 ( .A(n16752), .B(n16751), .Z(n16753) );
  NANDN U18508 ( .A(n16735), .B(n16734), .Z(n16739) );
  NAND U18509 ( .A(n16737), .B(n16736), .Z(n16738) );
  NAND U18510 ( .A(n16739), .B(n16738), .Z(n16754) );
  XNOR U18511 ( .A(n16753), .B(n16754), .Z(n16745) );
  XNOR U18512 ( .A(n16746), .B(n16745), .Z(n16747) );
  XNOR U18513 ( .A(n16748), .B(n16747), .Z(n16777) );
  XNOR U18514 ( .A(sreg[1358]), .B(n16777), .Z(n16779) );
  NANDN U18515 ( .A(sreg[1357]), .B(n16740), .Z(n16744) );
  NAND U18516 ( .A(n16742), .B(n16741), .Z(n16743) );
  NAND U18517 ( .A(n16744), .B(n16743), .Z(n16778) );
  XNOR U18518 ( .A(n16779), .B(n16778), .Z(c[1358]) );
  NANDN U18519 ( .A(n16746), .B(n16745), .Z(n16750) );
  NANDN U18520 ( .A(n16748), .B(n16747), .Z(n16749) );
  AND U18521 ( .A(n16750), .B(n16749), .Z(n16785) );
  NANDN U18522 ( .A(n16752), .B(n16751), .Z(n16756) );
  NANDN U18523 ( .A(n16754), .B(n16753), .Z(n16755) );
  AND U18524 ( .A(n16756), .B(n16755), .Z(n16783) );
  NAND U18525 ( .A(n42143), .B(n16757), .Z(n16759) );
  XNOR U18526 ( .A(a[337]), .B(n4120), .Z(n16794) );
  NAND U18527 ( .A(n42144), .B(n16794), .Z(n16758) );
  AND U18528 ( .A(n16759), .B(n16758), .Z(n16809) );
  XOR U18529 ( .A(a[341]), .B(n42012), .Z(n16797) );
  XNOR U18530 ( .A(n16809), .B(n16808), .Z(n16811) );
  AND U18531 ( .A(a[343]), .B(b[0]), .Z(n16761) );
  XNOR U18532 ( .A(n16761), .B(n4071), .Z(n16763) );
  NANDN U18533 ( .A(b[0]), .B(a[342]), .Z(n16762) );
  NAND U18534 ( .A(n16763), .B(n16762), .Z(n16805) );
  XOR U18535 ( .A(a[339]), .B(n42085), .Z(n16801) );
  AND U18536 ( .A(a[335]), .B(b[7]), .Z(n16802) );
  XNOR U18537 ( .A(n16803), .B(n16802), .Z(n16804) );
  XNOR U18538 ( .A(n16805), .B(n16804), .Z(n16810) );
  XOR U18539 ( .A(n16811), .B(n16810), .Z(n16789) );
  NANDN U18540 ( .A(n16766), .B(n16765), .Z(n16770) );
  NANDN U18541 ( .A(n16768), .B(n16767), .Z(n16769) );
  AND U18542 ( .A(n16770), .B(n16769), .Z(n16788) );
  XNOR U18543 ( .A(n16789), .B(n16788), .Z(n16790) );
  NANDN U18544 ( .A(n16772), .B(n16771), .Z(n16776) );
  NAND U18545 ( .A(n16774), .B(n16773), .Z(n16775) );
  NAND U18546 ( .A(n16776), .B(n16775), .Z(n16791) );
  XNOR U18547 ( .A(n16790), .B(n16791), .Z(n16782) );
  XNOR U18548 ( .A(n16783), .B(n16782), .Z(n16784) );
  XNOR U18549 ( .A(n16785), .B(n16784), .Z(n16814) );
  XNOR U18550 ( .A(sreg[1359]), .B(n16814), .Z(n16816) );
  NANDN U18551 ( .A(sreg[1358]), .B(n16777), .Z(n16781) );
  NAND U18552 ( .A(n16779), .B(n16778), .Z(n16780) );
  NAND U18553 ( .A(n16781), .B(n16780), .Z(n16815) );
  XNOR U18554 ( .A(n16816), .B(n16815), .Z(c[1359]) );
  NANDN U18555 ( .A(n16783), .B(n16782), .Z(n16787) );
  NANDN U18556 ( .A(n16785), .B(n16784), .Z(n16786) );
  AND U18557 ( .A(n16787), .B(n16786), .Z(n16822) );
  NANDN U18558 ( .A(n16789), .B(n16788), .Z(n16793) );
  NANDN U18559 ( .A(n16791), .B(n16790), .Z(n16792) );
  AND U18560 ( .A(n16793), .B(n16792), .Z(n16820) );
  NAND U18561 ( .A(n42143), .B(n16794), .Z(n16796) );
  XNOR U18562 ( .A(a[338]), .B(n4120), .Z(n16831) );
  NAND U18563 ( .A(n42144), .B(n16831), .Z(n16795) );
  AND U18564 ( .A(n16796), .B(n16795), .Z(n16846) );
  XOR U18565 ( .A(a[342]), .B(n42012), .Z(n16834) );
  XNOR U18566 ( .A(n16846), .B(n16845), .Z(n16848) );
  AND U18567 ( .A(a[344]), .B(b[0]), .Z(n16798) );
  XNOR U18568 ( .A(n16798), .B(n4071), .Z(n16800) );
  NANDN U18569 ( .A(b[0]), .B(a[343]), .Z(n16799) );
  NAND U18570 ( .A(n16800), .B(n16799), .Z(n16842) );
  XOR U18571 ( .A(a[340]), .B(n42085), .Z(n16838) );
  AND U18572 ( .A(a[336]), .B(b[7]), .Z(n16839) );
  XNOR U18573 ( .A(n16840), .B(n16839), .Z(n16841) );
  XNOR U18574 ( .A(n16842), .B(n16841), .Z(n16847) );
  XOR U18575 ( .A(n16848), .B(n16847), .Z(n16826) );
  NANDN U18576 ( .A(n16803), .B(n16802), .Z(n16807) );
  NANDN U18577 ( .A(n16805), .B(n16804), .Z(n16806) );
  AND U18578 ( .A(n16807), .B(n16806), .Z(n16825) );
  XNOR U18579 ( .A(n16826), .B(n16825), .Z(n16827) );
  NANDN U18580 ( .A(n16809), .B(n16808), .Z(n16813) );
  NAND U18581 ( .A(n16811), .B(n16810), .Z(n16812) );
  NAND U18582 ( .A(n16813), .B(n16812), .Z(n16828) );
  XNOR U18583 ( .A(n16827), .B(n16828), .Z(n16819) );
  XNOR U18584 ( .A(n16820), .B(n16819), .Z(n16821) );
  XNOR U18585 ( .A(n16822), .B(n16821), .Z(n16851) );
  XNOR U18586 ( .A(sreg[1360]), .B(n16851), .Z(n16853) );
  NANDN U18587 ( .A(sreg[1359]), .B(n16814), .Z(n16818) );
  NAND U18588 ( .A(n16816), .B(n16815), .Z(n16817) );
  NAND U18589 ( .A(n16818), .B(n16817), .Z(n16852) );
  XNOR U18590 ( .A(n16853), .B(n16852), .Z(c[1360]) );
  NANDN U18591 ( .A(n16820), .B(n16819), .Z(n16824) );
  NANDN U18592 ( .A(n16822), .B(n16821), .Z(n16823) );
  AND U18593 ( .A(n16824), .B(n16823), .Z(n16859) );
  NANDN U18594 ( .A(n16826), .B(n16825), .Z(n16830) );
  NANDN U18595 ( .A(n16828), .B(n16827), .Z(n16829) );
  AND U18596 ( .A(n16830), .B(n16829), .Z(n16857) );
  NAND U18597 ( .A(n42143), .B(n16831), .Z(n16833) );
  XNOR U18598 ( .A(a[339]), .B(n4120), .Z(n16868) );
  NAND U18599 ( .A(n42144), .B(n16868), .Z(n16832) );
  AND U18600 ( .A(n16833), .B(n16832), .Z(n16883) );
  XOR U18601 ( .A(a[343]), .B(n42012), .Z(n16871) );
  XNOR U18602 ( .A(n16883), .B(n16882), .Z(n16885) );
  AND U18603 ( .A(a[345]), .B(b[0]), .Z(n16835) );
  XNOR U18604 ( .A(n16835), .B(n4071), .Z(n16837) );
  NANDN U18605 ( .A(b[0]), .B(a[344]), .Z(n16836) );
  NAND U18606 ( .A(n16837), .B(n16836), .Z(n16879) );
  XOR U18607 ( .A(a[341]), .B(n42085), .Z(n16872) );
  AND U18608 ( .A(a[337]), .B(b[7]), .Z(n16876) );
  XNOR U18609 ( .A(n16877), .B(n16876), .Z(n16878) );
  XNOR U18610 ( .A(n16879), .B(n16878), .Z(n16884) );
  XOR U18611 ( .A(n16885), .B(n16884), .Z(n16863) );
  NANDN U18612 ( .A(n16840), .B(n16839), .Z(n16844) );
  NANDN U18613 ( .A(n16842), .B(n16841), .Z(n16843) );
  AND U18614 ( .A(n16844), .B(n16843), .Z(n16862) );
  XNOR U18615 ( .A(n16863), .B(n16862), .Z(n16864) );
  NANDN U18616 ( .A(n16846), .B(n16845), .Z(n16850) );
  NAND U18617 ( .A(n16848), .B(n16847), .Z(n16849) );
  NAND U18618 ( .A(n16850), .B(n16849), .Z(n16865) );
  XNOR U18619 ( .A(n16864), .B(n16865), .Z(n16856) );
  XNOR U18620 ( .A(n16857), .B(n16856), .Z(n16858) );
  XNOR U18621 ( .A(n16859), .B(n16858), .Z(n16888) );
  XNOR U18622 ( .A(sreg[1361]), .B(n16888), .Z(n16890) );
  NANDN U18623 ( .A(sreg[1360]), .B(n16851), .Z(n16855) );
  NAND U18624 ( .A(n16853), .B(n16852), .Z(n16854) );
  NAND U18625 ( .A(n16855), .B(n16854), .Z(n16889) );
  XNOR U18626 ( .A(n16890), .B(n16889), .Z(c[1361]) );
  NANDN U18627 ( .A(n16857), .B(n16856), .Z(n16861) );
  NANDN U18628 ( .A(n16859), .B(n16858), .Z(n16860) );
  AND U18629 ( .A(n16861), .B(n16860), .Z(n16896) );
  NANDN U18630 ( .A(n16863), .B(n16862), .Z(n16867) );
  NANDN U18631 ( .A(n16865), .B(n16864), .Z(n16866) );
  AND U18632 ( .A(n16867), .B(n16866), .Z(n16894) );
  NAND U18633 ( .A(n42143), .B(n16868), .Z(n16870) );
  XNOR U18634 ( .A(a[340]), .B(n4120), .Z(n16905) );
  NAND U18635 ( .A(n42144), .B(n16905), .Z(n16869) );
  AND U18636 ( .A(n16870), .B(n16869), .Z(n16920) );
  XOR U18637 ( .A(a[344]), .B(n42012), .Z(n16908) );
  XNOR U18638 ( .A(n16920), .B(n16919), .Z(n16922) );
  XOR U18639 ( .A(a[342]), .B(n42085), .Z(n16912) );
  AND U18640 ( .A(a[338]), .B(b[7]), .Z(n16913) );
  XNOR U18641 ( .A(n16914), .B(n16913), .Z(n16915) );
  AND U18642 ( .A(a[346]), .B(b[0]), .Z(n16873) );
  XNOR U18643 ( .A(n16873), .B(n4071), .Z(n16875) );
  NANDN U18644 ( .A(b[0]), .B(a[345]), .Z(n16874) );
  NAND U18645 ( .A(n16875), .B(n16874), .Z(n16916) );
  XNOR U18646 ( .A(n16915), .B(n16916), .Z(n16921) );
  XOR U18647 ( .A(n16922), .B(n16921), .Z(n16900) );
  NANDN U18648 ( .A(n16877), .B(n16876), .Z(n16881) );
  NANDN U18649 ( .A(n16879), .B(n16878), .Z(n16880) );
  AND U18650 ( .A(n16881), .B(n16880), .Z(n16899) );
  XNOR U18651 ( .A(n16900), .B(n16899), .Z(n16901) );
  NANDN U18652 ( .A(n16883), .B(n16882), .Z(n16887) );
  NAND U18653 ( .A(n16885), .B(n16884), .Z(n16886) );
  NAND U18654 ( .A(n16887), .B(n16886), .Z(n16902) );
  XNOR U18655 ( .A(n16901), .B(n16902), .Z(n16893) );
  XNOR U18656 ( .A(n16894), .B(n16893), .Z(n16895) );
  XNOR U18657 ( .A(n16896), .B(n16895), .Z(n16925) );
  XNOR U18658 ( .A(sreg[1362]), .B(n16925), .Z(n16927) );
  NANDN U18659 ( .A(sreg[1361]), .B(n16888), .Z(n16892) );
  NAND U18660 ( .A(n16890), .B(n16889), .Z(n16891) );
  NAND U18661 ( .A(n16892), .B(n16891), .Z(n16926) );
  XNOR U18662 ( .A(n16927), .B(n16926), .Z(c[1362]) );
  NANDN U18663 ( .A(n16894), .B(n16893), .Z(n16898) );
  NANDN U18664 ( .A(n16896), .B(n16895), .Z(n16897) );
  AND U18665 ( .A(n16898), .B(n16897), .Z(n16933) );
  NANDN U18666 ( .A(n16900), .B(n16899), .Z(n16904) );
  NANDN U18667 ( .A(n16902), .B(n16901), .Z(n16903) );
  AND U18668 ( .A(n16904), .B(n16903), .Z(n16931) );
  NAND U18669 ( .A(n42143), .B(n16905), .Z(n16907) );
  XNOR U18670 ( .A(a[341]), .B(n4120), .Z(n16942) );
  NAND U18671 ( .A(n42144), .B(n16942), .Z(n16906) );
  AND U18672 ( .A(n16907), .B(n16906), .Z(n16957) );
  XOR U18673 ( .A(a[345]), .B(n42012), .Z(n16945) );
  XNOR U18674 ( .A(n16957), .B(n16956), .Z(n16959) );
  AND U18675 ( .A(b[0]), .B(a[347]), .Z(n16909) );
  XOR U18676 ( .A(b[1]), .B(n16909), .Z(n16911) );
  NANDN U18677 ( .A(b[0]), .B(a[346]), .Z(n16910) );
  AND U18678 ( .A(n16911), .B(n16910), .Z(n16952) );
  XOR U18679 ( .A(a[343]), .B(n42085), .Z(n16949) );
  AND U18680 ( .A(a[339]), .B(b[7]), .Z(n16950) );
  XOR U18681 ( .A(n16951), .B(n16950), .Z(n16953) );
  XNOR U18682 ( .A(n16952), .B(n16953), .Z(n16958) );
  XOR U18683 ( .A(n16959), .B(n16958), .Z(n16937) );
  NANDN U18684 ( .A(n16914), .B(n16913), .Z(n16918) );
  NANDN U18685 ( .A(n16916), .B(n16915), .Z(n16917) );
  AND U18686 ( .A(n16918), .B(n16917), .Z(n16936) );
  XNOR U18687 ( .A(n16937), .B(n16936), .Z(n16938) );
  NANDN U18688 ( .A(n16920), .B(n16919), .Z(n16924) );
  NAND U18689 ( .A(n16922), .B(n16921), .Z(n16923) );
  NAND U18690 ( .A(n16924), .B(n16923), .Z(n16939) );
  XNOR U18691 ( .A(n16938), .B(n16939), .Z(n16930) );
  XNOR U18692 ( .A(n16931), .B(n16930), .Z(n16932) );
  XNOR U18693 ( .A(n16933), .B(n16932), .Z(n16962) );
  XNOR U18694 ( .A(sreg[1363]), .B(n16962), .Z(n16964) );
  NANDN U18695 ( .A(sreg[1362]), .B(n16925), .Z(n16929) );
  NAND U18696 ( .A(n16927), .B(n16926), .Z(n16928) );
  NAND U18697 ( .A(n16929), .B(n16928), .Z(n16963) );
  XNOR U18698 ( .A(n16964), .B(n16963), .Z(c[1363]) );
  NANDN U18699 ( .A(n16931), .B(n16930), .Z(n16935) );
  NANDN U18700 ( .A(n16933), .B(n16932), .Z(n16934) );
  AND U18701 ( .A(n16935), .B(n16934), .Z(n16970) );
  NANDN U18702 ( .A(n16937), .B(n16936), .Z(n16941) );
  NANDN U18703 ( .A(n16939), .B(n16938), .Z(n16940) );
  AND U18704 ( .A(n16941), .B(n16940), .Z(n16968) );
  NAND U18705 ( .A(n42143), .B(n16942), .Z(n16944) );
  XNOR U18706 ( .A(a[342]), .B(n4120), .Z(n16979) );
  NAND U18707 ( .A(n42144), .B(n16979), .Z(n16943) );
  AND U18708 ( .A(n16944), .B(n16943), .Z(n16994) );
  XOR U18709 ( .A(a[346]), .B(n42012), .Z(n16982) );
  XNOR U18710 ( .A(n16994), .B(n16993), .Z(n16996) );
  AND U18711 ( .A(a[348]), .B(b[0]), .Z(n16946) );
  XNOR U18712 ( .A(n16946), .B(n4071), .Z(n16948) );
  NANDN U18713 ( .A(b[0]), .B(a[347]), .Z(n16947) );
  NAND U18714 ( .A(n16948), .B(n16947), .Z(n16990) );
  XOR U18715 ( .A(a[344]), .B(n42085), .Z(n16986) );
  AND U18716 ( .A(a[340]), .B(b[7]), .Z(n16987) );
  XNOR U18717 ( .A(n16988), .B(n16987), .Z(n16989) );
  XNOR U18718 ( .A(n16990), .B(n16989), .Z(n16995) );
  XOR U18719 ( .A(n16996), .B(n16995), .Z(n16974) );
  NANDN U18720 ( .A(n16951), .B(n16950), .Z(n16955) );
  NANDN U18721 ( .A(n16953), .B(n16952), .Z(n16954) );
  AND U18722 ( .A(n16955), .B(n16954), .Z(n16973) );
  XNOR U18723 ( .A(n16974), .B(n16973), .Z(n16975) );
  NANDN U18724 ( .A(n16957), .B(n16956), .Z(n16961) );
  NAND U18725 ( .A(n16959), .B(n16958), .Z(n16960) );
  NAND U18726 ( .A(n16961), .B(n16960), .Z(n16976) );
  XNOR U18727 ( .A(n16975), .B(n16976), .Z(n16967) );
  XNOR U18728 ( .A(n16968), .B(n16967), .Z(n16969) );
  XNOR U18729 ( .A(n16970), .B(n16969), .Z(n16999) );
  XNOR U18730 ( .A(sreg[1364]), .B(n16999), .Z(n17001) );
  NANDN U18731 ( .A(sreg[1363]), .B(n16962), .Z(n16966) );
  NAND U18732 ( .A(n16964), .B(n16963), .Z(n16965) );
  NAND U18733 ( .A(n16966), .B(n16965), .Z(n17000) );
  XNOR U18734 ( .A(n17001), .B(n17000), .Z(c[1364]) );
  NANDN U18735 ( .A(n16968), .B(n16967), .Z(n16972) );
  NANDN U18736 ( .A(n16970), .B(n16969), .Z(n16971) );
  AND U18737 ( .A(n16972), .B(n16971), .Z(n17007) );
  NANDN U18738 ( .A(n16974), .B(n16973), .Z(n16978) );
  NANDN U18739 ( .A(n16976), .B(n16975), .Z(n16977) );
  AND U18740 ( .A(n16978), .B(n16977), .Z(n17005) );
  NAND U18741 ( .A(n42143), .B(n16979), .Z(n16981) );
  XNOR U18742 ( .A(a[343]), .B(n4120), .Z(n17016) );
  NAND U18743 ( .A(n42144), .B(n17016), .Z(n16980) );
  AND U18744 ( .A(n16981), .B(n16980), .Z(n17031) );
  XOR U18745 ( .A(a[347]), .B(n42012), .Z(n17019) );
  XNOR U18746 ( .A(n17031), .B(n17030), .Z(n17033) );
  AND U18747 ( .A(a[349]), .B(b[0]), .Z(n16983) );
  XNOR U18748 ( .A(n16983), .B(n4071), .Z(n16985) );
  NANDN U18749 ( .A(b[0]), .B(a[348]), .Z(n16984) );
  NAND U18750 ( .A(n16985), .B(n16984), .Z(n17027) );
  XOR U18751 ( .A(a[345]), .B(n42085), .Z(n17023) );
  AND U18752 ( .A(a[341]), .B(b[7]), .Z(n17024) );
  XNOR U18753 ( .A(n17025), .B(n17024), .Z(n17026) );
  XNOR U18754 ( .A(n17027), .B(n17026), .Z(n17032) );
  XOR U18755 ( .A(n17033), .B(n17032), .Z(n17011) );
  NANDN U18756 ( .A(n16988), .B(n16987), .Z(n16992) );
  NANDN U18757 ( .A(n16990), .B(n16989), .Z(n16991) );
  AND U18758 ( .A(n16992), .B(n16991), .Z(n17010) );
  XNOR U18759 ( .A(n17011), .B(n17010), .Z(n17012) );
  NANDN U18760 ( .A(n16994), .B(n16993), .Z(n16998) );
  NAND U18761 ( .A(n16996), .B(n16995), .Z(n16997) );
  NAND U18762 ( .A(n16998), .B(n16997), .Z(n17013) );
  XNOR U18763 ( .A(n17012), .B(n17013), .Z(n17004) );
  XNOR U18764 ( .A(n17005), .B(n17004), .Z(n17006) );
  XNOR U18765 ( .A(n17007), .B(n17006), .Z(n17036) );
  XNOR U18766 ( .A(sreg[1365]), .B(n17036), .Z(n17038) );
  NANDN U18767 ( .A(sreg[1364]), .B(n16999), .Z(n17003) );
  NAND U18768 ( .A(n17001), .B(n17000), .Z(n17002) );
  NAND U18769 ( .A(n17003), .B(n17002), .Z(n17037) );
  XNOR U18770 ( .A(n17038), .B(n17037), .Z(c[1365]) );
  NANDN U18771 ( .A(n17005), .B(n17004), .Z(n17009) );
  NANDN U18772 ( .A(n17007), .B(n17006), .Z(n17008) );
  AND U18773 ( .A(n17009), .B(n17008), .Z(n17044) );
  NANDN U18774 ( .A(n17011), .B(n17010), .Z(n17015) );
  NANDN U18775 ( .A(n17013), .B(n17012), .Z(n17014) );
  AND U18776 ( .A(n17015), .B(n17014), .Z(n17042) );
  NAND U18777 ( .A(n42143), .B(n17016), .Z(n17018) );
  XNOR U18778 ( .A(a[344]), .B(n4121), .Z(n17053) );
  NAND U18779 ( .A(n42144), .B(n17053), .Z(n17017) );
  AND U18780 ( .A(n17018), .B(n17017), .Z(n17068) );
  XOR U18781 ( .A(a[348]), .B(n42012), .Z(n17056) );
  XNOR U18782 ( .A(n17068), .B(n17067), .Z(n17070) );
  AND U18783 ( .A(a[350]), .B(b[0]), .Z(n17020) );
  XNOR U18784 ( .A(n17020), .B(n4071), .Z(n17022) );
  NANDN U18785 ( .A(b[0]), .B(a[349]), .Z(n17021) );
  NAND U18786 ( .A(n17022), .B(n17021), .Z(n17064) );
  XOR U18787 ( .A(a[346]), .B(n42085), .Z(n17060) );
  AND U18788 ( .A(a[342]), .B(b[7]), .Z(n17061) );
  XNOR U18789 ( .A(n17062), .B(n17061), .Z(n17063) );
  XNOR U18790 ( .A(n17064), .B(n17063), .Z(n17069) );
  XOR U18791 ( .A(n17070), .B(n17069), .Z(n17048) );
  NANDN U18792 ( .A(n17025), .B(n17024), .Z(n17029) );
  NANDN U18793 ( .A(n17027), .B(n17026), .Z(n17028) );
  AND U18794 ( .A(n17029), .B(n17028), .Z(n17047) );
  XNOR U18795 ( .A(n17048), .B(n17047), .Z(n17049) );
  NANDN U18796 ( .A(n17031), .B(n17030), .Z(n17035) );
  NAND U18797 ( .A(n17033), .B(n17032), .Z(n17034) );
  NAND U18798 ( .A(n17035), .B(n17034), .Z(n17050) );
  XNOR U18799 ( .A(n17049), .B(n17050), .Z(n17041) );
  XNOR U18800 ( .A(n17042), .B(n17041), .Z(n17043) );
  XNOR U18801 ( .A(n17044), .B(n17043), .Z(n17073) );
  XNOR U18802 ( .A(sreg[1366]), .B(n17073), .Z(n17075) );
  NANDN U18803 ( .A(sreg[1365]), .B(n17036), .Z(n17040) );
  NAND U18804 ( .A(n17038), .B(n17037), .Z(n17039) );
  NAND U18805 ( .A(n17040), .B(n17039), .Z(n17074) );
  XNOR U18806 ( .A(n17075), .B(n17074), .Z(c[1366]) );
  NANDN U18807 ( .A(n17042), .B(n17041), .Z(n17046) );
  NANDN U18808 ( .A(n17044), .B(n17043), .Z(n17045) );
  AND U18809 ( .A(n17046), .B(n17045), .Z(n17081) );
  NANDN U18810 ( .A(n17048), .B(n17047), .Z(n17052) );
  NANDN U18811 ( .A(n17050), .B(n17049), .Z(n17051) );
  AND U18812 ( .A(n17052), .B(n17051), .Z(n17079) );
  NAND U18813 ( .A(n42143), .B(n17053), .Z(n17055) );
  XNOR U18814 ( .A(a[345]), .B(n4121), .Z(n17090) );
  NAND U18815 ( .A(n42144), .B(n17090), .Z(n17054) );
  AND U18816 ( .A(n17055), .B(n17054), .Z(n17105) );
  XOR U18817 ( .A(a[349]), .B(n42012), .Z(n17093) );
  XNOR U18818 ( .A(n17105), .B(n17104), .Z(n17107) );
  AND U18819 ( .A(a[351]), .B(b[0]), .Z(n17057) );
  XNOR U18820 ( .A(n17057), .B(n4071), .Z(n17059) );
  NANDN U18821 ( .A(b[0]), .B(a[350]), .Z(n17058) );
  NAND U18822 ( .A(n17059), .B(n17058), .Z(n17101) );
  XOR U18823 ( .A(a[347]), .B(n42085), .Z(n17094) );
  AND U18824 ( .A(a[343]), .B(b[7]), .Z(n17098) );
  XNOR U18825 ( .A(n17099), .B(n17098), .Z(n17100) );
  XNOR U18826 ( .A(n17101), .B(n17100), .Z(n17106) );
  XOR U18827 ( .A(n17107), .B(n17106), .Z(n17085) );
  NANDN U18828 ( .A(n17062), .B(n17061), .Z(n17066) );
  NANDN U18829 ( .A(n17064), .B(n17063), .Z(n17065) );
  AND U18830 ( .A(n17066), .B(n17065), .Z(n17084) );
  XNOR U18831 ( .A(n17085), .B(n17084), .Z(n17086) );
  NANDN U18832 ( .A(n17068), .B(n17067), .Z(n17072) );
  NAND U18833 ( .A(n17070), .B(n17069), .Z(n17071) );
  NAND U18834 ( .A(n17072), .B(n17071), .Z(n17087) );
  XNOR U18835 ( .A(n17086), .B(n17087), .Z(n17078) );
  XNOR U18836 ( .A(n17079), .B(n17078), .Z(n17080) );
  XNOR U18837 ( .A(n17081), .B(n17080), .Z(n17110) );
  XNOR U18838 ( .A(sreg[1367]), .B(n17110), .Z(n17112) );
  NANDN U18839 ( .A(sreg[1366]), .B(n17073), .Z(n17077) );
  NAND U18840 ( .A(n17075), .B(n17074), .Z(n17076) );
  NAND U18841 ( .A(n17077), .B(n17076), .Z(n17111) );
  XNOR U18842 ( .A(n17112), .B(n17111), .Z(c[1367]) );
  NANDN U18843 ( .A(n17079), .B(n17078), .Z(n17083) );
  NANDN U18844 ( .A(n17081), .B(n17080), .Z(n17082) );
  AND U18845 ( .A(n17083), .B(n17082), .Z(n17118) );
  NANDN U18846 ( .A(n17085), .B(n17084), .Z(n17089) );
  NANDN U18847 ( .A(n17087), .B(n17086), .Z(n17088) );
  AND U18848 ( .A(n17089), .B(n17088), .Z(n17116) );
  NAND U18849 ( .A(n42143), .B(n17090), .Z(n17092) );
  XNOR U18850 ( .A(a[346]), .B(n4121), .Z(n17127) );
  NAND U18851 ( .A(n42144), .B(n17127), .Z(n17091) );
  AND U18852 ( .A(n17092), .B(n17091), .Z(n17142) );
  XOR U18853 ( .A(a[350]), .B(n42012), .Z(n17130) );
  XNOR U18854 ( .A(n17142), .B(n17141), .Z(n17144) );
  XOR U18855 ( .A(a[348]), .B(n42085), .Z(n17134) );
  AND U18856 ( .A(a[344]), .B(b[7]), .Z(n17135) );
  XNOR U18857 ( .A(n17136), .B(n17135), .Z(n17137) );
  AND U18858 ( .A(a[352]), .B(b[0]), .Z(n17095) );
  XNOR U18859 ( .A(n17095), .B(n4071), .Z(n17097) );
  NANDN U18860 ( .A(b[0]), .B(a[351]), .Z(n17096) );
  NAND U18861 ( .A(n17097), .B(n17096), .Z(n17138) );
  XNOR U18862 ( .A(n17137), .B(n17138), .Z(n17143) );
  XOR U18863 ( .A(n17144), .B(n17143), .Z(n17122) );
  NANDN U18864 ( .A(n17099), .B(n17098), .Z(n17103) );
  NANDN U18865 ( .A(n17101), .B(n17100), .Z(n17102) );
  AND U18866 ( .A(n17103), .B(n17102), .Z(n17121) );
  XNOR U18867 ( .A(n17122), .B(n17121), .Z(n17123) );
  NANDN U18868 ( .A(n17105), .B(n17104), .Z(n17109) );
  NAND U18869 ( .A(n17107), .B(n17106), .Z(n17108) );
  NAND U18870 ( .A(n17109), .B(n17108), .Z(n17124) );
  XNOR U18871 ( .A(n17123), .B(n17124), .Z(n17115) );
  XNOR U18872 ( .A(n17116), .B(n17115), .Z(n17117) );
  XNOR U18873 ( .A(n17118), .B(n17117), .Z(n17147) );
  XNOR U18874 ( .A(sreg[1368]), .B(n17147), .Z(n17149) );
  NANDN U18875 ( .A(sreg[1367]), .B(n17110), .Z(n17114) );
  NAND U18876 ( .A(n17112), .B(n17111), .Z(n17113) );
  NAND U18877 ( .A(n17114), .B(n17113), .Z(n17148) );
  XNOR U18878 ( .A(n17149), .B(n17148), .Z(c[1368]) );
  NANDN U18879 ( .A(n17116), .B(n17115), .Z(n17120) );
  NANDN U18880 ( .A(n17118), .B(n17117), .Z(n17119) );
  AND U18881 ( .A(n17120), .B(n17119), .Z(n17155) );
  NANDN U18882 ( .A(n17122), .B(n17121), .Z(n17126) );
  NANDN U18883 ( .A(n17124), .B(n17123), .Z(n17125) );
  AND U18884 ( .A(n17126), .B(n17125), .Z(n17153) );
  NAND U18885 ( .A(n42143), .B(n17127), .Z(n17129) );
  XNOR U18886 ( .A(a[347]), .B(n4121), .Z(n17164) );
  NAND U18887 ( .A(n42144), .B(n17164), .Z(n17128) );
  AND U18888 ( .A(n17129), .B(n17128), .Z(n17179) );
  XOR U18889 ( .A(a[351]), .B(n42012), .Z(n17167) );
  XNOR U18890 ( .A(n17179), .B(n17178), .Z(n17181) );
  AND U18891 ( .A(a[353]), .B(b[0]), .Z(n17131) );
  XNOR U18892 ( .A(n17131), .B(n4071), .Z(n17133) );
  NANDN U18893 ( .A(b[0]), .B(a[352]), .Z(n17132) );
  NAND U18894 ( .A(n17133), .B(n17132), .Z(n17175) );
  XOR U18895 ( .A(a[349]), .B(n42085), .Z(n17168) );
  AND U18896 ( .A(a[345]), .B(b[7]), .Z(n17172) );
  XNOR U18897 ( .A(n17173), .B(n17172), .Z(n17174) );
  XNOR U18898 ( .A(n17175), .B(n17174), .Z(n17180) );
  XOR U18899 ( .A(n17181), .B(n17180), .Z(n17159) );
  NANDN U18900 ( .A(n17136), .B(n17135), .Z(n17140) );
  NANDN U18901 ( .A(n17138), .B(n17137), .Z(n17139) );
  AND U18902 ( .A(n17140), .B(n17139), .Z(n17158) );
  XNOR U18903 ( .A(n17159), .B(n17158), .Z(n17160) );
  NANDN U18904 ( .A(n17142), .B(n17141), .Z(n17146) );
  NAND U18905 ( .A(n17144), .B(n17143), .Z(n17145) );
  NAND U18906 ( .A(n17146), .B(n17145), .Z(n17161) );
  XNOR U18907 ( .A(n17160), .B(n17161), .Z(n17152) );
  XNOR U18908 ( .A(n17153), .B(n17152), .Z(n17154) );
  XNOR U18909 ( .A(n17155), .B(n17154), .Z(n17184) );
  XNOR U18910 ( .A(sreg[1369]), .B(n17184), .Z(n17186) );
  NANDN U18911 ( .A(sreg[1368]), .B(n17147), .Z(n17151) );
  NAND U18912 ( .A(n17149), .B(n17148), .Z(n17150) );
  NAND U18913 ( .A(n17151), .B(n17150), .Z(n17185) );
  XNOR U18914 ( .A(n17186), .B(n17185), .Z(c[1369]) );
  NANDN U18915 ( .A(n17153), .B(n17152), .Z(n17157) );
  NANDN U18916 ( .A(n17155), .B(n17154), .Z(n17156) );
  AND U18917 ( .A(n17157), .B(n17156), .Z(n17192) );
  NANDN U18918 ( .A(n17159), .B(n17158), .Z(n17163) );
  NANDN U18919 ( .A(n17161), .B(n17160), .Z(n17162) );
  AND U18920 ( .A(n17163), .B(n17162), .Z(n17190) );
  NAND U18921 ( .A(n42143), .B(n17164), .Z(n17166) );
  XNOR U18922 ( .A(a[348]), .B(n4121), .Z(n17201) );
  NAND U18923 ( .A(n42144), .B(n17201), .Z(n17165) );
  AND U18924 ( .A(n17166), .B(n17165), .Z(n17216) );
  XOR U18925 ( .A(a[352]), .B(n42012), .Z(n17204) );
  XNOR U18926 ( .A(n17216), .B(n17215), .Z(n17218) );
  XOR U18927 ( .A(a[350]), .B(n42085), .Z(n17208) );
  AND U18928 ( .A(a[346]), .B(b[7]), .Z(n17209) );
  XNOR U18929 ( .A(n17210), .B(n17209), .Z(n17211) );
  AND U18930 ( .A(a[354]), .B(b[0]), .Z(n17169) );
  XNOR U18931 ( .A(n17169), .B(n4071), .Z(n17171) );
  NANDN U18932 ( .A(b[0]), .B(a[353]), .Z(n17170) );
  NAND U18933 ( .A(n17171), .B(n17170), .Z(n17212) );
  XNOR U18934 ( .A(n17211), .B(n17212), .Z(n17217) );
  XOR U18935 ( .A(n17218), .B(n17217), .Z(n17196) );
  NANDN U18936 ( .A(n17173), .B(n17172), .Z(n17177) );
  NANDN U18937 ( .A(n17175), .B(n17174), .Z(n17176) );
  AND U18938 ( .A(n17177), .B(n17176), .Z(n17195) );
  XNOR U18939 ( .A(n17196), .B(n17195), .Z(n17197) );
  NANDN U18940 ( .A(n17179), .B(n17178), .Z(n17183) );
  NAND U18941 ( .A(n17181), .B(n17180), .Z(n17182) );
  NAND U18942 ( .A(n17183), .B(n17182), .Z(n17198) );
  XNOR U18943 ( .A(n17197), .B(n17198), .Z(n17189) );
  XNOR U18944 ( .A(n17190), .B(n17189), .Z(n17191) );
  XNOR U18945 ( .A(n17192), .B(n17191), .Z(n17221) );
  XNOR U18946 ( .A(sreg[1370]), .B(n17221), .Z(n17223) );
  NANDN U18947 ( .A(sreg[1369]), .B(n17184), .Z(n17188) );
  NAND U18948 ( .A(n17186), .B(n17185), .Z(n17187) );
  NAND U18949 ( .A(n17188), .B(n17187), .Z(n17222) );
  XNOR U18950 ( .A(n17223), .B(n17222), .Z(c[1370]) );
  NANDN U18951 ( .A(n17190), .B(n17189), .Z(n17194) );
  NANDN U18952 ( .A(n17192), .B(n17191), .Z(n17193) );
  AND U18953 ( .A(n17194), .B(n17193), .Z(n17229) );
  NANDN U18954 ( .A(n17196), .B(n17195), .Z(n17200) );
  NANDN U18955 ( .A(n17198), .B(n17197), .Z(n17199) );
  AND U18956 ( .A(n17200), .B(n17199), .Z(n17227) );
  NAND U18957 ( .A(n42143), .B(n17201), .Z(n17203) );
  XNOR U18958 ( .A(a[349]), .B(n4121), .Z(n17238) );
  NAND U18959 ( .A(n42144), .B(n17238), .Z(n17202) );
  AND U18960 ( .A(n17203), .B(n17202), .Z(n17253) );
  XOR U18961 ( .A(a[353]), .B(n42012), .Z(n17241) );
  XNOR U18962 ( .A(n17253), .B(n17252), .Z(n17255) );
  AND U18963 ( .A(a[355]), .B(b[0]), .Z(n17205) );
  XNOR U18964 ( .A(n17205), .B(n4071), .Z(n17207) );
  NANDN U18965 ( .A(b[0]), .B(a[354]), .Z(n17206) );
  NAND U18966 ( .A(n17207), .B(n17206), .Z(n17249) );
  XOR U18967 ( .A(a[351]), .B(n42085), .Z(n17242) );
  AND U18968 ( .A(a[347]), .B(b[7]), .Z(n17246) );
  XNOR U18969 ( .A(n17247), .B(n17246), .Z(n17248) );
  XNOR U18970 ( .A(n17249), .B(n17248), .Z(n17254) );
  XOR U18971 ( .A(n17255), .B(n17254), .Z(n17233) );
  NANDN U18972 ( .A(n17210), .B(n17209), .Z(n17214) );
  NANDN U18973 ( .A(n17212), .B(n17211), .Z(n17213) );
  AND U18974 ( .A(n17214), .B(n17213), .Z(n17232) );
  XNOR U18975 ( .A(n17233), .B(n17232), .Z(n17234) );
  NANDN U18976 ( .A(n17216), .B(n17215), .Z(n17220) );
  NAND U18977 ( .A(n17218), .B(n17217), .Z(n17219) );
  NAND U18978 ( .A(n17220), .B(n17219), .Z(n17235) );
  XNOR U18979 ( .A(n17234), .B(n17235), .Z(n17226) );
  XNOR U18980 ( .A(n17227), .B(n17226), .Z(n17228) );
  XNOR U18981 ( .A(n17229), .B(n17228), .Z(n17258) );
  XNOR U18982 ( .A(sreg[1371]), .B(n17258), .Z(n17260) );
  NANDN U18983 ( .A(sreg[1370]), .B(n17221), .Z(n17225) );
  NAND U18984 ( .A(n17223), .B(n17222), .Z(n17224) );
  NAND U18985 ( .A(n17225), .B(n17224), .Z(n17259) );
  XNOR U18986 ( .A(n17260), .B(n17259), .Z(c[1371]) );
  NANDN U18987 ( .A(n17227), .B(n17226), .Z(n17231) );
  NANDN U18988 ( .A(n17229), .B(n17228), .Z(n17230) );
  AND U18989 ( .A(n17231), .B(n17230), .Z(n17266) );
  NANDN U18990 ( .A(n17233), .B(n17232), .Z(n17237) );
  NANDN U18991 ( .A(n17235), .B(n17234), .Z(n17236) );
  AND U18992 ( .A(n17237), .B(n17236), .Z(n17264) );
  NAND U18993 ( .A(n42143), .B(n17238), .Z(n17240) );
  XNOR U18994 ( .A(a[350]), .B(n4121), .Z(n17275) );
  NAND U18995 ( .A(n42144), .B(n17275), .Z(n17239) );
  AND U18996 ( .A(n17240), .B(n17239), .Z(n17290) );
  XOR U18997 ( .A(a[354]), .B(n42012), .Z(n17278) );
  XNOR U18998 ( .A(n17290), .B(n17289), .Z(n17292) );
  XOR U18999 ( .A(a[352]), .B(n42085), .Z(n17282) );
  AND U19000 ( .A(a[348]), .B(b[7]), .Z(n17283) );
  XNOR U19001 ( .A(n17284), .B(n17283), .Z(n17285) );
  AND U19002 ( .A(a[356]), .B(b[0]), .Z(n17243) );
  XNOR U19003 ( .A(n17243), .B(n4071), .Z(n17245) );
  NANDN U19004 ( .A(b[0]), .B(a[355]), .Z(n17244) );
  NAND U19005 ( .A(n17245), .B(n17244), .Z(n17286) );
  XNOR U19006 ( .A(n17285), .B(n17286), .Z(n17291) );
  XOR U19007 ( .A(n17292), .B(n17291), .Z(n17270) );
  NANDN U19008 ( .A(n17247), .B(n17246), .Z(n17251) );
  NANDN U19009 ( .A(n17249), .B(n17248), .Z(n17250) );
  AND U19010 ( .A(n17251), .B(n17250), .Z(n17269) );
  XNOR U19011 ( .A(n17270), .B(n17269), .Z(n17271) );
  NANDN U19012 ( .A(n17253), .B(n17252), .Z(n17257) );
  NAND U19013 ( .A(n17255), .B(n17254), .Z(n17256) );
  NAND U19014 ( .A(n17257), .B(n17256), .Z(n17272) );
  XNOR U19015 ( .A(n17271), .B(n17272), .Z(n17263) );
  XNOR U19016 ( .A(n17264), .B(n17263), .Z(n17265) );
  XNOR U19017 ( .A(n17266), .B(n17265), .Z(n17295) );
  XNOR U19018 ( .A(sreg[1372]), .B(n17295), .Z(n17297) );
  NANDN U19019 ( .A(sreg[1371]), .B(n17258), .Z(n17262) );
  NAND U19020 ( .A(n17260), .B(n17259), .Z(n17261) );
  NAND U19021 ( .A(n17262), .B(n17261), .Z(n17296) );
  XNOR U19022 ( .A(n17297), .B(n17296), .Z(c[1372]) );
  NANDN U19023 ( .A(n17264), .B(n17263), .Z(n17268) );
  NANDN U19024 ( .A(n17266), .B(n17265), .Z(n17267) );
  AND U19025 ( .A(n17268), .B(n17267), .Z(n17303) );
  NANDN U19026 ( .A(n17270), .B(n17269), .Z(n17274) );
  NANDN U19027 ( .A(n17272), .B(n17271), .Z(n17273) );
  AND U19028 ( .A(n17274), .B(n17273), .Z(n17301) );
  NAND U19029 ( .A(n42143), .B(n17275), .Z(n17277) );
  XNOR U19030 ( .A(a[351]), .B(n4122), .Z(n17312) );
  NAND U19031 ( .A(n42144), .B(n17312), .Z(n17276) );
  AND U19032 ( .A(n17277), .B(n17276), .Z(n17327) );
  XOR U19033 ( .A(a[355]), .B(n42012), .Z(n17315) );
  XNOR U19034 ( .A(n17327), .B(n17326), .Z(n17329) );
  AND U19035 ( .A(a[357]), .B(b[0]), .Z(n17279) );
  XNOR U19036 ( .A(n17279), .B(n4071), .Z(n17281) );
  NANDN U19037 ( .A(b[0]), .B(a[356]), .Z(n17280) );
  NAND U19038 ( .A(n17281), .B(n17280), .Z(n17323) );
  XOR U19039 ( .A(a[353]), .B(n42085), .Z(n17319) );
  AND U19040 ( .A(a[349]), .B(b[7]), .Z(n17320) );
  XNOR U19041 ( .A(n17321), .B(n17320), .Z(n17322) );
  XNOR U19042 ( .A(n17323), .B(n17322), .Z(n17328) );
  XOR U19043 ( .A(n17329), .B(n17328), .Z(n17307) );
  NANDN U19044 ( .A(n17284), .B(n17283), .Z(n17288) );
  NANDN U19045 ( .A(n17286), .B(n17285), .Z(n17287) );
  AND U19046 ( .A(n17288), .B(n17287), .Z(n17306) );
  XNOR U19047 ( .A(n17307), .B(n17306), .Z(n17308) );
  NANDN U19048 ( .A(n17290), .B(n17289), .Z(n17294) );
  NAND U19049 ( .A(n17292), .B(n17291), .Z(n17293) );
  NAND U19050 ( .A(n17294), .B(n17293), .Z(n17309) );
  XNOR U19051 ( .A(n17308), .B(n17309), .Z(n17300) );
  XNOR U19052 ( .A(n17301), .B(n17300), .Z(n17302) );
  XNOR U19053 ( .A(n17303), .B(n17302), .Z(n17332) );
  XNOR U19054 ( .A(sreg[1373]), .B(n17332), .Z(n17334) );
  NANDN U19055 ( .A(sreg[1372]), .B(n17295), .Z(n17299) );
  NAND U19056 ( .A(n17297), .B(n17296), .Z(n17298) );
  NAND U19057 ( .A(n17299), .B(n17298), .Z(n17333) );
  XNOR U19058 ( .A(n17334), .B(n17333), .Z(c[1373]) );
  NANDN U19059 ( .A(n17301), .B(n17300), .Z(n17305) );
  NANDN U19060 ( .A(n17303), .B(n17302), .Z(n17304) );
  AND U19061 ( .A(n17305), .B(n17304), .Z(n17340) );
  NANDN U19062 ( .A(n17307), .B(n17306), .Z(n17311) );
  NANDN U19063 ( .A(n17309), .B(n17308), .Z(n17310) );
  AND U19064 ( .A(n17311), .B(n17310), .Z(n17338) );
  NAND U19065 ( .A(n42143), .B(n17312), .Z(n17314) );
  XNOR U19066 ( .A(a[352]), .B(n4122), .Z(n17349) );
  NAND U19067 ( .A(n42144), .B(n17349), .Z(n17313) );
  AND U19068 ( .A(n17314), .B(n17313), .Z(n17364) );
  XOR U19069 ( .A(a[356]), .B(n42012), .Z(n17352) );
  XNOR U19070 ( .A(n17364), .B(n17363), .Z(n17366) );
  AND U19071 ( .A(a[358]), .B(b[0]), .Z(n17316) );
  XNOR U19072 ( .A(n17316), .B(n4071), .Z(n17318) );
  NANDN U19073 ( .A(b[0]), .B(a[357]), .Z(n17317) );
  NAND U19074 ( .A(n17318), .B(n17317), .Z(n17360) );
  XOR U19075 ( .A(a[354]), .B(n42085), .Z(n17356) );
  AND U19076 ( .A(a[350]), .B(b[7]), .Z(n17357) );
  XNOR U19077 ( .A(n17358), .B(n17357), .Z(n17359) );
  XNOR U19078 ( .A(n17360), .B(n17359), .Z(n17365) );
  XOR U19079 ( .A(n17366), .B(n17365), .Z(n17344) );
  NANDN U19080 ( .A(n17321), .B(n17320), .Z(n17325) );
  NANDN U19081 ( .A(n17323), .B(n17322), .Z(n17324) );
  AND U19082 ( .A(n17325), .B(n17324), .Z(n17343) );
  XNOR U19083 ( .A(n17344), .B(n17343), .Z(n17345) );
  NANDN U19084 ( .A(n17327), .B(n17326), .Z(n17331) );
  NAND U19085 ( .A(n17329), .B(n17328), .Z(n17330) );
  NAND U19086 ( .A(n17331), .B(n17330), .Z(n17346) );
  XNOR U19087 ( .A(n17345), .B(n17346), .Z(n17337) );
  XNOR U19088 ( .A(n17338), .B(n17337), .Z(n17339) );
  XNOR U19089 ( .A(n17340), .B(n17339), .Z(n17369) );
  XNOR U19090 ( .A(sreg[1374]), .B(n17369), .Z(n17371) );
  NANDN U19091 ( .A(sreg[1373]), .B(n17332), .Z(n17336) );
  NAND U19092 ( .A(n17334), .B(n17333), .Z(n17335) );
  NAND U19093 ( .A(n17336), .B(n17335), .Z(n17370) );
  XNOR U19094 ( .A(n17371), .B(n17370), .Z(c[1374]) );
  NANDN U19095 ( .A(n17338), .B(n17337), .Z(n17342) );
  NANDN U19096 ( .A(n17340), .B(n17339), .Z(n17341) );
  AND U19097 ( .A(n17342), .B(n17341), .Z(n17377) );
  NANDN U19098 ( .A(n17344), .B(n17343), .Z(n17348) );
  NANDN U19099 ( .A(n17346), .B(n17345), .Z(n17347) );
  AND U19100 ( .A(n17348), .B(n17347), .Z(n17375) );
  NAND U19101 ( .A(n42143), .B(n17349), .Z(n17351) );
  XNOR U19102 ( .A(a[353]), .B(n4122), .Z(n17386) );
  NAND U19103 ( .A(n42144), .B(n17386), .Z(n17350) );
  AND U19104 ( .A(n17351), .B(n17350), .Z(n17401) );
  XOR U19105 ( .A(a[357]), .B(n42012), .Z(n17389) );
  XNOR U19106 ( .A(n17401), .B(n17400), .Z(n17403) );
  AND U19107 ( .A(a[359]), .B(b[0]), .Z(n17353) );
  XNOR U19108 ( .A(n17353), .B(n4071), .Z(n17355) );
  NANDN U19109 ( .A(b[0]), .B(a[358]), .Z(n17354) );
  NAND U19110 ( .A(n17355), .B(n17354), .Z(n17397) );
  XOR U19111 ( .A(a[355]), .B(n42085), .Z(n17390) );
  AND U19112 ( .A(a[351]), .B(b[7]), .Z(n17394) );
  XNOR U19113 ( .A(n17395), .B(n17394), .Z(n17396) );
  XNOR U19114 ( .A(n17397), .B(n17396), .Z(n17402) );
  XOR U19115 ( .A(n17403), .B(n17402), .Z(n17381) );
  NANDN U19116 ( .A(n17358), .B(n17357), .Z(n17362) );
  NANDN U19117 ( .A(n17360), .B(n17359), .Z(n17361) );
  AND U19118 ( .A(n17362), .B(n17361), .Z(n17380) );
  XNOR U19119 ( .A(n17381), .B(n17380), .Z(n17382) );
  NANDN U19120 ( .A(n17364), .B(n17363), .Z(n17368) );
  NAND U19121 ( .A(n17366), .B(n17365), .Z(n17367) );
  NAND U19122 ( .A(n17368), .B(n17367), .Z(n17383) );
  XNOR U19123 ( .A(n17382), .B(n17383), .Z(n17374) );
  XNOR U19124 ( .A(n17375), .B(n17374), .Z(n17376) );
  XNOR U19125 ( .A(n17377), .B(n17376), .Z(n17406) );
  XNOR U19126 ( .A(sreg[1375]), .B(n17406), .Z(n17408) );
  NANDN U19127 ( .A(sreg[1374]), .B(n17369), .Z(n17373) );
  NAND U19128 ( .A(n17371), .B(n17370), .Z(n17372) );
  NAND U19129 ( .A(n17373), .B(n17372), .Z(n17407) );
  XNOR U19130 ( .A(n17408), .B(n17407), .Z(c[1375]) );
  NANDN U19131 ( .A(n17375), .B(n17374), .Z(n17379) );
  NANDN U19132 ( .A(n17377), .B(n17376), .Z(n17378) );
  AND U19133 ( .A(n17379), .B(n17378), .Z(n17414) );
  NANDN U19134 ( .A(n17381), .B(n17380), .Z(n17385) );
  NANDN U19135 ( .A(n17383), .B(n17382), .Z(n17384) );
  AND U19136 ( .A(n17385), .B(n17384), .Z(n17412) );
  NAND U19137 ( .A(n42143), .B(n17386), .Z(n17388) );
  XNOR U19138 ( .A(a[354]), .B(n4122), .Z(n17423) );
  NAND U19139 ( .A(n42144), .B(n17423), .Z(n17387) );
  AND U19140 ( .A(n17388), .B(n17387), .Z(n17438) );
  XOR U19141 ( .A(a[358]), .B(n42012), .Z(n17426) );
  XNOR U19142 ( .A(n17438), .B(n17437), .Z(n17440) );
  XOR U19143 ( .A(a[356]), .B(n42085), .Z(n17430) );
  AND U19144 ( .A(a[352]), .B(b[7]), .Z(n17431) );
  XNOR U19145 ( .A(n17432), .B(n17431), .Z(n17433) );
  AND U19146 ( .A(a[360]), .B(b[0]), .Z(n17391) );
  XNOR U19147 ( .A(n17391), .B(n4071), .Z(n17393) );
  NANDN U19148 ( .A(b[0]), .B(a[359]), .Z(n17392) );
  NAND U19149 ( .A(n17393), .B(n17392), .Z(n17434) );
  XNOR U19150 ( .A(n17433), .B(n17434), .Z(n17439) );
  XOR U19151 ( .A(n17440), .B(n17439), .Z(n17418) );
  NANDN U19152 ( .A(n17395), .B(n17394), .Z(n17399) );
  NANDN U19153 ( .A(n17397), .B(n17396), .Z(n17398) );
  AND U19154 ( .A(n17399), .B(n17398), .Z(n17417) );
  XNOR U19155 ( .A(n17418), .B(n17417), .Z(n17419) );
  NANDN U19156 ( .A(n17401), .B(n17400), .Z(n17405) );
  NAND U19157 ( .A(n17403), .B(n17402), .Z(n17404) );
  NAND U19158 ( .A(n17405), .B(n17404), .Z(n17420) );
  XNOR U19159 ( .A(n17419), .B(n17420), .Z(n17411) );
  XNOR U19160 ( .A(n17412), .B(n17411), .Z(n17413) );
  XNOR U19161 ( .A(n17414), .B(n17413), .Z(n17443) );
  XNOR U19162 ( .A(sreg[1376]), .B(n17443), .Z(n17445) );
  NANDN U19163 ( .A(sreg[1375]), .B(n17406), .Z(n17410) );
  NAND U19164 ( .A(n17408), .B(n17407), .Z(n17409) );
  NAND U19165 ( .A(n17410), .B(n17409), .Z(n17444) );
  XNOR U19166 ( .A(n17445), .B(n17444), .Z(c[1376]) );
  NANDN U19167 ( .A(n17412), .B(n17411), .Z(n17416) );
  NANDN U19168 ( .A(n17414), .B(n17413), .Z(n17415) );
  AND U19169 ( .A(n17416), .B(n17415), .Z(n17451) );
  NANDN U19170 ( .A(n17418), .B(n17417), .Z(n17422) );
  NANDN U19171 ( .A(n17420), .B(n17419), .Z(n17421) );
  AND U19172 ( .A(n17422), .B(n17421), .Z(n17449) );
  NAND U19173 ( .A(n42143), .B(n17423), .Z(n17425) );
  XNOR U19174 ( .A(a[355]), .B(n4122), .Z(n17460) );
  NAND U19175 ( .A(n42144), .B(n17460), .Z(n17424) );
  AND U19176 ( .A(n17425), .B(n17424), .Z(n17475) );
  XOR U19177 ( .A(a[359]), .B(n42012), .Z(n17463) );
  XNOR U19178 ( .A(n17475), .B(n17474), .Z(n17477) );
  AND U19179 ( .A(a[361]), .B(b[0]), .Z(n17427) );
  XNOR U19180 ( .A(n17427), .B(n4071), .Z(n17429) );
  NANDN U19181 ( .A(b[0]), .B(a[360]), .Z(n17428) );
  NAND U19182 ( .A(n17429), .B(n17428), .Z(n17471) );
  XOR U19183 ( .A(a[357]), .B(n42085), .Z(n17467) );
  AND U19184 ( .A(a[353]), .B(b[7]), .Z(n17468) );
  XNOR U19185 ( .A(n17469), .B(n17468), .Z(n17470) );
  XNOR U19186 ( .A(n17471), .B(n17470), .Z(n17476) );
  XOR U19187 ( .A(n17477), .B(n17476), .Z(n17455) );
  NANDN U19188 ( .A(n17432), .B(n17431), .Z(n17436) );
  NANDN U19189 ( .A(n17434), .B(n17433), .Z(n17435) );
  AND U19190 ( .A(n17436), .B(n17435), .Z(n17454) );
  XNOR U19191 ( .A(n17455), .B(n17454), .Z(n17456) );
  NANDN U19192 ( .A(n17438), .B(n17437), .Z(n17442) );
  NAND U19193 ( .A(n17440), .B(n17439), .Z(n17441) );
  NAND U19194 ( .A(n17442), .B(n17441), .Z(n17457) );
  XNOR U19195 ( .A(n17456), .B(n17457), .Z(n17448) );
  XNOR U19196 ( .A(n17449), .B(n17448), .Z(n17450) );
  XNOR U19197 ( .A(n17451), .B(n17450), .Z(n17480) );
  XNOR U19198 ( .A(sreg[1377]), .B(n17480), .Z(n17482) );
  NANDN U19199 ( .A(sreg[1376]), .B(n17443), .Z(n17447) );
  NAND U19200 ( .A(n17445), .B(n17444), .Z(n17446) );
  NAND U19201 ( .A(n17447), .B(n17446), .Z(n17481) );
  XNOR U19202 ( .A(n17482), .B(n17481), .Z(c[1377]) );
  NANDN U19203 ( .A(n17449), .B(n17448), .Z(n17453) );
  NANDN U19204 ( .A(n17451), .B(n17450), .Z(n17452) );
  AND U19205 ( .A(n17453), .B(n17452), .Z(n17488) );
  NANDN U19206 ( .A(n17455), .B(n17454), .Z(n17459) );
  NANDN U19207 ( .A(n17457), .B(n17456), .Z(n17458) );
  AND U19208 ( .A(n17459), .B(n17458), .Z(n17486) );
  NAND U19209 ( .A(n42143), .B(n17460), .Z(n17462) );
  XNOR U19210 ( .A(a[356]), .B(n4122), .Z(n17497) );
  NAND U19211 ( .A(n42144), .B(n17497), .Z(n17461) );
  AND U19212 ( .A(n17462), .B(n17461), .Z(n17512) );
  XOR U19213 ( .A(a[360]), .B(n42012), .Z(n17500) );
  XNOR U19214 ( .A(n17512), .B(n17511), .Z(n17514) );
  AND U19215 ( .A(a[362]), .B(b[0]), .Z(n17464) );
  XNOR U19216 ( .A(n17464), .B(n4071), .Z(n17466) );
  NANDN U19217 ( .A(b[0]), .B(a[361]), .Z(n17465) );
  NAND U19218 ( .A(n17466), .B(n17465), .Z(n17508) );
  XOR U19219 ( .A(a[358]), .B(n42085), .Z(n17504) );
  AND U19220 ( .A(a[354]), .B(b[7]), .Z(n17505) );
  XNOR U19221 ( .A(n17506), .B(n17505), .Z(n17507) );
  XNOR U19222 ( .A(n17508), .B(n17507), .Z(n17513) );
  XOR U19223 ( .A(n17514), .B(n17513), .Z(n17492) );
  NANDN U19224 ( .A(n17469), .B(n17468), .Z(n17473) );
  NANDN U19225 ( .A(n17471), .B(n17470), .Z(n17472) );
  AND U19226 ( .A(n17473), .B(n17472), .Z(n17491) );
  XNOR U19227 ( .A(n17492), .B(n17491), .Z(n17493) );
  NANDN U19228 ( .A(n17475), .B(n17474), .Z(n17479) );
  NAND U19229 ( .A(n17477), .B(n17476), .Z(n17478) );
  NAND U19230 ( .A(n17479), .B(n17478), .Z(n17494) );
  XNOR U19231 ( .A(n17493), .B(n17494), .Z(n17485) );
  XNOR U19232 ( .A(n17486), .B(n17485), .Z(n17487) );
  XNOR U19233 ( .A(n17488), .B(n17487), .Z(n17517) );
  XNOR U19234 ( .A(sreg[1378]), .B(n17517), .Z(n17519) );
  NANDN U19235 ( .A(sreg[1377]), .B(n17480), .Z(n17484) );
  NAND U19236 ( .A(n17482), .B(n17481), .Z(n17483) );
  NAND U19237 ( .A(n17484), .B(n17483), .Z(n17518) );
  XNOR U19238 ( .A(n17519), .B(n17518), .Z(c[1378]) );
  NANDN U19239 ( .A(n17486), .B(n17485), .Z(n17490) );
  NANDN U19240 ( .A(n17488), .B(n17487), .Z(n17489) );
  AND U19241 ( .A(n17490), .B(n17489), .Z(n17525) );
  NANDN U19242 ( .A(n17492), .B(n17491), .Z(n17496) );
  NANDN U19243 ( .A(n17494), .B(n17493), .Z(n17495) );
  AND U19244 ( .A(n17496), .B(n17495), .Z(n17523) );
  NAND U19245 ( .A(n42143), .B(n17497), .Z(n17499) );
  XNOR U19246 ( .A(a[357]), .B(n4122), .Z(n17534) );
  NAND U19247 ( .A(n42144), .B(n17534), .Z(n17498) );
  AND U19248 ( .A(n17499), .B(n17498), .Z(n17549) );
  XOR U19249 ( .A(a[361]), .B(n42012), .Z(n17537) );
  XNOR U19250 ( .A(n17549), .B(n17548), .Z(n17551) );
  AND U19251 ( .A(a[363]), .B(b[0]), .Z(n17501) );
  XNOR U19252 ( .A(n17501), .B(n4071), .Z(n17503) );
  NANDN U19253 ( .A(b[0]), .B(a[362]), .Z(n17502) );
  NAND U19254 ( .A(n17503), .B(n17502), .Z(n17545) );
  XOR U19255 ( .A(a[359]), .B(n42085), .Z(n17541) );
  AND U19256 ( .A(a[355]), .B(b[7]), .Z(n17542) );
  XNOR U19257 ( .A(n17543), .B(n17542), .Z(n17544) );
  XNOR U19258 ( .A(n17545), .B(n17544), .Z(n17550) );
  XOR U19259 ( .A(n17551), .B(n17550), .Z(n17529) );
  NANDN U19260 ( .A(n17506), .B(n17505), .Z(n17510) );
  NANDN U19261 ( .A(n17508), .B(n17507), .Z(n17509) );
  AND U19262 ( .A(n17510), .B(n17509), .Z(n17528) );
  XNOR U19263 ( .A(n17529), .B(n17528), .Z(n17530) );
  NANDN U19264 ( .A(n17512), .B(n17511), .Z(n17516) );
  NAND U19265 ( .A(n17514), .B(n17513), .Z(n17515) );
  NAND U19266 ( .A(n17516), .B(n17515), .Z(n17531) );
  XNOR U19267 ( .A(n17530), .B(n17531), .Z(n17522) );
  XNOR U19268 ( .A(n17523), .B(n17522), .Z(n17524) );
  XNOR U19269 ( .A(n17525), .B(n17524), .Z(n17554) );
  XNOR U19270 ( .A(sreg[1379]), .B(n17554), .Z(n17556) );
  NANDN U19271 ( .A(sreg[1378]), .B(n17517), .Z(n17521) );
  NAND U19272 ( .A(n17519), .B(n17518), .Z(n17520) );
  NAND U19273 ( .A(n17521), .B(n17520), .Z(n17555) );
  XNOR U19274 ( .A(n17556), .B(n17555), .Z(c[1379]) );
  NANDN U19275 ( .A(n17523), .B(n17522), .Z(n17527) );
  NANDN U19276 ( .A(n17525), .B(n17524), .Z(n17526) );
  AND U19277 ( .A(n17527), .B(n17526), .Z(n17562) );
  NANDN U19278 ( .A(n17529), .B(n17528), .Z(n17533) );
  NANDN U19279 ( .A(n17531), .B(n17530), .Z(n17532) );
  AND U19280 ( .A(n17533), .B(n17532), .Z(n17560) );
  NAND U19281 ( .A(n42143), .B(n17534), .Z(n17536) );
  XNOR U19282 ( .A(a[358]), .B(n4123), .Z(n17571) );
  NAND U19283 ( .A(n42144), .B(n17571), .Z(n17535) );
  AND U19284 ( .A(n17536), .B(n17535), .Z(n17586) );
  XOR U19285 ( .A(a[362]), .B(n42012), .Z(n17574) );
  XNOR U19286 ( .A(n17586), .B(n17585), .Z(n17588) );
  AND U19287 ( .A(a[364]), .B(b[0]), .Z(n17538) );
  XNOR U19288 ( .A(n17538), .B(n4071), .Z(n17540) );
  NANDN U19289 ( .A(b[0]), .B(a[363]), .Z(n17539) );
  NAND U19290 ( .A(n17540), .B(n17539), .Z(n17582) );
  XOR U19291 ( .A(a[360]), .B(n42085), .Z(n17578) );
  AND U19292 ( .A(a[356]), .B(b[7]), .Z(n17579) );
  XNOR U19293 ( .A(n17580), .B(n17579), .Z(n17581) );
  XNOR U19294 ( .A(n17582), .B(n17581), .Z(n17587) );
  XOR U19295 ( .A(n17588), .B(n17587), .Z(n17566) );
  NANDN U19296 ( .A(n17543), .B(n17542), .Z(n17547) );
  NANDN U19297 ( .A(n17545), .B(n17544), .Z(n17546) );
  AND U19298 ( .A(n17547), .B(n17546), .Z(n17565) );
  XNOR U19299 ( .A(n17566), .B(n17565), .Z(n17567) );
  NANDN U19300 ( .A(n17549), .B(n17548), .Z(n17553) );
  NAND U19301 ( .A(n17551), .B(n17550), .Z(n17552) );
  NAND U19302 ( .A(n17553), .B(n17552), .Z(n17568) );
  XNOR U19303 ( .A(n17567), .B(n17568), .Z(n17559) );
  XNOR U19304 ( .A(n17560), .B(n17559), .Z(n17561) );
  XNOR U19305 ( .A(n17562), .B(n17561), .Z(n17591) );
  XNOR U19306 ( .A(sreg[1380]), .B(n17591), .Z(n17593) );
  NANDN U19307 ( .A(sreg[1379]), .B(n17554), .Z(n17558) );
  NAND U19308 ( .A(n17556), .B(n17555), .Z(n17557) );
  NAND U19309 ( .A(n17558), .B(n17557), .Z(n17592) );
  XNOR U19310 ( .A(n17593), .B(n17592), .Z(c[1380]) );
  NANDN U19311 ( .A(n17560), .B(n17559), .Z(n17564) );
  NANDN U19312 ( .A(n17562), .B(n17561), .Z(n17563) );
  AND U19313 ( .A(n17564), .B(n17563), .Z(n17599) );
  NANDN U19314 ( .A(n17566), .B(n17565), .Z(n17570) );
  NANDN U19315 ( .A(n17568), .B(n17567), .Z(n17569) );
  AND U19316 ( .A(n17570), .B(n17569), .Z(n17597) );
  NAND U19317 ( .A(n42143), .B(n17571), .Z(n17573) );
  XNOR U19318 ( .A(a[359]), .B(n4123), .Z(n17608) );
  NAND U19319 ( .A(n42144), .B(n17608), .Z(n17572) );
  AND U19320 ( .A(n17573), .B(n17572), .Z(n17623) );
  XOR U19321 ( .A(a[363]), .B(n42012), .Z(n17611) );
  XNOR U19322 ( .A(n17623), .B(n17622), .Z(n17625) );
  AND U19323 ( .A(b[0]), .B(a[365]), .Z(n17575) );
  XOR U19324 ( .A(b[1]), .B(n17575), .Z(n17577) );
  NANDN U19325 ( .A(b[0]), .B(a[364]), .Z(n17576) );
  AND U19326 ( .A(n17577), .B(n17576), .Z(n17618) );
  XOR U19327 ( .A(a[361]), .B(n42085), .Z(n17615) );
  AND U19328 ( .A(a[357]), .B(b[7]), .Z(n17616) );
  XOR U19329 ( .A(n17617), .B(n17616), .Z(n17619) );
  XNOR U19330 ( .A(n17618), .B(n17619), .Z(n17624) );
  XOR U19331 ( .A(n17625), .B(n17624), .Z(n17603) );
  NANDN U19332 ( .A(n17580), .B(n17579), .Z(n17584) );
  NANDN U19333 ( .A(n17582), .B(n17581), .Z(n17583) );
  AND U19334 ( .A(n17584), .B(n17583), .Z(n17602) );
  XNOR U19335 ( .A(n17603), .B(n17602), .Z(n17604) );
  NANDN U19336 ( .A(n17586), .B(n17585), .Z(n17590) );
  NAND U19337 ( .A(n17588), .B(n17587), .Z(n17589) );
  NAND U19338 ( .A(n17590), .B(n17589), .Z(n17605) );
  XNOR U19339 ( .A(n17604), .B(n17605), .Z(n17596) );
  XNOR U19340 ( .A(n17597), .B(n17596), .Z(n17598) );
  XNOR U19341 ( .A(n17599), .B(n17598), .Z(n17628) );
  XNOR U19342 ( .A(sreg[1381]), .B(n17628), .Z(n17630) );
  NANDN U19343 ( .A(sreg[1380]), .B(n17591), .Z(n17595) );
  NAND U19344 ( .A(n17593), .B(n17592), .Z(n17594) );
  NAND U19345 ( .A(n17595), .B(n17594), .Z(n17629) );
  XNOR U19346 ( .A(n17630), .B(n17629), .Z(c[1381]) );
  NANDN U19347 ( .A(n17597), .B(n17596), .Z(n17601) );
  NANDN U19348 ( .A(n17599), .B(n17598), .Z(n17600) );
  AND U19349 ( .A(n17601), .B(n17600), .Z(n17636) );
  NANDN U19350 ( .A(n17603), .B(n17602), .Z(n17607) );
  NANDN U19351 ( .A(n17605), .B(n17604), .Z(n17606) );
  AND U19352 ( .A(n17607), .B(n17606), .Z(n17634) );
  NAND U19353 ( .A(n42143), .B(n17608), .Z(n17610) );
  XNOR U19354 ( .A(a[360]), .B(n4123), .Z(n17645) );
  NAND U19355 ( .A(n42144), .B(n17645), .Z(n17609) );
  AND U19356 ( .A(n17610), .B(n17609), .Z(n17660) );
  XOR U19357 ( .A(a[364]), .B(n42012), .Z(n17648) );
  XNOR U19358 ( .A(n17660), .B(n17659), .Z(n17662) );
  AND U19359 ( .A(a[366]), .B(b[0]), .Z(n17612) );
  XNOR U19360 ( .A(n17612), .B(n4071), .Z(n17614) );
  NANDN U19361 ( .A(b[0]), .B(a[365]), .Z(n17613) );
  NAND U19362 ( .A(n17614), .B(n17613), .Z(n17656) );
  XOR U19363 ( .A(a[362]), .B(n42085), .Z(n17649) );
  AND U19364 ( .A(a[358]), .B(b[7]), .Z(n17653) );
  XNOR U19365 ( .A(n17654), .B(n17653), .Z(n17655) );
  XNOR U19366 ( .A(n17656), .B(n17655), .Z(n17661) );
  XOR U19367 ( .A(n17662), .B(n17661), .Z(n17640) );
  NANDN U19368 ( .A(n17617), .B(n17616), .Z(n17621) );
  NANDN U19369 ( .A(n17619), .B(n17618), .Z(n17620) );
  AND U19370 ( .A(n17621), .B(n17620), .Z(n17639) );
  XNOR U19371 ( .A(n17640), .B(n17639), .Z(n17641) );
  NANDN U19372 ( .A(n17623), .B(n17622), .Z(n17627) );
  NAND U19373 ( .A(n17625), .B(n17624), .Z(n17626) );
  NAND U19374 ( .A(n17627), .B(n17626), .Z(n17642) );
  XNOR U19375 ( .A(n17641), .B(n17642), .Z(n17633) );
  XNOR U19376 ( .A(n17634), .B(n17633), .Z(n17635) );
  XNOR U19377 ( .A(n17636), .B(n17635), .Z(n17665) );
  XNOR U19378 ( .A(sreg[1382]), .B(n17665), .Z(n17667) );
  NANDN U19379 ( .A(sreg[1381]), .B(n17628), .Z(n17632) );
  NAND U19380 ( .A(n17630), .B(n17629), .Z(n17631) );
  NAND U19381 ( .A(n17632), .B(n17631), .Z(n17666) );
  XNOR U19382 ( .A(n17667), .B(n17666), .Z(c[1382]) );
  NANDN U19383 ( .A(n17634), .B(n17633), .Z(n17638) );
  NANDN U19384 ( .A(n17636), .B(n17635), .Z(n17637) );
  AND U19385 ( .A(n17638), .B(n17637), .Z(n17673) );
  NANDN U19386 ( .A(n17640), .B(n17639), .Z(n17644) );
  NANDN U19387 ( .A(n17642), .B(n17641), .Z(n17643) );
  AND U19388 ( .A(n17644), .B(n17643), .Z(n17671) );
  NAND U19389 ( .A(n42143), .B(n17645), .Z(n17647) );
  XNOR U19390 ( .A(a[361]), .B(n4123), .Z(n17682) );
  NAND U19391 ( .A(n42144), .B(n17682), .Z(n17646) );
  AND U19392 ( .A(n17647), .B(n17646), .Z(n17697) );
  XOR U19393 ( .A(a[365]), .B(n42012), .Z(n17685) );
  XNOR U19394 ( .A(n17697), .B(n17696), .Z(n17699) );
  XOR U19395 ( .A(a[363]), .B(n42085), .Z(n17689) );
  AND U19396 ( .A(a[359]), .B(b[7]), .Z(n17690) );
  XNOR U19397 ( .A(n17691), .B(n17690), .Z(n17692) );
  AND U19398 ( .A(a[367]), .B(b[0]), .Z(n17650) );
  XNOR U19399 ( .A(n17650), .B(n4071), .Z(n17652) );
  NANDN U19400 ( .A(b[0]), .B(a[366]), .Z(n17651) );
  NAND U19401 ( .A(n17652), .B(n17651), .Z(n17693) );
  XNOR U19402 ( .A(n17692), .B(n17693), .Z(n17698) );
  XOR U19403 ( .A(n17699), .B(n17698), .Z(n17677) );
  NANDN U19404 ( .A(n17654), .B(n17653), .Z(n17658) );
  NANDN U19405 ( .A(n17656), .B(n17655), .Z(n17657) );
  AND U19406 ( .A(n17658), .B(n17657), .Z(n17676) );
  XNOR U19407 ( .A(n17677), .B(n17676), .Z(n17678) );
  NANDN U19408 ( .A(n17660), .B(n17659), .Z(n17664) );
  NAND U19409 ( .A(n17662), .B(n17661), .Z(n17663) );
  NAND U19410 ( .A(n17664), .B(n17663), .Z(n17679) );
  XNOR U19411 ( .A(n17678), .B(n17679), .Z(n17670) );
  XNOR U19412 ( .A(n17671), .B(n17670), .Z(n17672) );
  XNOR U19413 ( .A(n17673), .B(n17672), .Z(n17702) );
  XNOR U19414 ( .A(sreg[1383]), .B(n17702), .Z(n17704) );
  NANDN U19415 ( .A(sreg[1382]), .B(n17665), .Z(n17669) );
  NAND U19416 ( .A(n17667), .B(n17666), .Z(n17668) );
  NAND U19417 ( .A(n17669), .B(n17668), .Z(n17703) );
  XNOR U19418 ( .A(n17704), .B(n17703), .Z(c[1383]) );
  NANDN U19419 ( .A(n17671), .B(n17670), .Z(n17675) );
  NANDN U19420 ( .A(n17673), .B(n17672), .Z(n17674) );
  AND U19421 ( .A(n17675), .B(n17674), .Z(n17710) );
  NANDN U19422 ( .A(n17677), .B(n17676), .Z(n17681) );
  NANDN U19423 ( .A(n17679), .B(n17678), .Z(n17680) );
  AND U19424 ( .A(n17681), .B(n17680), .Z(n17708) );
  NAND U19425 ( .A(n42143), .B(n17682), .Z(n17684) );
  XNOR U19426 ( .A(a[362]), .B(n4123), .Z(n17719) );
  NAND U19427 ( .A(n42144), .B(n17719), .Z(n17683) );
  AND U19428 ( .A(n17684), .B(n17683), .Z(n17734) );
  XOR U19429 ( .A(a[366]), .B(n42012), .Z(n17722) );
  XNOR U19430 ( .A(n17734), .B(n17733), .Z(n17736) );
  AND U19431 ( .A(a[368]), .B(b[0]), .Z(n17686) );
  XNOR U19432 ( .A(n17686), .B(n4071), .Z(n17688) );
  NANDN U19433 ( .A(b[0]), .B(a[367]), .Z(n17687) );
  NAND U19434 ( .A(n17688), .B(n17687), .Z(n17730) );
  XOR U19435 ( .A(a[364]), .B(n42085), .Z(n17726) );
  AND U19436 ( .A(a[360]), .B(b[7]), .Z(n17727) );
  XNOR U19437 ( .A(n17728), .B(n17727), .Z(n17729) );
  XNOR U19438 ( .A(n17730), .B(n17729), .Z(n17735) );
  XOR U19439 ( .A(n17736), .B(n17735), .Z(n17714) );
  NANDN U19440 ( .A(n17691), .B(n17690), .Z(n17695) );
  NANDN U19441 ( .A(n17693), .B(n17692), .Z(n17694) );
  AND U19442 ( .A(n17695), .B(n17694), .Z(n17713) );
  XNOR U19443 ( .A(n17714), .B(n17713), .Z(n17715) );
  NANDN U19444 ( .A(n17697), .B(n17696), .Z(n17701) );
  NAND U19445 ( .A(n17699), .B(n17698), .Z(n17700) );
  NAND U19446 ( .A(n17701), .B(n17700), .Z(n17716) );
  XNOR U19447 ( .A(n17715), .B(n17716), .Z(n17707) );
  XNOR U19448 ( .A(n17708), .B(n17707), .Z(n17709) );
  XNOR U19449 ( .A(n17710), .B(n17709), .Z(n17739) );
  XNOR U19450 ( .A(sreg[1384]), .B(n17739), .Z(n17741) );
  NANDN U19451 ( .A(sreg[1383]), .B(n17702), .Z(n17706) );
  NAND U19452 ( .A(n17704), .B(n17703), .Z(n17705) );
  NAND U19453 ( .A(n17706), .B(n17705), .Z(n17740) );
  XNOR U19454 ( .A(n17741), .B(n17740), .Z(c[1384]) );
  NANDN U19455 ( .A(n17708), .B(n17707), .Z(n17712) );
  NANDN U19456 ( .A(n17710), .B(n17709), .Z(n17711) );
  AND U19457 ( .A(n17712), .B(n17711), .Z(n17747) );
  NANDN U19458 ( .A(n17714), .B(n17713), .Z(n17718) );
  NANDN U19459 ( .A(n17716), .B(n17715), .Z(n17717) );
  AND U19460 ( .A(n17718), .B(n17717), .Z(n17745) );
  NAND U19461 ( .A(n42143), .B(n17719), .Z(n17721) );
  XNOR U19462 ( .A(a[363]), .B(n4123), .Z(n17756) );
  NAND U19463 ( .A(n42144), .B(n17756), .Z(n17720) );
  AND U19464 ( .A(n17721), .B(n17720), .Z(n17771) );
  XOR U19465 ( .A(a[367]), .B(n42012), .Z(n17759) );
  XNOR U19466 ( .A(n17771), .B(n17770), .Z(n17773) );
  AND U19467 ( .A(a[369]), .B(b[0]), .Z(n17723) );
  XNOR U19468 ( .A(n17723), .B(n4071), .Z(n17725) );
  NANDN U19469 ( .A(b[0]), .B(a[368]), .Z(n17724) );
  NAND U19470 ( .A(n17725), .B(n17724), .Z(n17767) );
  XOR U19471 ( .A(a[365]), .B(n42085), .Z(n17763) );
  AND U19472 ( .A(a[361]), .B(b[7]), .Z(n17764) );
  XNOR U19473 ( .A(n17765), .B(n17764), .Z(n17766) );
  XNOR U19474 ( .A(n17767), .B(n17766), .Z(n17772) );
  XOR U19475 ( .A(n17773), .B(n17772), .Z(n17751) );
  NANDN U19476 ( .A(n17728), .B(n17727), .Z(n17732) );
  NANDN U19477 ( .A(n17730), .B(n17729), .Z(n17731) );
  AND U19478 ( .A(n17732), .B(n17731), .Z(n17750) );
  XNOR U19479 ( .A(n17751), .B(n17750), .Z(n17752) );
  NANDN U19480 ( .A(n17734), .B(n17733), .Z(n17738) );
  NAND U19481 ( .A(n17736), .B(n17735), .Z(n17737) );
  NAND U19482 ( .A(n17738), .B(n17737), .Z(n17753) );
  XNOR U19483 ( .A(n17752), .B(n17753), .Z(n17744) );
  XNOR U19484 ( .A(n17745), .B(n17744), .Z(n17746) );
  XNOR U19485 ( .A(n17747), .B(n17746), .Z(n17776) );
  XNOR U19486 ( .A(sreg[1385]), .B(n17776), .Z(n17778) );
  NANDN U19487 ( .A(sreg[1384]), .B(n17739), .Z(n17743) );
  NAND U19488 ( .A(n17741), .B(n17740), .Z(n17742) );
  NAND U19489 ( .A(n17743), .B(n17742), .Z(n17777) );
  XNOR U19490 ( .A(n17778), .B(n17777), .Z(c[1385]) );
  NANDN U19491 ( .A(n17745), .B(n17744), .Z(n17749) );
  NANDN U19492 ( .A(n17747), .B(n17746), .Z(n17748) );
  AND U19493 ( .A(n17749), .B(n17748), .Z(n17784) );
  NANDN U19494 ( .A(n17751), .B(n17750), .Z(n17755) );
  NANDN U19495 ( .A(n17753), .B(n17752), .Z(n17754) );
  AND U19496 ( .A(n17755), .B(n17754), .Z(n17782) );
  NAND U19497 ( .A(n42143), .B(n17756), .Z(n17758) );
  XNOR U19498 ( .A(a[364]), .B(n4123), .Z(n17793) );
  NAND U19499 ( .A(n42144), .B(n17793), .Z(n17757) );
  AND U19500 ( .A(n17758), .B(n17757), .Z(n17808) );
  XOR U19501 ( .A(a[368]), .B(n42012), .Z(n17796) );
  XNOR U19502 ( .A(n17808), .B(n17807), .Z(n17810) );
  AND U19503 ( .A(a[370]), .B(b[0]), .Z(n17760) );
  XNOR U19504 ( .A(n17760), .B(n4071), .Z(n17762) );
  NANDN U19505 ( .A(b[0]), .B(a[369]), .Z(n17761) );
  NAND U19506 ( .A(n17762), .B(n17761), .Z(n17804) );
  XOR U19507 ( .A(a[366]), .B(n42085), .Z(n17797) );
  AND U19508 ( .A(a[362]), .B(b[7]), .Z(n17801) );
  XNOR U19509 ( .A(n17802), .B(n17801), .Z(n17803) );
  XNOR U19510 ( .A(n17804), .B(n17803), .Z(n17809) );
  XOR U19511 ( .A(n17810), .B(n17809), .Z(n17788) );
  NANDN U19512 ( .A(n17765), .B(n17764), .Z(n17769) );
  NANDN U19513 ( .A(n17767), .B(n17766), .Z(n17768) );
  AND U19514 ( .A(n17769), .B(n17768), .Z(n17787) );
  XNOR U19515 ( .A(n17788), .B(n17787), .Z(n17789) );
  NANDN U19516 ( .A(n17771), .B(n17770), .Z(n17775) );
  NAND U19517 ( .A(n17773), .B(n17772), .Z(n17774) );
  NAND U19518 ( .A(n17775), .B(n17774), .Z(n17790) );
  XNOR U19519 ( .A(n17789), .B(n17790), .Z(n17781) );
  XNOR U19520 ( .A(n17782), .B(n17781), .Z(n17783) );
  XNOR U19521 ( .A(n17784), .B(n17783), .Z(n17813) );
  XNOR U19522 ( .A(sreg[1386]), .B(n17813), .Z(n17815) );
  NANDN U19523 ( .A(sreg[1385]), .B(n17776), .Z(n17780) );
  NAND U19524 ( .A(n17778), .B(n17777), .Z(n17779) );
  NAND U19525 ( .A(n17780), .B(n17779), .Z(n17814) );
  XNOR U19526 ( .A(n17815), .B(n17814), .Z(c[1386]) );
  NANDN U19527 ( .A(n17782), .B(n17781), .Z(n17786) );
  NANDN U19528 ( .A(n17784), .B(n17783), .Z(n17785) );
  AND U19529 ( .A(n17786), .B(n17785), .Z(n17821) );
  NANDN U19530 ( .A(n17788), .B(n17787), .Z(n17792) );
  NANDN U19531 ( .A(n17790), .B(n17789), .Z(n17791) );
  AND U19532 ( .A(n17792), .B(n17791), .Z(n17819) );
  NAND U19533 ( .A(n42143), .B(n17793), .Z(n17795) );
  XNOR U19534 ( .A(a[365]), .B(n4124), .Z(n17830) );
  NAND U19535 ( .A(n42144), .B(n17830), .Z(n17794) );
  AND U19536 ( .A(n17795), .B(n17794), .Z(n17845) );
  XOR U19537 ( .A(a[369]), .B(n42012), .Z(n17833) );
  XNOR U19538 ( .A(n17845), .B(n17844), .Z(n17847) );
  XOR U19539 ( .A(a[367]), .B(n42085), .Z(n17837) );
  AND U19540 ( .A(a[363]), .B(b[7]), .Z(n17838) );
  XNOR U19541 ( .A(n17839), .B(n17838), .Z(n17840) );
  AND U19542 ( .A(a[371]), .B(b[0]), .Z(n17798) );
  XNOR U19543 ( .A(n17798), .B(n4071), .Z(n17800) );
  NANDN U19544 ( .A(b[0]), .B(a[370]), .Z(n17799) );
  NAND U19545 ( .A(n17800), .B(n17799), .Z(n17841) );
  XNOR U19546 ( .A(n17840), .B(n17841), .Z(n17846) );
  XOR U19547 ( .A(n17847), .B(n17846), .Z(n17825) );
  NANDN U19548 ( .A(n17802), .B(n17801), .Z(n17806) );
  NANDN U19549 ( .A(n17804), .B(n17803), .Z(n17805) );
  AND U19550 ( .A(n17806), .B(n17805), .Z(n17824) );
  XNOR U19551 ( .A(n17825), .B(n17824), .Z(n17826) );
  NANDN U19552 ( .A(n17808), .B(n17807), .Z(n17812) );
  NAND U19553 ( .A(n17810), .B(n17809), .Z(n17811) );
  NAND U19554 ( .A(n17812), .B(n17811), .Z(n17827) );
  XNOR U19555 ( .A(n17826), .B(n17827), .Z(n17818) );
  XNOR U19556 ( .A(n17819), .B(n17818), .Z(n17820) );
  XNOR U19557 ( .A(n17821), .B(n17820), .Z(n17850) );
  XNOR U19558 ( .A(sreg[1387]), .B(n17850), .Z(n17852) );
  NANDN U19559 ( .A(sreg[1386]), .B(n17813), .Z(n17817) );
  NAND U19560 ( .A(n17815), .B(n17814), .Z(n17816) );
  NAND U19561 ( .A(n17817), .B(n17816), .Z(n17851) );
  XNOR U19562 ( .A(n17852), .B(n17851), .Z(c[1387]) );
  NANDN U19563 ( .A(n17819), .B(n17818), .Z(n17823) );
  NANDN U19564 ( .A(n17821), .B(n17820), .Z(n17822) );
  AND U19565 ( .A(n17823), .B(n17822), .Z(n17858) );
  NANDN U19566 ( .A(n17825), .B(n17824), .Z(n17829) );
  NANDN U19567 ( .A(n17827), .B(n17826), .Z(n17828) );
  AND U19568 ( .A(n17829), .B(n17828), .Z(n17856) );
  NAND U19569 ( .A(n42143), .B(n17830), .Z(n17832) );
  XNOR U19570 ( .A(a[366]), .B(n4124), .Z(n17867) );
  NAND U19571 ( .A(n42144), .B(n17867), .Z(n17831) );
  AND U19572 ( .A(n17832), .B(n17831), .Z(n17882) );
  XOR U19573 ( .A(a[370]), .B(n42012), .Z(n17870) );
  XNOR U19574 ( .A(n17882), .B(n17881), .Z(n17884) );
  AND U19575 ( .A(a[372]), .B(b[0]), .Z(n17834) );
  XNOR U19576 ( .A(n17834), .B(n4071), .Z(n17836) );
  NANDN U19577 ( .A(b[0]), .B(a[371]), .Z(n17835) );
  NAND U19578 ( .A(n17836), .B(n17835), .Z(n17878) );
  XOR U19579 ( .A(a[368]), .B(n42085), .Z(n17874) );
  AND U19580 ( .A(a[364]), .B(b[7]), .Z(n17875) );
  XNOR U19581 ( .A(n17876), .B(n17875), .Z(n17877) );
  XNOR U19582 ( .A(n17878), .B(n17877), .Z(n17883) );
  XOR U19583 ( .A(n17884), .B(n17883), .Z(n17862) );
  NANDN U19584 ( .A(n17839), .B(n17838), .Z(n17843) );
  NANDN U19585 ( .A(n17841), .B(n17840), .Z(n17842) );
  AND U19586 ( .A(n17843), .B(n17842), .Z(n17861) );
  XNOR U19587 ( .A(n17862), .B(n17861), .Z(n17863) );
  NANDN U19588 ( .A(n17845), .B(n17844), .Z(n17849) );
  NAND U19589 ( .A(n17847), .B(n17846), .Z(n17848) );
  NAND U19590 ( .A(n17849), .B(n17848), .Z(n17864) );
  XNOR U19591 ( .A(n17863), .B(n17864), .Z(n17855) );
  XNOR U19592 ( .A(n17856), .B(n17855), .Z(n17857) );
  XNOR U19593 ( .A(n17858), .B(n17857), .Z(n17887) );
  XNOR U19594 ( .A(sreg[1388]), .B(n17887), .Z(n17889) );
  NANDN U19595 ( .A(sreg[1387]), .B(n17850), .Z(n17854) );
  NAND U19596 ( .A(n17852), .B(n17851), .Z(n17853) );
  NAND U19597 ( .A(n17854), .B(n17853), .Z(n17888) );
  XNOR U19598 ( .A(n17889), .B(n17888), .Z(c[1388]) );
  NANDN U19599 ( .A(n17856), .B(n17855), .Z(n17860) );
  NANDN U19600 ( .A(n17858), .B(n17857), .Z(n17859) );
  AND U19601 ( .A(n17860), .B(n17859), .Z(n17895) );
  NANDN U19602 ( .A(n17862), .B(n17861), .Z(n17866) );
  NANDN U19603 ( .A(n17864), .B(n17863), .Z(n17865) );
  AND U19604 ( .A(n17866), .B(n17865), .Z(n17893) );
  NAND U19605 ( .A(n42143), .B(n17867), .Z(n17869) );
  XNOR U19606 ( .A(a[367]), .B(n4124), .Z(n17904) );
  NAND U19607 ( .A(n42144), .B(n17904), .Z(n17868) );
  AND U19608 ( .A(n17869), .B(n17868), .Z(n17919) );
  XOR U19609 ( .A(a[371]), .B(n42012), .Z(n17907) );
  XNOR U19610 ( .A(n17919), .B(n17918), .Z(n17921) );
  AND U19611 ( .A(a[373]), .B(b[0]), .Z(n17871) );
  XNOR U19612 ( .A(n17871), .B(n4071), .Z(n17873) );
  NANDN U19613 ( .A(b[0]), .B(a[372]), .Z(n17872) );
  NAND U19614 ( .A(n17873), .B(n17872), .Z(n17915) );
  XOR U19615 ( .A(a[369]), .B(n42085), .Z(n17911) );
  AND U19616 ( .A(a[365]), .B(b[7]), .Z(n17912) );
  XNOR U19617 ( .A(n17913), .B(n17912), .Z(n17914) );
  XNOR U19618 ( .A(n17915), .B(n17914), .Z(n17920) );
  XOR U19619 ( .A(n17921), .B(n17920), .Z(n17899) );
  NANDN U19620 ( .A(n17876), .B(n17875), .Z(n17880) );
  NANDN U19621 ( .A(n17878), .B(n17877), .Z(n17879) );
  AND U19622 ( .A(n17880), .B(n17879), .Z(n17898) );
  XNOR U19623 ( .A(n17899), .B(n17898), .Z(n17900) );
  NANDN U19624 ( .A(n17882), .B(n17881), .Z(n17886) );
  NAND U19625 ( .A(n17884), .B(n17883), .Z(n17885) );
  NAND U19626 ( .A(n17886), .B(n17885), .Z(n17901) );
  XNOR U19627 ( .A(n17900), .B(n17901), .Z(n17892) );
  XNOR U19628 ( .A(n17893), .B(n17892), .Z(n17894) );
  XNOR U19629 ( .A(n17895), .B(n17894), .Z(n17924) );
  XNOR U19630 ( .A(sreg[1389]), .B(n17924), .Z(n17926) );
  NANDN U19631 ( .A(sreg[1388]), .B(n17887), .Z(n17891) );
  NAND U19632 ( .A(n17889), .B(n17888), .Z(n17890) );
  NAND U19633 ( .A(n17891), .B(n17890), .Z(n17925) );
  XNOR U19634 ( .A(n17926), .B(n17925), .Z(c[1389]) );
  NANDN U19635 ( .A(n17893), .B(n17892), .Z(n17897) );
  NANDN U19636 ( .A(n17895), .B(n17894), .Z(n17896) );
  AND U19637 ( .A(n17897), .B(n17896), .Z(n17932) );
  NANDN U19638 ( .A(n17899), .B(n17898), .Z(n17903) );
  NANDN U19639 ( .A(n17901), .B(n17900), .Z(n17902) );
  AND U19640 ( .A(n17903), .B(n17902), .Z(n17930) );
  NAND U19641 ( .A(n42143), .B(n17904), .Z(n17906) );
  XNOR U19642 ( .A(a[368]), .B(n4124), .Z(n17941) );
  NAND U19643 ( .A(n42144), .B(n17941), .Z(n17905) );
  AND U19644 ( .A(n17906), .B(n17905), .Z(n17956) );
  XOR U19645 ( .A(a[372]), .B(n42012), .Z(n17944) );
  XNOR U19646 ( .A(n17956), .B(n17955), .Z(n17958) );
  AND U19647 ( .A(a[374]), .B(b[0]), .Z(n17908) );
  XNOR U19648 ( .A(n17908), .B(n4071), .Z(n17910) );
  NANDN U19649 ( .A(b[0]), .B(a[373]), .Z(n17909) );
  NAND U19650 ( .A(n17910), .B(n17909), .Z(n17952) );
  XOR U19651 ( .A(a[370]), .B(n42085), .Z(n17948) );
  AND U19652 ( .A(a[366]), .B(b[7]), .Z(n17949) );
  XNOR U19653 ( .A(n17950), .B(n17949), .Z(n17951) );
  XNOR U19654 ( .A(n17952), .B(n17951), .Z(n17957) );
  XOR U19655 ( .A(n17958), .B(n17957), .Z(n17936) );
  NANDN U19656 ( .A(n17913), .B(n17912), .Z(n17917) );
  NANDN U19657 ( .A(n17915), .B(n17914), .Z(n17916) );
  AND U19658 ( .A(n17917), .B(n17916), .Z(n17935) );
  XNOR U19659 ( .A(n17936), .B(n17935), .Z(n17937) );
  NANDN U19660 ( .A(n17919), .B(n17918), .Z(n17923) );
  NAND U19661 ( .A(n17921), .B(n17920), .Z(n17922) );
  NAND U19662 ( .A(n17923), .B(n17922), .Z(n17938) );
  XNOR U19663 ( .A(n17937), .B(n17938), .Z(n17929) );
  XNOR U19664 ( .A(n17930), .B(n17929), .Z(n17931) );
  XNOR U19665 ( .A(n17932), .B(n17931), .Z(n17961) );
  XNOR U19666 ( .A(sreg[1390]), .B(n17961), .Z(n17963) );
  NANDN U19667 ( .A(sreg[1389]), .B(n17924), .Z(n17928) );
  NAND U19668 ( .A(n17926), .B(n17925), .Z(n17927) );
  NAND U19669 ( .A(n17928), .B(n17927), .Z(n17962) );
  XNOR U19670 ( .A(n17963), .B(n17962), .Z(c[1390]) );
  NANDN U19671 ( .A(n17930), .B(n17929), .Z(n17934) );
  NANDN U19672 ( .A(n17932), .B(n17931), .Z(n17933) );
  AND U19673 ( .A(n17934), .B(n17933), .Z(n17969) );
  NANDN U19674 ( .A(n17936), .B(n17935), .Z(n17940) );
  NANDN U19675 ( .A(n17938), .B(n17937), .Z(n17939) );
  AND U19676 ( .A(n17940), .B(n17939), .Z(n17967) );
  NAND U19677 ( .A(n42143), .B(n17941), .Z(n17943) );
  XNOR U19678 ( .A(a[369]), .B(n4124), .Z(n17978) );
  NAND U19679 ( .A(n42144), .B(n17978), .Z(n17942) );
  AND U19680 ( .A(n17943), .B(n17942), .Z(n17993) );
  XOR U19681 ( .A(a[373]), .B(n42012), .Z(n17981) );
  XNOR U19682 ( .A(n17993), .B(n17992), .Z(n17995) );
  AND U19683 ( .A(a[375]), .B(b[0]), .Z(n17945) );
  XNOR U19684 ( .A(n17945), .B(n4071), .Z(n17947) );
  NANDN U19685 ( .A(b[0]), .B(a[374]), .Z(n17946) );
  NAND U19686 ( .A(n17947), .B(n17946), .Z(n17989) );
  XOR U19687 ( .A(a[371]), .B(n42085), .Z(n17985) );
  AND U19688 ( .A(a[367]), .B(b[7]), .Z(n17986) );
  XNOR U19689 ( .A(n17987), .B(n17986), .Z(n17988) );
  XNOR U19690 ( .A(n17989), .B(n17988), .Z(n17994) );
  XOR U19691 ( .A(n17995), .B(n17994), .Z(n17973) );
  NANDN U19692 ( .A(n17950), .B(n17949), .Z(n17954) );
  NANDN U19693 ( .A(n17952), .B(n17951), .Z(n17953) );
  AND U19694 ( .A(n17954), .B(n17953), .Z(n17972) );
  XNOR U19695 ( .A(n17973), .B(n17972), .Z(n17974) );
  NANDN U19696 ( .A(n17956), .B(n17955), .Z(n17960) );
  NAND U19697 ( .A(n17958), .B(n17957), .Z(n17959) );
  NAND U19698 ( .A(n17960), .B(n17959), .Z(n17975) );
  XNOR U19699 ( .A(n17974), .B(n17975), .Z(n17966) );
  XNOR U19700 ( .A(n17967), .B(n17966), .Z(n17968) );
  XNOR U19701 ( .A(n17969), .B(n17968), .Z(n17998) );
  XNOR U19702 ( .A(sreg[1391]), .B(n17998), .Z(n18000) );
  NANDN U19703 ( .A(sreg[1390]), .B(n17961), .Z(n17965) );
  NAND U19704 ( .A(n17963), .B(n17962), .Z(n17964) );
  NAND U19705 ( .A(n17965), .B(n17964), .Z(n17999) );
  XNOR U19706 ( .A(n18000), .B(n17999), .Z(c[1391]) );
  NANDN U19707 ( .A(n17967), .B(n17966), .Z(n17971) );
  NANDN U19708 ( .A(n17969), .B(n17968), .Z(n17970) );
  AND U19709 ( .A(n17971), .B(n17970), .Z(n18006) );
  NANDN U19710 ( .A(n17973), .B(n17972), .Z(n17977) );
  NANDN U19711 ( .A(n17975), .B(n17974), .Z(n17976) );
  AND U19712 ( .A(n17977), .B(n17976), .Z(n18004) );
  NAND U19713 ( .A(n42143), .B(n17978), .Z(n17980) );
  XNOR U19714 ( .A(a[370]), .B(n4124), .Z(n18015) );
  NAND U19715 ( .A(n42144), .B(n18015), .Z(n17979) );
  AND U19716 ( .A(n17980), .B(n17979), .Z(n18030) );
  XOR U19717 ( .A(a[374]), .B(n42012), .Z(n18018) );
  XNOR U19718 ( .A(n18030), .B(n18029), .Z(n18032) );
  AND U19719 ( .A(a[376]), .B(b[0]), .Z(n17982) );
  XNOR U19720 ( .A(n17982), .B(n4071), .Z(n17984) );
  NANDN U19721 ( .A(b[0]), .B(a[375]), .Z(n17983) );
  NAND U19722 ( .A(n17984), .B(n17983), .Z(n18026) );
  XOR U19723 ( .A(a[372]), .B(n42085), .Z(n18022) );
  AND U19724 ( .A(a[368]), .B(b[7]), .Z(n18023) );
  XNOR U19725 ( .A(n18024), .B(n18023), .Z(n18025) );
  XNOR U19726 ( .A(n18026), .B(n18025), .Z(n18031) );
  XOR U19727 ( .A(n18032), .B(n18031), .Z(n18010) );
  NANDN U19728 ( .A(n17987), .B(n17986), .Z(n17991) );
  NANDN U19729 ( .A(n17989), .B(n17988), .Z(n17990) );
  AND U19730 ( .A(n17991), .B(n17990), .Z(n18009) );
  XNOR U19731 ( .A(n18010), .B(n18009), .Z(n18011) );
  NANDN U19732 ( .A(n17993), .B(n17992), .Z(n17997) );
  NAND U19733 ( .A(n17995), .B(n17994), .Z(n17996) );
  NAND U19734 ( .A(n17997), .B(n17996), .Z(n18012) );
  XNOR U19735 ( .A(n18011), .B(n18012), .Z(n18003) );
  XNOR U19736 ( .A(n18004), .B(n18003), .Z(n18005) );
  XNOR U19737 ( .A(n18006), .B(n18005), .Z(n18035) );
  XNOR U19738 ( .A(sreg[1392]), .B(n18035), .Z(n18037) );
  NANDN U19739 ( .A(sreg[1391]), .B(n17998), .Z(n18002) );
  NAND U19740 ( .A(n18000), .B(n17999), .Z(n18001) );
  NAND U19741 ( .A(n18002), .B(n18001), .Z(n18036) );
  XNOR U19742 ( .A(n18037), .B(n18036), .Z(c[1392]) );
  NANDN U19743 ( .A(n18004), .B(n18003), .Z(n18008) );
  NANDN U19744 ( .A(n18006), .B(n18005), .Z(n18007) );
  AND U19745 ( .A(n18008), .B(n18007), .Z(n18043) );
  NANDN U19746 ( .A(n18010), .B(n18009), .Z(n18014) );
  NANDN U19747 ( .A(n18012), .B(n18011), .Z(n18013) );
  AND U19748 ( .A(n18014), .B(n18013), .Z(n18041) );
  NAND U19749 ( .A(n42143), .B(n18015), .Z(n18017) );
  XNOR U19750 ( .A(a[371]), .B(n4124), .Z(n18052) );
  NAND U19751 ( .A(n42144), .B(n18052), .Z(n18016) );
  AND U19752 ( .A(n18017), .B(n18016), .Z(n18067) );
  XOR U19753 ( .A(a[375]), .B(n42012), .Z(n18055) );
  XNOR U19754 ( .A(n18067), .B(n18066), .Z(n18069) );
  AND U19755 ( .A(a[377]), .B(b[0]), .Z(n18019) );
  XNOR U19756 ( .A(n18019), .B(n4071), .Z(n18021) );
  NANDN U19757 ( .A(b[0]), .B(a[376]), .Z(n18020) );
  NAND U19758 ( .A(n18021), .B(n18020), .Z(n18063) );
  XOR U19759 ( .A(a[373]), .B(n42085), .Z(n18059) );
  AND U19760 ( .A(a[369]), .B(b[7]), .Z(n18060) );
  XNOR U19761 ( .A(n18061), .B(n18060), .Z(n18062) );
  XNOR U19762 ( .A(n18063), .B(n18062), .Z(n18068) );
  XOR U19763 ( .A(n18069), .B(n18068), .Z(n18047) );
  NANDN U19764 ( .A(n18024), .B(n18023), .Z(n18028) );
  NANDN U19765 ( .A(n18026), .B(n18025), .Z(n18027) );
  AND U19766 ( .A(n18028), .B(n18027), .Z(n18046) );
  XNOR U19767 ( .A(n18047), .B(n18046), .Z(n18048) );
  NANDN U19768 ( .A(n18030), .B(n18029), .Z(n18034) );
  NAND U19769 ( .A(n18032), .B(n18031), .Z(n18033) );
  NAND U19770 ( .A(n18034), .B(n18033), .Z(n18049) );
  XNOR U19771 ( .A(n18048), .B(n18049), .Z(n18040) );
  XNOR U19772 ( .A(n18041), .B(n18040), .Z(n18042) );
  XNOR U19773 ( .A(n18043), .B(n18042), .Z(n18072) );
  XNOR U19774 ( .A(sreg[1393]), .B(n18072), .Z(n18074) );
  NANDN U19775 ( .A(sreg[1392]), .B(n18035), .Z(n18039) );
  NAND U19776 ( .A(n18037), .B(n18036), .Z(n18038) );
  NAND U19777 ( .A(n18039), .B(n18038), .Z(n18073) );
  XNOR U19778 ( .A(n18074), .B(n18073), .Z(c[1393]) );
  NANDN U19779 ( .A(n18041), .B(n18040), .Z(n18045) );
  NANDN U19780 ( .A(n18043), .B(n18042), .Z(n18044) );
  AND U19781 ( .A(n18045), .B(n18044), .Z(n18080) );
  NANDN U19782 ( .A(n18047), .B(n18046), .Z(n18051) );
  NANDN U19783 ( .A(n18049), .B(n18048), .Z(n18050) );
  AND U19784 ( .A(n18051), .B(n18050), .Z(n18078) );
  NAND U19785 ( .A(n42143), .B(n18052), .Z(n18054) );
  XNOR U19786 ( .A(a[372]), .B(n4125), .Z(n18089) );
  NAND U19787 ( .A(n42144), .B(n18089), .Z(n18053) );
  AND U19788 ( .A(n18054), .B(n18053), .Z(n18104) );
  XOR U19789 ( .A(a[376]), .B(n42012), .Z(n18092) );
  XNOR U19790 ( .A(n18104), .B(n18103), .Z(n18106) );
  AND U19791 ( .A(a[378]), .B(b[0]), .Z(n18056) );
  XNOR U19792 ( .A(n18056), .B(n4071), .Z(n18058) );
  NANDN U19793 ( .A(b[0]), .B(a[377]), .Z(n18057) );
  NAND U19794 ( .A(n18058), .B(n18057), .Z(n18100) );
  XOR U19795 ( .A(a[374]), .B(n42085), .Z(n18096) );
  AND U19796 ( .A(a[370]), .B(b[7]), .Z(n18097) );
  XNOR U19797 ( .A(n18098), .B(n18097), .Z(n18099) );
  XNOR U19798 ( .A(n18100), .B(n18099), .Z(n18105) );
  XOR U19799 ( .A(n18106), .B(n18105), .Z(n18084) );
  NANDN U19800 ( .A(n18061), .B(n18060), .Z(n18065) );
  NANDN U19801 ( .A(n18063), .B(n18062), .Z(n18064) );
  AND U19802 ( .A(n18065), .B(n18064), .Z(n18083) );
  XNOR U19803 ( .A(n18084), .B(n18083), .Z(n18085) );
  NANDN U19804 ( .A(n18067), .B(n18066), .Z(n18071) );
  NAND U19805 ( .A(n18069), .B(n18068), .Z(n18070) );
  NAND U19806 ( .A(n18071), .B(n18070), .Z(n18086) );
  XNOR U19807 ( .A(n18085), .B(n18086), .Z(n18077) );
  XNOR U19808 ( .A(n18078), .B(n18077), .Z(n18079) );
  XNOR U19809 ( .A(n18080), .B(n18079), .Z(n18109) );
  XNOR U19810 ( .A(sreg[1394]), .B(n18109), .Z(n18111) );
  NANDN U19811 ( .A(sreg[1393]), .B(n18072), .Z(n18076) );
  NAND U19812 ( .A(n18074), .B(n18073), .Z(n18075) );
  NAND U19813 ( .A(n18076), .B(n18075), .Z(n18110) );
  XNOR U19814 ( .A(n18111), .B(n18110), .Z(c[1394]) );
  NANDN U19815 ( .A(n18078), .B(n18077), .Z(n18082) );
  NANDN U19816 ( .A(n18080), .B(n18079), .Z(n18081) );
  AND U19817 ( .A(n18082), .B(n18081), .Z(n18117) );
  NANDN U19818 ( .A(n18084), .B(n18083), .Z(n18088) );
  NANDN U19819 ( .A(n18086), .B(n18085), .Z(n18087) );
  AND U19820 ( .A(n18088), .B(n18087), .Z(n18115) );
  NAND U19821 ( .A(n42143), .B(n18089), .Z(n18091) );
  XNOR U19822 ( .A(a[373]), .B(n4125), .Z(n18126) );
  NAND U19823 ( .A(n42144), .B(n18126), .Z(n18090) );
  AND U19824 ( .A(n18091), .B(n18090), .Z(n18141) );
  XOR U19825 ( .A(a[377]), .B(n42012), .Z(n18129) );
  XNOR U19826 ( .A(n18141), .B(n18140), .Z(n18143) );
  AND U19827 ( .A(a[379]), .B(b[0]), .Z(n18093) );
  XNOR U19828 ( .A(n18093), .B(n4071), .Z(n18095) );
  NANDN U19829 ( .A(b[0]), .B(a[378]), .Z(n18094) );
  NAND U19830 ( .A(n18095), .B(n18094), .Z(n18137) );
  XOR U19831 ( .A(a[375]), .B(n42085), .Z(n18133) );
  AND U19832 ( .A(a[371]), .B(b[7]), .Z(n18134) );
  XNOR U19833 ( .A(n18135), .B(n18134), .Z(n18136) );
  XNOR U19834 ( .A(n18137), .B(n18136), .Z(n18142) );
  XOR U19835 ( .A(n18143), .B(n18142), .Z(n18121) );
  NANDN U19836 ( .A(n18098), .B(n18097), .Z(n18102) );
  NANDN U19837 ( .A(n18100), .B(n18099), .Z(n18101) );
  AND U19838 ( .A(n18102), .B(n18101), .Z(n18120) );
  XNOR U19839 ( .A(n18121), .B(n18120), .Z(n18122) );
  NANDN U19840 ( .A(n18104), .B(n18103), .Z(n18108) );
  NAND U19841 ( .A(n18106), .B(n18105), .Z(n18107) );
  NAND U19842 ( .A(n18108), .B(n18107), .Z(n18123) );
  XNOR U19843 ( .A(n18122), .B(n18123), .Z(n18114) );
  XNOR U19844 ( .A(n18115), .B(n18114), .Z(n18116) );
  XNOR U19845 ( .A(n18117), .B(n18116), .Z(n18146) );
  XNOR U19846 ( .A(sreg[1395]), .B(n18146), .Z(n18148) );
  NANDN U19847 ( .A(sreg[1394]), .B(n18109), .Z(n18113) );
  NAND U19848 ( .A(n18111), .B(n18110), .Z(n18112) );
  NAND U19849 ( .A(n18113), .B(n18112), .Z(n18147) );
  XNOR U19850 ( .A(n18148), .B(n18147), .Z(c[1395]) );
  NANDN U19851 ( .A(n18115), .B(n18114), .Z(n18119) );
  NANDN U19852 ( .A(n18117), .B(n18116), .Z(n18118) );
  AND U19853 ( .A(n18119), .B(n18118), .Z(n18154) );
  NANDN U19854 ( .A(n18121), .B(n18120), .Z(n18125) );
  NANDN U19855 ( .A(n18123), .B(n18122), .Z(n18124) );
  AND U19856 ( .A(n18125), .B(n18124), .Z(n18152) );
  NAND U19857 ( .A(n42143), .B(n18126), .Z(n18128) );
  XNOR U19858 ( .A(a[374]), .B(n4125), .Z(n18163) );
  NAND U19859 ( .A(n42144), .B(n18163), .Z(n18127) );
  AND U19860 ( .A(n18128), .B(n18127), .Z(n18178) );
  XOR U19861 ( .A(a[378]), .B(n42012), .Z(n18166) );
  XNOR U19862 ( .A(n18178), .B(n18177), .Z(n18180) );
  AND U19863 ( .A(a[380]), .B(b[0]), .Z(n18130) );
  XNOR U19864 ( .A(n18130), .B(n4071), .Z(n18132) );
  NANDN U19865 ( .A(b[0]), .B(a[379]), .Z(n18131) );
  NAND U19866 ( .A(n18132), .B(n18131), .Z(n18174) );
  XOR U19867 ( .A(a[376]), .B(n42085), .Z(n18167) );
  AND U19868 ( .A(a[372]), .B(b[7]), .Z(n18171) );
  XNOR U19869 ( .A(n18172), .B(n18171), .Z(n18173) );
  XNOR U19870 ( .A(n18174), .B(n18173), .Z(n18179) );
  XOR U19871 ( .A(n18180), .B(n18179), .Z(n18158) );
  NANDN U19872 ( .A(n18135), .B(n18134), .Z(n18139) );
  NANDN U19873 ( .A(n18137), .B(n18136), .Z(n18138) );
  AND U19874 ( .A(n18139), .B(n18138), .Z(n18157) );
  XNOR U19875 ( .A(n18158), .B(n18157), .Z(n18159) );
  NANDN U19876 ( .A(n18141), .B(n18140), .Z(n18145) );
  NAND U19877 ( .A(n18143), .B(n18142), .Z(n18144) );
  NAND U19878 ( .A(n18145), .B(n18144), .Z(n18160) );
  XNOR U19879 ( .A(n18159), .B(n18160), .Z(n18151) );
  XNOR U19880 ( .A(n18152), .B(n18151), .Z(n18153) );
  XNOR U19881 ( .A(n18154), .B(n18153), .Z(n18183) );
  XNOR U19882 ( .A(sreg[1396]), .B(n18183), .Z(n18185) );
  NANDN U19883 ( .A(sreg[1395]), .B(n18146), .Z(n18150) );
  NAND U19884 ( .A(n18148), .B(n18147), .Z(n18149) );
  NAND U19885 ( .A(n18150), .B(n18149), .Z(n18184) );
  XNOR U19886 ( .A(n18185), .B(n18184), .Z(c[1396]) );
  NANDN U19887 ( .A(n18152), .B(n18151), .Z(n18156) );
  NANDN U19888 ( .A(n18154), .B(n18153), .Z(n18155) );
  AND U19889 ( .A(n18156), .B(n18155), .Z(n18191) );
  NANDN U19890 ( .A(n18158), .B(n18157), .Z(n18162) );
  NANDN U19891 ( .A(n18160), .B(n18159), .Z(n18161) );
  AND U19892 ( .A(n18162), .B(n18161), .Z(n18189) );
  NAND U19893 ( .A(n42143), .B(n18163), .Z(n18165) );
  XNOR U19894 ( .A(a[375]), .B(n4125), .Z(n18200) );
  NAND U19895 ( .A(n42144), .B(n18200), .Z(n18164) );
  AND U19896 ( .A(n18165), .B(n18164), .Z(n18215) );
  XOR U19897 ( .A(a[379]), .B(n42012), .Z(n18203) );
  XNOR U19898 ( .A(n18215), .B(n18214), .Z(n18217) );
  XOR U19899 ( .A(a[377]), .B(n42085), .Z(n18207) );
  AND U19900 ( .A(a[373]), .B(b[7]), .Z(n18208) );
  XNOR U19901 ( .A(n18209), .B(n18208), .Z(n18210) );
  AND U19902 ( .A(a[381]), .B(b[0]), .Z(n18168) );
  XNOR U19903 ( .A(n18168), .B(n4071), .Z(n18170) );
  NANDN U19904 ( .A(b[0]), .B(a[380]), .Z(n18169) );
  NAND U19905 ( .A(n18170), .B(n18169), .Z(n18211) );
  XNOR U19906 ( .A(n18210), .B(n18211), .Z(n18216) );
  XOR U19907 ( .A(n18217), .B(n18216), .Z(n18195) );
  NANDN U19908 ( .A(n18172), .B(n18171), .Z(n18176) );
  NANDN U19909 ( .A(n18174), .B(n18173), .Z(n18175) );
  AND U19910 ( .A(n18176), .B(n18175), .Z(n18194) );
  XNOR U19911 ( .A(n18195), .B(n18194), .Z(n18196) );
  NANDN U19912 ( .A(n18178), .B(n18177), .Z(n18182) );
  NAND U19913 ( .A(n18180), .B(n18179), .Z(n18181) );
  NAND U19914 ( .A(n18182), .B(n18181), .Z(n18197) );
  XNOR U19915 ( .A(n18196), .B(n18197), .Z(n18188) );
  XNOR U19916 ( .A(n18189), .B(n18188), .Z(n18190) );
  XNOR U19917 ( .A(n18191), .B(n18190), .Z(n18220) );
  XNOR U19918 ( .A(sreg[1397]), .B(n18220), .Z(n18222) );
  NANDN U19919 ( .A(sreg[1396]), .B(n18183), .Z(n18187) );
  NAND U19920 ( .A(n18185), .B(n18184), .Z(n18186) );
  NAND U19921 ( .A(n18187), .B(n18186), .Z(n18221) );
  XNOR U19922 ( .A(n18222), .B(n18221), .Z(c[1397]) );
  NANDN U19923 ( .A(n18189), .B(n18188), .Z(n18193) );
  NANDN U19924 ( .A(n18191), .B(n18190), .Z(n18192) );
  AND U19925 ( .A(n18193), .B(n18192), .Z(n18228) );
  NANDN U19926 ( .A(n18195), .B(n18194), .Z(n18199) );
  NANDN U19927 ( .A(n18197), .B(n18196), .Z(n18198) );
  AND U19928 ( .A(n18199), .B(n18198), .Z(n18226) );
  NAND U19929 ( .A(n42143), .B(n18200), .Z(n18202) );
  XNOR U19930 ( .A(a[376]), .B(n4125), .Z(n18237) );
  NAND U19931 ( .A(n42144), .B(n18237), .Z(n18201) );
  AND U19932 ( .A(n18202), .B(n18201), .Z(n18252) );
  XOR U19933 ( .A(a[380]), .B(n42012), .Z(n18240) );
  XNOR U19934 ( .A(n18252), .B(n18251), .Z(n18254) );
  AND U19935 ( .A(a[382]), .B(b[0]), .Z(n18204) );
  XNOR U19936 ( .A(n18204), .B(n4071), .Z(n18206) );
  NANDN U19937 ( .A(b[0]), .B(a[381]), .Z(n18205) );
  NAND U19938 ( .A(n18206), .B(n18205), .Z(n18248) );
  XOR U19939 ( .A(a[378]), .B(n42085), .Z(n18244) );
  AND U19940 ( .A(a[374]), .B(b[7]), .Z(n18245) );
  XNOR U19941 ( .A(n18246), .B(n18245), .Z(n18247) );
  XNOR U19942 ( .A(n18248), .B(n18247), .Z(n18253) );
  XOR U19943 ( .A(n18254), .B(n18253), .Z(n18232) );
  NANDN U19944 ( .A(n18209), .B(n18208), .Z(n18213) );
  NANDN U19945 ( .A(n18211), .B(n18210), .Z(n18212) );
  AND U19946 ( .A(n18213), .B(n18212), .Z(n18231) );
  XNOR U19947 ( .A(n18232), .B(n18231), .Z(n18233) );
  NANDN U19948 ( .A(n18215), .B(n18214), .Z(n18219) );
  NAND U19949 ( .A(n18217), .B(n18216), .Z(n18218) );
  NAND U19950 ( .A(n18219), .B(n18218), .Z(n18234) );
  XNOR U19951 ( .A(n18233), .B(n18234), .Z(n18225) );
  XNOR U19952 ( .A(n18226), .B(n18225), .Z(n18227) );
  XNOR U19953 ( .A(n18228), .B(n18227), .Z(n18257) );
  XNOR U19954 ( .A(sreg[1398]), .B(n18257), .Z(n18259) );
  NANDN U19955 ( .A(sreg[1397]), .B(n18220), .Z(n18224) );
  NAND U19956 ( .A(n18222), .B(n18221), .Z(n18223) );
  NAND U19957 ( .A(n18224), .B(n18223), .Z(n18258) );
  XNOR U19958 ( .A(n18259), .B(n18258), .Z(c[1398]) );
  NANDN U19959 ( .A(n18226), .B(n18225), .Z(n18230) );
  NANDN U19960 ( .A(n18228), .B(n18227), .Z(n18229) );
  AND U19961 ( .A(n18230), .B(n18229), .Z(n18265) );
  NANDN U19962 ( .A(n18232), .B(n18231), .Z(n18236) );
  NANDN U19963 ( .A(n18234), .B(n18233), .Z(n18235) );
  AND U19964 ( .A(n18236), .B(n18235), .Z(n18263) );
  NAND U19965 ( .A(n42143), .B(n18237), .Z(n18239) );
  XNOR U19966 ( .A(a[377]), .B(n4125), .Z(n18274) );
  NAND U19967 ( .A(n42144), .B(n18274), .Z(n18238) );
  AND U19968 ( .A(n18239), .B(n18238), .Z(n18289) );
  XOR U19969 ( .A(a[381]), .B(n42012), .Z(n18277) );
  XNOR U19970 ( .A(n18289), .B(n18288), .Z(n18291) );
  AND U19971 ( .A(a[383]), .B(b[0]), .Z(n18241) );
  XNOR U19972 ( .A(n18241), .B(n4071), .Z(n18243) );
  NANDN U19973 ( .A(b[0]), .B(a[382]), .Z(n18242) );
  NAND U19974 ( .A(n18243), .B(n18242), .Z(n18285) );
  XOR U19975 ( .A(a[379]), .B(n42085), .Z(n18281) );
  AND U19976 ( .A(a[375]), .B(b[7]), .Z(n18282) );
  XNOR U19977 ( .A(n18283), .B(n18282), .Z(n18284) );
  XNOR U19978 ( .A(n18285), .B(n18284), .Z(n18290) );
  XOR U19979 ( .A(n18291), .B(n18290), .Z(n18269) );
  NANDN U19980 ( .A(n18246), .B(n18245), .Z(n18250) );
  NANDN U19981 ( .A(n18248), .B(n18247), .Z(n18249) );
  AND U19982 ( .A(n18250), .B(n18249), .Z(n18268) );
  XNOR U19983 ( .A(n18269), .B(n18268), .Z(n18270) );
  NANDN U19984 ( .A(n18252), .B(n18251), .Z(n18256) );
  NAND U19985 ( .A(n18254), .B(n18253), .Z(n18255) );
  NAND U19986 ( .A(n18256), .B(n18255), .Z(n18271) );
  XNOR U19987 ( .A(n18270), .B(n18271), .Z(n18262) );
  XNOR U19988 ( .A(n18263), .B(n18262), .Z(n18264) );
  XNOR U19989 ( .A(n18265), .B(n18264), .Z(n18294) );
  XNOR U19990 ( .A(sreg[1399]), .B(n18294), .Z(n18296) );
  NANDN U19991 ( .A(sreg[1398]), .B(n18257), .Z(n18261) );
  NAND U19992 ( .A(n18259), .B(n18258), .Z(n18260) );
  NAND U19993 ( .A(n18261), .B(n18260), .Z(n18295) );
  XNOR U19994 ( .A(n18296), .B(n18295), .Z(c[1399]) );
  NANDN U19995 ( .A(n18263), .B(n18262), .Z(n18267) );
  NANDN U19996 ( .A(n18265), .B(n18264), .Z(n18266) );
  AND U19997 ( .A(n18267), .B(n18266), .Z(n18302) );
  NANDN U19998 ( .A(n18269), .B(n18268), .Z(n18273) );
  NANDN U19999 ( .A(n18271), .B(n18270), .Z(n18272) );
  AND U20000 ( .A(n18273), .B(n18272), .Z(n18300) );
  NAND U20001 ( .A(n42143), .B(n18274), .Z(n18276) );
  XNOR U20002 ( .A(a[378]), .B(n4125), .Z(n18311) );
  NAND U20003 ( .A(n42144), .B(n18311), .Z(n18275) );
  AND U20004 ( .A(n18276), .B(n18275), .Z(n18326) );
  XOR U20005 ( .A(a[382]), .B(n42012), .Z(n18314) );
  XNOR U20006 ( .A(n18326), .B(n18325), .Z(n18328) );
  AND U20007 ( .A(a[384]), .B(b[0]), .Z(n18278) );
  XNOR U20008 ( .A(n18278), .B(n4071), .Z(n18280) );
  NANDN U20009 ( .A(b[0]), .B(a[383]), .Z(n18279) );
  NAND U20010 ( .A(n18280), .B(n18279), .Z(n18322) );
  XOR U20011 ( .A(a[380]), .B(n42085), .Z(n18318) );
  AND U20012 ( .A(a[376]), .B(b[7]), .Z(n18319) );
  XNOR U20013 ( .A(n18320), .B(n18319), .Z(n18321) );
  XNOR U20014 ( .A(n18322), .B(n18321), .Z(n18327) );
  XOR U20015 ( .A(n18328), .B(n18327), .Z(n18306) );
  NANDN U20016 ( .A(n18283), .B(n18282), .Z(n18287) );
  NANDN U20017 ( .A(n18285), .B(n18284), .Z(n18286) );
  AND U20018 ( .A(n18287), .B(n18286), .Z(n18305) );
  XNOR U20019 ( .A(n18306), .B(n18305), .Z(n18307) );
  NANDN U20020 ( .A(n18289), .B(n18288), .Z(n18293) );
  NAND U20021 ( .A(n18291), .B(n18290), .Z(n18292) );
  NAND U20022 ( .A(n18293), .B(n18292), .Z(n18308) );
  XNOR U20023 ( .A(n18307), .B(n18308), .Z(n18299) );
  XNOR U20024 ( .A(n18300), .B(n18299), .Z(n18301) );
  XNOR U20025 ( .A(n18302), .B(n18301), .Z(n18331) );
  XNOR U20026 ( .A(sreg[1400]), .B(n18331), .Z(n18333) );
  NANDN U20027 ( .A(sreg[1399]), .B(n18294), .Z(n18298) );
  NAND U20028 ( .A(n18296), .B(n18295), .Z(n18297) );
  NAND U20029 ( .A(n18298), .B(n18297), .Z(n18332) );
  XNOR U20030 ( .A(n18333), .B(n18332), .Z(c[1400]) );
  NANDN U20031 ( .A(n18300), .B(n18299), .Z(n18304) );
  NANDN U20032 ( .A(n18302), .B(n18301), .Z(n18303) );
  AND U20033 ( .A(n18304), .B(n18303), .Z(n18339) );
  NANDN U20034 ( .A(n18306), .B(n18305), .Z(n18310) );
  NANDN U20035 ( .A(n18308), .B(n18307), .Z(n18309) );
  AND U20036 ( .A(n18310), .B(n18309), .Z(n18337) );
  NAND U20037 ( .A(n42143), .B(n18311), .Z(n18313) );
  XNOR U20038 ( .A(a[379]), .B(n4126), .Z(n18348) );
  NAND U20039 ( .A(n42144), .B(n18348), .Z(n18312) );
  AND U20040 ( .A(n18313), .B(n18312), .Z(n18363) );
  XOR U20041 ( .A(a[383]), .B(n42012), .Z(n18351) );
  XNOR U20042 ( .A(n18363), .B(n18362), .Z(n18365) );
  AND U20043 ( .A(a[385]), .B(b[0]), .Z(n18315) );
  XNOR U20044 ( .A(n18315), .B(n4071), .Z(n18317) );
  NANDN U20045 ( .A(b[0]), .B(a[384]), .Z(n18316) );
  NAND U20046 ( .A(n18317), .B(n18316), .Z(n18359) );
  XOR U20047 ( .A(a[381]), .B(n42085), .Z(n18355) );
  AND U20048 ( .A(a[377]), .B(b[7]), .Z(n18356) );
  XNOR U20049 ( .A(n18357), .B(n18356), .Z(n18358) );
  XNOR U20050 ( .A(n18359), .B(n18358), .Z(n18364) );
  XOR U20051 ( .A(n18365), .B(n18364), .Z(n18343) );
  NANDN U20052 ( .A(n18320), .B(n18319), .Z(n18324) );
  NANDN U20053 ( .A(n18322), .B(n18321), .Z(n18323) );
  AND U20054 ( .A(n18324), .B(n18323), .Z(n18342) );
  XNOR U20055 ( .A(n18343), .B(n18342), .Z(n18344) );
  NANDN U20056 ( .A(n18326), .B(n18325), .Z(n18330) );
  NAND U20057 ( .A(n18328), .B(n18327), .Z(n18329) );
  NAND U20058 ( .A(n18330), .B(n18329), .Z(n18345) );
  XNOR U20059 ( .A(n18344), .B(n18345), .Z(n18336) );
  XNOR U20060 ( .A(n18337), .B(n18336), .Z(n18338) );
  XNOR U20061 ( .A(n18339), .B(n18338), .Z(n18368) );
  XNOR U20062 ( .A(sreg[1401]), .B(n18368), .Z(n18370) );
  NANDN U20063 ( .A(sreg[1400]), .B(n18331), .Z(n18335) );
  NAND U20064 ( .A(n18333), .B(n18332), .Z(n18334) );
  NAND U20065 ( .A(n18335), .B(n18334), .Z(n18369) );
  XNOR U20066 ( .A(n18370), .B(n18369), .Z(c[1401]) );
  NANDN U20067 ( .A(n18337), .B(n18336), .Z(n18341) );
  NANDN U20068 ( .A(n18339), .B(n18338), .Z(n18340) );
  AND U20069 ( .A(n18341), .B(n18340), .Z(n18376) );
  NANDN U20070 ( .A(n18343), .B(n18342), .Z(n18347) );
  NANDN U20071 ( .A(n18345), .B(n18344), .Z(n18346) );
  AND U20072 ( .A(n18347), .B(n18346), .Z(n18374) );
  NAND U20073 ( .A(n42143), .B(n18348), .Z(n18350) );
  XNOR U20074 ( .A(a[380]), .B(n4126), .Z(n18385) );
  NAND U20075 ( .A(n42144), .B(n18385), .Z(n18349) );
  AND U20076 ( .A(n18350), .B(n18349), .Z(n18400) );
  XOR U20077 ( .A(a[384]), .B(n42012), .Z(n18388) );
  XNOR U20078 ( .A(n18400), .B(n18399), .Z(n18402) );
  AND U20079 ( .A(a[386]), .B(b[0]), .Z(n18352) );
  XNOR U20080 ( .A(n18352), .B(n4071), .Z(n18354) );
  NANDN U20081 ( .A(b[0]), .B(a[385]), .Z(n18353) );
  NAND U20082 ( .A(n18354), .B(n18353), .Z(n18396) );
  XOR U20083 ( .A(a[382]), .B(n42085), .Z(n18392) );
  AND U20084 ( .A(a[378]), .B(b[7]), .Z(n18393) );
  XNOR U20085 ( .A(n18394), .B(n18393), .Z(n18395) );
  XNOR U20086 ( .A(n18396), .B(n18395), .Z(n18401) );
  XOR U20087 ( .A(n18402), .B(n18401), .Z(n18380) );
  NANDN U20088 ( .A(n18357), .B(n18356), .Z(n18361) );
  NANDN U20089 ( .A(n18359), .B(n18358), .Z(n18360) );
  AND U20090 ( .A(n18361), .B(n18360), .Z(n18379) );
  XNOR U20091 ( .A(n18380), .B(n18379), .Z(n18381) );
  NANDN U20092 ( .A(n18363), .B(n18362), .Z(n18367) );
  NAND U20093 ( .A(n18365), .B(n18364), .Z(n18366) );
  NAND U20094 ( .A(n18367), .B(n18366), .Z(n18382) );
  XNOR U20095 ( .A(n18381), .B(n18382), .Z(n18373) );
  XNOR U20096 ( .A(n18374), .B(n18373), .Z(n18375) );
  XNOR U20097 ( .A(n18376), .B(n18375), .Z(n18405) );
  XNOR U20098 ( .A(sreg[1402]), .B(n18405), .Z(n18407) );
  NANDN U20099 ( .A(sreg[1401]), .B(n18368), .Z(n18372) );
  NAND U20100 ( .A(n18370), .B(n18369), .Z(n18371) );
  NAND U20101 ( .A(n18372), .B(n18371), .Z(n18406) );
  XNOR U20102 ( .A(n18407), .B(n18406), .Z(c[1402]) );
  NANDN U20103 ( .A(n18374), .B(n18373), .Z(n18378) );
  NANDN U20104 ( .A(n18376), .B(n18375), .Z(n18377) );
  AND U20105 ( .A(n18378), .B(n18377), .Z(n18413) );
  NANDN U20106 ( .A(n18380), .B(n18379), .Z(n18384) );
  NANDN U20107 ( .A(n18382), .B(n18381), .Z(n18383) );
  AND U20108 ( .A(n18384), .B(n18383), .Z(n18411) );
  NAND U20109 ( .A(n42143), .B(n18385), .Z(n18387) );
  XNOR U20110 ( .A(a[381]), .B(n4126), .Z(n18422) );
  NAND U20111 ( .A(n42144), .B(n18422), .Z(n18386) );
  AND U20112 ( .A(n18387), .B(n18386), .Z(n18437) );
  XOR U20113 ( .A(a[385]), .B(n42012), .Z(n18425) );
  XNOR U20114 ( .A(n18437), .B(n18436), .Z(n18439) );
  AND U20115 ( .A(a[387]), .B(b[0]), .Z(n18389) );
  XNOR U20116 ( .A(n18389), .B(n4071), .Z(n18391) );
  NANDN U20117 ( .A(b[0]), .B(a[386]), .Z(n18390) );
  NAND U20118 ( .A(n18391), .B(n18390), .Z(n18433) );
  XOR U20119 ( .A(a[383]), .B(n42085), .Z(n18429) );
  AND U20120 ( .A(a[379]), .B(b[7]), .Z(n18430) );
  XNOR U20121 ( .A(n18431), .B(n18430), .Z(n18432) );
  XNOR U20122 ( .A(n18433), .B(n18432), .Z(n18438) );
  XOR U20123 ( .A(n18439), .B(n18438), .Z(n18417) );
  NANDN U20124 ( .A(n18394), .B(n18393), .Z(n18398) );
  NANDN U20125 ( .A(n18396), .B(n18395), .Z(n18397) );
  AND U20126 ( .A(n18398), .B(n18397), .Z(n18416) );
  XNOR U20127 ( .A(n18417), .B(n18416), .Z(n18418) );
  NANDN U20128 ( .A(n18400), .B(n18399), .Z(n18404) );
  NAND U20129 ( .A(n18402), .B(n18401), .Z(n18403) );
  NAND U20130 ( .A(n18404), .B(n18403), .Z(n18419) );
  XNOR U20131 ( .A(n18418), .B(n18419), .Z(n18410) );
  XNOR U20132 ( .A(n18411), .B(n18410), .Z(n18412) );
  XNOR U20133 ( .A(n18413), .B(n18412), .Z(n18442) );
  XNOR U20134 ( .A(sreg[1403]), .B(n18442), .Z(n18444) );
  NANDN U20135 ( .A(sreg[1402]), .B(n18405), .Z(n18409) );
  NAND U20136 ( .A(n18407), .B(n18406), .Z(n18408) );
  NAND U20137 ( .A(n18409), .B(n18408), .Z(n18443) );
  XNOR U20138 ( .A(n18444), .B(n18443), .Z(c[1403]) );
  NANDN U20139 ( .A(n18411), .B(n18410), .Z(n18415) );
  NANDN U20140 ( .A(n18413), .B(n18412), .Z(n18414) );
  AND U20141 ( .A(n18415), .B(n18414), .Z(n18450) );
  NANDN U20142 ( .A(n18417), .B(n18416), .Z(n18421) );
  NANDN U20143 ( .A(n18419), .B(n18418), .Z(n18420) );
  AND U20144 ( .A(n18421), .B(n18420), .Z(n18448) );
  NAND U20145 ( .A(n42143), .B(n18422), .Z(n18424) );
  XNOR U20146 ( .A(a[382]), .B(n4126), .Z(n18459) );
  NAND U20147 ( .A(n42144), .B(n18459), .Z(n18423) );
  AND U20148 ( .A(n18424), .B(n18423), .Z(n18474) );
  XOR U20149 ( .A(a[386]), .B(n42012), .Z(n18462) );
  XNOR U20150 ( .A(n18474), .B(n18473), .Z(n18476) );
  AND U20151 ( .A(a[388]), .B(b[0]), .Z(n18426) );
  XNOR U20152 ( .A(n18426), .B(n4071), .Z(n18428) );
  NANDN U20153 ( .A(b[0]), .B(a[387]), .Z(n18427) );
  NAND U20154 ( .A(n18428), .B(n18427), .Z(n18470) );
  XOR U20155 ( .A(a[384]), .B(n42085), .Z(n18463) );
  AND U20156 ( .A(a[380]), .B(b[7]), .Z(n18467) );
  XNOR U20157 ( .A(n18468), .B(n18467), .Z(n18469) );
  XNOR U20158 ( .A(n18470), .B(n18469), .Z(n18475) );
  XOR U20159 ( .A(n18476), .B(n18475), .Z(n18454) );
  NANDN U20160 ( .A(n18431), .B(n18430), .Z(n18435) );
  NANDN U20161 ( .A(n18433), .B(n18432), .Z(n18434) );
  AND U20162 ( .A(n18435), .B(n18434), .Z(n18453) );
  XNOR U20163 ( .A(n18454), .B(n18453), .Z(n18455) );
  NANDN U20164 ( .A(n18437), .B(n18436), .Z(n18441) );
  NAND U20165 ( .A(n18439), .B(n18438), .Z(n18440) );
  NAND U20166 ( .A(n18441), .B(n18440), .Z(n18456) );
  XNOR U20167 ( .A(n18455), .B(n18456), .Z(n18447) );
  XNOR U20168 ( .A(n18448), .B(n18447), .Z(n18449) );
  XNOR U20169 ( .A(n18450), .B(n18449), .Z(n18479) );
  XNOR U20170 ( .A(sreg[1404]), .B(n18479), .Z(n18481) );
  NANDN U20171 ( .A(sreg[1403]), .B(n18442), .Z(n18446) );
  NAND U20172 ( .A(n18444), .B(n18443), .Z(n18445) );
  NAND U20173 ( .A(n18446), .B(n18445), .Z(n18480) );
  XNOR U20174 ( .A(n18481), .B(n18480), .Z(c[1404]) );
  NANDN U20175 ( .A(n18448), .B(n18447), .Z(n18452) );
  NANDN U20176 ( .A(n18450), .B(n18449), .Z(n18451) );
  AND U20177 ( .A(n18452), .B(n18451), .Z(n18487) );
  NANDN U20178 ( .A(n18454), .B(n18453), .Z(n18458) );
  NANDN U20179 ( .A(n18456), .B(n18455), .Z(n18457) );
  AND U20180 ( .A(n18458), .B(n18457), .Z(n18485) );
  NAND U20181 ( .A(n42143), .B(n18459), .Z(n18461) );
  XNOR U20182 ( .A(a[383]), .B(n4126), .Z(n18496) );
  NAND U20183 ( .A(n42144), .B(n18496), .Z(n18460) );
  AND U20184 ( .A(n18461), .B(n18460), .Z(n18511) );
  XOR U20185 ( .A(a[387]), .B(n42012), .Z(n18499) );
  XNOR U20186 ( .A(n18511), .B(n18510), .Z(n18513) );
  XOR U20187 ( .A(a[385]), .B(n42085), .Z(n18503) );
  AND U20188 ( .A(a[381]), .B(b[7]), .Z(n18504) );
  XNOR U20189 ( .A(n18505), .B(n18504), .Z(n18506) );
  AND U20190 ( .A(a[389]), .B(b[0]), .Z(n18464) );
  XNOR U20191 ( .A(n18464), .B(n4071), .Z(n18466) );
  NANDN U20192 ( .A(b[0]), .B(a[388]), .Z(n18465) );
  NAND U20193 ( .A(n18466), .B(n18465), .Z(n18507) );
  XNOR U20194 ( .A(n18506), .B(n18507), .Z(n18512) );
  XOR U20195 ( .A(n18513), .B(n18512), .Z(n18491) );
  NANDN U20196 ( .A(n18468), .B(n18467), .Z(n18472) );
  NANDN U20197 ( .A(n18470), .B(n18469), .Z(n18471) );
  AND U20198 ( .A(n18472), .B(n18471), .Z(n18490) );
  XNOR U20199 ( .A(n18491), .B(n18490), .Z(n18492) );
  NANDN U20200 ( .A(n18474), .B(n18473), .Z(n18478) );
  NAND U20201 ( .A(n18476), .B(n18475), .Z(n18477) );
  NAND U20202 ( .A(n18478), .B(n18477), .Z(n18493) );
  XNOR U20203 ( .A(n18492), .B(n18493), .Z(n18484) );
  XNOR U20204 ( .A(n18485), .B(n18484), .Z(n18486) );
  XNOR U20205 ( .A(n18487), .B(n18486), .Z(n18516) );
  XNOR U20206 ( .A(sreg[1405]), .B(n18516), .Z(n18518) );
  NANDN U20207 ( .A(sreg[1404]), .B(n18479), .Z(n18483) );
  NAND U20208 ( .A(n18481), .B(n18480), .Z(n18482) );
  NAND U20209 ( .A(n18483), .B(n18482), .Z(n18517) );
  XNOR U20210 ( .A(n18518), .B(n18517), .Z(c[1405]) );
  NANDN U20211 ( .A(n18485), .B(n18484), .Z(n18489) );
  NANDN U20212 ( .A(n18487), .B(n18486), .Z(n18488) );
  AND U20213 ( .A(n18489), .B(n18488), .Z(n18524) );
  NANDN U20214 ( .A(n18491), .B(n18490), .Z(n18495) );
  NANDN U20215 ( .A(n18493), .B(n18492), .Z(n18494) );
  AND U20216 ( .A(n18495), .B(n18494), .Z(n18522) );
  NAND U20217 ( .A(n42143), .B(n18496), .Z(n18498) );
  XNOR U20218 ( .A(a[384]), .B(n4126), .Z(n18533) );
  NAND U20219 ( .A(n42144), .B(n18533), .Z(n18497) );
  AND U20220 ( .A(n18498), .B(n18497), .Z(n18548) );
  XOR U20221 ( .A(a[388]), .B(n42012), .Z(n18536) );
  XNOR U20222 ( .A(n18548), .B(n18547), .Z(n18550) );
  AND U20223 ( .A(a[390]), .B(b[0]), .Z(n18500) );
  XNOR U20224 ( .A(n18500), .B(n4071), .Z(n18502) );
  NANDN U20225 ( .A(b[0]), .B(a[389]), .Z(n18501) );
  NAND U20226 ( .A(n18502), .B(n18501), .Z(n18544) );
  XOR U20227 ( .A(a[386]), .B(n42085), .Z(n18540) );
  AND U20228 ( .A(a[382]), .B(b[7]), .Z(n18541) );
  XNOR U20229 ( .A(n18542), .B(n18541), .Z(n18543) );
  XNOR U20230 ( .A(n18544), .B(n18543), .Z(n18549) );
  XOR U20231 ( .A(n18550), .B(n18549), .Z(n18528) );
  NANDN U20232 ( .A(n18505), .B(n18504), .Z(n18509) );
  NANDN U20233 ( .A(n18507), .B(n18506), .Z(n18508) );
  AND U20234 ( .A(n18509), .B(n18508), .Z(n18527) );
  XNOR U20235 ( .A(n18528), .B(n18527), .Z(n18529) );
  NANDN U20236 ( .A(n18511), .B(n18510), .Z(n18515) );
  NAND U20237 ( .A(n18513), .B(n18512), .Z(n18514) );
  NAND U20238 ( .A(n18515), .B(n18514), .Z(n18530) );
  XNOR U20239 ( .A(n18529), .B(n18530), .Z(n18521) );
  XNOR U20240 ( .A(n18522), .B(n18521), .Z(n18523) );
  XNOR U20241 ( .A(n18524), .B(n18523), .Z(n18553) );
  XNOR U20242 ( .A(sreg[1406]), .B(n18553), .Z(n18555) );
  NANDN U20243 ( .A(sreg[1405]), .B(n18516), .Z(n18520) );
  NAND U20244 ( .A(n18518), .B(n18517), .Z(n18519) );
  NAND U20245 ( .A(n18520), .B(n18519), .Z(n18554) );
  XNOR U20246 ( .A(n18555), .B(n18554), .Z(c[1406]) );
  NANDN U20247 ( .A(n18522), .B(n18521), .Z(n18526) );
  NANDN U20248 ( .A(n18524), .B(n18523), .Z(n18525) );
  AND U20249 ( .A(n18526), .B(n18525), .Z(n18561) );
  NANDN U20250 ( .A(n18528), .B(n18527), .Z(n18532) );
  NANDN U20251 ( .A(n18530), .B(n18529), .Z(n18531) );
  AND U20252 ( .A(n18532), .B(n18531), .Z(n18559) );
  NAND U20253 ( .A(n42143), .B(n18533), .Z(n18535) );
  XNOR U20254 ( .A(a[385]), .B(n4126), .Z(n18570) );
  NAND U20255 ( .A(n42144), .B(n18570), .Z(n18534) );
  AND U20256 ( .A(n18535), .B(n18534), .Z(n18585) );
  XOR U20257 ( .A(a[389]), .B(n42012), .Z(n18573) );
  XNOR U20258 ( .A(n18585), .B(n18584), .Z(n18587) );
  AND U20259 ( .A(a[391]), .B(b[0]), .Z(n18537) );
  XNOR U20260 ( .A(n18537), .B(n4071), .Z(n18539) );
  NANDN U20261 ( .A(b[0]), .B(a[390]), .Z(n18538) );
  NAND U20262 ( .A(n18539), .B(n18538), .Z(n18581) );
  XOR U20263 ( .A(a[387]), .B(n42085), .Z(n18577) );
  AND U20264 ( .A(a[383]), .B(b[7]), .Z(n18578) );
  XNOR U20265 ( .A(n18579), .B(n18578), .Z(n18580) );
  XNOR U20266 ( .A(n18581), .B(n18580), .Z(n18586) );
  XOR U20267 ( .A(n18587), .B(n18586), .Z(n18565) );
  NANDN U20268 ( .A(n18542), .B(n18541), .Z(n18546) );
  NANDN U20269 ( .A(n18544), .B(n18543), .Z(n18545) );
  AND U20270 ( .A(n18546), .B(n18545), .Z(n18564) );
  XNOR U20271 ( .A(n18565), .B(n18564), .Z(n18566) );
  NANDN U20272 ( .A(n18548), .B(n18547), .Z(n18552) );
  NAND U20273 ( .A(n18550), .B(n18549), .Z(n18551) );
  NAND U20274 ( .A(n18552), .B(n18551), .Z(n18567) );
  XNOR U20275 ( .A(n18566), .B(n18567), .Z(n18558) );
  XNOR U20276 ( .A(n18559), .B(n18558), .Z(n18560) );
  XNOR U20277 ( .A(n18561), .B(n18560), .Z(n18590) );
  XNOR U20278 ( .A(sreg[1407]), .B(n18590), .Z(n18592) );
  NANDN U20279 ( .A(sreg[1406]), .B(n18553), .Z(n18557) );
  NAND U20280 ( .A(n18555), .B(n18554), .Z(n18556) );
  NAND U20281 ( .A(n18557), .B(n18556), .Z(n18591) );
  XNOR U20282 ( .A(n18592), .B(n18591), .Z(c[1407]) );
  NANDN U20283 ( .A(n18559), .B(n18558), .Z(n18563) );
  NANDN U20284 ( .A(n18561), .B(n18560), .Z(n18562) );
  AND U20285 ( .A(n18563), .B(n18562), .Z(n18598) );
  NANDN U20286 ( .A(n18565), .B(n18564), .Z(n18569) );
  NANDN U20287 ( .A(n18567), .B(n18566), .Z(n18568) );
  AND U20288 ( .A(n18569), .B(n18568), .Z(n18596) );
  NAND U20289 ( .A(n42143), .B(n18570), .Z(n18572) );
  XNOR U20290 ( .A(a[386]), .B(n4127), .Z(n18607) );
  NAND U20291 ( .A(n42144), .B(n18607), .Z(n18571) );
  AND U20292 ( .A(n18572), .B(n18571), .Z(n18622) );
  XOR U20293 ( .A(a[390]), .B(n42012), .Z(n18610) );
  XNOR U20294 ( .A(n18622), .B(n18621), .Z(n18624) );
  AND U20295 ( .A(a[392]), .B(b[0]), .Z(n18574) );
  XNOR U20296 ( .A(n18574), .B(n4071), .Z(n18576) );
  NANDN U20297 ( .A(b[0]), .B(a[391]), .Z(n18575) );
  NAND U20298 ( .A(n18576), .B(n18575), .Z(n18618) );
  XOR U20299 ( .A(a[388]), .B(n42085), .Z(n18611) );
  AND U20300 ( .A(a[384]), .B(b[7]), .Z(n18615) );
  XNOR U20301 ( .A(n18616), .B(n18615), .Z(n18617) );
  XNOR U20302 ( .A(n18618), .B(n18617), .Z(n18623) );
  XOR U20303 ( .A(n18624), .B(n18623), .Z(n18602) );
  NANDN U20304 ( .A(n18579), .B(n18578), .Z(n18583) );
  NANDN U20305 ( .A(n18581), .B(n18580), .Z(n18582) );
  AND U20306 ( .A(n18583), .B(n18582), .Z(n18601) );
  XNOR U20307 ( .A(n18602), .B(n18601), .Z(n18603) );
  NANDN U20308 ( .A(n18585), .B(n18584), .Z(n18589) );
  NAND U20309 ( .A(n18587), .B(n18586), .Z(n18588) );
  NAND U20310 ( .A(n18589), .B(n18588), .Z(n18604) );
  XNOR U20311 ( .A(n18603), .B(n18604), .Z(n18595) );
  XNOR U20312 ( .A(n18596), .B(n18595), .Z(n18597) );
  XNOR U20313 ( .A(n18598), .B(n18597), .Z(n18627) );
  XNOR U20314 ( .A(sreg[1408]), .B(n18627), .Z(n18629) );
  NANDN U20315 ( .A(sreg[1407]), .B(n18590), .Z(n18594) );
  NAND U20316 ( .A(n18592), .B(n18591), .Z(n18593) );
  NAND U20317 ( .A(n18594), .B(n18593), .Z(n18628) );
  XNOR U20318 ( .A(n18629), .B(n18628), .Z(c[1408]) );
  NANDN U20319 ( .A(n18596), .B(n18595), .Z(n18600) );
  NANDN U20320 ( .A(n18598), .B(n18597), .Z(n18599) );
  AND U20321 ( .A(n18600), .B(n18599), .Z(n18635) );
  NANDN U20322 ( .A(n18602), .B(n18601), .Z(n18606) );
  NANDN U20323 ( .A(n18604), .B(n18603), .Z(n18605) );
  AND U20324 ( .A(n18606), .B(n18605), .Z(n18633) );
  NAND U20325 ( .A(n42143), .B(n18607), .Z(n18609) );
  XNOR U20326 ( .A(a[387]), .B(n4127), .Z(n18644) );
  NAND U20327 ( .A(n42144), .B(n18644), .Z(n18608) );
  AND U20328 ( .A(n18609), .B(n18608), .Z(n18659) );
  XOR U20329 ( .A(a[391]), .B(n42012), .Z(n18647) );
  XNOR U20330 ( .A(n18659), .B(n18658), .Z(n18661) );
  XOR U20331 ( .A(a[389]), .B(n42085), .Z(n18648) );
  AND U20332 ( .A(a[385]), .B(b[7]), .Z(n18652) );
  XNOR U20333 ( .A(n18653), .B(n18652), .Z(n18654) );
  AND U20334 ( .A(a[393]), .B(b[0]), .Z(n18612) );
  XNOR U20335 ( .A(n18612), .B(n4071), .Z(n18614) );
  NANDN U20336 ( .A(b[0]), .B(a[392]), .Z(n18613) );
  NAND U20337 ( .A(n18614), .B(n18613), .Z(n18655) );
  XNOR U20338 ( .A(n18654), .B(n18655), .Z(n18660) );
  XOR U20339 ( .A(n18661), .B(n18660), .Z(n18639) );
  NANDN U20340 ( .A(n18616), .B(n18615), .Z(n18620) );
  NANDN U20341 ( .A(n18618), .B(n18617), .Z(n18619) );
  AND U20342 ( .A(n18620), .B(n18619), .Z(n18638) );
  XNOR U20343 ( .A(n18639), .B(n18638), .Z(n18640) );
  NANDN U20344 ( .A(n18622), .B(n18621), .Z(n18626) );
  NAND U20345 ( .A(n18624), .B(n18623), .Z(n18625) );
  NAND U20346 ( .A(n18626), .B(n18625), .Z(n18641) );
  XNOR U20347 ( .A(n18640), .B(n18641), .Z(n18632) );
  XNOR U20348 ( .A(n18633), .B(n18632), .Z(n18634) );
  XNOR U20349 ( .A(n18635), .B(n18634), .Z(n18664) );
  XNOR U20350 ( .A(sreg[1409]), .B(n18664), .Z(n18666) );
  NANDN U20351 ( .A(sreg[1408]), .B(n18627), .Z(n18631) );
  NAND U20352 ( .A(n18629), .B(n18628), .Z(n18630) );
  NAND U20353 ( .A(n18631), .B(n18630), .Z(n18665) );
  XNOR U20354 ( .A(n18666), .B(n18665), .Z(c[1409]) );
  NANDN U20355 ( .A(n18633), .B(n18632), .Z(n18637) );
  NANDN U20356 ( .A(n18635), .B(n18634), .Z(n18636) );
  AND U20357 ( .A(n18637), .B(n18636), .Z(n18672) );
  NANDN U20358 ( .A(n18639), .B(n18638), .Z(n18643) );
  NANDN U20359 ( .A(n18641), .B(n18640), .Z(n18642) );
  AND U20360 ( .A(n18643), .B(n18642), .Z(n18670) );
  NAND U20361 ( .A(n42143), .B(n18644), .Z(n18646) );
  XNOR U20362 ( .A(a[388]), .B(n4127), .Z(n18681) );
  NAND U20363 ( .A(n42144), .B(n18681), .Z(n18645) );
  AND U20364 ( .A(n18646), .B(n18645), .Z(n18696) );
  XOR U20365 ( .A(a[392]), .B(n42012), .Z(n18684) );
  XNOR U20366 ( .A(n18696), .B(n18695), .Z(n18698) );
  XOR U20367 ( .A(a[390]), .B(n42085), .Z(n18688) );
  AND U20368 ( .A(a[386]), .B(b[7]), .Z(n18689) );
  XNOR U20369 ( .A(n18690), .B(n18689), .Z(n18691) );
  AND U20370 ( .A(a[394]), .B(b[0]), .Z(n18649) );
  XNOR U20371 ( .A(n18649), .B(n4071), .Z(n18651) );
  NANDN U20372 ( .A(b[0]), .B(a[393]), .Z(n18650) );
  NAND U20373 ( .A(n18651), .B(n18650), .Z(n18692) );
  XNOR U20374 ( .A(n18691), .B(n18692), .Z(n18697) );
  XOR U20375 ( .A(n18698), .B(n18697), .Z(n18676) );
  NANDN U20376 ( .A(n18653), .B(n18652), .Z(n18657) );
  NANDN U20377 ( .A(n18655), .B(n18654), .Z(n18656) );
  AND U20378 ( .A(n18657), .B(n18656), .Z(n18675) );
  XNOR U20379 ( .A(n18676), .B(n18675), .Z(n18677) );
  NANDN U20380 ( .A(n18659), .B(n18658), .Z(n18663) );
  NAND U20381 ( .A(n18661), .B(n18660), .Z(n18662) );
  NAND U20382 ( .A(n18663), .B(n18662), .Z(n18678) );
  XNOR U20383 ( .A(n18677), .B(n18678), .Z(n18669) );
  XNOR U20384 ( .A(n18670), .B(n18669), .Z(n18671) );
  XNOR U20385 ( .A(n18672), .B(n18671), .Z(n18701) );
  XNOR U20386 ( .A(sreg[1410]), .B(n18701), .Z(n18703) );
  NANDN U20387 ( .A(sreg[1409]), .B(n18664), .Z(n18668) );
  NAND U20388 ( .A(n18666), .B(n18665), .Z(n18667) );
  NAND U20389 ( .A(n18668), .B(n18667), .Z(n18702) );
  XNOR U20390 ( .A(n18703), .B(n18702), .Z(c[1410]) );
  NANDN U20391 ( .A(n18670), .B(n18669), .Z(n18674) );
  NANDN U20392 ( .A(n18672), .B(n18671), .Z(n18673) );
  AND U20393 ( .A(n18674), .B(n18673), .Z(n18709) );
  NANDN U20394 ( .A(n18676), .B(n18675), .Z(n18680) );
  NANDN U20395 ( .A(n18678), .B(n18677), .Z(n18679) );
  AND U20396 ( .A(n18680), .B(n18679), .Z(n18707) );
  NAND U20397 ( .A(n42143), .B(n18681), .Z(n18683) );
  XNOR U20398 ( .A(a[389]), .B(n4127), .Z(n18718) );
  NAND U20399 ( .A(n42144), .B(n18718), .Z(n18682) );
  AND U20400 ( .A(n18683), .B(n18682), .Z(n18733) );
  XOR U20401 ( .A(a[393]), .B(n42012), .Z(n18721) );
  XNOR U20402 ( .A(n18733), .B(n18732), .Z(n18735) );
  AND U20403 ( .A(a[395]), .B(b[0]), .Z(n18685) );
  XNOR U20404 ( .A(n18685), .B(n4071), .Z(n18687) );
  NANDN U20405 ( .A(b[0]), .B(a[394]), .Z(n18686) );
  NAND U20406 ( .A(n18687), .B(n18686), .Z(n18729) );
  XOR U20407 ( .A(a[391]), .B(n42085), .Z(n18725) );
  AND U20408 ( .A(a[387]), .B(b[7]), .Z(n18726) );
  XNOR U20409 ( .A(n18727), .B(n18726), .Z(n18728) );
  XNOR U20410 ( .A(n18729), .B(n18728), .Z(n18734) );
  XOR U20411 ( .A(n18735), .B(n18734), .Z(n18713) );
  NANDN U20412 ( .A(n18690), .B(n18689), .Z(n18694) );
  NANDN U20413 ( .A(n18692), .B(n18691), .Z(n18693) );
  AND U20414 ( .A(n18694), .B(n18693), .Z(n18712) );
  XNOR U20415 ( .A(n18713), .B(n18712), .Z(n18714) );
  NANDN U20416 ( .A(n18696), .B(n18695), .Z(n18700) );
  NAND U20417 ( .A(n18698), .B(n18697), .Z(n18699) );
  NAND U20418 ( .A(n18700), .B(n18699), .Z(n18715) );
  XNOR U20419 ( .A(n18714), .B(n18715), .Z(n18706) );
  XNOR U20420 ( .A(n18707), .B(n18706), .Z(n18708) );
  XNOR U20421 ( .A(n18709), .B(n18708), .Z(n18738) );
  XNOR U20422 ( .A(sreg[1411]), .B(n18738), .Z(n18740) );
  NANDN U20423 ( .A(sreg[1410]), .B(n18701), .Z(n18705) );
  NAND U20424 ( .A(n18703), .B(n18702), .Z(n18704) );
  NAND U20425 ( .A(n18705), .B(n18704), .Z(n18739) );
  XNOR U20426 ( .A(n18740), .B(n18739), .Z(c[1411]) );
  NANDN U20427 ( .A(n18707), .B(n18706), .Z(n18711) );
  NANDN U20428 ( .A(n18709), .B(n18708), .Z(n18710) );
  AND U20429 ( .A(n18711), .B(n18710), .Z(n18746) );
  NANDN U20430 ( .A(n18713), .B(n18712), .Z(n18717) );
  NANDN U20431 ( .A(n18715), .B(n18714), .Z(n18716) );
  AND U20432 ( .A(n18717), .B(n18716), .Z(n18744) );
  NAND U20433 ( .A(n42143), .B(n18718), .Z(n18720) );
  XNOR U20434 ( .A(a[390]), .B(n4127), .Z(n18755) );
  NAND U20435 ( .A(n42144), .B(n18755), .Z(n18719) );
  AND U20436 ( .A(n18720), .B(n18719), .Z(n18770) );
  XOR U20437 ( .A(a[394]), .B(n42012), .Z(n18758) );
  XNOR U20438 ( .A(n18770), .B(n18769), .Z(n18772) );
  AND U20439 ( .A(a[396]), .B(b[0]), .Z(n18722) );
  XNOR U20440 ( .A(n18722), .B(n4071), .Z(n18724) );
  NANDN U20441 ( .A(b[0]), .B(a[395]), .Z(n18723) );
  NAND U20442 ( .A(n18724), .B(n18723), .Z(n18766) );
  XOR U20443 ( .A(a[392]), .B(n42085), .Z(n18759) );
  AND U20444 ( .A(a[388]), .B(b[7]), .Z(n18763) );
  XNOR U20445 ( .A(n18764), .B(n18763), .Z(n18765) );
  XNOR U20446 ( .A(n18766), .B(n18765), .Z(n18771) );
  XOR U20447 ( .A(n18772), .B(n18771), .Z(n18750) );
  NANDN U20448 ( .A(n18727), .B(n18726), .Z(n18731) );
  NANDN U20449 ( .A(n18729), .B(n18728), .Z(n18730) );
  AND U20450 ( .A(n18731), .B(n18730), .Z(n18749) );
  XNOR U20451 ( .A(n18750), .B(n18749), .Z(n18751) );
  NANDN U20452 ( .A(n18733), .B(n18732), .Z(n18737) );
  NAND U20453 ( .A(n18735), .B(n18734), .Z(n18736) );
  NAND U20454 ( .A(n18737), .B(n18736), .Z(n18752) );
  XNOR U20455 ( .A(n18751), .B(n18752), .Z(n18743) );
  XNOR U20456 ( .A(n18744), .B(n18743), .Z(n18745) );
  XNOR U20457 ( .A(n18746), .B(n18745), .Z(n18775) );
  XNOR U20458 ( .A(sreg[1412]), .B(n18775), .Z(n18777) );
  NANDN U20459 ( .A(sreg[1411]), .B(n18738), .Z(n18742) );
  NAND U20460 ( .A(n18740), .B(n18739), .Z(n18741) );
  NAND U20461 ( .A(n18742), .B(n18741), .Z(n18776) );
  XNOR U20462 ( .A(n18777), .B(n18776), .Z(c[1412]) );
  NANDN U20463 ( .A(n18744), .B(n18743), .Z(n18748) );
  NANDN U20464 ( .A(n18746), .B(n18745), .Z(n18747) );
  AND U20465 ( .A(n18748), .B(n18747), .Z(n18783) );
  NANDN U20466 ( .A(n18750), .B(n18749), .Z(n18754) );
  NANDN U20467 ( .A(n18752), .B(n18751), .Z(n18753) );
  AND U20468 ( .A(n18754), .B(n18753), .Z(n18781) );
  NAND U20469 ( .A(n42143), .B(n18755), .Z(n18757) );
  XNOR U20470 ( .A(a[391]), .B(n4127), .Z(n18792) );
  NAND U20471 ( .A(n42144), .B(n18792), .Z(n18756) );
  AND U20472 ( .A(n18757), .B(n18756), .Z(n18807) );
  XOR U20473 ( .A(a[395]), .B(n42012), .Z(n18795) );
  XNOR U20474 ( .A(n18807), .B(n18806), .Z(n18809) );
  XOR U20475 ( .A(a[393]), .B(n42085), .Z(n18796) );
  AND U20476 ( .A(a[389]), .B(b[7]), .Z(n18800) );
  XNOR U20477 ( .A(n18801), .B(n18800), .Z(n18802) );
  AND U20478 ( .A(a[397]), .B(b[0]), .Z(n18760) );
  XNOR U20479 ( .A(n18760), .B(n4071), .Z(n18762) );
  NANDN U20480 ( .A(b[0]), .B(a[396]), .Z(n18761) );
  NAND U20481 ( .A(n18762), .B(n18761), .Z(n18803) );
  XNOR U20482 ( .A(n18802), .B(n18803), .Z(n18808) );
  XOR U20483 ( .A(n18809), .B(n18808), .Z(n18787) );
  NANDN U20484 ( .A(n18764), .B(n18763), .Z(n18768) );
  NANDN U20485 ( .A(n18766), .B(n18765), .Z(n18767) );
  AND U20486 ( .A(n18768), .B(n18767), .Z(n18786) );
  XNOR U20487 ( .A(n18787), .B(n18786), .Z(n18788) );
  NANDN U20488 ( .A(n18770), .B(n18769), .Z(n18774) );
  NAND U20489 ( .A(n18772), .B(n18771), .Z(n18773) );
  NAND U20490 ( .A(n18774), .B(n18773), .Z(n18789) );
  XNOR U20491 ( .A(n18788), .B(n18789), .Z(n18780) );
  XNOR U20492 ( .A(n18781), .B(n18780), .Z(n18782) );
  XNOR U20493 ( .A(n18783), .B(n18782), .Z(n18812) );
  XNOR U20494 ( .A(sreg[1413]), .B(n18812), .Z(n18814) );
  NANDN U20495 ( .A(sreg[1412]), .B(n18775), .Z(n18779) );
  NAND U20496 ( .A(n18777), .B(n18776), .Z(n18778) );
  NAND U20497 ( .A(n18779), .B(n18778), .Z(n18813) );
  XNOR U20498 ( .A(n18814), .B(n18813), .Z(c[1413]) );
  NANDN U20499 ( .A(n18781), .B(n18780), .Z(n18785) );
  NANDN U20500 ( .A(n18783), .B(n18782), .Z(n18784) );
  AND U20501 ( .A(n18785), .B(n18784), .Z(n18820) );
  NANDN U20502 ( .A(n18787), .B(n18786), .Z(n18791) );
  NANDN U20503 ( .A(n18789), .B(n18788), .Z(n18790) );
  AND U20504 ( .A(n18791), .B(n18790), .Z(n18818) );
  NAND U20505 ( .A(n42143), .B(n18792), .Z(n18794) );
  XNOR U20506 ( .A(a[392]), .B(n4127), .Z(n18829) );
  NAND U20507 ( .A(n42144), .B(n18829), .Z(n18793) );
  AND U20508 ( .A(n18794), .B(n18793), .Z(n18844) );
  XOR U20509 ( .A(a[396]), .B(n42012), .Z(n18832) );
  XNOR U20510 ( .A(n18844), .B(n18843), .Z(n18846) );
  XOR U20511 ( .A(a[394]), .B(n42085), .Z(n18833) );
  AND U20512 ( .A(a[390]), .B(b[7]), .Z(n18837) );
  XNOR U20513 ( .A(n18838), .B(n18837), .Z(n18839) );
  AND U20514 ( .A(a[398]), .B(b[0]), .Z(n18797) );
  XNOR U20515 ( .A(n18797), .B(n4071), .Z(n18799) );
  NANDN U20516 ( .A(b[0]), .B(a[397]), .Z(n18798) );
  NAND U20517 ( .A(n18799), .B(n18798), .Z(n18840) );
  XNOR U20518 ( .A(n18839), .B(n18840), .Z(n18845) );
  XOR U20519 ( .A(n18846), .B(n18845), .Z(n18824) );
  NANDN U20520 ( .A(n18801), .B(n18800), .Z(n18805) );
  NANDN U20521 ( .A(n18803), .B(n18802), .Z(n18804) );
  AND U20522 ( .A(n18805), .B(n18804), .Z(n18823) );
  XNOR U20523 ( .A(n18824), .B(n18823), .Z(n18825) );
  NANDN U20524 ( .A(n18807), .B(n18806), .Z(n18811) );
  NAND U20525 ( .A(n18809), .B(n18808), .Z(n18810) );
  NAND U20526 ( .A(n18811), .B(n18810), .Z(n18826) );
  XNOR U20527 ( .A(n18825), .B(n18826), .Z(n18817) );
  XNOR U20528 ( .A(n18818), .B(n18817), .Z(n18819) );
  XNOR U20529 ( .A(n18820), .B(n18819), .Z(n18849) );
  XNOR U20530 ( .A(sreg[1414]), .B(n18849), .Z(n18851) );
  NANDN U20531 ( .A(sreg[1413]), .B(n18812), .Z(n18816) );
  NAND U20532 ( .A(n18814), .B(n18813), .Z(n18815) );
  NAND U20533 ( .A(n18816), .B(n18815), .Z(n18850) );
  XNOR U20534 ( .A(n18851), .B(n18850), .Z(c[1414]) );
  NANDN U20535 ( .A(n18818), .B(n18817), .Z(n18822) );
  NANDN U20536 ( .A(n18820), .B(n18819), .Z(n18821) );
  AND U20537 ( .A(n18822), .B(n18821), .Z(n18857) );
  NANDN U20538 ( .A(n18824), .B(n18823), .Z(n18828) );
  NANDN U20539 ( .A(n18826), .B(n18825), .Z(n18827) );
  AND U20540 ( .A(n18828), .B(n18827), .Z(n18855) );
  NAND U20541 ( .A(n42143), .B(n18829), .Z(n18831) );
  XNOR U20542 ( .A(a[393]), .B(n4128), .Z(n18866) );
  NAND U20543 ( .A(n42144), .B(n18866), .Z(n18830) );
  AND U20544 ( .A(n18831), .B(n18830), .Z(n18881) );
  XOR U20545 ( .A(a[397]), .B(n42012), .Z(n18869) );
  XNOR U20546 ( .A(n18881), .B(n18880), .Z(n18883) );
  XOR U20547 ( .A(a[395]), .B(n42085), .Z(n18873) );
  AND U20548 ( .A(a[391]), .B(b[7]), .Z(n18874) );
  XNOR U20549 ( .A(n18875), .B(n18874), .Z(n18876) );
  AND U20550 ( .A(a[399]), .B(b[0]), .Z(n18834) );
  XNOR U20551 ( .A(n18834), .B(n4071), .Z(n18836) );
  NANDN U20552 ( .A(b[0]), .B(a[398]), .Z(n18835) );
  NAND U20553 ( .A(n18836), .B(n18835), .Z(n18877) );
  XNOR U20554 ( .A(n18876), .B(n18877), .Z(n18882) );
  XOR U20555 ( .A(n18883), .B(n18882), .Z(n18861) );
  NANDN U20556 ( .A(n18838), .B(n18837), .Z(n18842) );
  NANDN U20557 ( .A(n18840), .B(n18839), .Z(n18841) );
  AND U20558 ( .A(n18842), .B(n18841), .Z(n18860) );
  XNOR U20559 ( .A(n18861), .B(n18860), .Z(n18862) );
  NANDN U20560 ( .A(n18844), .B(n18843), .Z(n18848) );
  NAND U20561 ( .A(n18846), .B(n18845), .Z(n18847) );
  NAND U20562 ( .A(n18848), .B(n18847), .Z(n18863) );
  XNOR U20563 ( .A(n18862), .B(n18863), .Z(n18854) );
  XNOR U20564 ( .A(n18855), .B(n18854), .Z(n18856) );
  XNOR U20565 ( .A(n18857), .B(n18856), .Z(n18886) );
  XNOR U20566 ( .A(sreg[1415]), .B(n18886), .Z(n18888) );
  NANDN U20567 ( .A(sreg[1414]), .B(n18849), .Z(n18853) );
  NAND U20568 ( .A(n18851), .B(n18850), .Z(n18852) );
  NAND U20569 ( .A(n18853), .B(n18852), .Z(n18887) );
  XNOR U20570 ( .A(n18888), .B(n18887), .Z(c[1415]) );
  NANDN U20571 ( .A(n18855), .B(n18854), .Z(n18859) );
  NANDN U20572 ( .A(n18857), .B(n18856), .Z(n18858) );
  AND U20573 ( .A(n18859), .B(n18858), .Z(n18894) );
  NANDN U20574 ( .A(n18861), .B(n18860), .Z(n18865) );
  NANDN U20575 ( .A(n18863), .B(n18862), .Z(n18864) );
  AND U20576 ( .A(n18865), .B(n18864), .Z(n18892) );
  NAND U20577 ( .A(n42143), .B(n18866), .Z(n18868) );
  XNOR U20578 ( .A(a[394]), .B(n4128), .Z(n18903) );
  NAND U20579 ( .A(n42144), .B(n18903), .Z(n18867) );
  AND U20580 ( .A(n18868), .B(n18867), .Z(n18918) );
  XOR U20581 ( .A(a[398]), .B(n42012), .Z(n18906) );
  XNOR U20582 ( .A(n18918), .B(n18917), .Z(n18920) );
  AND U20583 ( .A(a[400]), .B(b[0]), .Z(n18870) );
  XNOR U20584 ( .A(n18870), .B(n4071), .Z(n18872) );
  NANDN U20585 ( .A(b[0]), .B(a[399]), .Z(n18871) );
  NAND U20586 ( .A(n18872), .B(n18871), .Z(n18914) );
  XOR U20587 ( .A(a[396]), .B(n42085), .Z(n18907) );
  AND U20588 ( .A(a[392]), .B(b[7]), .Z(n18911) );
  XNOR U20589 ( .A(n18912), .B(n18911), .Z(n18913) );
  XNOR U20590 ( .A(n18914), .B(n18913), .Z(n18919) );
  XOR U20591 ( .A(n18920), .B(n18919), .Z(n18898) );
  NANDN U20592 ( .A(n18875), .B(n18874), .Z(n18879) );
  NANDN U20593 ( .A(n18877), .B(n18876), .Z(n18878) );
  AND U20594 ( .A(n18879), .B(n18878), .Z(n18897) );
  XNOR U20595 ( .A(n18898), .B(n18897), .Z(n18899) );
  NANDN U20596 ( .A(n18881), .B(n18880), .Z(n18885) );
  NAND U20597 ( .A(n18883), .B(n18882), .Z(n18884) );
  NAND U20598 ( .A(n18885), .B(n18884), .Z(n18900) );
  XNOR U20599 ( .A(n18899), .B(n18900), .Z(n18891) );
  XNOR U20600 ( .A(n18892), .B(n18891), .Z(n18893) );
  XNOR U20601 ( .A(n18894), .B(n18893), .Z(n18923) );
  XNOR U20602 ( .A(sreg[1416]), .B(n18923), .Z(n18925) );
  NANDN U20603 ( .A(sreg[1415]), .B(n18886), .Z(n18890) );
  NAND U20604 ( .A(n18888), .B(n18887), .Z(n18889) );
  NAND U20605 ( .A(n18890), .B(n18889), .Z(n18924) );
  XNOR U20606 ( .A(n18925), .B(n18924), .Z(c[1416]) );
  NANDN U20607 ( .A(n18892), .B(n18891), .Z(n18896) );
  NANDN U20608 ( .A(n18894), .B(n18893), .Z(n18895) );
  AND U20609 ( .A(n18896), .B(n18895), .Z(n18931) );
  NANDN U20610 ( .A(n18898), .B(n18897), .Z(n18902) );
  NANDN U20611 ( .A(n18900), .B(n18899), .Z(n18901) );
  AND U20612 ( .A(n18902), .B(n18901), .Z(n18929) );
  NAND U20613 ( .A(n42143), .B(n18903), .Z(n18905) );
  XNOR U20614 ( .A(a[395]), .B(n4128), .Z(n18940) );
  NAND U20615 ( .A(n42144), .B(n18940), .Z(n18904) );
  AND U20616 ( .A(n18905), .B(n18904), .Z(n18955) );
  XOR U20617 ( .A(a[399]), .B(n42012), .Z(n18943) );
  XNOR U20618 ( .A(n18955), .B(n18954), .Z(n18957) );
  XOR U20619 ( .A(a[397]), .B(n42085), .Z(n18944) );
  AND U20620 ( .A(a[393]), .B(b[7]), .Z(n18948) );
  XNOR U20621 ( .A(n18949), .B(n18948), .Z(n18950) );
  AND U20622 ( .A(a[401]), .B(b[0]), .Z(n18908) );
  XNOR U20623 ( .A(n18908), .B(n4071), .Z(n18910) );
  NANDN U20624 ( .A(b[0]), .B(a[400]), .Z(n18909) );
  NAND U20625 ( .A(n18910), .B(n18909), .Z(n18951) );
  XNOR U20626 ( .A(n18950), .B(n18951), .Z(n18956) );
  XOR U20627 ( .A(n18957), .B(n18956), .Z(n18935) );
  NANDN U20628 ( .A(n18912), .B(n18911), .Z(n18916) );
  NANDN U20629 ( .A(n18914), .B(n18913), .Z(n18915) );
  AND U20630 ( .A(n18916), .B(n18915), .Z(n18934) );
  XNOR U20631 ( .A(n18935), .B(n18934), .Z(n18936) );
  NANDN U20632 ( .A(n18918), .B(n18917), .Z(n18922) );
  NAND U20633 ( .A(n18920), .B(n18919), .Z(n18921) );
  NAND U20634 ( .A(n18922), .B(n18921), .Z(n18937) );
  XNOR U20635 ( .A(n18936), .B(n18937), .Z(n18928) );
  XNOR U20636 ( .A(n18929), .B(n18928), .Z(n18930) );
  XNOR U20637 ( .A(n18931), .B(n18930), .Z(n18960) );
  XNOR U20638 ( .A(sreg[1417]), .B(n18960), .Z(n18962) );
  NANDN U20639 ( .A(sreg[1416]), .B(n18923), .Z(n18927) );
  NAND U20640 ( .A(n18925), .B(n18924), .Z(n18926) );
  NAND U20641 ( .A(n18927), .B(n18926), .Z(n18961) );
  XNOR U20642 ( .A(n18962), .B(n18961), .Z(c[1417]) );
  NANDN U20643 ( .A(n18929), .B(n18928), .Z(n18933) );
  NANDN U20644 ( .A(n18931), .B(n18930), .Z(n18932) );
  AND U20645 ( .A(n18933), .B(n18932), .Z(n18968) );
  NANDN U20646 ( .A(n18935), .B(n18934), .Z(n18939) );
  NANDN U20647 ( .A(n18937), .B(n18936), .Z(n18938) );
  AND U20648 ( .A(n18939), .B(n18938), .Z(n18966) );
  NAND U20649 ( .A(n42143), .B(n18940), .Z(n18942) );
  XNOR U20650 ( .A(a[396]), .B(n4128), .Z(n18977) );
  NAND U20651 ( .A(n42144), .B(n18977), .Z(n18941) );
  AND U20652 ( .A(n18942), .B(n18941), .Z(n18992) );
  XOR U20653 ( .A(a[400]), .B(n42012), .Z(n18980) );
  XNOR U20654 ( .A(n18992), .B(n18991), .Z(n18994) );
  XOR U20655 ( .A(a[398]), .B(n42085), .Z(n18984) );
  AND U20656 ( .A(a[394]), .B(b[7]), .Z(n18985) );
  XNOR U20657 ( .A(n18986), .B(n18985), .Z(n18987) );
  AND U20658 ( .A(a[402]), .B(b[0]), .Z(n18945) );
  XNOR U20659 ( .A(n18945), .B(n4071), .Z(n18947) );
  NANDN U20660 ( .A(b[0]), .B(a[401]), .Z(n18946) );
  NAND U20661 ( .A(n18947), .B(n18946), .Z(n18988) );
  XNOR U20662 ( .A(n18987), .B(n18988), .Z(n18993) );
  XOR U20663 ( .A(n18994), .B(n18993), .Z(n18972) );
  NANDN U20664 ( .A(n18949), .B(n18948), .Z(n18953) );
  NANDN U20665 ( .A(n18951), .B(n18950), .Z(n18952) );
  AND U20666 ( .A(n18953), .B(n18952), .Z(n18971) );
  XNOR U20667 ( .A(n18972), .B(n18971), .Z(n18973) );
  NANDN U20668 ( .A(n18955), .B(n18954), .Z(n18959) );
  NAND U20669 ( .A(n18957), .B(n18956), .Z(n18958) );
  NAND U20670 ( .A(n18959), .B(n18958), .Z(n18974) );
  XNOR U20671 ( .A(n18973), .B(n18974), .Z(n18965) );
  XNOR U20672 ( .A(n18966), .B(n18965), .Z(n18967) );
  XNOR U20673 ( .A(n18968), .B(n18967), .Z(n18997) );
  XNOR U20674 ( .A(sreg[1418]), .B(n18997), .Z(n18999) );
  NANDN U20675 ( .A(sreg[1417]), .B(n18960), .Z(n18964) );
  NAND U20676 ( .A(n18962), .B(n18961), .Z(n18963) );
  NAND U20677 ( .A(n18964), .B(n18963), .Z(n18998) );
  XNOR U20678 ( .A(n18999), .B(n18998), .Z(c[1418]) );
  NANDN U20679 ( .A(n18966), .B(n18965), .Z(n18970) );
  NANDN U20680 ( .A(n18968), .B(n18967), .Z(n18969) );
  AND U20681 ( .A(n18970), .B(n18969), .Z(n19005) );
  NANDN U20682 ( .A(n18972), .B(n18971), .Z(n18976) );
  NANDN U20683 ( .A(n18974), .B(n18973), .Z(n18975) );
  AND U20684 ( .A(n18976), .B(n18975), .Z(n19003) );
  NAND U20685 ( .A(n42143), .B(n18977), .Z(n18979) );
  XNOR U20686 ( .A(a[397]), .B(n4128), .Z(n19014) );
  NAND U20687 ( .A(n42144), .B(n19014), .Z(n18978) );
  AND U20688 ( .A(n18979), .B(n18978), .Z(n19029) );
  XOR U20689 ( .A(a[401]), .B(n42012), .Z(n19017) );
  XNOR U20690 ( .A(n19029), .B(n19028), .Z(n19031) );
  AND U20691 ( .A(a[403]), .B(b[0]), .Z(n18981) );
  XNOR U20692 ( .A(n18981), .B(n4071), .Z(n18983) );
  NANDN U20693 ( .A(b[0]), .B(a[402]), .Z(n18982) );
  NAND U20694 ( .A(n18983), .B(n18982), .Z(n19025) );
  XOR U20695 ( .A(a[399]), .B(n42085), .Z(n19018) );
  AND U20696 ( .A(a[395]), .B(b[7]), .Z(n19022) );
  XNOR U20697 ( .A(n19023), .B(n19022), .Z(n19024) );
  XNOR U20698 ( .A(n19025), .B(n19024), .Z(n19030) );
  XOR U20699 ( .A(n19031), .B(n19030), .Z(n19009) );
  NANDN U20700 ( .A(n18986), .B(n18985), .Z(n18990) );
  NANDN U20701 ( .A(n18988), .B(n18987), .Z(n18989) );
  AND U20702 ( .A(n18990), .B(n18989), .Z(n19008) );
  XNOR U20703 ( .A(n19009), .B(n19008), .Z(n19010) );
  NANDN U20704 ( .A(n18992), .B(n18991), .Z(n18996) );
  NAND U20705 ( .A(n18994), .B(n18993), .Z(n18995) );
  NAND U20706 ( .A(n18996), .B(n18995), .Z(n19011) );
  XNOR U20707 ( .A(n19010), .B(n19011), .Z(n19002) );
  XNOR U20708 ( .A(n19003), .B(n19002), .Z(n19004) );
  XNOR U20709 ( .A(n19005), .B(n19004), .Z(n19034) );
  XNOR U20710 ( .A(sreg[1419]), .B(n19034), .Z(n19036) );
  NANDN U20711 ( .A(sreg[1418]), .B(n18997), .Z(n19001) );
  NAND U20712 ( .A(n18999), .B(n18998), .Z(n19000) );
  NAND U20713 ( .A(n19001), .B(n19000), .Z(n19035) );
  XNOR U20714 ( .A(n19036), .B(n19035), .Z(c[1419]) );
  NANDN U20715 ( .A(n19003), .B(n19002), .Z(n19007) );
  NANDN U20716 ( .A(n19005), .B(n19004), .Z(n19006) );
  AND U20717 ( .A(n19007), .B(n19006), .Z(n19042) );
  NANDN U20718 ( .A(n19009), .B(n19008), .Z(n19013) );
  NANDN U20719 ( .A(n19011), .B(n19010), .Z(n19012) );
  AND U20720 ( .A(n19013), .B(n19012), .Z(n19040) );
  NAND U20721 ( .A(n42143), .B(n19014), .Z(n19016) );
  XNOR U20722 ( .A(a[398]), .B(n4128), .Z(n19051) );
  NAND U20723 ( .A(n42144), .B(n19051), .Z(n19015) );
  AND U20724 ( .A(n19016), .B(n19015), .Z(n19066) );
  XOR U20725 ( .A(a[402]), .B(n42012), .Z(n19054) );
  XNOR U20726 ( .A(n19066), .B(n19065), .Z(n19068) );
  XOR U20727 ( .A(a[400]), .B(n42085), .Z(n19058) );
  AND U20728 ( .A(a[396]), .B(b[7]), .Z(n19059) );
  XNOR U20729 ( .A(n19060), .B(n19059), .Z(n19061) );
  AND U20730 ( .A(a[404]), .B(b[0]), .Z(n19019) );
  XNOR U20731 ( .A(n19019), .B(n4071), .Z(n19021) );
  NANDN U20732 ( .A(b[0]), .B(a[403]), .Z(n19020) );
  NAND U20733 ( .A(n19021), .B(n19020), .Z(n19062) );
  XNOR U20734 ( .A(n19061), .B(n19062), .Z(n19067) );
  XOR U20735 ( .A(n19068), .B(n19067), .Z(n19046) );
  NANDN U20736 ( .A(n19023), .B(n19022), .Z(n19027) );
  NANDN U20737 ( .A(n19025), .B(n19024), .Z(n19026) );
  AND U20738 ( .A(n19027), .B(n19026), .Z(n19045) );
  XNOR U20739 ( .A(n19046), .B(n19045), .Z(n19047) );
  NANDN U20740 ( .A(n19029), .B(n19028), .Z(n19033) );
  NAND U20741 ( .A(n19031), .B(n19030), .Z(n19032) );
  NAND U20742 ( .A(n19033), .B(n19032), .Z(n19048) );
  XNOR U20743 ( .A(n19047), .B(n19048), .Z(n19039) );
  XNOR U20744 ( .A(n19040), .B(n19039), .Z(n19041) );
  XNOR U20745 ( .A(n19042), .B(n19041), .Z(n19071) );
  XNOR U20746 ( .A(sreg[1420]), .B(n19071), .Z(n19073) );
  NANDN U20747 ( .A(sreg[1419]), .B(n19034), .Z(n19038) );
  NAND U20748 ( .A(n19036), .B(n19035), .Z(n19037) );
  NAND U20749 ( .A(n19038), .B(n19037), .Z(n19072) );
  XNOR U20750 ( .A(n19073), .B(n19072), .Z(c[1420]) );
  NANDN U20751 ( .A(n19040), .B(n19039), .Z(n19044) );
  NANDN U20752 ( .A(n19042), .B(n19041), .Z(n19043) );
  AND U20753 ( .A(n19044), .B(n19043), .Z(n19079) );
  NANDN U20754 ( .A(n19046), .B(n19045), .Z(n19050) );
  NANDN U20755 ( .A(n19048), .B(n19047), .Z(n19049) );
  AND U20756 ( .A(n19050), .B(n19049), .Z(n19077) );
  NAND U20757 ( .A(n42143), .B(n19051), .Z(n19053) );
  XNOR U20758 ( .A(a[399]), .B(n4128), .Z(n19088) );
  NAND U20759 ( .A(n42144), .B(n19088), .Z(n19052) );
  AND U20760 ( .A(n19053), .B(n19052), .Z(n19103) );
  XOR U20761 ( .A(a[403]), .B(n42012), .Z(n19091) );
  XNOR U20762 ( .A(n19103), .B(n19102), .Z(n19105) );
  AND U20763 ( .A(a[405]), .B(b[0]), .Z(n19055) );
  XNOR U20764 ( .A(n19055), .B(n4071), .Z(n19057) );
  NANDN U20765 ( .A(b[0]), .B(a[404]), .Z(n19056) );
  NAND U20766 ( .A(n19057), .B(n19056), .Z(n19099) );
  XOR U20767 ( .A(a[401]), .B(n42085), .Z(n19092) );
  AND U20768 ( .A(a[397]), .B(b[7]), .Z(n19096) );
  XNOR U20769 ( .A(n19097), .B(n19096), .Z(n19098) );
  XNOR U20770 ( .A(n19099), .B(n19098), .Z(n19104) );
  XOR U20771 ( .A(n19105), .B(n19104), .Z(n19083) );
  NANDN U20772 ( .A(n19060), .B(n19059), .Z(n19064) );
  NANDN U20773 ( .A(n19062), .B(n19061), .Z(n19063) );
  AND U20774 ( .A(n19064), .B(n19063), .Z(n19082) );
  XNOR U20775 ( .A(n19083), .B(n19082), .Z(n19084) );
  NANDN U20776 ( .A(n19066), .B(n19065), .Z(n19070) );
  NAND U20777 ( .A(n19068), .B(n19067), .Z(n19069) );
  NAND U20778 ( .A(n19070), .B(n19069), .Z(n19085) );
  XNOR U20779 ( .A(n19084), .B(n19085), .Z(n19076) );
  XNOR U20780 ( .A(n19077), .B(n19076), .Z(n19078) );
  XNOR U20781 ( .A(n19079), .B(n19078), .Z(n19108) );
  XNOR U20782 ( .A(sreg[1421]), .B(n19108), .Z(n19110) );
  NANDN U20783 ( .A(sreg[1420]), .B(n19071), .Z(n19075) );
  NAND U20784 ( .A(n19073), .B(n19072), .Z(n19074) );
  NAND U20785 ( .A(n19075), .B(n19074), .Z(n19109) );
  XNOR U20786 ( .A(n19110), .B(n19109), .Z(c[1421]) );
  NANDN U20787 ( .A(n19077), .B(n19076), .Z(n19081) );
  NANDN U20788 ( .A(n19079), .B(n19078), .Z(n19080) );
  AND U20789 ( .A(n19081), .B(n19080), .Z(n19116) );
  NANDN U20790 ( .A(n19083), .B(n19082), .Z(n19087) );
  NANDN U20791 ( .A(n19085), .B(n19084), .Z(n19086) );
  AND U20792 ( .A(n19087), .B(n19086), .Z(n19114) );
  NAND U20793 ( .A(n42143), .B(n19088), .Z(n19090) );
  XNOR U20794 ( .A(a[400]), .B(n4129), .Z(n19125) );
  NAND U20795 ( .A(n42144), .B(n19125), .Z(n19089) );
  AND U20796 ( .A(n19090), .B(n19089), .Z(n19140) );
  XOR U20797 ( .A(a[404]), .B(n42012), .Z(n19128) );
  XNOR U20798 ( .A(n19140), .B(n19139), .Z(n19142) );
  XOR U20799 ( .A(a[402]), .B(n42085), .Z(n19132) );
  AND U20800 ( .A(a[398]), .B(b[7]), .Z(n19133) );
  XNOR U20801 ( .A(n19134), .B(n19133), .Z(n19135) );
  AND U20802 ( .A(a[406]), .B(b[0]), .Z(n19093) );
  XNOR U20803 ( .A(n19093), .B(n4071), .Z(n19095) );
  NANDN U20804 ( .A(b[0]), .B(a[405]), .Z(n19094) );
  NAND U20805 ( .A(n19095), .B(n19094), .Z(n19136) );
  XNOR U20806 ( .A(n19135), .B(n19136), .Z(n19141) );
  XOR U20807 ( .A(n19142), .B(n19141), .Z(n19120) );
  NANDN U20808 ( .A(n19097), .B(n19096), .Z(n19101) );
  NANDN U20809 ( .A(n19099), .B(n19098), .Z(n19100) );
  AND U20810 ( .A(n19101), .B(n19100), .Z(n19119) );
  XNOR U20811 ( .A(n19120), .B(n19119), .Z(n19121) );
  NANDN U20812 ( .A(n19103), .B(n19102), .Z(n19107) );
  NAND U20813 ( .A(n19105), .B(n19104), .Z(n19106) );
  NAND U20814 ( .A(n19107), .B(n19106), .Z(n19122) );
  XNOR U20815 ( .A(n19121), .B(n19122), .Z(n19113) );
  XNOR U20816 ( .A(n19114), .B(n19113), .Z(n19115) );
  XNOR U20817 ( .A(n19116), .B(n19115), .Z(n19145) );
  XNOR U20818 ( .A(sreg[1422]), .B(n19145), .Z(n19147) );
  NANDN U20819 ( .A(sreg[1421]), .B(n19108), .Z(n19112) );
  NAND U20820 ( .A(n19110), .B(n19109), .Z(n19111) );
  NAND U20821 ( .A(n19112), .B(n19111), .Z(n19146) );
  XNOR U20822 ( .A(n19147), .B(n19146), .Z(c[1422]) );
  NANDN U20823 ( .A(n19114), .B(n19113), .Z(n19118) );
  NANDN U20824 ( .A(n19116), .B(n19115), .Z(n19117) );
  AND U20825 ( .A(n19118), .B(n19117), .Z(n19153) );
  NANDN U20826 ( .A(n19120), .B(n19119), .Z(n19124) );
  NANDN U20827 ( .A(n19122), .B(n19121), .Z(n19123) );
  AND U20828 ( .A(n19124), .B(n19123), .Z(n19151) );
  NAND U20829 ( .A(n42143), .B(n19125), .Z(n19127) );
  XNOR U20830 ( .A(a[401]), .B(n4129), .Z(n19162) );
  NAND U20831 ( .A(n42144), .B(n19162), .Z(n19126) );
  AND U20832 ( .A(n19127), .B(n19126), .Z(n19177) );
  XOR U20833 ( .A(a[405]), .B(n42012), .Z(n19165) );
  XNOR U20834 ( .A(n19177), .B(n19176), .Z(n19179) );
  AND U20835 ( .A(a[407]), .B(b[0]), .Z(n19129) );
  XNOR U20836 ( .A(n19129), .B(n4071), .Z(n19131) );
  NANDN U20837 ( .A(b[0]), .B(a[406]), .Z(n19130) );
  NAND U20838 ( .A(n19131), .B(n19130), .Z(n19173) );
  XOR U20839 ( .A(a[403]), .B(n42085), .Z(n19166) );
  AND U20840 ( .A(a[399]), .B(b[7]), .Z(n19170) );
  XNOR U20841 ( .A(n19171), .B(n19170), .Z(n19172) );
  XNOR U20842 ( .A(n19173), .B(n19172), .Z(n19178) );
  XOR U20843 ( .A(n19179), .B(n19178), .Z(n19157) );
  NANDN U20844 ( .A(n19134), .B(n19133), .Z(n19138) );
  NANDN U20845 ( .A(n19136), .B(n19135), .Z(n19137) );
  AND U20846 ( .A(n19138), .B(n19137), .Z(n19156) );
  XNOR U20847 ( .A(n19157), .B(n19156), .Z(n19158) );
  NANDN U20848 ( .A(n19140), .B(n19139), .Z(n19144) );
  NAND U20849 ( .A(n19142), .B(n19141), .Z(n19143) );
  NAND U20850 ( .A(n19144), .B(n19143), .Z(n19159) );
  XNOR U20851 ( .A(n19158), .B(n19159), .Z(n19150) );
  XNOR U20852 ( .A(n19151), .B(n19150), .Z(n19152) );
  XNOR U20853 ( .A(n19153), .B(n19152), .Z(n19182) );
  XNOR U20854 ( .A(sreg[1423]), .B(n19182), .Z(n19184) );
  NANDN U20855 ( .A(sreg[1422]), .B(n19145), .Z(n19149) );
  NAND U20856 ( .A(n19147), .B(n19146), .Z(n19148) );
  NAND U20857 ( .A(n19149), .B(n19148), .Z(n19183) );
  XNOR U20858 ( .A(n19184), .B(n19183), .Z(c[1423]) );
  NANDN U20859 ( .A(n19151), .B(n19150), .Z(n19155) );
  NANDN U20860 ( .A(n19153), .B(n19152), .Z(n19154) );
  AND U20861 ( .A(n19155), .B(n19154), .Z(n19190) );
  NANDN U20862 ( .A(n19157), .B(n19156), .Z(n19161) );
  NANDN U20863 ( .A(n19159), .B(n19158), .Z(n19160) );
  AND U20864 ( .A(n19161), .B(n19160), .Z(n19188) );
  NAND U20865 ( .A(n42143), .B(n19162), .Z(n19164) );
  XNOR U20866 ( .A(a[402]), .B(n4129), .Z(n19199) );
  NAND U20867 ( .A(n42144), .B(n19199), .Z(n19163) );
  AND U20868 ( .A(n19164), .B(n19163), .Z(n19214) );
  XOR U20869 ( .A(a[406]), .B(n42012), .Z(n19202) );
  XNOR U20870 ( .A(n19214), .B(n19213), .Z(n19216) );
  XOR U20871 ( .A(a[404]), .B(n42085), .Z(n19206) );
  AND U20872 ( .A(a[400]), .B(b[7]), .Z(n19207) );
  XNOR U20873 ( .A(n19208), .B(n19207), .Z(n19209) );
  AND U20874 ( .A(a[408]), .B(b[0]), .Z(n19167) );
  XNOR U20875 ( .A(n19167), .B(n4071), .Z(n19169) );
  NANDN U20876 ( .A(b[0]), .B(a[407]), .Z(n19168) );
  NAND U20877 ( .A(n19169), .B(n19168), .Z(n19210) );
  XNOR U20878 ( .A(n19209), .B(n19210), .Z(n19215) );
  XOR U20879 ( .A(n19216), .B(n19215), .Z(n19194) );
  NANDN U20880 ( .A(n19171), .B(n19170), .Z(n19175) );
  NANDN U20881 ( .A(n19173), .B(n19172), .Z(n19174) );
  AND U20882 ( .A(n19175), .B(n19174), .Z(n19193) );
  XNOR U20883 ( .A(n19194), .B(n19193), .Z(n19195) );
  NANDN U20884 ( .A(n19177), .B(n19176), .Z(n19181) );
  NAND U20885 ( .A(n19179), .B(n19178), .Z(n19180) );
  NAND U20886 ( .A(n19181), .B(n19180), .Z(n19196) );
  XNOR U20887 ( .A(n19195), .B(n19196), .Z(n19187) );
  XNOR U20888 ( .A(n19188), .B(n19187), .Z(n19189) );
  XNOR U20889 ( .A(n19190), .B(n19189), .Z(n19219) );
  XNOR U20890 ( .A(sreg[1424]), .B(n19219), .Z(n19221) );
  NANDN U20891 ( .A(sreg[1423]), .B(n19182), .Z(n19186) );
  NAND U20892 ( .A(n19184), .B(n19183), .Z(n19185) );
  NAND U20893 ( .A(n19186), .B(n19185), .Z(n19220) );
  XNOR U20894 ( .A(n19221), .B(n19220), .Z(c[1424]) );
  NANDN U20895 ( .A(n19188), .B(n19187), .Z(n19192) );
  NANDN U20896 ( .A(n19190), .B(n19189), .Z(n19191) );
  AND U20897 ( .A(n19192), .B(n19191), .Z(n19227) );
  NANDN U20898 ( .A(n19194), .B(n19193), .Z(n19198) );
  NANDN U20899 ( .A(n19196), .B(n19195), .Z(n19197) );
  AND U20900 ( .A(n19198), .B(n19197), .Z(n19225) );
  NAND U20901 ( .A(n42143), .B(n19199), .Z(n19201) );
  XNOR U20902 ( .A(a[403]), .B(n4129), .Z(n19236) );
  NAND U20903 ( .A(n42144), .B(n19236), .Z(n19200) );
  AND U20904 ( .A(n19201), .B(n19200), .Z(n19251) );
  XOR U20905 ( .A(a[407]), .B(n42012), .Z(n19239) );
  XNOR U20906 ( .A(n19251), .B(n19250), .Z(n19253) );
  AND U20907 ( .A(a[409]), .B(b[0]), .Z(n19203) );
  XNOR U20908 ( .A(n19203), .B(n4071), .Z(n19205) );
  NANDN U20909 ( .A(b[0]), .B(a[408]), .Z(n19204) );
  NAND U20910 ( .A(n19205), .B(n19204), .Z(n19247) );
  XOR U20911 ( .A(a[405]), .B(n42085), .Z(n19243) );
  AND U20912 ( .A(a[401]), .B(b[7]), .Z(n19244) );
  XNOR U20913 ( .A(n19245), .B(n19244), .Z(n19246) );
  XNOR U20914 ( .A(n19247), .B(n19246), .Z(n19252) );
  XOR U20915 ( .A(n19253), .B(n19252), .Z(n19231) );
  NANDN U20916 ( .A(n19208), .B(n19207), .Z(n19212) );
  NANDN U20917 ( .A(n19210), .B(n19209), .Z(n19211) );
  AND U20918 ( .A(n19212), .B(n19211), .Z(n19230) );
  XNOR U20919 ( .A(n19231), .B(n19230), .Z(n19232) );
  NANDN U20920 ( .A(n19214), .B(n19213), .Z(n19218) );
  NAND U20921 ( .A(n19216), .B(n19215), .Z(n19217) );
  NAND U20922 ( .A(n19218), .B(n19217), .Z(n19233) );
  XNOR U20923 ( .A(n19232), .B(n19233), .Z(n19224) );
  XNOR U20924 ( .A(n19225), .B(n19224), .Z(n19226) );
  XNOR U20925 ( .A(n19227), .B(n19226), .Z(n19256) );
  XNOR U20926 ( .A(sreg[1425]), .B(n19256), .Z(n19258) );
  NANDN U20927 ( .A(sreg[1424]), .B(n19219), .Z(n19223) );
  NAND U20928 ( .A(n19221), .B(n19220), .Z(n19222) );
  NAND U20929 ( .A(n19223), .B(n19222), .Z(n19257) );
  XNOR U20930 ( .A(n19258), .B(n19257), .Z(c[1425]) );
  NANDN U20931 ( .A(n19225), .B(n19224), .Z(n19229) );
  NANDN U20932 ( .A(n19227), .B(n19226), .Z(n19228) );
  AND U20933 ( .A(n19229), .B(n19228), .Z(n19264) );
  NANDN U20934 ( .A(n19231), .B(n19230), .Z(n19235) );
  NANDN U20935 ( .A(n19233), .B(n19232), .Z(n19234) );
  AND U20936 ( .A(n19235), .B(n19234), .Z(n19262) );
  NAND U20937 ( .A(n42143), .B(n19236), .Z(n19238) );
  XNOR U20938 ( .A(a[404]), .B(n4129), .Z(n19273) );
  NAND U20939 ( .A(n42144), .B(n19273), .Z(n19237) );
  AND U20940 ( .A(n19238), .B(n19237), .Z(n19288) );
  XOR U20941 ( .A(a[408]), .B(n42012), .Z(n19276) );
  XNOR U20942 ( .A(n19288), .B(n19287), .Z(n19290) );
  AND U20943 ( .A(a[410]), .B(b[0]), .Z(n19240) );
  XNOR U20944 ( .A(n19240), .B(n4071), .Z(n19242) );
  NANDN U20945 ( .A(b[0]), .B(a[409]), .Z(n19241) );
  NAND U20946 ( .A(n19242), .B(n19241), .Z(n19284) );
  XOR U20947 ( .A(a[406]), .B(n42085), .Z(n19280) );
  AND U20948 ( .A(a[402]), .B(b[7]), .Z(n19281) );
  XNOR U20949 ( .A(n19282), .B(n19281), .Z(n19283) );
  XNOR U20950 ( .A(n19284), .B(n19283), .Z(n19289) );
  XOR U20951 ( .A(n19290), .B(n19289), .Z(n19268) );
  NANDN U20952 ( .A(n19245), .B(n19244), .Z(n19249) );
  NANDN U20953 ( .A(n19247), .B(n19246), .Z(n19248) );
  AND U20954 ( .A(n19249), .B(n19248), .Z(n19267) );
  XNOR U20955 ( .A(n19268), .B(n19267), .Z(n19269) );
  NANDN U20956 ( .A(n19251), .B(n19250), .Z(n19255) );
  NAND U20957 ( .A(n19253), .B(n19252), .Z(n19254) );
  NAND U20958 ( .A(n19255), .B(n19254), .Z(n19270) );
  XNOR U20959 ( .A(n19269), .B(n19270), .Z(n19261) );
  XNOR U20960 ( .A(n19262), .B(n19261), .Z(n19263) );
  XNOR U20961 ( .A(n19264), .B(n19263), .Z(n19293) );
  XNOR U20962 ( .A(sreg[1426]), .B(n19293), .Z(n19295) );
  NANDN U20963 ( .A(sreg[1425]), .B(n19256), .Z(n19260) );
  NAND U20964 ( .A(n19258), .B(n19257), .Z(n19259) );
  NAND U20965 ( .A(n19260), .B(n19259), .Z(n19294) );
  XNOR U20966 ( .A(n19295), .B(n19294), .Z(c[1426]) );
  NANDN U20967 ( .A(n19262), .B(n19261), .Z(n19266) );
  NANDN U20968 ( .A(n19264), .B(n19263), .Z(n19265) );
  AND U20969 ( .A(n19266), .B(n19265), .Z(n19301) );
  NANDN U20970 ( .A(n19268), .B(n19267), .Z(n19272) );
  NANDN U20971 ( .A(n19270), .B(n19269), .Z(n19271) );
  AND U20972 ( .A(n19272), .B(n19271), .Z(n19299) );
  NAND U20973 ( .A(n42143), .B(n19273), .Z(n19275) );
  XNOR U20974 ( .A(a[405]), .B(n4129), .Z(n19310) );
  NAND U20975 ( .A(n42144), .B(n19310), .Z(n19274) );
  AND U20976 ( .A(n19275), .B(n19274), .Z(n19325) );
  XOR U20977 ( .A(a[409]), .B(n42012), .Z(n19313) );
  XNOR U20978 ( .A(n19325), .B(n19324), .Z(n19327) );
  AND U20979 ( .A(a[411]), .B(b[0]), .Z(n19277) );
  XNOR U20980 ( .A(n19277), .B(n4071), .Z(n19279) );
  NANDN U20981 ( .A(b[0]), .B(a[410]), .Z(n19278) );
  NAND U20982 ( .A(n19279), .B(n19278), .Z(n19321) );
  XOR U20983 ( .A(a[407]), .B(n42085), .Z(n19317) );
  AND U20984 ( .A(a[403]), .B(b[7]), .Z(n19318) );
  XNOR U20985 ( .A(n19319), .B(n19318), .Z(n19320) );
  XNOR U20986 ( .A(n19321), .B(n19320), .Z(n19326) );
  XOR U20987 ( .A(n19327), .B(n19326), .Z(n19305) );
  NANDN U20988 ( .A(n19282), .B(n19281), .Z(n19286) );
  NANDN U20989 ( .A(n19284), .B(n19283), .Z(n19285) );
  AND U20990 ( .A(n19286), .B(n19285), .Z(n19304) );
  XNOR U20991 ( .A(n19305), .B(n19304), .Z(n19306) );
  NANDN U20992 ( .A(n19288), .B(n19287), .Z(n19292) );
  NAND U20993 ( .A(n19290), .B(n19289), .Z(n19291) );
  NAND U20994 ( .A(n19292), .B(n19291), .Z(n19307) );
  XNOR U20995 ( .A(n19306), .B(n19307), .Z(n19298) );
  XNOR U20996 ( .A(n19299), .B(n19298), .Z(n19300) );
  XNOR U20997 ( .A(n19301), .B(n19300), .Z(n19330) );
  XNOR U20998 ( .A(sreg[1427]), .B(n19330), .Z(n19332) );
  NANDN U20999 ( .A(sreg[1426]), .B(n19293), .Z(n19297) );
  NAND U21000 ( .A(n19295), .B(n19294), .Z(n19296) );
  NAND U21001 ( .A(n19297), .B(n19296), .Z(n19331) );
  XNOR U21002 ( .A(n19332), .B(n19331), .Z(c[1427]) );
  NANDN U21003 ( .A(n19299), .B(n19298), .Z(n19303) );
  NANDN U21004 ( .A(n19301), .B(n19300), .Z(n19302) );
  AND U21005 ( .A(n19303), .B(n19302), .Z(n19338) );
  NANDN U21006 ( .A(n19305), .B(n19304), .Z(n19309) );
  NANDN U21007 ( .A(n19307), .B(n19306), .Z(n19308) );
  AND U21008 ( .A(n19309), .B(n19308), .Z(n19336) );
  NAND U21009 ( .A(n42143), .B(n19310), .Z(n19312) );
  XNOR U21010 ( .A(a[406]), .B(n4129), .Z(n19347) );
  NAND U21011 ( .A(n42144), .B(n19347), .Z(n19311) );
  AND U21012 ( .A(n19312), .B(n19311), .Z(n19362) );
  XOR U21013 ( .A(a[410]), .B(n42012), .Z(n19350) );
  XNOR U21014 ( .A(n19362), .B(n19361), .Z(n19364) );
  AND U21015 ( .A(a[412]), .B(b[0]), .Z(n19314) );
  XNOR U21016 ( .A(n19314), .B(n4071), .Z(n19316) );
  NANDN U21017 ( .A(b[0]), .B(a[411]), .Z(n19315) );
  NAND U21018 ( .A(n19316), .B(n19315), .Z(n19358) );
  XOR U21019 ( .A(a[408]), .B(n42085), .Z(n19354) );
  AND U21020 ( .A(a[404]), .B(b[7]), .Z(n19355) );
  XNOR U21021 ( .A(n19356), .B(n19355), .Z(n19357) );
  XNOR U21022 ( .A(n19358), .B(n19357), .Z(n19363) );
  XOR U21023 ( .A(n19364), .B(n19363), .Z(n19342) );
  NANDN U21024 ( .A(n19319), .B(n19318), .Z(n19323) );
  NANDN U21025 ( .A(n19321), .B(n19320), .Z(n19322) );
  AND U21026 ( .A(n19323), .B(n19322), .Z(n19341) );
  XNOR U21027 ( .A(n19342), .B(n19341), .Z(n19343) );
  NANDN U21028 ( .A(n19325), .B(n19324), .Z(n19329) );
  NAND U21029 ( .A(n19327), .B(n19326), .Z(n19328) );
  NAND U21030 ( .A(n19329), .B(n19328), .Z(n19344) );
  XNOR U21031 ( .A(n19343), .B(n19344), .Z(n19335) );
  XNOR U21032 ( .A(n19336), .B(n19335), .Z(n19337) );
  XNOR U21033 ( .A(n19338), .B(n19337), .Z(n19367) );
  XNOR U21034 ( .A(sreg[1428]), .B(n19367), .Z(n19369) );
  NANDN U21035 ( .A(sreg[1427]), .B(n19330), .Z(n19334) );
  NAND U21036 ( .A(n19332), .B(n19331), .Z(n19333) );
  NAND U21037 ( .A(n19334), .B(n19333), .Z(n19368) );
  XNOR U21038 ( .A(n19369), .B(n19368), .Z(c[1428]) );
  NANDN U21039 ( .A(n19336), .B(n19335), .Z(n19340) );
  NANDN U21040 ( .A(n19338), .B(n19337), .Z(n19339) );
  AND U21041 ( .A(n19340), .B(n19339), .Z(n19375) );
  NANDN U21042 ( .A(n19342), .B(n19341), .Z(n19346) );
  NANDN U21043 ( .A(n19344), .B(n19343), .Z(n19345) );
  AND U21044 ( .A(n19346), .B(n19345), .Z(n19373) );
  NAND U21045 ( .A(n42143), .B(n19347), .Z(n19349) );
  XNOR U21046 ( .A(a[407]), .B(n4130), .Z(n19384) );
  NAND U21047 ( .A(n42144), .B(n19384), .Z(n19348) );
  AND U21048 ( .A(n19349), .B(n19348), .Z(n19399) );
  XOR U21049 ( .A(a[411]), .B(n42012), .Z(n19387) );
  XNOR U21050 ( .A(n19399), .B(n19398), .Z(n19401) );
  AND U21051 ( .A(a[413]), .B(b[0]), .Z(n19351) );
  XNOR U21052 ( .A(n19351), .B(n4071), .Z(n19353) );
  NANDN U21053 ( .A(b[0]), .B(a[412]), .Z(n19352) );
  NAND U21054 ( .A(n19353), .B(n19352), .Z(n19395) );
  XOR U21055 ( .A(a[409]), .B(n42085), .Z(n19391) );
  AND U21056 ( .A(a[405]), .B(b[7]), .Z(n19392) );
  XNOR U21057 ( .A(n19393), .B(n19392), .Z(n19394) );
  XNOR U21058 ( .A(n19395), .B(n19394), .Z(n19400) );
  XOR U21059 ( .A(n19401), .B(n19400), .Z(n19379) );
  NANDN U21060 ( .A(n19356), .B(n19355), .Z(n19360) );
  NANDN U21061 ( .A(n19358), .B(n19357), .Z(n19359) );
  AND U21062 ( .A(n19360), .B(n19359), .Z(n19378) );
  XNOR U21063 ( .A(n19379), .B(n19378), .Z(n19380) );
  NANDN U21064 ( .A(n19362), .B(n19361), .Z(n19366) );
  NAND U21065 ( .A(n19364), .B(n19363), .Z(n19365) );
  NAND U21066 ( .A(n19366), .B(n19365), .Z(n19381) );
  XNOR U21067 ( .A(n19380), .B(n19381), .Z(n19372) );
  XNOR U21068 ( .A(n19373), .B(n19372), .Z(n19374) );
  XNOR U21069 ( .A(n19375), .B(n19374), .Z(n19404) );
  XNOR U21070 ( .A(sreg[1429]), .B(n19404), .Z(n19406) );
  NANDN U21071 ( .A(sreg[1428]), .B(n19367), .Z(n19371) );
  NAND U21072 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U21073 ( .A(n19371), .B(n19370), .Z(n19405) );
  XNOR U21074 ( .A(n19406), .B(n19405), .Z(c[1429]) );
  NANDN U21075 ( .A(n19373), .B(n19372), .Z(n19377) );
  NANDN U21076 ( .A(n19375), .B(n19374), .Z(n19376) );
  AND U21077 ( .A(n19377), .B(n19376), .Z(n19412) );
  NANDN U21078 ( .A(n19379), .B(n19378), .Z(n19383) );
  NANDN U21079 ( .A(n19381), .B(n19380), .Z(n19382) );
  AND U21080 ( .A(n19383), .B(n19382), .Z(n19410) );
  NAND U21081 ( .A(n42143), .B(n19384), .Z(n19386) );
  XNOR U21082 ( .A(a[408]), .B(n4130), .Z(n19421) );
  NAND U21083 ( .A(n42144), .B(n19421), .Z(n19385) );
  AND U21084 ( .A(n19386), .B(n19385), .Z(n19436) );
  XOR U21085 ( .A(a[412]), .B(n42012), .Z(n19424) );
  XNOR U21086 ( .A(n19436), .B(n19435), .Z(n19438) );
  AND U21087 ( .A(a[414]), .B(b[0]), .Z(n19388) );
  XNOR U21088 ( .A(n19388), .B(n4071), .Z(n19390) );
  NANDN U21089 ( .A(b[0]), .B(a[413]), .Z(n19389) );
  NAND U21090 ( .A(n19390), .B(n19389), .Z(n19432) );
  XOR U21091 ( .A(a[410]), .B(n42085), .Z(n19425) );
  AND U21092 ( .A(a[406]), .B(b[7]), .Z(n19429) );
  XNOR U21093 ( .A(n19430), .B(n19429), .Z(n19431) );
  XNOR U21094 ( .A(n19432), .B(n19431), .Z(n19437) );
  XOR U21095 ( .A(n19438), .B(n19437), .Z(n19416) );
  NANDN U21096 ( .A(n19393), .B(n19392), .Z(n19397) );
  NANDN U21097 ( .A(n19395), .B(n19394), .Z(n19396) );
  AND U21098 ( .A(n19397), .B(n19396), .Z(n19415) );
  XNOR U21099 ( .A(n19416), .B(n19415), .Z(n19417) );
  NANDN U21100 ( .A(n19399), .B(n19398), .Z(n19403) );
  NAND U21101 ( .A(n19401), .B(n19400), .Z(n19402) );
  NAND U21102 ( .A(n19403), .B(n19402), .Z(n19418) );
  XNOR U21103 ( .A(n19417), .B(n19418), .Z(n19409) );
  XNOR U21104 ( .A(n19410), .B(n19409), .Z(n19411) );
  XNOR U21105 ( .A(n19412), .B(n19411), .Z(n19441) );
  XNOR U21106 ( .A(sreg[1430]), .B(n19441), .Z(n19443) );
  NANDN U21107 ( .A(sreg[1429]), .B(n19404), .Z(n19408) );
  NAND U21108 ( .A(n19406), .B(n19405), .Z(n19407) );
  NAND U21109 ( .A(n19408), .B(n19407), .Z(n19442) );
  XNOR U21110 ( .A(n19443), .B(n19442), .Z(c[1430]) );
  NANDN U21111 ( .A(n19410), .B(n19409), .Z(n19414) );
  NANDN U21112 ( .A(n19412), .B(n19411), .Z(n19413) );
  AND U21113 ( .A(n19414), .B(n19413), .Z(n19449) );
  NANDN U21114 ( .A(n19416), .B(n19415), .Z(n19420) );
  NANDN U21115 ( .A(n19418), .B(n19417), .Z(n19419) );
  AND U21116 ( .A(n19420), .B(n19419), .Z(n19447) );
  NAND U21117 ( .A(n42143), .B(n19421), .Z(n19423) );
  XNOR U21118 ( .A(a[409]), .B(n4130), .Z(n19458) );
  NAND U21119 ( .A(n42144), .B(n19458), .Z(n19422) );
  AND U21120 ( .A(n19423), .B(n19422), .Z(n19473) );
  XOR U21121 ( .A(a[413]), .B(n42012), .Z(n19461) );
  XNOR U21122 ( .A(n19473), .B(n19472), .Z(n19475) );
  XOR U21123 ( .A(a[411]), .B(n42085), .Z(n19465) );
  AND U21124 ( .A(a[407]), .B(b[7]), .Z(n19466) );
  XNOR U21125 ( .A(n19467), .B(n19466), .Z(n19468) );
  AND U21126 ( .A(a[415]), .B(b[0]), .Z(n19426) );
  XNOR U21127 ( .A(n19426), .B(n4071), .Z(n19428) );
  NANDN U21128 ( .A(b[0]), .B(a[414]), .Z(n19427) );
  NAND U21129 ( .A(n19428), .B(n19427), .Z(n19469) );
  XNOR U21130 ( .A(n19468), .B(n19469), .Z(n19474) );
  XOR U21131 ( .A(n19475), .B(n19474), .Z(n19453) );
  NANDN U21132 ( .A(n19430), .B(n19429), .Z(n19434) );
  NANDN U21133 ( .A(n19432), .B(n19431), .Z(n19433) );
  AND U21134 ( .A(n19434), .B(n19433), .Z(n19452) );
  XNOR U21135 ( .A(n19453), .B(n19452), .Z(n19454) );
  NANDN U21136 ( .A(n19436), .B(n19435), .Z(n19440) );
  NAND U21137 ( .A(n19438), .B(n19437), .Z(n19439) );
  NAND U21138 ( .A(n19440), .B(n19439), .Z(n19455) );
  XNOR U21139 ( .A(n19454), .B(n19455), .Z(n19446) );
  XNOR U21140 ( .A(n19447), .B(n19446), .Z(n19448) );
  XNOR U21141 ( .A(n19449), .B(n19448), .Z(n19478) );
  XNOR U21142 ( .A(sreg[1431]), .B(n19478), .Z(n19480) );
  NANDN U21143 ( .A(sreg[1430]), .B(n19441), .Z(n19445) );
  NAND U21144 ( .A(n19443), .B(n19442), .Z(n19444) );
  NAND U21145 ( .A(n19445), .B(n19444), .Z(n19479) );
  XNOR U21146 ( .A(n19480), .B(n19479), .Z(c[1431]) );
  NANDN U21147 ( .A(n19447), .B(n19446), .Z(n19451) );
  NANDN U21148 ( .A(n19449), .B(n19448), .Z(n19450) );
  AND U21149 ( .A(n19451), .B(n19450), .Z(n19486) );
  NANDN U21150 ( .A(n19453), .B(n19452), .Z(n19457) );
  NANDN U21151 ( .A(n19455), .B(n19454), .Z(n19456) );
  AND U21152 ( .A(n19457), .B(n19456), .Z(n19484) );
  NAND U21153 ( .A(n42143), .B(n19458), .Z(n19460) );
  XNOR U21154 ( .A(a[410]), .B(n4130), .Z(n19495) );
  NAND U21155 ( .A(n42144), .B(n19495), .Z(n19459) );
  AND U21156 ( .A(n19460), .B(n19459), .Z(n19510) );
  XOR U21157 ( .A(a[414]), .B(n42012), .Z(n19498) );
  XNOR U21158 ( .A(n19510), .B(n19509), .Z(n19512) );
  AND U21159 ( .A(a[416]), .B(b[0]), .Z(n19462) );
  XNOR U21160 ( .A(n19462), .B(n4071), .Z(n19464) );
  NANDN U21161 ( .A(b[0]), .B(a[415]), .Z(n19463) );
  NAND U21162 ( .A(n19464), .B(n19463), .Z(n19506) );
  XOR U21163 ( .A(a[412]), .B(n42085), .Z(n19502) );
  AND U21164 ( .A(a[408]), .B(b[7]), .Z(n19503) );
  XNOR U21165 ( .A(n19504), .B(n19503), .Z(n19505) );
  XNOR U21166 ( .A(n19506), .B(n19505), .Z(n19511) );
  XOR U21167 ( .A(n19512), .B(n19511), .Z(n19490) );
  NANDN U21168 ( .A(n19467), .B(n19466), .Z(n19471) );
  NANDN U21169 ( .A(n19469), .B(n19468), .Z(n19470) );
  AND U21170 ( .A(n19471), .B(n19470), .Z(n19489) );
  XNOR U21171 ( .A(n19490), .B(n19489), .Z(n19491) );
  NANDN U21172 ( .A(n19473), .B(n19472), .Z(n19477) );
  NAND U21173 ( .A(n19475), .B(n19474), .Z(n19476) );
  NAND U21174 ( .A(n19477), .B(n19476), .Z(n19492) );
  XNOR U21175 ( .A(n19491), .B(n19492), .Z(n19483) );
  XNOR U21176 ( .A(n19484), .B(n19483), .Z(n19485) );
  XNOR U21177 ( .A(n19486), .B(n19485), .Z(n19515) );
  XNOR U21178 ( .A(sreg[1432]), .B(n19515), .Z(n19517) );
  NANDN U21179 ( .A(sreg[1431]), .B(n19478), .Z(n19482) );
  NAND U21180 ( .A(n19480), .B(n19479), .Z(n19481) );
  NAND U21181 ( .A(n19482), .B(n19481), .Z(n19516) );
  XNOR U21182 ( .A(n19517), .B(n19516), .Z(c[1432]) );
  NANDN U21183 ( .A(n19484), .B(n19483), .Z(n19488) );
  NANDN U21184 ( .A(n19486), .B(n19485), .Z(n19487) );
  AND U21185 ( .A(n19488), .B(n19487), .Z(n19523) );
  NANDN U21186 ( .A(n19490), .B(n19489), .Z(n19494) );
  NANDN U21187 ( .A(n19492), .B(n19491), .Z(n19493) );
  AND U21188 ( .A(n19494), .B(n19493), .Z(n19521) );
  NAND U21189 ( .A(n42143), .B(n19495), .Z(n19497) );
  XNOR U21190 ( .A(a[411]), .B(n4130), .Z(n19532) );
  NAND U21191 ( .A(n42144), .B(n19532), .Z(n19496) );
  AND U21192 ( .A(n19497), .B(n19496), .Z(n19547) );
  XOR U21193 ( .A(a[415]), .B(n42012), .Z(n19535) );
  XNOR U21194 ( .A(n19547), .B(n19546), .Z(n19549) );
  AND U21195 ( .A(a[417]), .B(b[0]), .Z(n19499) );
  XNOR U21196 ( .A(n19499), .B(n4071), .Z(n19501) );
  NANDN U21197 ( .A(b[0]), .B(a[416]), .Z(n19500) );
  NAND U21198 ( .A(n19501), .B(n19500), .Z(n19543) );
  XOR U21199 ( .A(a[413]), .B(n42085), .Z(n19539) );
  AND U21200 ( .A(a[409]), .B(b[7]), .Z(n19540) );
  XNOR U21201 ( .A(n19541), .B(n19540), .Z(n19542) );
  XNOR U21202 ( .A(n19543), .B(n19542), .Z(n19548) );
  XOR U21203 ( .A(n19549), .B(n19548), .Z(n19527) );
  NANDN U21204 ( .A(n19504), .B(n19503), .Z(n19508) );
  NANDN U21205 ( .A(n19506), .B(n19505), .Z(n19507) );
  AND U21206 ( .A(n19508), .B(n19507), .Z(n19526) );
  XNOR U21207 ( .A(n19527), .B(n19526), .Z(n19528) );
  NANDN U21208 ( .A(n19510), .B(n19509), .Z(n19514) );
  NAND U21209 ( .A(n19512), .B(n19511), .Z(n19513) );
  NAND U21210 ( .A(n19514), .B(n19513), .Z(n19529) );
  XNOR U21211 ( .A(n19528), .B(n19529), .Z(n19520) );
  XNOR U21212 ( .A(n19521), .B(n19520), .Z(n19522) );
  XNOR U21213 ( .A(n19523), .B(n19522), .Z(n19552) );
  XNOR U21214 ( .A(sreg[1433]), .B(n19552), .Z(n19554) );
  NANDN U21215 ( .A(sreg[1432]), .B(n19515), .Z(n19519) );
  NAND U21216 ( .A(n19517), .B(n19516), .Z(n19518) );
  NAND U21217 ( .A(n19519), .B(n19518), .Z(n19553) );
  XNOR U21218 ( .A(n19554), .B(n19553), .Z(c[1433]) );
  NANDN U21219 ( .A(n19521), .B(n19520), .Z(n19525) );
  NANDN U21220 ( .A(n19523), .B(n19522), .Z(n19524) );
  AND U21221 ( .A(n19525), .B(n19524), .Z(n19560) );
  NANDN U21222 ( .A(n19527), .B(n19526), .Z(n19531) );
  NANDN U21223 ( .A(n19529), .B(n19528), .Z(n19530) );
  AND U21224 ( .A(n19531), .B(n19530), .Z(n19558) );
  NAND U21225 ( .A(n42143), .B(n19532), .Z(n19534) );
  XNOR U21226 ( .A(a[412]), .B(n4130), .Z(n19569) );
  NAND U21227 ( .A(n42144), .B(n19569), .Z(n19533) );
  AND U21228 ( .A(n19534), .B(n19533), .Z(n19584) );
  XOR U21229 ( .A(a[416]), .B(n42012), .Z(n19572) );
  XNOR U21230 ( .A(n19584), .B(n19583), .Z(n19586) );
  AND U21231 ( .A(a[418]), .B(b[0]), .Z(n19536) );
  XNOR U21232 ( .A(n19536), .B(n4071), .Z(n19538) );
  NANDN U21233 ( .A(b[0]), .B(a[417]), .Z(n19537) );
  NAND U21234 ( .A(n19538), .B(n19537), .Z(n19580) );
  XOR U21235 ( .A(a[414]), .B(n42085), .Z(n19576) );
  AND U21236 ( .A(a[410]), .B(b[7]), .Z(n19577) );
  XNOR U21237 ( .A(n19578), .B(n19577), .Z(n19579) );
  XNOR U21238 ( .A(n19580), .B(n19579), .Z(n19585) );
  XOR U21239 ( .A(n19586), .B(n19585), .Z(n19564) );
  NANDN U21240 ( .A(n19541), .B(n19540), .Z(n19545) );
  NANDN U21241 ( .A(n19543), .B(n19542), .Z(n19544) );
  AND U21242 ( .A(n19545), .B(n19544), .Z(n19563) );
  XNOR U21243 ( .A(n19564), .B(n19563), .Z(n19565) );
  NANDN U21244 ( .A(n19547), .B(n19546), .Z(n19551) );
  NAND U21245 ( .A(n19549), .B(n19548), .Z(n19550) );
  NAND U21246 ( .A(n19551), .B(n19550), .Z(n19566) );
  XNOR U21247 ( .A(n19565), .B(n19566), .Z(n19557) );
  XNOR U21248 ( .A(n19558), .B(n19557), .Z(n19559) );
  XNOR U21249 ( .A(n19560), .B(n19559), .Z(n19589) );
  XNOR U21250 ( .A(sreg[1434]), .B(n19589), .Z(n19591) );
  NANDN U21251 ( .A(sreg[1433]), .B(n19552), .Z(n19556) );
  NAND U21252 ( .A(n19554), .B(n19553), .Z(n19555) );
  NAND U21253 ( .A(n19556), .B(n19555), .Z(n19590) );
  XNOR U21254 ( .A(n19591), .B(n19590), .Z(c[1434]) );
  NANDN U21255 ( .A(n19558), .B(n19557), .Z(n19562) );
  NANDN U21256 ( .A(n19560), .B(n19559), .Z(n19561) );
  AND U21257 ( .A(n19562), .B(n19561), .Z(n19597) );
  NANDN U21258 ( .A(n19564), .B(n19563), .Z(n19568) );
  NANDN U21259 ( .A(n19566), .B(n19565), .Z(n19567) );
  AND U21260 ( .A(n19568), .B(n19567), .Z(n19595) );
  NAND U21261 ( .A(n42143), .B(n19569), .Z(n19571) );
  XNOR U21262 ( .A(a[413]), .B(n4130), .Z(n19606) );
  NAND U21263 ( .A(n42144), .B(n19606), .Z(n19570) );
  AND U21264 ( .A(n19571), .B(n19570), .Z(n19621) );
  XOR U21265 ( .A(a[417]), .B(n42012), .Z(n19609) );
  XNOR U21266 ( .A(n19621), .B(n19620), .Z(n19623) );
  AND U21267 ( .A(a[419]), .B(b[0]), .Z(n19573) );
  XNOR U21268 ( .A(n19573), .B(n4071), .Z(n19575) );
  NANDN U21269 ( .A(b[0]), .B(a[418]), .Z(n19574) );
  NAND U21270 ( .A(n19575), .B(n19574), .Z(n19617) );
  XOR U21271 ( .A(a[415]), .B(n42085), .Z(n19613) );
  AND U21272 ( .A(a[411]), .B(b[7]), .Z(n19614) );
  XNOR U21273 ( .A(n19615), .B(n19614), .Z(n19616) );
  XNOR U21274 ( .A(n19617), .B(n19616), .Z(n19622) );
  XOR U21275 ( .A(n19623), .B(n19622), .Z(n19601) );
  NANDN U21276 ( .A(n19578), .B(n19577), .Z(n19582) );
  NANDN U21277 ( .A(n19580), .B(n19579), .Z(n19581) );
  AND U21278 ( .A(n19582), .B(n19581), .Z(n19600) );
  XNOR U21279 ( .A(n19601), .B(n19600), .Z(n19602) );
  NANDN U21280 ( .A(n19584), .B(n19583), .Z(n19588) );
  NAND U21281 ( .A(n19586), .B(n19585), .Z(n19587) );
  NAND U21282 ( .A(n19588), .B(n19587), .Z(n19603) );
  XNOR U21283 ( .A(n19602), .B(n19603), .Z(n19594) );
  XNOR U21284 ( .A(n19595), .B(n19594), .Z(n19596) );
  XNOR U21285 ( .A(n19597), .B(n19596), .Z(n19626) );
  XNOR U21286 ( .A(sreg[1435]), .B(n19626), .Z(n19628) );
  NANDN U21287 ( .A(sreg[1434]), .B(n19589), .Z(n19593) );
  NAND U21288 ( .A(n19591), .B(n19590), .Z(n19592) );
  NAND U21289 ( .A(n19593), .B(n19592), .Z(n19627) );
  XNOR U21290 ( .A(n19628), .B(n19627), .Z(c[1435]) );
  NANDN U21291 ( .A(n19595), .B(n19594), .Z(n19599) );
  NANDN U21292 ( .A(n19597), .B(n19596), .Z(n19598) );
  AND U21293 ( .A(n19599), .B(n19598), .Z(n19634) );
  NANDN U21294 ( .A(n19601), .B(n19600), .Z(n19605) );
  NANDN U21295 ( .A(n19603), .B(n19602), .Z(n19604) );
  AND U21296 ( .A(n19605), .B(n19604), .Z(n19632) );
  NAND U21297 ( .A(n42143), .B(n19606), .Z(n19608) );
  XNOR U21298 ( .A(a[414]), .B(n4131), .Z(n19643) );
  NAND U21299 ( .A(n42144), .B(n19643), .Z(n19607) );
  AND U21300 ( .A(n19608), .B(n19607), .Z(n19658) );
  XOR U21301 ( .A(a[418]), .B(n42012), .Z(n19646) );
  XNOR U21302 ( .A(n19658), .B(n19657), .Z(n19660) );
  AND U21303 ( .A(a[420]), .B(b[0]), .Z(n19610) );
  XNOR U21304 ( .A(n19610), .B(n4071), .Z(n19612) );
  NANDN U21305 ( .A(b[0]), .B(a[419]), .Z(n19611) );
  NAND U21306 ( .A(n19612), .B(n19611), .Z(n19654) );
  XOR U21307 ( .A(a[416]), .B(n42085), .Z(n19650) );
  AND U21308 ( .A(a[412]), .B(b[7]), .Z(n19651) );
  XNOR U21309 ( .A(n19652), .B(n19651), .Z(n19653) );
  XNOR U21310 ( .A(n19654), .B(n19653), .Z(n19659) );
  XOR U21311 ( .A(n19660), .B(n19659), .Z(n19638) );
  NANDN U21312 ( .A(n19615), .B(n19614), .Z(n19619) );
  NANDN U21313 ( .A(n19617), .B(n19616), .Z(n19618) );
  AND U21314 ( .A(n19619), .B(n19618), .Z(n19637) );
  XNOR U21315 ( .A(n19638), .B(n19637), .Z(n19639) );
  NANDN U21316 ( .A(n19621), .B(n19620), .Z(n19625) );
  NAND U21317 ( .A(n19623), .B(n19622), .Z(n19624) );
  NAND U21318 ( .A(n19625), .B(n19624), .Z(n19640) );
  XNOR U21319 ( .A(n19639), .B(n19640), .Z(n19631) );
  XNOR U21320 ( .A(n19632), .B(n19631), .Z(n19633) );
  XNOR U21321 ( .A(n19634), .B(n19633), .Z(n19663) );
  XNOR U21322 ( .A(sreg[1436]), .B(n19663), .Z(n19665) );
  NANDN U21323 ( .A(sreg[1435]), .B(n19626), .Z(n19630) );
  NAND U21324 ( .A(n19628), .B(n19627), .Z(n19629) );
  NAND U21325 ( .A(n19630), .B(n19629), .Z(n19664) );
  XNOR U21326 ( .A(n19665), .B(n19664), .Z(c[1436]) );
  NANDN U21327 ( .A(n19632), .B(n19631), .Z(n19636) );
  NANDN U21328 ( .A(n19634), .B(n19633), .Z(n19635) );
  AND U21329 ( .A(n19636), .B(n19635), .Z(n19671) );
  NANDN U21330 ( .A(n19638), .B(n19637), .Z(n19642) );
  NANDN U21331 ( .A(n19640), .B(n19639), .Z(n19641) );
  AND U21332 ( .A(n19642), .B(n19641), .Z(n19669) );
  NAND U21333 ( .A(n42143), .B(n19643), .Z(n19645) );
  XNOR U21334 ( .A(a[415]), .B(n4131), .Z(n19680) );
  NAND U21335 ( .A(n42144), .B(n19680), .Z(n19644) );
  AND U21336 ( .A(n19645), .B(n19644), .Z(n19695) );
  XOR U21337 ( .A(a[419]), .B(n42012), .Z(n19683) );
  XNOR U21338 ( .A(n19695), .B(n19694), .Z(n19697) );
  AND U21339 ( .A(a[421]), .B(b[0]), .Z(n19647) );
  XNOR U21340 ( .A(n19647), .B(n4071), .Z(n19649) );
  NANDN U21341 ( .A(b[0]), .B(a[420]), .Z(n19648) );
  NAND U21342 ( .A(n19649), .B(n19648), .Z(n19691) );
  XOR U21343 ( .A(a[417]), .B(n42085), .Z(n19687) );
  AND U21344 ( .A(a[413]), .B(b[7]), .Z(n19688) );
  XNOR U21345 ( .A(n19689), .B(n19688), .Z(n19690) );
  XNOR U21346 ( .A(n19691), .B(n19690), .Z(n19696) );
  XOR U21347 ( .A(n19697), .B(n19696), .Z(n19675) );
  NANDN U21348 ( .A(n19652), .B(n19651), .Z(n19656) );
  NANDN U21349 ( .A(n19654), .B(n19653), .Z(n19655) );
  AND U21350 ( .A(n19656), .B(n19655), .Z(n19674) );
  XNOR U21351 ( .A(n19675), .B(n19674), .Z(n19676) );
  NANDN U21352 ( .A(n19658), .B(n19657), .Z(n19662) );
  NAND U21353 ( .A(n19660), .B(n19659), .Z(n19661) );
  NAND U21354 ( .A(n19662), .B(n19661), .Z(n19677) );
  XNOR U21355 ( .A(n19676), .B(n19677), .Z(n19668) );
  XNOR U21356 ( .A(n19669), .B(n19668), .Z(n19670) );
  XNOR U21357 ( .A(n19671), .B(n19670), .Z(n19700) );
  XNOR U21358 ( .A(sreg[1437]), .B(n19700), .Z(n19702) );
  NANDN U21359 ( .A(sreg[1436]), .B(n19663), .Z(n19667) );
  NAND U21360 ( .A(n19665), .B(n19664), .Z(n19666) );
  NAND U21361 ( .A(n19667), .B(n19666), .Z(n19701) );
  XNOR U21362 ( .A(n19702), .B(n19701), .Z(c[1437]) );
  NANDN U21363 ( .A(n19669), .B(n19668), .Z(n19673) );
  NANDN U21364 ( .A(n19671), .B(n19670), .Z(n19672) );
  AND U21365 ( .A(n19673), .B(n19672), .Z(n19708) );
  NANDN U21366 ( .A(n19675), .B(n19674), .Z(n19679) );
  NANDN U21367 ( .A(n19677), .B(n19676), .Z(n19678) );
  AND U21368 ( .A(n19679), .B(n19678), .Z(n19706) );
  NAND U21369 ( .A(n42143), .B(n19680), .Z(n19682) );
  XNOR U21370 ( .A(a[416]), .B(n4131), .Z(n19717) );
  NAND U21371 ( .A(n42144), .B(n19717), .Z(n19681) );
  AND U21372 ( .A(n19682), .B(n19681), .Z(n19732) );
  XOR U21373 ( .A(a[420]), .B(n42012), .Z(n19720) );
  XNOR U21374 ( .A(n19732), .B(n19731), .Z(n19734) );
  AND U21375 ( .A(a[422]), .B(b[0]), .Z(n19684) );
  XNOR U21376 ( .A(n19684), .B(n4071), .Z(n19686) );
  NANDN U21377 ( .A(b[0]), .B(a[421]), .Z(n19685) );
  NAND U21378 ( .A(n19686), .B(n19685), .Z(n19728) );
  XOR U21379 ( .A(a[418]), .B(n42085), .Z(n19721) );
  AND U21380 ( .A(a[414]), .B(b[7]), .Z(n19725) );
  XNOR U21381 ( .A(n19726), .B(n19725), .Z(n19727) );
  XNOR U21382 ( .A(n19728), .B(n19727), .Z(n19733) );
  XOR U21383 ( .A(n19734), .B(n19733), .Z(n19712) );
  NANDN U21384 ( .A(n19689), .B(n19688), .Z(n19693) );
  NANDN U21385 ( .A(n19691), .B(n19690), .Z(n19692) );
  AND U21386 ( .A(n19693), .B(n19692), .Z(n19711) );
  XNOR U21387 ( .A(n19712), .B(n19711), .Z(n19713) );
  NANDN U21388 ( .A(n19695), .B(n19694), .Z(n19699) );
  NAND U21389 ( .A(n19697), .B(n19696), .Z(n19698) );
  NAND U21390 ( .A(n19699), .B(n19698), .Z(n19714) );
  XNOR U21391 ( .A(n19713), .B(n19714), .Z(n19705) );
  XNOR U21392 ( .A(n19706), .B(n19705), .Z(n19707) );
  XNOR U21393 ( .A(n19708), .B(n19707), .Z(n19737) );
  XNOR U21394 ( .A(sreg[1438]), .B(n19737), .Z(n19739) );
  NANDN U21395 ( .A(sreg[1437]), .B(n19700), .Z(n19704) );
  NAND U21396 ( .A(n19702), .B(n19701), .Z(n19703) );
  NAND U21397 ( .A(n19704), .B(n19703), .Z(n19738) );
  XNOR U21398 ( .A(n19739), .B(n19738), .Z(c[1438]) );
  NANDN U21399 ( .A(n19706), .B(n19705), .Z(n19710) );
  NANDN U21400 ( .A(n19708), .B(n19707), .Z(n19709) );
  AND U21401 ( .A(n19710), .B(n19709), .Z(n19745) );
  NANDN U21402 ( .A(n19712), .B(n19711), .Z(n19716) );
  NANDN U21403 ( .A(n19714), .B(n19713), .Z(n19715) );
  AND U21404 ( .A(n19716), .B(n19715), .Z(n19743) );
  NAND U21405 ( .A(n42143), .B(n19717), .Z(n19719) );
  XNOR U21406 ( .A(a[417]), .B(n4131), .Z(n19754) );
  NAND U21407 ( .A(n42144), .B(n19754), .Z(n19718) );
  AND U21408 ( .A(n19719), .B(n19718), .Z(n19769) );
  XOR U21409 ( .A(a[421]), .B(n42012), .Z(n19757) );
  XNOR U21410 ( .A(n19769), .B(n19768), .Z(n19771) );
  XOR U21411 ( .A(a[419]), .B(n42085), .Z(n19761) );
  AND U21412 ( .A(a[415]), .B(b[7]), .Z(n19762) );
  XNOR U21413 ( .A(n19763), .B(n19762), .Z(n19764) );
  AND U21414 ( .A(a[423]), .B(b[0]), .Z(n19722) );
  XNOR U21415 ( .A(n19722), .B(n4071), .Z(n19724) );
  NANDN U21416 ( .A(b[0]), .B(a[422]), .Z(n19723) );
  NAND U21417 ( .A(n19724), .B(n19723), .Z(n19765) );
  XNOR U21418 ( .A(n19764), .B(n19765), .Z(n19770) );
  XOR U21419 ( .A(n19771), .B(n19770), .Z(n19749) );
  NANDN U21420 ( .A(n19726), .B(n19725), .Z(n19730) );
  NANDN U21421 ( .A(n19728), .B(n19727), .Z(n19729) );
  AND U21422 ( .A(n19730), .B(n19729), .Z(n19748) );
  XNOR U21423 ( .A(n19749), .B(n19748), .Z(n19750) );
  NANDN U21424 ( .A(n19732), .B(n19731), .Z(n19736) );
  NAND U21425 ( .A(n19734), .B(n19733), .Z(n19735) );
  NAND U21426 ( .A(n19736), .B(n19735), .Z(n19751) );
  XNOR U21427 ( .A(n19750), .B(n19751), .Z(n19742) );
  XNOR U21428 ( .A(n19743), .B(n19742), .Z(n19744) );
  XNOR U21429 ( .A(n19745), .B(n19744), .Z(n19774) );
  XNOR U21430 ( .A(sreg[1439]), .B(n19774), .Z(n19776) );
  NANDN U21431 ( .A(sreg[1438]), .B(n19737), .Z(n19741) );
  NAND U21432 ( .A(n19739), .B(n19738), .Z(n19740) );
  NAND U21433 ( .A(n19741), .B(n19740), .Z(n19775) );
  XNOR U21434 ( .A(n19776), .B(n19775), .Z(c[1439]) );
  NANDN U21435 ( .A(n19743), .B(n19742), .Z(n19747) );
  NANDN U21436 ( .A(n19745), .B(n19744), .Z(n19746) );
  AND U21437 ( .A(n19747), .B(n19746), .Z(n19782) );
  NANDN U21438 ( .A(n19749), .B(n19748), .Z(n19753) );
  NANDN U21439 ( .A(n19751), .B(n19750), .Z(n19752) );
  AND U21440 ( .A(n19753), .B(n19752), .Z(n19780) );
  NAND U21441 ( .A(n42143), .B(n19754), .Z(n19756) );
  XNOR U21442 ( .A(a[418]), .B(n4131), .Z(n19791) );
  NAND U21443 ( .A(n42144), .B(n19791), .Z(n19755) );
  AND U21444 ( .A(n19756), .B(n19755), .Z(n19806) );
  XOR U21445 ( .A(a[422]), .B(n42012), .Z(n19794) );
  XNOR U21446 ( .A(n19806), .B(n19805), .Z(n19808) );
  AND U21447 ( .A(a[424]), .B(b[0]), .Z(n19758) );
  XNOR U21448 ( .A(n19758), .B(n4071), .Z(n19760) );
  NANDN U21449 ( .A(b[0]), .B(a[423]), .Z(n19759) );
  NAND U21450 ( .A(n19760), .B(n19759), .Z(n19802) );
  XOR U21451 ( .A(a[420]), .B(n42085), .Z(n19798) );
  AND U21452 ( .A(a[416]), .B(b[7]), .Z(n19799) );
  XNOR U21453 ( .A(n19800), .B(n19799), .Z(n19801) );
  XNOR U21454 ( .A(n19802), .B(n19801), .Z(n19807) );
  XOR U21455 ( .A(n19808), .B(n19807), .Z(n19786) );
  NANDN U21456 ( .A(n19763), .B(n19762), .Z(n19767) );
  NANDN U21457 ( .A(n19765), .B(n19764), .Z(n19766) );
  AND U21458 ( .A(n19767), .B(n19766), .Z(n19785) );
  XNOR U21459 ( .A(n19786), .B(n19785), .Z(n19787) );
  NANDN U21460 ( .A(n19769), .B(n19768), .Z(n19773) );
  NAND U21461 ( .A(n19771), .B(n19770), .Z(n19772) );
  NAND U21462 ( .A(n19773), .B(n19772), .Z(n19788) );
  XNOR U21463 ( .A(n19787), .B(n19788), .Z(n19779) );
  XNOR U21464 ( .A(n19780), .B(n19779), .Z(n19781) );
  XNOR U21465 ( .A(n19782), .B(n19781), .Z(n19811) );
  XNOR U21466 ( .A(sreg[1440]), .B(n19811), .Z(n19813) );
  NANDN U21467 ( .A(sreg[1439]), .B(n19774), .Z(n19778) );
  NAND U21468 ( .A(n19776), .B(n19775), .Z(n19777) );
  NAND U21469 ( .A(n19778), .B(n19777), .Z(n19812) );
  XNOR U21470 ( .A(n19813), .B(n19812), .Z(c[1440]) );
  NANDN U21471 ( .A(n19780), .B(n19779), .Z(n19784) );
  NANDN U21472 ( .A(n19782), .B(n19781), .Z(n19783) );
  AND U21473 ( .A(n19784), .B(n19783), .Z(n19819) );
  NANDN U21474 ( .A(n19786), .B(n19785), .Z(n19790) );
  NANDN U21475 ( .A(n19788), .B(n19787), .Z(n19789) );
  AND U21476 ( .A(n19790), .B(n19789), .Z(n19817) );
  NAND U21477 ( .A(n42143), .B(n19791), .Z(n19793) );
  XNOR U21478 ( .A(a[419]), .B(n4131), .Z(n19828) );
  NAND U21479 ( .A(n42144), .B(n19828), .Z(n19792) );
  AND U21480 ( .A(n19793), .B(n19792), .Z(n19843) );
  XOR U21481 ( .A(a[423]), .B(n42012), .Z(n19831) );
  XNOR U21482 ( .A(n19843), .B(n19842), .Z(n19845) );
  AND U21483 ( .A(a[425]), .B(b[0]), .Z(n19795) );
  XNOR U21484 ( .A(n19795), .B(n4071), .Z(n19797) );
  NANDN U21485 ( .A(b[0]), .B(a[424]), .Z(n19796) );
  NAND U21486 ( .A(n19797), .B(n19796), .Z(n19839) );
  XOR U21487 ( .A(a[421]), .B(n42085), .Z(n19832) );
  AND U21488 ( .A(a[417]), .B(b[7]), .Z(n19836) );
  XNOR U21489 ( .A(n19837), .B(n19836), .Z(n19838) );
  XNOR U21490 ( .A(n19839), .B(n19838), .Z(n19844) );
  XOR U21491 ( .A(n19845), .B(n19844), .Z(n19823) );
  NANDN U21492 ( .A(n19800), .B(n19799), .Z(n19804) );
  NANDN U21493 ( .A(n19802), .B(n19801), .Z(n19803) );
  AND U21494 ( .A(n19804), .B(n19803), .Z(n19822) );
  XNOR U21495 ( .A(n19823), .B(n19822), .Z(n19824) );
  NANDN U21496 ( .A(n19806), .B(n19805), .Z(n19810) );
  NAND U21497 ( .A(n19808), .B(n19807), .Z(n19809) );
  NAND U21498 ( .A(n19810), .B(n19809), .Z(n19825) );
  XNOR U21499 ( .A(n19824), .B(n19825), .Z(n19816) );
  XNOR U21500 ( .A(n19817), .B(n19816), .Z(n19818) );
  XNOR U21501 ( .A(n19819), .B(n19818), .Z(n19848) );
  XNOR U21502 ( .A(sreg[1441]), .B(n19848), .Z(n19850) );
  NANDN U21503 ( .A(sreg[1440]), .B(n19811), .Z(n19815) );
  NAND U21504 ( .A(n19813), .B(n19812), .Z(n19814) );
  NAND U21505 ( .A(n19815), .B(n19814), .Z(n19849) );
  XNOR U21506 ( .A(n19850), .B(n19849), .Z(c[1441]) );
  NANDN U21507 ( .A(n19817), .B(n19816), .Z(n19821) );
  NANDN U21508 ( .A(n19819), .B(n19818), .Z(n19820) );
  AND U21509 ( .A(n19821), .B(n19820), .Z(n19856) );
  NANDN U21510 ( .A(n19823), .B(n19822), .Z(n19827) );
  NANDN U21511 ( .A(n19825), .B(n19824), .Z(n19826) );
  AND U21512 ( .A(n19827), .B(n19826), .Z(n19854) );
  NAND U21513 ( .A(n42143), .B(n19828), .Z(n19830) );
  XNOR U21514 ( .A(a[420]), .B(n4131), .Z(n19865) );
  NAND U21515 ( .A(n42144), .B(n19865), .Z(n19829) );
  AND U21516 ( .A(n19830), .B(n19829), .Z(n19880) );
  XOR U21517 ( .A(a[424]), .B(n42012), .Z(n19868) );
  XNOR U21518 ( .A(n19880), .B(n19879), .Z(n19882) );
  XOR U21519 ( .A(a[422]), .B(n42085), .Z(n19872) );
  AND U21520 ( .A(a[418]), .B(b[7]), .Z(n19873) );
  XNOR U21521 ( .A(n19874), .B(n19873), .Z(n19875) );
  AND U21522 ( .A(a[426]), .B(b[0]), .Z(n19833) );
  XNOR U21523 ( .A(n19833), .B(n4071), .Z(n19835) );
  NANDN U21524 ( .A(b[0]), .B(a[425]), .Z(n19834) );
  NAND U21525 ( .A(n19835), .B(n19834), .Z(n19876) );
  XNOR U21526 ( .A(n19875), .B(n19876), .Z(n19881) );
  XOR U21527 ( .A(n19882), .B(n19881), .Z(n19860) );
  NANDN U21528 ( .A(n19837), .B(n19836), .Z(n19841) );
  NANDN U21529 ( .A(n19839), .B(n19838), .Z(n19840) );
  AND U21530 ( .A(n19841), .B(n19840), .Z(n19859) );
  XNOR U21531 ( .A(n19860), .B(n19859), .Z(n19861) );
  NANDN U21532 ( .A(n19843), .B(n19842), .Z(n19847) );
  NAND U21533 ( .A(n19845), .B(n19844), .Z(n19846) );
  NAND U21534 ( .A(n19847), .B(n19846), .Z(n19862) );
  XNOR U21535 ( .A(n19861), .B(n19862), .Z(n19853) );
  XNOR U21536 ( .A(n19854), .B(n19853), .Z(n19855) );
  XNOR U21537 ( .A(n19856), .B(n19855), .Z(n19885) );
  XNOR U21538 ( .A(sreg[1442]), .B(n19885), .Z(n19887) );
  NANDN U21539 ( .A(sreg[1441]), .B(n19848), .Z(n19852) );
  NAND U21540 ( .A(n19850), .B(n19849), .Z(n19851) );
  NAND U21541 ( .A(n19852), .B(n19851), .Z(n19886) );
  XNOR U21542 ( .A(n19887), .B(n19886), .Z(c[1442]) );
  NANDN U21543 ( .A(n19854), .B(n19853), .Z(n19858) );
  NANDN U21544 ( .A(n19856), .B(n19855), .Z(n19857) );
  AND U21545 ( .A(n19858), .B(n19857), .Z(n19893) );
  NANDN U21546 ( .A(n19860), .B(n19859), .Z(n19864) );
  NANDN U21547 ( .A(n19862), .B(n19861), .Z(n19863) );
  AND U21548 ( .A(n19864), .B(n19863), .Z(n19891) );
  NAND U21549 ( .A(n42143), .B(n19865), .Z(n19867) );
  XNOR U21550 ( .A(a[421]), .B(n4132), .Z(n19902) );
  NAND U21551 ( .A(n42144), .B(n19902), .Z(n19866) );
  AND U21552 ( .A(n19867), .B(n19866), .Z(n19917) );
  XOR U21553 ( .A(a[425]), .B(n42012), .Z(n19905) );
  XNOR U21554 ( .A(n19917), .B(n19916), .Z(n19919) );
  AND U21555 ( .A(a[427]), .B(b[0]), .Z(n19869) );
  XNOR U21556 ( .A(n19869), .B(n4071), .Z(n19871) );
  NANDN U21557 ( .A(b[0]), .B(a[426]), .Z(n19870) );
  NAND U21558 ( .A(n19871), .B(n19870), .Z(n19913) );
  XOR U21559 ( .A(a[423]), .B(n42085), .Z(n19909) );
  AND U21560 ( .A(a[419]), .B(b[7]), .Z(n19910) );
  XNOR U21561 ( .A(n19911), .B(n19910), .Z(n19912) );
  XNOR U21562 ( .A(n19913), .B(n19912), .Z(n19918) );
  XOR U21563 ( .A(n19919), .B(n19918), .Z(n19897) );
  NANDN U21564 ( .A(n19874), .B(n19873), .Z(n19878) );
  NANDN U21565 ( .A(n19876), .B(n19875), .Z(n19877) );
  AND U21566 ( .A(n19878), .B(n19877), .Z(n19896) );
  XNOR U21567 ( .A(n19897), .B(n19896), .Z(n19898) );
  NANDN U21568 ( .A(n19880), .B(n19879), .Z(n19884) );
  NAND U21569 ( .A(n19882), .B(n19881), .Z(n19883) );
  NAND U21570 ( .A(n19884), .B(n19883), .Z(n19899) );
  XNOR U21571 ( .A(n19898), .B(n19899), .Z(n19890) );
  XNOR U21572 ( .A(n19891), .B(n19890), .Z(n19892) );
  XNOR U21573 ( .A(n19893), .B(n19892), .Z(n19922) );
  XNOR U21574 ( .A(sreg[1443]), .B(n19922), .Z(n19924) );
  NANDN U21575 ( .A(sreg[1442]), .B(n19885), .Z(n19889) );
  NAND U21576 ( .A(n19887), .B(n19886), .Z(n19888) );
  NAND U21577 ( .A(n19889), .B(n19888), .Z(n19923) );
  XNOR U21578 ( .A(n19924), .B(n19923), .Z(c[1443]) );
  NANDN U21579 ( .A(n19891), .B(n19890), .Z(n19895) );
  NANDN U21580 ( .A(n19893), .B(n19892), .Z(n19894) );
  AND U21581 ( .A(n19895), .B(n19894), .Z(n19930) );
  NANDN U21582 ( .A(n19897), .B(n19896), .Z(n19901) );
  NANDN U21583 ( .A(n19899), .B(n19898), .Z(n19900) );
  AND U21584 ( .A(n19901), .B(n19900), .Z(n19928) );
  NAND U21585 ( .A(n42143), .B(n19902), .Z(n19904) );
  XNOR U21586 ( .A(a[422]), .B(n4132), .Z(n19939) );
  NAND U21587 ( .A(n42144), .B(n19939), .Z(n19903) );
  AND U21588 ( .A(n19904), .B(n19903), .Z(n19954) );
  XOR U21589 ( .A(a[426]), .B(n42012), .Z(n19942) );
  XNOR U21590 ( .A(n19954), .B(n19953), .Z(n19956) );
  AND U21591 ( .A(a[428]), .B(b[0]), .Z(n19906) );
  XNOR U21592 ( .A(n19906), .B(n4071), .Z(n19908) );
  NANDN U21593 ( .A(b[0]), .B(a[427]), .Z(n19907) );
  NAND U21594 ( .A(n19908), .B(n19907), .Z(n19950) );
  XOR U21595 ( .A(a[424]), .B(n42085), .Z(n19946) );
  AND U21596 ( .A(a[420]), .B(b[7]), .Z(n19947) );
  XNOR U21597 ( .A(n19948), .B(n19947), .Z(n19949) );
  XNOR U21598 ( .A(n19950), .B(n19949), .Z(n19955) );
  XOR U21599 ( .A(n19956), .B(n19955), .Z(n19934) );
  NANDN U21600 ( .A(n19911), .B(n19910), .Z(n19915) );
  NANDN U21601 ( .A(n19913), .B(n19912), .Z(n19914) );
  AND U21602 ( .A(n19915), .B(n19914), .Z(n19933) );
  XNOR U21603 ( .A(n19934), .B(n19933), .Z(n19935) );
  NANDN U21604 ( .A(n19917), .B(n19916), .Z(n19921) );
  NAND U21605 ( .A(n19919), .B(n19918), .Z(n19920) );
  NAND U21606 ( .A(n19921), .B(n19920), .Z(n19936) );
  XNOR U21607 ( .A(n19935), .B(n19936), .Z(n19927) );
  XNOR U21608 ( .A(n19928), .B(n19927), .Z(n19929) );
  XNOR U21609 ( .A(n19930), .B(n19929), .Z(n19959) );
  XNOR U21610 ( .A(sreg[1444]), .B(n19959), .Z(n19961) );
  NANDN U21611 ( .A(sreg[1443]), .B(n19922), .Z(n19926) );
  NAND U21612 ( .A(n19924), .B(n19923), .Z(n19925) );
  NAND U21613 ( .A(n19926), .B(n19925), .Z(n19960) );
  XNOR U21614 ( .A(n19961), .B(n19960), .Z(c[1444]) );
  NANDN U21615 ( .A(n19928), .B(n19927), .Z(n19932) );
  NANDN U21616 ( .A(n19930), .B(n19929), .Z(n19931) );
  AND U21617 ( .A(n19932), .B(n19931), .Z(n19967) );
  NANDN U21618 ( .A(n19934), .B(n19933), .Z(n19938) );
  NANDN U21619 ( .A(n19936), .B(n19935), .Z(n19937) );
  AND U21620 ( .A(n19938), .B(n19937), .Z(n19965) );
  NAND U21621 ( .A(n42143), .B(n19939), .Z(n19941) );
  XNOR U21622 ( .A(a[423]), .B(n4132), .Z(n19976) );
  NAND U21623 ( .A(n42144), .B(n19976), .Z(n19940) );
  AND U21624 ( .A(n19941), .B(n19940), .Z(n19991) );
  XOR U21625 ( .A(a[427]), .B(n42012), .Z(n19979) );
  XNOR U21626 ( .A(n19991), .B(n19990), .Z(n19993) );
  AND U21627 ( .A(a[429]), .B(b[0]), .Z(n19943) );
  XNOR U21628 ( .A(n19943), .B(n4071), .Z(n19945) );
  NANDN U21629 ( .A(b[0]), .B(a[428]), .Z(n19944) );
  NAND U21630 ( .A(n19945), .B(n19944), .Z(n19987) );
  XOR U21631 ( .A(a[425]), .B(n42085), .Z(n19980) );
  AND U21632 ( .A(a[421]), .B(b[7]), .Z(n19984) );
  XNOR U21633 ( .A(n19985), .B(n19984), .Z(n19986) );
  XNOR U21634 ( .A(n19987), .B(n19986), .Z(n19992) );
  XOR U21635 ( .A(n19993), .B(n19992), .Z(n19971) );
  NANDN U21636 ( .A(n19948), .B(n19947), .Z(n19952) );
  NANDN U21637 ( .A(n19950), .B(n19949), .Z(n19951) );
  AND U21638 ( .A(n19952), .B(n19951), .Z(n19970) );
  XNOR U21639 ( .A(n19971), .B(n19970), .Z(n19972) );
  NANDN U21640 ( .A(n19954), .B(n19953), .Z(n19958) );
  NAND U21641 ( .A(n19956), .B(n19955), .Z(n19957) );
  NAND U21642 ( .A(n19958), .B(n19957), .Z(n19973) );
  XNOR U21643 ( .A(n19972), .B(n19973), .Z(n19964) );
  XNOR U21644 ( .A(n19965), .B(n19964), .Z(n19966) );
  XNOR U21645 ( .A(n19967), .B(n19966), .Z(n19996) );
  XNOR U21646 ( .A(sreg[1445]), .B(n19996), .Z(n19998) );
  NANDN U21647 ( .A(sreg[1444]), .B(n19959), .Z(n19963) );
  NAND U21648 ( .A(n19961), .B(n19960), .Z(n19962) );
  NAND U21649 ( .A(n19963), .B(n19962), .Z(n19997) );
  XNOR U21650 ( .A(n19998), .B(n19997), .Z(c[1445]) );
  NANDN U21651 ( .A(n19965), .B(n19964), .Z(n19969) );
  NANDN U21652 ( .A(n19967), .B(n19966), .Z(n19968) );
  AND U21653 ( .A(n19969), .B(n19968), .Z(n20004) );
  NANDN U21654 ( .A(n19971), .B(n19970), .Z(n19975) );
  NANDN U21655 ( .A(n19973), .B(n19972), .Z(n19974) );
  AND U21656 ( .A(n19975), .B(n19974), .Z(n20002) );
  NAND U21657 ( .A(n42143), .B(n19976), .Z(n19978) );
  XNOR U21658 ( .A(a[424]), .B(n4132), .Z(n20013) );
  NAND U21659 ( .A(n42144), .B(n20013), .Z(n19977) );
  AND U21660 ( .A(n19978), .B(n19977), .Z(n20028) );
  XOR U21661 ( .A(a[428]), .B(n42012), .Z(n20016) );
  XNOR U21662 ( .A(n20028), .B(n20027), .Z(n20030) );
  XOR U21663 ( .A(a[426]), .B(n42085), .Z(n20020) );
  AND U21664 ( .A(a[422]), .B(b[7]), .Z(n20021) );
  XNOR U21665 ( .A(n20022), .B(n20021), .Z(n20023) );
  AND U21666 ( .A(a[430]), .B(b[0]), .Z(n19981) );
  XNOR U21667 ( .A(n19981), .B(n4071), .Z(n19983) );
  NANDN U21668 ( .A(b[0]), .B(a[429]), .Z(n19982) );
  NAND U21669 ( .A(n19983), .B(n19982), .Z(n20024) );
  XNOR U21670 ( .A(n20023), .B(n20024), .Z(n20029) );
  XOR U21671 ( .A(n20030), .B(n20029), .Z(n20008) );
  NANDN U21672 ( .A(n19985), .B(n19984), .Z(n19989) );
  NANDN U21673 ( .A(n19987), .B(n19986), .Z(n19988) );
  AND U21674 ( .A(n19989), .B(n19988), .Z(n20007) );
  XNOR U21675 ( .A(n20008), .B(n20007), .Z(n20009) );
  NANDN U21676 ( .A(n19991), .B(n19990), .Z(n19995) );
  NAND U21677 ( .A(n19993), .B(n19992), .Z(n19994) );
  NAND U21678 ( .A(n19995), .B(n19994), .Z(n20010) );
  XNOR U21679 ( .A(n20009), .B(n20010), .Z(n20001) );
  XNOR U21680 ( .A(n20002), .B(n20001), .Z(n20003) );
  XNOR U21681 ( .A(n20004), .B(n20003), .Z(n20033) );
  XNOR U21682 ( .A(sreg[1446]), .B(n20033), .Z(n20035) );
  NANDN U21683 ( .A(sreg[1445]), .B(n19996), .Z(n20000) );
  NAND U21684 ( .A(n19998), .B(n19997), .Z(n19999) );
  NAND U21685 ( .A(n20000), .B(n19999), .Z(n20034) );
  XNOR U21686 ( .A(n20035), .B(n20034), .Z(c[1446]) );
  NANDN U21687 ( .A(n20002), .B(n20001), .Z(n20006) );
  NANDN U21688 ( .A(n20004), .B(n20003), .Z(n20005) );
  AND U21689 ( .A(n20006), .B(n20005), .Z(n20041) );
  NANDN U21690 ( .A(n20008), .B(n20007), .Z(n20012) );
  NANDN U21691 ( .A(n20010), .B(n20009), .Z(n20011) );
  AND U21692 ( .A(n20012), .B(n20011), .Z(n20039) );
  NAND U21693 ( .A(n42143), .B(n20013), .Z(n20015) );
  XNOR U21694 ( .A(a[425]), .B(n4132), .Z(n20050) );
  NAND U21695 ( .A(n42144), .B(n20050), .Z(n20014) );
  AND U21696 ( .A(n20015), .B(n20014), .Z(n20065) );
  XOR U21697 ( .A(a[429]), .B(n42012), .Z(n20053) );
  XNOR U21698 ( .A(n20065), .B(n20064), .Z(n20067) );
  AND U21699 ( .A(a[431]), .B(b[0]), .Z(n20017) );
  XNOR U21700 ( .A(n20017), .B(n4071), .Z(n20019) );
  NANDN U21701 ( .A(b[0]), .B(a[430]), .Z(n20018) );
  NAND U21702 ( .A(n20019), .B(n20018), .Z(n20061) );
  XOR U21703 ( .A(a[427]), .B(n42085), .Z(n20057) );
  AND U21704 ( .A(a[423]), .B(b[7]), .Z(n20058) );
  XNOR U21705 ( .A(n20059), .B(n20058), .Z(n20060) );
  XNOR U21706 ( .A(n20061), .B(n20060), .Z(n20066) );
  XOR U21707 ( .A(n20067), .B(n20066), .Z(n20045) );
  NANDN U21708 ( .A(n20022), .B(n20021), .Z(n20026) );
  NANDN U21709 ( .A(n20024), .B(n20023), .Z(n20025) );
  AND U21710 ( .A(n20026), .B(n20025), .Z(n20044) );
  XNOR U21711 ( .A(n20045), .B(n20044), .Z(n20046) );
  NANDN U21712 ( .A(n20028), .B(n20027), .Z(n20032) );
  NAND U21713 ( .A(n20030), .B(n20029), .Z(n20031) );
  NAND U21714 ( .A(n20032), .B(n20031), .Z(n20047) );
  XNOR U21715 ( .A(n20046), .B(n20047), .Z(n20038) );
  XNOR U21716 ( .A(n20039), .B(n20038), .Z(n20040) );
  XNOR U21717 ( .A(n20041), .B(n20040), .Z(n20070) );
  XNOR U21718 ( .A(sreg[1447]), .B(n20070), .Z(n20072) );
  NANDN U21719 ( .A(sreg[1446]), .B(n20033), .Z(n20037) );
  NAND U21720 ( .A(n20035), .B(n20034), .Z(n20036) );
  NAND U21721 ( .A(n20037), .B(n20036), .Z(n20071) );
  XNOR U21722 ( .A(n20072), .B(n20071), .Z(c[1447]) );
  NANDN U21723 ( .A(n20039), .B(n20038), .Z(n20043) );
  NANDN U21724 ( .A(n20041), .B(n20040), .Z(n20042) );
  AND U21725 ( .A(n20043), .B(n20042), .Z(n20078) );
  NANDN U21726 ( .A(n20045), .B(n20044), .Z(n20049) );
  NANDN U21727 ( .A(n20047), .B(n20046), .Z(n20048) );
  AND U21728 ( .A(n20049), .B(n20048), .Z(n20076) );
  NAND U21729 ( .A(n42143), .B(n20050), .Z(n20052) );
  XNOR U21730 ( .A(a[426]), .B(n4132), .Z(n20087) );
  NAND U21731 ( .A(n42144), .B(n20087), .Z(n20051) );
  AND U21732 ( .A(n20052), .B(n20051), .Z(n20102) );
  XOR U21733 ( .A(a[430]), .B(n42012), .Z(n20090) );
  XNOR U21734 ( .A(n20102), .B(n20101), .Z(n20104) );
  AND U21735 ( .A(b[0]), .B(a[432]), .Z(n20054) );
  XOR U21736 ( .A(b[1]), .B(n20054), .Z(n20056) );
  NANDN U21737 ( .A(b[0]), .B(a[431]), .Z(n20055) );
  AND U21738 ( .A(n20056), .B(n20055), .Z(n20097) );
  XOR U21739 ( .A(a[428]), .B(n42085), .Z(n20094) );
  AND U21740 ( .A(a[424]), .B(b[7]), .Z(n20095) );
  XOR U21741 ( .A(n20096), .B(n20095), .Z(n20098) );
  XNOR U21742 ( .A(n20097), .B(n20098), .Z(n20103) );
  XOR U21743 ( .A(n20104), .B(n20103), .Z(n20082) );
  NANDN U21744 ( .A(n20059), .B(n20058), .Z(n20063) );
  NANDN U21745 ( .A(n20061), .B(n20060), .Z(n20062) );
  AND U21746 ( .A(n20063), .B(n20062), .Z(n20081) );
  XNOR U21747 ( .A(n20082), .B(n20081), .Z(n20083) );
  NANDN U21748 ( .A(n20065), .B(n20064), .Z(n20069) );
  NAND U21749 ( .A(n20067), .B(n20066), .Z(n20068) );
  NAND U21750 ( .A(n20069), .B(n20068), .Z(n20084) );
  XNOR U21751 ( .A(n20083), .B(n20084), .Z(n20075) );
  XNOR U21752 ( .A(n20076), .B(n20075), .Z(n20077) );
  XNOR U21753 ( .A(n20078), .B(n20077), .Z(n20107) );
  XNOR U21754 ( .A(sreg[1448]), .B(n20107), .Z(n20109) );
  NANDN U21755 ( .A(sreg[1447]), .B(n20070), .Z(n20074) );
  NAND U21756 ( .A(n20072), .B(n20071), .Z(n20073) );
  NAND U21757 ( .A(n20074), .B(n20073), .Z(n20108) );
  XNOR U21758 ( .A(n20109), .B(n20108), .Z(c[1448]) );
  NANDN U21759 ( .A(n20076), .B(n20075), .Z(n20080) );
  NANDN U21760 ( .A(n20078), .B(n20077), .Z(n20079) );
  AND U21761 ( .A(n20080), .B(n20079), .Z(n20115) );
  NANDN U21762 ( .A(n20082), .B(n20081), .Z(n20086) );
  NANDN U21763 ( .A(n20084), .B(n20083), .Z(n20085) );
  AND U21764 ( .A(n20086), .B(n20085), .Z(n20113) );
  NAND U21765 ( .A(n42143), .B(n20087), .Z(n20089) );
  XNOR U21766 ( .A(a[427]), .B(n4132), .Z(n20124) );
  NAND U21767 ( .A(n42144), .B(n20124), .Z(n20088) );
  AND U21768 ( .A(n20089), .B(n20088), .Z(n20139) );
  XOR U21769 ( .A(a[431]), .B(n42012), .Z(n20127) );
  XNOR U21770 ( .A(n20139), .B(n20138), .Z(n20141) );
  AND U21771 ( .A(a[433]), .B(b[0]), .Z(n20091) );
  XNOR U21772 ( .A(n20091), .B(n4071), .Z(n20093) );
  NANDN U21773 ( .A(b[0]), .B(a[432]), .Z(n20092) );
  NAND U21774 ( .A(n20093), .B(n20092), .Z(n20135) );
  XOR U21775 ( .A(a[429]), .B(n42085), .Z(n20131) );
  AND U21776 ( .A(a[425]), .B(b[7]), .Z(n20132) );
  XNOR U21777 ( .A(n20133), .B(n20132), .Z(n20134) );
  XNOR U21778 ( .A(n20135), .B(n20134), .Z(n20140) );
  XOR U21779 ( .A(n20141), .B(n20140), .Z(n20119) );
  NANDN U21780 ( .A(n20096), .B(n20095), .Z(n20100) );
  NANDN U21781 ( .A(n20098), .B(n20097), .Z(n20099) );
  AND U21782 ( .A(n20100), .B(n20099), .Z(n20118) );
  XNOR U21783 ( .A(n20119), .B(n20118), .Z(n20120) );
  NANDN U21784 ( .A(n20102), .B(n20101), .Z(n20106) );
  NAND U21785 ( .A(n20104), .B(n20103), .Z(n20105) );
  NAND U21786 ( .A(n20106), .B(n20105), .Z(n20121) );
  XNOR U21787 ( .A(n20120), .B(n20121), .Z(n20112) );
  XNOR U21788 ( .A(n20113), .B(n20112), .Z(n20114) );
  XNOR U21789 ( .A(n20115), .B(n20114), .Z(n20144) );
  XNOR U21790 ( .A(sreg[1449]), .B(n20144), .Z(n20146) );
  NANDN U21791 ( .A(sreg[1448]), .B(n20107), .Z(n20111) );
  NAND U21792 ( .A(n20109), .B(n20108), .Z(n20110) );
  NAND U21793 ( .A(n20111), .B(n20110), .Z(n20145) );
  XNOR U21794 ( .A(n20146), .B(n20145), .Z(c[1449]) );
  NANDN U21795 ( .A(n20113), .B(n20112), .Z(n20117) );
  NANDN U21796 ( .A(n20115), .B(n20114), .Z(n20116) );
  AND U21797 ( .A(n20117), .B(n20116), .Z(n20152) );
  NANDN U21798 ( .A(n20119), .B(n20118), .Z(n20123) );
  NANDN U21799 ( .A(n20121), .B(n20120), .Z(n20122) );
  AND U21800 ( .A(n20123), .B(n20122), .Z(n20150) );
  NAND U21801 ( .A(n42143), .B(n20124), .Z(n20126) );
  XNOR U21802 ( .A(a[428]), .B(n4133), .Z(n20161) );
  NAND U21803 ( .A(n42144), .B(n20161), .Z(n20125) );
  AND U21804 ( .A(n20126), .B(n20125), .Z(n20176) );
  XOR U21805 ( .A(a[432]), .B(n42012), .Z(n20164) );
  XNOR U21806 ( .A(n20176), .B(n20175), .Z(n20178) );
  AND U21807 ( .A(a[434]), .B(b[0]), .Z(n20128) );
  XNOR U21808 ( .A(n20128), .B(n4071), .Z(n20130) );
  NANDN U21809 ( .A(b[0]), .B(a[433]), .Z(n20129) );
  NAND U21810 ( .A(n20130), .B(n20129), .Z(n20172) );
  XOR U21811 ( .A(a[430]), .B(n42085), .Z(n20165) );
  AND U21812 ( .A(a[426]), .B(b[7]), .Z(n20169) );
  XNOR U21813 ( .A(n20170), .B(n20169), .Z(n20171) );
  XNOR U21814 ( .A(n20172), .B(n20171), .Z(n20177) );
  XOR U21815 ( .A(n20178), .B(n20177), .Z(n20156) );
  NANDN U21816 ( .A(n20133), .B(n20132), .Z(n20137) );
  NANDN U21817 ( .A(n20135), .B(n20134), .Z(n20136) );
  AND U21818 ( .A(n20137), .B(n20136), .Z(n20155) );
  XNOR U21819 ( .A(n20156), .B(n20155), .Z(n20157) );
  NANDN U21820 ( .A(n20139), .B(n20138), .Z(n20143) );
  NAND U21821 ( .A(n20141), .B(n20140), .Z(n20142) );
  NAND U21822 ( .A(n20143), .B(n20142), .Z(n20158) );
  XNOR U21823 ( .A(n20157), .B(n20158), .Z(n20149) );
  XNOR U21824 ( .A(n20150), .B(n20149), .Z(n20151) );
  XNOR U21825 ( .A(n20152), .B(n20151), .Z(n20181) );
  XNOR U21826 ( .A(sreg[1450]), .B(n20181), .Z(n20183) );
  NANDN U21827 ( .A(sreg[1449]), .B(n20144), .Z(n20148) );
  NAND U21828 ( .A(n20146), .B(n20145), .Z(n20147) );
  NAND U21829 ( .A(n20148), .B(n20147), .Z(n20182) );
  XNOR U21830 ( .A(n20183), .B(n20182), .Z(c[1450]) );
  NANDN U21831 ( .A(n20150), .B(n20149), .Z(n20154) );
  NANDN U21832 ( .A(n20152), .B(n20151), .Z(n20153) );
  AND U21833 ( .A(n20154), .B(n20153), .Z(n20189) );
  NANDN U21834 ( .A(n20156), .B(n20155), .Z(n20160) );
  NANDN U21835 ( .A(n20158), .B(n20157), .Z(n20159) );
  AND U21836 ( .A(n20160), .B(n20159), .Z(n20187) );
  NAND U21837 ( .A(n42143), .B(n20161), .Z(n20163) );
  XNOR U21838 ( .A(a[429]), .B(n4133), .Z(n20198) );
  NAND U21839 ( .A(n42144), .B(n20198), .Z(n20162) );
  AND U21840 ( .A(n20163), .B(n20162), .Z(n20213) );
  XOR U21841 ( .A(a[433]), .B(n42012), .Z(n20201) );
  XNOR U21842 ( .A(n20213), .B(n20212), .Z(n20215) );
  XOR U21843 ( .A(a[431]), .B(n42085), .Z(n20205) );
  AND U21844 ( .A(a[427]), .B(b[7]), .Z(n20206) );
  XNOR U21845 ( .A(n20207), .B(n20206), .Z(n20208) );
  AND U21846 ( .A(a[435]), .B(b[0]), .Z(n20166) );
  XNOR U21847 ( .A(n20166), .B(n4071), .Z(n20168) );
  NANDN U21848 ( .A(b[0]), .B(a[434]), .Z(n20167) );
  NAND U21849 ( .A(n20168), .B(n20167), .Z(n20209) );
  XNOR U21850 ( .A(n20208), .B(n20209), .Z(n20214) );
  XOR U21851 ( .A(n20215), .B(n20214), .Z(n20193) );
  NANDN U21852 ( .A(n20170), .B(n20169), .Z(n20174) );
  NANDN U21853 ( .A(n20172), .B(n20171), .Z(n20173) );
  AND U21854 ( .A(n20174), .B(n20173), .Z(n20192) );
  XNOR U21855 ( .A(n20193), .B(n20192), .Z(n20194) );
  NANDN U21856 ( .A(n20176), .B(n20175), .Z(n20180) );
  NAND U21857 ( .A(n20178), .B(n20177), .Z(n20179) );
  NAND U21858 ( .A(n20180), .B(n20179), .Z(n20195) );
  XNOR U21859 ( .A(n20194), .B(n20195), .Z(n20186) );
  XNOR U21860 ( .A(n20187), .B(n20186), .Z(n20188) );
  XNOR U21861 ( .A(n20189), .B(n20188), .Z(n20218) );
  XNOR U21862 ( .A(sreg[1451]), .B(n20218), .Z(n20220) );
  NANDN U21863 ( .A(sreg[1450]), .B(n20181), .Z(n20185) );
  NAND U21864 ( .A(n20183), .B(n20182), .Z(n20184) );
  NAND U21865 ( .A(n20185), .B(n20184), .Z(n20219) );
  XNOR U21866 ( .A(n20220), .B(n20219), .Z(c[1451]) );
  NANDN U21867 ( .A(n20187), .B(n20186), .Z(n20191) );
  NANDN U21868 ( .A(n20189), .B(n20188), .Z(n20190) );
  AND U21869 ( .A(n20191), .B(n20190), .Z(n20226) );
  NANDN U21870 ( .A(n20193), .B(n20192), .Z(n20197) );
  NANDN U21871 ( .A(n20195), .B(n20194), .Z(n20196) );
  AND U21872 ( .A(n20197), .B(n20196), .Z(n20224) );
  NAND U21873 ( .A(n42143), .B(n20198), .Z(n20200) );
  XNOR U21874 ( .A(a[430]), .B(n4133), .Z(n20235) );
  NAND U21875 ( .A(n42144), .B(n20235), .Z(n20199) );
  AND U21876 ( .A(n20200), .B(n20199), .Z(n20250) );
  XOR U21877 ( .A(a[434]), .B(n42012), .Z(n20238) );
  XNOR U21878 ( .A(n20250), .B(n20249), .Z(n20252) );
  AND U21879 ( .A(a[436]), .B(b[0]), .Z(n20202) );
  XNOR U21880 ( .A(n20202), .B(n4071), .Z(n20204) );
  NANDN U21881 ( .A(b[0]), .B(a[435]), .Z(n20203) );
  NAND U21882 ( .A(n20204), .B(n20203), .Z(n20246) );
  XOR U21883 ( .A(a[432]), .B(n42085), .Z(n20242) );
  AND U21884 ( .A(a[428]), .B(b[7]), .Z(n20243) );
  XNOR U21885 ( .A(n20244), .B(n20243), .Z(n20245) );
  XNOR U21886 ( .A(n20246), .B(n20245), .Z(n20251) );
  XOR U21887 ( .A(n20252), .B(n20251), .Z(n20230) );
  NANDN U21888 ( .A(n20207), .B(n20206), .Z(n20211) );
  NANDN U21889 ( .A(n20209), .B(n20208), .Z(n20210) );
  AND U21890 ( .A(n20211), .B(n20210), .Z(n20229) );
  XNOR U21891 ( .A(n20230), .B(n20229), .Z(n20231) );
  NANDN U21892 ( .A(n20213), .B(n20212), .Z(n20217) );
  NAND U21893 ( .A(n20215), .B(n20214), .Z(n20216) );
  NAND U21894 ( .A(n20217), .B(n20216), .Z(n20232) );
  XNOR U21895 ( .A(n20231), .B(n20232), .Z(n20223) );
  XNOR U21896 ( .A(n20224), .B(n20223), .Z(n20225) );
  XNOR U21897 ( .A(n20226), .B(n20225), .Z(n20255) );
  XNOR U21898 ( .A(sreg[1452]), .B(n20255), .Z(n20257) );
  NANDN U21899 ( .A(sreg[1451]), .B(n20218), .Z(n20222) );
  NAND U21900 ( .A(n20220), .B(n20219), .Z(n20221) );
  NAND U21901 ( .A(n20222), .B(n20221), .Z(n20256) );
  XNOR U21902 ( .A(n20257), .B(n20256), .Z(c[1452]) );
  NANDN U21903 ( .A(n20224), .B(n20223), .Z(n20228) );
  NANDN U21904 ( .A(n20226), .B(n20225), .Z(n20227) );
  AND U21905 ( .A(n20228), .B(n20227), .Z(n20263) );
  NANDN U21906 ( .A(n20230), .B(n20229), .Z(n20234) );
  NANDN U21907 ( .A(n20232), .B(n20231), .Z(n20233) );
  AND U21908 ( .A(n20234), .B(n20233), .Z(n20261) );
  NAND U21909 ( .A(n42143), .B(n20235), .Z(n20237) );
  XNOR U21910 ( .A(a[431]), .B(n4133), .Z(n20272) );
  NAND U21911 ( .A(n42144), .B(n20272), .Z(n20236) );
  AND U21912 ( .A(n20237), .B(n20236), .Z(n20287) );
  XOR U21913 ( .A(a[435]), .B(n42012), .Z(n20275) );
  XNOR U21914 ( .A(n20287), .B(n20286), .Z(n20289) );
  AND U21915 ( .A(a[437]), .B(b[0]), .Z(n20239) );
  XNOR U21916 ( .A(n20239), .B(n4071), .Z(n20241) );
  NANDN U21917 ( .A(b[0]), .B(a[436]), .Z(n20240) );
  NAND U21918 ( .A(n20241), .B(n20240), .Z(n20283) );
  XOR U21919 ( .A(a[433]), .B(n42085), .Z(n20279) );
  AND U21920 ( .A(a[429]), .B(b[7]), .Z(n20280) );
  XNOR U21921 ( .A(n20281), .B(n20280), .Z(n20282) );
  XNOR U21922 ( .A(n20283), .B(n20282), .Z(n20288) );
  XOR U21923 ( .A(n20289), .B(n20288), .Z(n20267) );
  NANDN U21924 ( .A(n20244), .B(n20243), .Z(n20248) );
  NANDN U21925 ( .A(n20246), .B(n20245), .Z(n20247) );
  AND U21926 ( .A(n20248), .B(n20247), .Z(n20266) );
  XNOR U21927 ( .A(n20267), .B(n20266), .Z(n20268) );
  NANDN U21928 ( .A(n20250), .B(n20249), .Z(n20254) );
  NAND U21929 ( .A(n20252), .B(n20251), .Z(n20253) );
  NAND U21930 ( .A(n20254), .B(n20253), .Z(n20269) );
  XNOR U21931 ( .A(n20268), .B(n20269), .Z(n20260) );
  XNOR U21932 ( .A(n20261), .B(n20260), .Z(n20262) );
  XNOR U21933 ( .A(n20263), .B(n20262), .Z(n20292) );
  XNOR U21934 ( .A(sreg[1453]), .B(n20292), .Z(n20294) );
  NANDN U21935 ( .A(sreg[1452]), .B(n20255), .Z(n20259) );
  NAND U21936 ( .A(n20257), .B(n20256), .Z(n20258) );
  NAND U21937 ( .A(n20259), .B(n20258), .Z(n20293) );
  XNOR U21938 ( .A(n20294), .B(n20293), .Z(c[1453]) );
  NANDN U21939 ( .A(n20261), .B(n20260), .Z(n20265) );
  NANDN U21940 ( .A(n20263), .B(n20262), .Z(n20264) );
  AND U21941 ( .A(n20265), .B(n20264), .Z(n20300) );
  NANDN U21942 ( .A(n20267), .B(n20266), .Z(n20271) );
  NANDN U21943 ( .A(n20269), .B(n20268), .Z(n20270) );
  AND U21944 ( .A(n20271), .B(n20270), .Z(n20298) );
  NAND U21945 ( .A(n42143), .B(n20272), .Z(n20274) );
  XNOR U21946 ( .A(a[432]), .B(n4133), .Z(n20309) );
  NAND U21947 ( .A(n42144), .B(n20309), .Z(n20273) );
  AND U21948 ( .A(n20274), .B(n20273), .Z(n20324) );
  XOR U21949 ( .A(a[436]), .B(n42012), .Z(n20312) );
  XNOR U21950 ( .A(n20324), .B(n20323), .Z(n20326) );
  AND U21951 ( .A(a[438]), .B(b[0]), .Z(n20276) );
  XNOR U21952 ( .A(n20276), .B(n4071), .Z(n20278) );
  NANDN U21953 ( .A(b[0]), .B(a[437]), .Z(n20277) );
  NAND U21954 ( .A(n20278), .B(n20277), .Z(n20320) );
  XOR U21955 ( .A(a[434]), .B(n42085), .Z(n20316) );
  AND U21956 ( .A(a[430]), .B(b[7]), .Z(n20317) );
  XNOR U21957 ( .A(n20318), .B(n20317), .Z(n20319) );
  XNOR U21958 ( .A(n20320), .B(n20319), .Z(n20325) );
  XOR U21959 ( .A(n20326), .B(n20325), .Z(n20304) );
  NANDN U21960 ( .A(n20281), .B(n20280), .Z(n20285) );
  NANDN U21961 ( .A(n20283), .B(n20282), .Z(n20284) );
  AND U21962 ( .A(n20285), .B(n20284), .Z(n20303) );
  XNOR U21963 ( .A(n20304), .B(n20303), .Z(n20305) );
  NANDN U21964 ( .A(n20287), .B(n20286), .Z(n20291) );
  NAND U21965 ( .A(n20289), .B(n20288), .Z(n20290) );
  NAND U21966 ( .A(n20291), .B(n20290), .Z(n20306) );
  XNOR U21967 ( .A(n20305), .B(n20306), .Z(n20297) );
  XNOR U21968 ( .A(n20298), .B(n20297), .Z(n20299) );
  XNOR U21969 ( .A(n20300), .B(n20299), .Z(n20329) );
  XNOR U21970 ( .A(sreg[1454]), .B(n20329), .Z(n20331) );
  NANDN U21971 ( .A(sreg[1453]), .B(n20292), .Z(n20296) );
  NAND U21972 ( .A(n20294), .B(n20293), .Z(n20295) );
  NAND U21973 ( .A(n20296), .B(n20295), .Z(n20330) );
  XNOR U21974 ( .A(n20331), .B(n20330), .Z(c[1454]) );
  NANDN U21975 ( .A(n20298), .B(n20297), .Z(n20302) );
  NANDN U21976 ( .A(n20300), .B(n20299), .Z(n20301) );
  AND U21977 ( .A(n20302), .B(n20301), .Z(n20337) );
  NANDN U21978 ( .A(n20304), .B(n20303), .Z(n20308) );
  NANDN U21979 ( .A(n20306), .B(n20305), .Z(n20307) );
  AND U21980 ( .A(n20308), .B(n20307), .Z(n20335) );
  NAND U21981 ( .A(n42143), .B(n20309), .Z(n20311) );
  XNOR U21982 ( .A(a[433]), .B(n4133), .Z(n20346) );
  NAND U21983 ( .A(n42144), .B(n20346), .Z(n20310) );
  AND U21984 ( .A(n20311), .B(n20310), .Z(n20361) );
  XOR U21985 ( .A(a[437]), .B(n42012), .Z(n20349) );
  XNOR U21986 ( .A(n20361), .B(n20360), .Z(n20363) );
  AND U21987 ( .A(a[439]), .B(b[0]), .Z(n20313) );
  XNOR U21988 ( .A(n20313), .B(n4071), .Z(n20315) );
  NANDN U21989 ( .A(b[0]), .B(a[438]), .Z(n20314) );
  NAND U21990 ( .A(n20315), .B(n20314), .Z(n20357) );
  XOR U21991 ( .A(a[435]), .B(n42085), .Z(n20353) );
  AND U21992 ( .A(a[431]), .B(b[7]), .Z(n20354) );
  XNOR U21993 ( .A(n20355), .B(n20354), .Z(n20356) );
  XNOR U21994 ( .A(n20357), .B(n20356), .Z(n20362) );
  XOR U21995 ( .A(n20363), .B(n20362), .Z(n20341) );
  NANDN U21996 ( .A(n20318), .B(n20317), .Z(n20322) );
  NANDN U21997 ( .A(n20320), .B(n20319), .Z(n20321) );
  AND U21998 ( .A(n20322), .B(n20321), .Z(n20340) );
  XNOR U21999 ( .A(n20341), .B(n20340), .Z(n20342) );
  NANDN U22000 ( .A(n20324), .B(n20323), .Z(n20328) );
  NAND U22001 ( .A(n20326), .B(n20325), .Z(n20327) );
  NAND U22002 ( .A(n20328), .B(n20327), .Z(n20343) );
  XNOR U22003 ( .A(n20342), .B(n20343), .Z(n20334) );
  XNOR U22004 ( .A(n20335), .B(n20334), .Z(n20336) );
  XNOR U22005 ( .A(n20337), .B(n20336), .Z(n20366) );
  XNOR U22006 ( .A(sreg[1455]), .B(n20366), .Z(n20368) );
  NANDN U22007 ( .A(sreg[1454]), .B(n20329), .Z(n20333) );
  NAND U22008 ( .A(n20331), .B(n20330), .Z(n20332) );
  NAND U22009 ( .A(n20333), .B(n20332), .Z(n20367) );
  XNOR U22010 ( .A(n20368), .B(n20367), .Z(c[1455]) );
  NANDN U22011 ( .A(n20335), .B(n20334), .Z(n20339) );
  NANDN U22012 ( .A(n20337), .B(n20336), .Z(n20338) );
  AND U22013 ( .A(n20339), .B(n20338), .Z(n20374) );
  NANDN U22014 ( .A(n20341), .B(n20340), .Z(n20345) );
  NANDN U22015 ( .A(n20343), .B(n20342), .Z(n20344) );
  AND U22016 ( .A(n20345), .B(n20344), .Z(n20372) );
  NAND U22017 ( .A(n42143), .B(n20346), .Z(n20348) );
  XNOR U22018 ( .A(a[434]), .B(n4133), .Z(n20383) );
  NAND U22019 ( .A(n42144), .B(n20383), .Z(n20347) );
  AND U22020 ( .A(n20348), .B(n20347), .Z(n20398) );
  XOR U22021 ( .A(a[438]), .B(n42012), .Z(n20386) );
  XNOR U22022 ( .A(n20398), .B(n20397), .Z(n20400) );
  AND U22023 ( .A(a[440]), .B(b[0]), .Z(n20350) );
  XNOR U22024 ( .A(n20350), .B(n4071), .Z(n20352) );
  NANDN U22025 ( .A(b[0]), .B(a[439]), .Z(n20351) );
  NAND U22026 ( .A(n20352), .B(n20351), .Z(n20394) );
  XOR U22027 ( .A(a[436]), .B(n42085), .Z(n20390) );
  AND U22028 ( .A(a[432]), .B(b[7]), .Z(n20391) );
  XNOR U22029 ( .A(n20392), .B(n20391), .Z(n20393) );
  XNOR U22030 ( .A(n20394), .B(n20393), .Z(n20399) );
  XOR U22031 ( .A(n20400), .B(n20399), .Z(n20378) );
  NANDN U22032 ( .A(n20355), .B(n20354), .Z(n20359) );
  NANDN U22033 ( .A(n20357), .B(n20356), .Z(n20358) );
  AND U22034 ( .A(n20359), .B(n20358), .Z(n20377) );
  XNOR U22035 ( .A(n20378), .B(n20377), .Z(n20379) );
  NANDN U22036 ( .A(n20361), .B(n20360), .Z(n20365) );
  NAND U22037 ( .A(n20363), .B(n20362), .Z(n20364) );
  NAND U22038 ( .A(n20365), .B(n20364), .Z(n20380) );
  XNOR U22039 ( .A(n20379), .B(n20380), .Z(n20371) );
  XNOR U22040 ( .A(n20372), .B(n20371), .Z(n20373) );
  XNOR U22041 ( .A(n20374), .B(n20373), .Z(n20403) );
  XNOR U22042 ( .A(sreg[1456]), .B(n20403), .Z(n20405) );
  NANDN U22043 ( .A(sreg[1455]), .B(n20366), .Z(n20370) );
  NAND U22044 ( .A(n20368), .B(n20367), .Z(n20369) );
  NAND U22045 ( .A(n20370), .B(n20369), .Z(n20404) );
  XNOR U22046 ( .A(n20405), .B(n20404), .Z(c[1456]) );
  NANDN U22047 ( .A(n20372), .B(n20371), .Z(n20376) );
  NANDN U22048 ( .A(n20374), .B(n20373), .Z(n20375) );
  AND U22049 ( .A(n20376), .B(n20375), .Z(n20411) );
  NANDN U22050 ( .A(n20378), .B(n20377), .Z(n20382) );
  NANDN U22051 ( .A(n20380), .B(n20379), .Z(n20381) );
  AND U22052 ( .A(n20382), .B(n20381), .Z(n20409) );
  NAND U22053 ( .A(n42143), .B(n20383), .Z(n20385) );
  XNOR U22054 ( .A(a[435]), .B(n4134), .Z(n20420) );
  NAND U22055 ( .A(n42144), .B(n20420), .Z(n20384) );
  AND U22056 ( .A(n20385), .B(n20384), .Z(n20435) );
  XOR U22057 ( .A(a[439]), .B(n42012), .Z(n20423) );
  XNOR U22058 ( .A(n20435), .B(n20434), .Z(n20437) );
  AND U22059 ( .A(a[441]), .B(b[0]), .Z(n20387) );
  XNOR U22060 ( .A(n20387), .B(n4071), .Z(n20389) );
  NANDN U22061 ( .A(b[0]), .B(a[440]), .Z(n20388) );
  NAND U22062 ( .A(n20389), .B(n20388), .Z(n20431) );
  XOR U22063 ( .A(a[437]), .B(n42085), .Z(n20424) );
  AND U22064 ( .A(a[433]), .B(b[7]), .Z(n20428) );
  XNOR U22065 ( .A(n20429), .B(n20428), .Z(n20430) );
  XNOR U22066 ( .A(n20431), .B(n20430), .Z(n20436) );
  XOR U22067 ( .A(n20437), .B(n20436), .Z(n20415) );
  NANDN U22068 ( .A(n20392), .B(n20391), .Z(n20396) );
  NANDN U22069 ( .A(n20394), .B(n20393), .Z(n20395) );
  AND U22070 ( .A(n20396), .B(n20395), .Z(n20414) );
  XNOR U22071 ( .A(n20415), .B(n20414), .Z(n20416) );
  NANDN U22072 ( .A(n20398), .B(n20397), .Z(n20402) );
  NAND U22073 ( .A(n20400), .B(n20399), .Z(n20401) );
  NAND U22074 ( .A(n20402), .B(n20401), .Z(n20417) );
  XNOR U22075 ( .A(n20416), .B(n20417), .Z(n20408) );
  XNOR U22076 ( .A(n20409), .B(n20408), .Z(n20410) );
  XNOR U22077 ( .A(n20411), .B(n20410), .Z(n20440) );
  XNOR U22078 ( .A(sreg[1457]), .B(n20440), .Z(n20442) );
  NANDN U22079 ( .A(sreg[1456]), .B(n20403), .Z(n20407) );
  NAND U22080 ( .A(n20405), .B(n20404), .Z(n20406) );
  NAND U22081 ( .A(n20407), .B(n20406), .Z(n20441) );
  XNOR U22082 ( .A(n20442), .B(n20441), .Z(c[1457]) );
  NANDN U22083 ( .A(n20409), .B(n20408), .Z(n20413) );
  NANDN U22084 ( .A(n20411), .B(n20410), .Z(n20412) );
  AND U22085 ( .A(n20413), .B(n20412), .Z(n20448) );
  NANDN U22086 ( .A(n20415), .B(n20414), .Z(n20419) );
  NANDN U22087 ( .A(n20417), .B(n20416), .Z(n20418) );
  AND U22088 ( .A(n20419), .B(n20418), .Z(n20446) );
  NAND U22089 ( .A(n42143), .B(n20420), .Z(n20422) );
  XNOR U22090 ( .A(a[436]), .B(n4134), .Z(n20457) );
  NAND U22091 ( .A(n42144), .B(n20457), .Z(n20421) );
  AND U22092 ( .A(n20422), .B(n20421), .Z(n20472) );
  XOR U22093 ( .A(a[440]), .B(n42012), .Z(n20460) );
  XNOR U22094 ( .A(n20472), .B(n20471), .Z(n20474) );
  XOR U22095 ( .A(a[438]), .B(n42085), .Z(n20464) );
  AND U22096 ( .A(a[434]), .B(b[7]), .Z(n20465) );
  XNOR U22097 ( .A(n20466), .B(n20465), .Z(n20467) );
  AND U22098 ( .A(a[442]), .B(b[0]), .Z(n20425) );
  XNOR U22099 ( .A(n20425), .B(n4071), .Z(n20427) );
  NANDN U22100 ( .A(b[0]), .B(a[441]), .Z(n20426) );
  NAND U22101 ( .A(n20427), .B(n20426), .Z(n20468) );
  XNOR U22102 ( .A(n20467), .B(n20468), .Z(n20473) );
  XOR U22103 ( .A(n20474), .B(n20473), .Z(n20452) );
  NANDN U22104 ( .A(n20429), .B(n20428), .Z(n20433) );
  NANDN U22105 ( .A(n20431), .B(n20430), .Z(n20432) );
  AND U22106 ( .A(n20433), .B(n20432), .Z(n20451) );
  XNOR U22107 ( .A(n20452), .B(n20451), .Z(n20453) );
  NANDN U22108 ( .A(n20435), .B(n20434), .Z(n20439) );
  NAND U22109 ( .A(n20437), .B(n20436), .Z(n20438) );
  NAND U22110 ( .A(n20439), .B(n20438), .Z(n20454) );
  XNOR U22111 ( .A(n20453), .B(n20454), .Z(n20445) );
  XNOR U22112 ( .A(n20446), .B(n20445), .Z(n20447) );
  XNOR U22113 ( .A(n20448), .B(n20447), .Z(n20477) );
  XNOR U22114 ( .A(sreg[1458]), .B(n20477), .Z(n20479) );
  NANDN U22115 ( .A(sreg[1457]), .B(n20440), .Z(n20444) );
  NAND U22116 ( .A(n20442), .B(n20441), .Z(n20443) );
  NAND U22117 ( .A(n20444), .B(n20443), .Z(n20478) );
  XNOR U22118 ( .A(n20479), .B(n20478), .Z(c[1458]) );
  NANDN U22119 ( .A(n20446), .B(n20445), .Z(n20450) );
  NANDN U22120 ( .A(n20448), .B(n20447), .Z(n20449) );
  AND U22121 ( .A(n20450), .B(n20449), .Z(n20485) );
  NANDN U22122 ( .A(n20452), .B(n20451), .Z(n20456) );
  NANDN U22123 ( .A(n20454), .B(n20453), .Z(n20455) );
  AND U22124 ( .A(n20456), .B(n20455), .Z(n20483) );
  NAND U22125 ( .A(n42143), .B(n20457), .Z(n20459) );
  XNOR U22126 ( .A(a[437]), .B(n4134), .Z(n20494) );
  NAND U22127 ( .A(n42144), .B(n20494), .Z(n20458) );
  AND U22128 ( .A(n20459), .B(n20458), .Z(n20509) );
  XOR U22129 ( .A(a[441]), .B(n42012), .Z(n20497) );
  XNOR U22130 ( .A(n20509), .B(n20508), .Z(n20511) );
  AND U22131 ( .A(a[443]), .B(b[0]), .Z(n20461) );
  XNOR U22132 ( .A(n20461), .B(n4071), .Z(n20463) );
  NANDN U22133 ( .A(b[0]), .B(a[442]), .Z(n20462) );
  NAND U22134 ( .A(n20463), .B(n20462), .Z(n20505) );
  XOR U22135 ( .A(a[439]), .B(n42085), .Z(n20501) );
  AND U22136 ( .A(a[435]), .B(b[7]), .Z(n20502) );
  XNOR U22137 ( .A(n20503), .B(n20502), .Z(n20504) );
  XNOR U22138 ( .A(n20505), .B(n20504), .Z(n20510) );
  XOR U22139 ( .A(n20511), .B(n20510), .Z(n20489) );
  NANDN U22140 ( .A(n20466), .B(n20465), .Z(n20470) );
  NANDN U22141 ( .A(n20468), .B(n20467), .Z(n20469) );
  AND U22142 ( .A(n20470), .B(n20469), .Z(n20488) );
  XNOR U22143 ( .A(n20489), .B(n20488), .Z(n20490) );
  NANDN U22144 ( .A(n20472), .B(n20471), .Z(n20476) );
  NAND U22145 ( .A(n20474), .B(n20473), .Z(n20475) );
  NAND U22146 ( .A(n20476), .B(n20475), .Z(n20491) );
  XNOR U22147 ( .A(n20490), .B(n20491), .Z(n20482) );
  XNOR U22148 ( .A(n20483), .B(n20482), .Z(n20484) );
  XNOR U22149 ( .A(n20485), .B(n20484), .Z(n20514) );
  XNOR U22150 ( .A(sreg[1459]), .B(n20514), .Z(n20516) );
  NANDN U22151 ( .A(sreg[1458]), .B(n20477), .Z(n20481) );
  NAND U22152 ( .A(n20479), .B(n20478), .Z(n20480) );
  NAND U22153 ( .A(n20481), .B(n20480), .Z(n20515) );
  XNOR U22154 ( .A(n20516), .B(n20515), .Z(c[1459]) );
  NANDN U22155 ( .A(n20483), .B(n20482), .Z(n20487) );
  NANDN U22156 ( .A(n20485), .B(n20484), .Z(n20486) );
  AND U22157 ( .A(n20487), .B(n20486), .Z(n20522) );
  NANDN U22158 ( .A(n20489), .B(n20488), .Z(n20493) );
  NANDN U22159 ( .A(n20491), .B(n20490), .Z(n20492) );
  AND U22160 ( .A(n20493), .B(n20492), .Z(n20520) );
  NAND U22161 ( .A(n42143), .B(n20494), .Z(n20496) );
  XNOR U22162 ( .A(a[438]), .B(n4134), .Z(n20531) );
  NAND U22163 ( .A(n42144), .B(n20531), .Z(n20495) );
  AND U22164 ( .A(n20496), .B(n20495), .Z(n20546) );
  XOR U22165 ( .A(a[442]), .B(n42012), .Z(n20534) );
  XNOR U22166 ( .A(n20546), .B(n20545), .Z(n20548) );
  AND U22167 ( .A(a[444]), .B(b[0]), .Z(n20498) );
  XNOR U22168 ( .A(n20498), .B(n4071), .Z(n20500) );
  NANDN U22169 ( .A(b[0]), .B(a[443]), .Z(n20499) );
  NAND U22170 ( .A(n20500), .B(n20499), .Z(n20542) );
  XOR U22171 ( .A(a[440]), .B(n42085), .Z(n20538) );
  AND U22172 ( .A(a[436]), .B(b[7]), .Z(n20539) );
  XNOR U22173 ( .A(n20540), .B(n20539), .Z(n20541) );
  XNOR U22174 ( .A(n20542), .B(n20541), .Z(n20547) );
  XOR U22175 ( .A(n20548), .B(n20547), .Z(n20526) );
  NANDN U22176 ( .A(n20503), .B(n20502), .Z(n20507) );
  NANDN U22177 ( .A(n20505), .B(n20504), .Z(n20506) );
  AND U22178 ( .A(n20507), .B(n20506), .Z(n20525) );
  XNOR U22179 ( .A(n20526), .B(n20525), .Z(n20527) );
  NANDN U22180 ( .A(n20509), .B(n20508), .Z(n20513) );
  NAND U22181 ( .A(n20511), .B(n20510), .Z(n20512) );
  NAND U22182 ( .A(n20513), .B(n20512), .Z(n20528) );
  XNOR U22183 ( .A(n20527), .B(n20528), .Z(n20519) );
  XNOR U22184 ( .A(n20520), .B(n20519), .Z(n20521) );
  XNOR U22185 ( .A(n20522), .B(n20521), .Z(n20551) );
  XNOR U22186 ( .A(sreg[1460]), .B(n20551), .Z(n20553) );
  NANDN U22187 ( .A(sreg[1459]), .B(n20514), .Z(n20518) );
  NAND U22188 ( .A(n20516), .B(n20515), .Z(n20517) );
  NAND U22189 ( .A(n20518), .B(n20517), .Z(n20552) );
  XNOR U22190 ( .A(n20553), .B(n20552), .Z(c[1460]) );
  NANDN U22191 ( .A(n20520), .B(n20519), .Z(n20524) );
  NANDN U22192 ( .A(n20522), .B(n20521), .Z(n20523) );
  AND U22193 ( .A(n20524), .B(n20523), .Z(n20559) );
  NANDN U22194 ( .A(n20526), .B(n20525), .Z(n20530) );
  NANDN U22195 ( .A(n20528), .B(n20527), .Z(n20529) );
  AND U22196 ( .A(n20530), .B(n20529), .Z(n20557) );
  NAND U22197 ( .A(n42143), .B(n20531), .Z(n20533) );
  XNOR U22198 ( .A(a[439]), .B(n4134), .Z(n20568) );
  NAND U22199 ( .A(n42144), .B(n20568), .Z(n20532) );
  AND U22200 ( .A(n20533), .B(n20532), .Z(n20583) );
  XOR U22201 ( .A(a[443]), .B(n42012), .Z(n20571) );
  XNOR U22202 ( .A(n20583), .B(n20582), .Z(n20585) );
  AND U22203 ( .A(a[445]), .B(b[0]), .Z(n20535) );
  XNOR U22204 ( .A(n20535), .B(n4071), .Z(n20537) );
  NANDN U22205 ( .A(b[0]), .B(a[444]), .Z(n20536) );
  NAND U22206 ( .A(n20537), .B(n20536), .Z(n20579) );
  XOR U22207 ( .A(a[441]), .B(n42085), .Z(n20572) );
  AND U22208 ( .A(a[437]), .B(b[7]), .Z(n20576) );
  XNOR U22209 ( .A(n20577), .B(n20576), .Z(n20578) );
  XNOR U22210 ( .A(n20579), .B(n20578), .Z(n20584) );
  XOR U22211 ( .A(n20585), .B(n20584), .Z(n20563) );
  NANDN U22212 ( .A(n20540), .B(n20539), .Z(n20544) );
  NANDN U22213 ( .A(n20542), .B(n20541), .Z(n20543) );
  AND U22214 ( .A(n20544), .B(n20543), .Z(n20562) );
  XNOR U22215 ( .A(n20563), .B(n20562), .Z(n20564) );
  NANDN U22216 ( .A(n20546), .B(n20545), .Z(n20550) );
  NAND U22217 ( .A(n20548), .B(n20547), .Z(n20549) );
  NAND U22218 ( .A(n20550), .B(n20549), .Z(n20565) );
  XNOR U22219 ( .A(n20564), .B(n20565), .Z(n20556) );
  XNOR U22220 ( .A(n20557), .B(n20556), .Z(n20558) );
  XNOR U22221 ( .A(n20559), .B(n20558), .Z(n20588) );
  XNOR U22222 ( .A(sreg[1461]), .B(n20588), .Z(n20590) );
  NANDN U22223 ( .A(sreg[1460]), .B(n20551), .Z(n20555) );
  NAND U22224 ( .A(n20553), .B(n20552), .Z(n20554) );
  NAND U22225 ( .A(n20555), .B(n20554), .Z(n20589) );
  XNOR U22226 ( .A(n20590), .B(n20589), .Z(c[1461]) );
  NANDN U22227 ( .A(n20557), .B(n20556), .Z(n20561) );
  NANDN U22228 ( .A(n20559), .B(n20558), .Z(n20560) );
  AND U22229 ( .A(n20561), .B(n20560), .Z(n20596) );
  NANDN U22230 ( .A(n20563), .B(n20562), .Z(n20567) );
  NANDN U22231 ( .A(n20565), .B(n20564), .Z(n20566) );
  AND U22232 ( .A(n20567), .B(n20566), .Z(n20594) );
  NAND U22233 ( .A(n42143), .B(n20568), .Z(n20570) );
  XNOR U22234 ( .A(a[440]), .B(n4134), .Z(n20605) );
  NAND U22235 ( .A(n42144), .B(n20605), .Z(n20569) );
  AND U22236 ( .A(n20570), .B(n20569), .Z(n20620) );
  XOR U22237 ( .A(a[444]), .B(n42012), .Z(n20608) );
  XNOR U22238 ( .A(n20620), .B(n20619), .Z(n20622) );
  XOR U22239 ( .A(a[442]), .B(n42085), .Z(n20612) );
  AND U22240 ( .A(a[438]), .B(b[7]), .Z(n20613) );
  XNOR U22241 ( .A(n20614), .B(n20613), .Z(n20615) );
  AND U22242 ( .A(a[446]), .B(b[0]), .Z(n20573) );
  XNOR U22243 ( .A(n20573), .B(n4071), .Z(n20575) );
  NANDN U22244 ( .A(b[0]), .B(a[445]), .Z(n20574) );
  NAND U22245 ( .A(n20575), .B(n20574), .Z(n20616) );
  XNOR U22246 ( .A(n20615), .B(n20616), .Z(n20621) );
  XOR U22247 ( .A(n20622), .B(n20621), .Z(n20600) );
  NANDN U22248 ( .A(n20577), .B(n20576), .Z(n20581) );
  NANDN U22249 ( .A(n20579), .B(n20578), .Z(n20580) );
  AND U22250 ( .A(n20581), .B(n20580), .Z(n20599) );
  XNOR U22251 ( .A(n20600), .B(n20599), .Z(n20601) );
  NANDN U22252 ( .A(n20583), .B(n20582), .Z(n20587) );
  NAND U22253 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U22254 ( .A(n20587), .B(n20586), .Z(n20602) );
  XNOR U22255 ( .A(n20601), .B(n20602), .Z(n20593) );
  XNOR U22256 ( .A(n20594), .B(n20593), .Z(n20595) );
  XNOR U22257 ( .A(n20596), .B(n20595), .Z(n20625) );
  XNOR U22258 ( .A(sreg[1462]), .B(n20625), .Z(n20627) );
  NANDN U22259 ( .A(sreg[1461]), .B(n20588), .Z(n20592) );
  NAND U22260 ( .A(n20590), .B(n20589), .Z(n20591) );
  NAND U22261 ( .A(n20592), .B(n20591), .Z(n20626) );
  XNOR U22262 ( .A(n20627), .B(n20626), .Z(c[1462]) );
  NANDN U22263 ( .A(n20594), .B(n20593), .Z(n20598) );
  NANDN U22264 ( .A(n20596), .B(n20595), .Z(n20597) );
  AND U22265 ( .A(n20598), .B(n20597), .Z(n20633) );
  NANDN U22266 ( .A(n20600), .B(n20599), .Z(n20604) );
  NANDN U22267 ( .A(n20602), .B(n20601), .Z(n20603) );
  AND U22268 ( .A(n20604), .B(n20603), .Z(n20631) );
  NAND U22269 ( .A(n42143), .B(n20605), .Z(n20607) );
  XNOR U22270 ( .A(a[441]), .B(n4134), .Z(n20642) );
  NAND U22271 ( .A(n42144), .B(n20642), .Z(n20606) );
  AND U22272 ( .A(n20607), .B(n20606), .Z(n20657) );
  XOR U22273 ( .A(a[445]), .B(n42012), .Z(n20645) );
  XNOR U22274 ( .A(n20657), .B(n20656), .Z(n20659) );
  AND U22275 ( .A(a[447]), .B(b[0]), .Z(n20609) );
  XNOR U22276 ( .A(n20609), .B(n4071), .Z(n20611) );
  NANDN U22277 ( .A(b[0]), .B(a[446]), .Z(n20610) );
  NAND U22278 ( .A(n20611), .B(n20610), .Z(n20653) );
  XOR U22279 ( .A(a[443]), .B(n42085), .Z(n20649) );
  AND U22280 ( .A(a[439]), .B(b[7]), .Z(n20650) );
  XNOR U22281 ( .A(n20651), .B(n20650), .Z(n20652) );
  XNOR U22282 ( .A(n20653), .B(n20652), .Z(n20658) );
  XOR U22283 ( .A(n20659), .B(n20658), .Z(n20637) );
  NANDN U22284 ( .A(n20614), .B(n20613), .Z(n20618) );
  NANDN U22285 ( .A(n20616), .B(n20615), .Z(n20617) );
  AND U22286 ( .A(n20618), .B(n20617), .Z(n20636) );
  XNOR U22287 ( .A(n20637), .B(n20636), .Z(n20638) );
  NANDN U22288 ( .A(n20620), .B(n20619), .Z(n20624) );
  NAND U22289 ( .A(n20622), .B(n20621), .Z(n20623) );
  NAND U22290 ( .A(n20624), .B(n20623), .Z(n20639) );
  XNOR U22291 ( .A(n20638), .B(n20639), .Z(n20630) );
  XNOR U22292 ( .A(n20631), .B(n20630), .Z(n20632) );
  XNOR U22293 ( .A(n20633), .B(n20632), .Z(n20662) );
  XNOR U22294 ( .A(sreg[1463]), .B(n20662), .Z(n20664) );
  NANDN U22295 ( .A(sreg[1462]), .B(n20625), .Z(n20629) );
  NAND U22296 ( .A(n20627), .B(n20626), .Z(n20628) );
  NAND U22297 ( .A(n20629), .B(n20628), .Z(n20663) );
  XNOR U22298 ( .A(n20664), .B(n20663), .Z(c[1463]) );
  NANDN U22299 ( .A(n20631), .B(n20630), .Z(n20635) );
  NANDN U22300 ( .A(n20633), .B(n20632), .Z(n20634) );
  AND U22301 ( .A(n20635), .B(n20634), .Z(n20670) );
  NANDN U22302 ( .A(n20637), .B(n20636), .Z(n20641) );
  NANDN U22303 ( .A(n20639), .B(n20638), .Z(n20640) );
  AND U22304 ( .A(n20641), .B(n20640), .Z(n20668) );
  NAND U22305 ( .A(n42143), .B(n20642), .Z(n20644) );
  XNOR U22306 ( .A(a[442]), .B(n4135), .Z(n20679) );
  NAND U22307 ( .A(n42144), .B(n20679), .Z(n20643) );
  AND U22308 ( .A(n20644), .B(n20643), .Z(n20694) );
  XOR U22309 ( .A(a[446]), .B(n42012), .Z(n20682) );
  XNOR U22310 ( .A(n20694), .B(n20693), .Z(n20696) );
  AND U22311 ( .A(a[448]), .B(b[0]), .Z(n20646) );
  XNOR U22312 ( .A(n20646), .B(n4071), .Z(n20648) );
  NANDN U22313 ( .A(b[0]), .B(a[447]), .Z(n20647) );
  NAND U22314 ( .A(n20648), .B(n20647), .Z(n20690) );
  XOR U22315 ( .A(a[444]), .B(n42085), .Z(n20686) );
  AND U22316 ( .A(a[440]), .B(b[7]), .Z(n20687) );
  XNOR U22317 ( .A(n20688), .B(n20687), .Z(n20689) );
  XNOR U22318 ( .A(n20690), .B(n20689), .Z(n20695) );
  XOR U22319 ( .A(n20696), .B(n20695), .Z(n20674) );
  NANDN U22320 ( .A(n20651), .B(n20650), .Z(n20655) );
  NANDN U22321 ( .A(n20653), .B(n20652), .Z(n20654) );
  AND U22322 ( .A(n20655), .B(n20654), .Z(n20673) );
  XNOR U22323 ( .A(n20674), .B(n20673), .Z(n20675) );
  NANDN U22324 ( .A(n20657), .B(n20656), .Z(n20661) );
  NAND U22325 ( .A(n20659), .B(n20658), .Z(n20660) );
  NAND U22326 ( .A(n20661), .B(n20660), .Z(n20676) );
  XNOR U22327 ( .A(n20675), .B(n20676), .Z(n20667) );
  XNOR U22328 ( .A(n20668), .B(n20667), .Z(n20669) );
  XNOR U22329 ( .A(n20670), .B(n20669), .Z(n20699) );
  XNOR U22330 ( .A(sreg[1464]), .B(n20699), .Z(n20701) );
  NANDN U22331 ( .A(sreg[1463]), .B(n20662), .Z(n20666) );
  NAND U22332 ( .A(n20664), .B(n20663), .Z(n20665) );
  NAND U22333 ( .A(n20666), .B(n20665), .Z(n20700) );
  XNOR U22334 ( .A(n20701), .B(n20700), .Z(c[1464]) );
  NANDN U22335 ( .A(n20668), .B(n20667), .Z(n20672) );
  NANDN U22336 ( .A(n20670), .B(n20669), .Z(n20671) );
  AND U22337 ( .A(n20672), .B(n20671), .Z(n20707) );
  NANDN U22338 ( .A(n20674), .B(n20673), .Z(n20678) );
  NANDN U22339 ( .A(n20676), .B(n20675), .Z(n20677) );
  AND U22340 ( .A(n20678), .B(n20677), .Z(n20705) );
  NAND U22341 ( .A(n42143), .B(n20679), .Z(n20681) );
  XNOR U22342 ( .A(a[443]), .B(n4135), .Z(n20716) );
  NAND U22343 ( .A(n42144), .B(n20716), .Z(n20680) );
  AND U22344 ( .A(n20681), .B(n20680), .Z(n20731) );
  XOR U22345 ( .A(a[447]), .B(n42012), .Z(n20719) );
  XNOR U22346 ( .A(n20731), .B(n20730), .Z(n20733) );
  AND U22347 ( .A(a[449]), .B(b[0]), .Z(n20683) );
  XNOR U22348 ( .A(n20683), .B(n4071), .Z(n20685) );
  NANDN U22349 ( .A(b[0]), .B(a[448]), .Z(n20684) );
  NAND U22350 ( .A(n20685), .B(n20684), .Z(n20727) );
  XOR U22351 ( .A(a[445]), .B(n42085), .Z(n20723) );
  AND U22352 ( .A(a[441]), .B(b[7]), .Z(n20724) );
  XNOR U22353 ( .A(n20725), .B(n20724), .Z(n20726) );
  XNOR U22354 ( .A(n20727), .B(n20726), .Z(n20732) );
  XOR U22355 ( .A(n20733), .B(n20732), .Z(n20711) );
  NANDN U22356 ( .A(n20688), .B(n20687), .Z(n20692) );
  NANDN U22357 ( .A(n20690), .B(n20689), .Z(n20691) );
  AND U22358 ( .A(n20692), .B(n20691), .Z(n20710) );
  XNOR U22359 ( .A(n20711), .B(n20710), .Z(n20712) );
  NANDN U22360 ( .A(n20694), .B(n20693), .Z(n20698) );
  NAND U22361 ( .A(n20696), .B(n20695), .Z(n20697) );
  NAND U22362 ( .A(n20698), .B(n20697), .Z(n20713) );
  XNOR U22363 ( .A(n20712), .B(n20713), .Z(n20704) );
  XNOR U22364 ( .A(n20705), .B(n20704), .Z(n20706) );
  XNOR U22365 ( .A(n20707), .B(n20706), .Z(n20736) );
  XNOR U22366 ( .A(sreg[1465]), .B(n20736), .Z(n20738) );
  NANDN U22367 ( .A(sreg[1464]), .B(n20699), .Z(n20703) );
  NAND U22368 ( .A(n20701), .B(n20700), .Z(n20702) );
  NAND U22369 ( .A(n20703), .B(n20702), .Z(n20737) );
  XNOR U22370 ( .A(n20738), .B(n20737), .Z(c[1465]) );
  NANDN U22371 ( .A(n20705), .B(n20704), .Z(n20709) );
  NANDN U22372 ( .A(n20707), .B(n20706), .Z(n20708) );
  AND U22373 ( .A(n20709), .B(n20708), .Z(n20744) );
  NANDN U22374 ( .A(n20711), .B(n20710), .Z(n20715) );
  NANDN U22375 ( .A(n20713), .B(n20712), .Z(n20714) );
  AND U22376 ( .A(n20715), .B(n20714), .Z(n20742) );
  NAND U22377 ( .A(n42143), .B(n20716), .Z(n20718) );
  XNOR U22378 ( .A(a[444]), .B(n4135), .Z(n20753) );
  NAND U22379 ( .A(n42144), .B(n20753), .Z(n20717) );
  AND U22380 ( .A(n20718), .B(n20717), .Z(n20768) );
  XOR U22381 ( .A(a[448]), .B(n42012), .Z(n20756) );
  XNOR U22382 ( .A(n20768), .B(n20767), .Z(n20770) );
  AND U22383 ( .A(a[450]), .B(b[0]), .Z(n20720) );
  XNOR U22384 ( .A(n20720), .B(n4071), .Z(n20722) );
  NANDN U22385 ( .A(b[0]), .B(a[449]), .Z(n20721) );
  NAND U22386 ( .A(n20722), .B(n20721), .Z(n20764) );
  XOR U22387 ( .A(a[446]), .B(n42085), .Z(n20760) );
  AND U22388 ( .A(a[442]), .B(b[7]), .Z(n20761) );
  XNOR U22389 ( .A(n20762), .B(n20761), .Z(n20763) );
  XNOR U22390 ( .A(n20764), .B(n20763), .Z(n20769) );
  XOR U22391 ( .A(n20770), .B(n20769), .Z(n20748) );
  NANDN U22392 ( .A(n20725), .B(n20724), .Z(n20729) );
  NANDN U22393 ( .A(n20727), .B(n20726), .Z(n20728) );
  AND U22394 ( .A(n20729), .B(n20728), .Z(n20747) );
  XNOR U22395 ( .A(n20748), .B(n20747), .Z(n20749) );
  NANDN U22396 ( .A(n20731), .B(n20730), .Z(n20735) );
  NAND U22397 ( .A(n20733), .B(n20732), .Z(n20734) );
  NAND U22398 ( .A(n20735), .B(n20734), .Z(n20750) );
  XNOR U22399 ( .A(n20749), .B(n20750), .Z(n20741) );
  XNOR U22400 ( .A(n20742), .B(n20741), .Z(n20743) );
  XNOR U22401 ( .A(n20744), .B(n20743), .Z(n20773) );
  XNOR U22402 ( .A(sreg[1466]), .B(n20773), .Z(n20775) );
  NANDN U22403 ( .A(sreg[1465]), .B(n20736), .Z(n20740) );
  NAND U22404 ( .A(n20738), .B(n20737), .Z(n20739) );
  NAND U22405 ( .A(n20740), .B(n20739), .Z(n20774) );
  XNOR U22406 ( .A(n20775), .B(n20774), .Z(c[1466]) );
  NANDN U22407 ( .A(n20742), .B(n20741), .Z(n20746) );
  NANDN U22408 ( .A(n20744), .B(n20743), .Z(n20745) );
  AND U22409 ( .A(n20746), .B(n20745), .Z(n20781) );
  NANDN U22410 ( .A(n20748), .B(n20747), .Z(n20752) );
  NANDN U22411 ( .A(n20750), .B(n20749), .Z(n20751) );
  AND U22412 ( .A(n20752), .B(n20751), .Z(n20779) );
  NAND U22413 ( .A(n42143), .B(n20753), .Z(n20755) );
  XNOR U22414 ( .A(a[445]), .B(n4135), .Z(n20790) );
  NAND U22415 ( .A(n42144), .B(n20790), .Z(n20754) );
  AND U22416 ( .A(n20755), .B(n20754), .Z(n20805) );
  XOR U22417 ( .A(a[449]), .B(n42012), .Z(n20793) );
  XNOR U22418 ( .A(n20805), .B(n20804), .Z(n20807) );
  AND U22419 ( .A(a[451]), .B(b[0]), .Z(n20757) );
  XNOR U22420 ( .A(n20757), .B(n4071), .Z(n20759) );
  NANDN U22421 ( .A(b[0]), .B(a[450]), .Z(n20758) );
  NAND U22422 ( .A(n20759), .B(n20758), .Z(n20801) );
  XOR U22423 ( .A(a[447]), .B(n42085), .Z(n20797) );
  AND U22424 ( .A(a[443]), .B(b[7]), .Z(n20798) );
  XNOR U22425 ( .A(n20799), .B(n20798), .Z(n20800) );
  XNOR U22426 ( .A(n20801), .B(n20800), .Z(n20806) );
  XOR U22427 ( .A(n20807), .B(n20806), .Z(n20785) );
  NANDN U22428 ( .A(n20762), .B(n20761), .Z(n20766) );
  NANDN U22429 ( .A(n20764), .B(n20763), .Z(n20765) );
  AND U22430 ( .A(n20766), .B(n20765), .Z(n20784) );
  XNOR U22431 ( .A(n20785), .B(n20784), .Z(n20786) );
  NANDN U22432 ( .A(n20768), .B(n20767), .Z(n20772) );
  NAND U22433 ( .A(n20770), .B(n20769), .Z(n20771) );
  NAND U22434 ( .A(n20772), .B(n20771), .Z(n20787) );
  XNOR U22435 ( .A(n20786), .B(n20787), .Z(n20778) );
  XNOR U22436 ( .A(n20779), .B(n20778), .Z(n20780) );
  XNOR U22437 ( .A(n20781), .B(n20780), .Z(n20810) );
  XNOR U22438 ( .A(sreg[1467]), .B(n20810), .Z(n20812) );
  NANDN U22439 ( .A(sreg[1466]), .B(n20773), .Z(n20777) );
  NAND U22440 ( .A(n20775), .B(n20774), .Z(n20776) );
  NAND U22441 ( .A(n20777), .B(n20776), .Z(n20811) );
  XNOR U22442 ( .A(n20812), .B(n20811), .Z(c[1467]) );
  NANDN U22443 ( .A(n20779), .B(n20778), .Z(n20783) );
  NANDN U22444 ( .A(n20781), .B(n20780), .Z(n20782) );
  AND U22445 ( .A(n20783), .B(n20782), .Z(n20818) );
  NANDN U22446 ( .A(n20785), .B(n20784), .Z(n20789) );
  NANDN U22447 ( .A(n20787), .B(n20786), .Z(n20788) );
  AND U22448 ( .A(n20789), .B(n20788), .Z(n20816) );
  NAND U22449 ( .A(n42143), .B(n20790), .Z(n20792) );
  XNOR U22450 ( .A(a[446]), .B(n4135), .Z(n20827) );
  NAND U22451 ( .A(n42144), .B(n20827), .Z(n20791) );
  AND U22452 ( .A(n20792), .B(n20791), .Z(n20842) );
  XOR U22453 ( .A(a[450]), .B(n42012), .Z(n20830) );
  XNOR U22454 ( .A(n20842), .B(n20841), .Z(n20844) );
  AND U22455 ( .A(a[452]), .B(b[0]), .Z(n20794) );
  XNOR U22456 ( .A(n20794), .B(n4071), .Z(n20796) );
  NANDN U22457 ( .A(b[0]), .B(a[451]), .Z(n20795) );
  NAND U22458 ( .A(n20796), .B(n20795), .Z(n20838) );
  XOR U22459 ( .A(a[448]), .B(n42085), .Z(n20834) );
  AND U22460 ( .A(a[444]), .B(b[7]), .Z(n20835) );
  XNOR U22461 ( .A(n20836), .B(n20835), .Z(n20837) );
  XNOR U22462 ( .A(n20838), .B(n20837), .Z(n20843) );
  XOR U22463 ( .A(n20844), .B(n20843), .Z(n20822) );
  NANDN U22464 ( .A(n20799), .B(n20798), .Z(n20803) );
  NANDN U22465 ( .A(n20801), .B(n20800), .Z(n20802) );
  AND U22466 ( .A(n20803), .B(n20802), .Z(n20821) );
  XNOR U22467 ( .A(n20822), .B(n20821), .Z(n20823) );
  NANDN U22468 ( .A(n20805), .B(n20804), .Z(n20809) );
  NAND U22469 ( .A(n20807), .B(n20806), .Z(n20808) );
  NAND U22470 ( .A(n20809), .B(n20808), .Z(n20824) );
  XNOR U22471 ( .A(n20823), .B(n20824), .Z(n20815) );
  XNOR U22472 ( .A(n20816), .B(n20815), .Z(n20817) );
  XNOR U22473 ( .A(n20818), .B(n20817), .Z(n20847) );
  XNOR U22474 ( .A(sreg[1468]), .B(n20847), .Z(n20849) );
  NANDN U22475 ( .A(sreg[1467]), .B(n20810), .Z(n20814) );
  NAND U22476 ( .A(n20812), .B(n20811), .Z(n20813) );
  NAND U22477 ( .A(n20814), .B(n20813), .Z(n20848) );
  XNOR U22478 ( .A(n20849), .B(n20848), .Z(c[1468]) );
  NANDN U22479 ( .A(n20816), .B(n20815), .Z(n20820) );
  NANDN U22480 ( .A(n20818), .B(n20817), .Z(n20819) );
  AND U22481 ( .A(n20820), .B(n20819), .Z(n20855) );
  NANDN U22482 ( .A(n20822), .B(n20821), .Z(n20826) );
  NANDN U22483 ( .A(n20824), .B(n20823), .Z(n20825) );
  AND U22484 ( .A(n20826), .B(n20825), .Z(n20853) );
  NAND U22485 ( .A(n42143), .B(n20827), .Z(n20829) );
  XNOR U22486 ( .A(a[447]), .B(n4135), .Z(n20864) );
  NAND U22487 ( .A(n42144), .B(n20864), .Z(n20828) );
  AND U22488 ( .A(n20829), .B(n20828), .Z(n20879) );
  XOR U22489 ( .A(a[451]), .B(n42012), .Z(n20867) );
  XNOR U22490 ( .A(n20879), .B(n20878), .Z(n20881) );
  AND U22491 ( .A(a[453]), .B(b[0]), .Z(n20831) );
  XNOR U22492 ( .A(n20831), .B(n4071), .Z(n20833) );
  NANDN U22493 ( .A(b[0]), .B(a[452]), .Z(n20832) );
  NAND U22494 ( .A(n20833), .B(n20832), .Z(n20875) );
  XOR U22495 ( .A(a[449]), .B(n42085), .Z(n20871) );
  AND U22496 ( .A(a[445]), .B(b[7]), .Z(n20872) );
  XNOR U22497 ( .A(n20873), .B(n20872), .Z(n20874) );
  XNOR U22498 ( .A(n20875), .B(n20874), .Z(n20880) );
  XOR U22499 ( .A(n20881), .B(n20880), .Z(n20859) );
  NANDN U22500 ( .A(n20836), .B(n20835), .Z(n20840) );
  NANDN U22501 ( .A(n20838), .B(n20837), .Z(n20839) );
  AND U22502 ( .A(n20840), .B(n20839), .Z(n20858) );
  XNOR U22503 ( .A(n20859), .B(n20858), .Z(n20860) );
  NANDN U22504 ( .A(n20842), .B(n20841), .Z(n20846) );
  NAND U22505 ( .A(n20844), .B(n20843), .Z(n20845) );
  NAND U22506 ( .A(n20846), .B(n20845), .Z(n20861) );
  XNOR U22507 ( .A(n20860), .B(n20861), .Z(n20852) );
  XNOR U22508 ( .A(n20853), .B(n20852), .Z(n20854) );
  XNOR U22509 ( .A(n20855), .B(n20854), .Z(n20884) );
  XNOR U22510 ( .A(sreg[1469]), .B(n20884), .Z(n20886) );
  NANDN U22511 ( .A(sreg[1468]), .B(n20847), .Z(n20851) );
  NAND U22512 ( .A(n20849), .B(n20848), .Z(n20850) );
  NAND U22513 ( .A(n20851), .B(n20850), .Z(n20885) );
  XNOR U22514 ( .A(n20886), .B(n20885), .Z(c[1469]) );
  NANDN U22515 ( .A(n20853), .B(n20852), .Z(n20857) );
  NANDN U22516 ( .A(n20855), .B(n20854), .Z(n20856) );
  AND U22517 ( .A(n20857), .B(n20856), .Z(n20892) );
  NANDN U22518 ( .A(n20859), .B(n20858), .Z(n20863) );
  NANDN U22519 ( .A(n20861), .B(n20860), .Z(n20862) );
  AND U22520 ( .A(n20863), .B(n20862), .Z(n20890) );
  NAND U22521 ( .A(n42143), .B(n20864), .Z(n20866) );
  XNOR U22522 ( .A(a[448]), .B(n4135), .Z(n20901) );
  NAND U22523 ( .A(n42144), .B(n20901), .Z(n20865) );
  AND U22524 ( .A(n20866), .B(n20865), .Z(n20916) );
  XOR U22525 ( .A(a[452]), .B(n42012), .Z(n20904) );
  XNOR U22526 ( .A(n20916), .B(n20915), .Z(n20918) );
  AND U22527 ( .A(a[454]), .B(b[0]), .Z(n20868) );
  XNOR U22528 ( .A(n20868), .B(n4071), .Z(n20870) );
  NANDN U22529 ( .A(b[0]), .B(a[453]), .Z(n20869) );
  NAND U22530 ( .A(n20870), .B(n20869), .Z(n20912) );
  XOR U22531 ( .A(a[450]), .B(n42085), .Z(n20908) );
  AND U22532 ( .A(a[446]), .B(b[7]), .Z(n20909) );
  XNOR U22533 ( .A(n20910), .B(n20909), .Z(n20911) );
  XNOR U22534 ( .A(n20912), .B(n20911), .Z(n20917) );
  XOR U22535 ( .A(n20918), .B(n20917), .Z(n20896) );
  NANDN U22536 ( .A(n20873), .B(n20872), .Z(n20877) );
  NANDN U22537 ( .A(n20875), .B(n20874), .Z(n20876) );
  AND U22538 ( .A(n20877), .B(n20876), .Z(n20895) );
  XNOR U22539 ( .A(n20896), .B(n20895), .Z(n20897) );
  NANDN U22540 ( .A(n20879), .B(n20878), .Z(n20883) );
  NAND U22541 ( .A(n20881), .B(n20880), .Z(n20882) );
  NAND U22542 ( .A(n20883), .B(n20882), .Z(n20898) );
  XNOR U22543 ( .A(n20897), .B(n20898), .Z(n20889) );
  XNOR U22544 ( .A(n20890), .B(n20889), .Z(n20891) );
  XNOR U22545 ( .A(n20892), .B(n20891), .Z(n20921) );
  XNOR U22546 ( .A(sreg[1470]), .B(n20921), .Z(n20923) );
  NANDN U22547 ( .A(sreg[1469]), .B(n20884), .Z(n20888) );
  NAND U22548 ( .A(n20886), .B(n20885), .Z(n20887) );
  NAND U22549 ( .A(n20888), .B(n20887), .Z(n20922) );
  XNOR U22550 ( .A(n20923), .B(n20922), .Z(c[1470]) );
  NANDN U22551 ( .A(n20890), .B(n20889), .Z(n20894) );
  NANDN U22552 ( .A(n20892), .B(n20891), .Z(n20893) );
  AND U22553 ( .A(n20894), .B(n20893), .Z(n20929) );
  NANDN U22554 ( .A(n20896), .B(n20895), .Z(n20900) );
  NANDN U22555 ( .A(n20898), .B(n20897), .Z(n20899) );
  AND U22556 ( .A(n20900), .B(n20899), .Z(n20927) );
  NAND U22557 ( .A(n42143), .B(n20901), .Z(n20903) );
  XNOR U22558 ( .A(a[449]), .B(n4136), .Z(n20938) );
  NAND U22559 ( .A(n42144), .B(n20938), .Z(n20902) );
  AND U22560 ( .A(n20903), .B(n20902), .Z(n20953) );
  XOR U22561 ( .A(a[453]), .B(n42012), .Z(n20941) );
  XNOR U22562 ( .A(n20953), .B(n20952), .Z(n20955) );
  AND U22563 ( .A(a[455]), .B(b[0]), .Z(n20905) );
  XNOR U22564 ( .A(n20905), .B(n4071), .Z(n20907) );
  NANDN U22565 ( .A(b[0]), .B(a[454]), .Z(n20906) );
  NAND U22566 ( .A(n20907), .B(n20906), .Z(n20949) );
  XOR U22567 ( .A(a[451]), .B(n42085), .Z(n20945) );
  AND U22568 ( .A(a[447]), .B(b[7]), .Z(n20946) );
  XNOR U22569 ( .A(n20947), .B(n20946), .Z(n20948) );
  XNOR U22570 ( .A(n20949), .B(n20948), .Z(n20954) );
  XOR U22571 ( .A(n20955), .B(n20954), .Z(n20933) );
  NANDN U22572 ( .A(n20910), .B(n20909), .Z(n20914) );
  NANDN U22573 ( .A(n20912), .B(n20911), .Z(n20913) );
  AND U22574 ( .A(n20914), .B(n20913), .Z(n20932) );
  XNOR U22575 ( .A(n20933), .B(n20932), .Z(n20934) );
  NANDN U22576 ( .A(n20916), .B(n20915), .Z(n20920) );
  NAND U22577 ( .A(n20918), .B(n20917), .Z(n20919) );
  NAND U22578 ( .A(n20920), .B(n20919), .Z(n20935) );
  XNOR U22579 ( .A(n20934), .B(n20935), .Z(n20926) );
  XNOR U22580 ( .A(n20927), .B(n20926), .Z(n20928) );
  XNOR U22581 ( .A(n20929), .B(n20928), .Z(n20958) );
  XNOR U22582 ( .A(sreg[1471]), .B(n20958), .Z(n20960) );
  NANDN U22583 ( .A(sreg[1470]), .B(n20921), .Z(n20925) );
  NAND U22584 ( .A(n20923), .B(n20922), .Z(n20924) );
  NAND U22585 ( .A(n20925), .B(n20924), .Z(n20959) );
  XNOR U22586 ( .A(n20960), .B(n20959), .Z(c[1471]) );
  NANDN U22587 ( .A(n20927), .B(n20926), .Z(n20931) );
  NANDN U22588 ( .A(n20929), .B(n20928), .Z(n20930) );
  AND U22589 ( .A(n20931), .B(n20930), .Z(n20966) );
  NANDN U22590 ( .A(n20933), .B(n20932), .Z(n20937) );
  NANDN U22591 ( .A(n20935), .B(n20934), .Z(n20936) );
  AND U22592 ( .A(n20937), .B(n20936), .Z(n20964) );
  NAND U22593 ( .A(n42143), .B(n20938), .Z(n20940) );
  XNOR U22594 ( .A(a[450]), .B(n4136), .Z(n20975) );
  NAND U22595 ( .A(n42144), .B(n20975), .Z(n20939) );
  AND U22596 ( .A(n20940), .B(n20939), .Z(n20990) );
  XOR U22597 ( .A(a[454]), .B(n42012), .Z(n20978) );
  XNOR U22598 ( .A(n20990), .B(n20989), .Z(n20992) );
  AND U22599 ( .A(a[456]), .B(b[0]), .Z(n20942) );
  XNOR U22600 ( .A(n20942), .B(n4071), .Z(n20944) );
  NANDN U22601 ( .A(b[0]), .B(a[455]), .Z(n20943) );
  NAND U22602 ( .A(n20944), .B(n20943), .Z(n20986) );
  XOR U22603 ( .A(a[452]), .B(n42085), .Z(n20982) );
  AND U22604 ( .A(a[448]), .B(b[7]), .Z(n20983) );
  XNOR U22605 ( .A(n20984), .B(n20983), .Z(n20985) );
  XNOR U22606 ( .A(n20986), .B(n20985), .Z(n20991) );
  XOR U22607 ( .A(n20992), .B(n20991), .Z(n20970) );
  NANDN U22608 ( .A(n20947), .B(n20946), .Z(n20951) );
  NANDN U22609 ( .A(n20949), .B(n20948), .Z(n20950) );
  AND U22610 ( .A(n20951), .B(n20950), .Z(n20969) );
  XNOR U22611 ( .A(n20970), .B(n20969), .Z(n20971) );
  NANDN U22612 ( .A(n20953), .B(n20952), .Z(n20957) );
  NAND U22613 ( .A(n20955), .B(n20954), .Z(n20956) );
  NAND U22614 ( .A(n20957), .B(n20956), .Z(n20972) );
  XNOR U22615 ( .A(n20971), .B(n20972), .Z(n20963) );
  XNOR U22616 ( .A(n20964), .B(n20963), .Z(n20965) );
  XNOR U22617 ( .A(n20966), .B(n20965), .Z(n20995) );
  XNOR U22618 ( .A(sreg[1472]), .B(n20995), .Z(n20997) );
  NANDN U22619 ( .A(sreg[1471]), .B(n20958), .Z(n20962) );
  NAND U22620 ( .A(n20960), .B(n20959), .Z(n20961) );
  NAND U22621 ( .A(n20962), .B(n20961), .Z(n20996) );
  XNOR U22622 ( .A(n20997), .B(n20996), .Z(c[1472]) );
  NANDN U22623 ( .A(n20964), .B(n20963), .Z(n20968) );
  NANDN U22624 ( .A(n20966), .B(n20965), .Z(n20967) );
  AND U22625 ( .A(n20968), .B(n20967), .Z(n21003) );
  NANDN U22626 ( .A(n20970), .B(n20969), .Z(n20974) );
  NANDN U22627 ( .A(n20972), .B(n20971), .Z(n20973) );
  AND U22628 ( .A(n20974), .B(n20973), .Z(n21001) );
  NAND U22629 ( .A(n42143), .B(n20975), .Z(n20977) );
  XNOR U22630 ( .A(a[451]), .B(n4136), .Z(n21012) );
  NAND U22631 ( .A(n42144), .B(n21012), .Z(n20976) );
  AND U22632 ( .A(n20977), .B(n20976), .Z(n21027) );
  XOR U22633 ( .A(a[455]), .B(n42012), .Z(n21015) );
  XNOR U22634 ( .A(n21027), .B(n21026), .Z(n21029) );
  AND U22635 ( .A(a[457]), .B(b[0]), .Z(n20979) );
  XNOR U22636 ( .A(n20979), .B(n4071), .Z(n20981) );
  NANDN U22637 ( .A(b[0]), .B(a[456]), .Z(n20980) );
  NAND U22638 ( .A(n20981), .B(n20980), .Z(n21023) );
  XOR U22639 ( .A(a[453]), .B(n42085), .Z(n21019) );
  AND U22640 ( .A(a[449]), .B(b[7]), .Z(n21020) );
  XNOR U22641 ( .A(n21021), .B(n21020), .Z(n21022) );
  XNOR U22642 ( .A(n21023), .B(n21022), .Z(n21028) );
  XOR U22643 ( .A(n21029), .B(n21028), .Z(n21007) );
  NANDN U22644 ( .A(n20984), .B(n20983), .Z(n20988) );
  NANDN U22645 ( .A(n20986), .B(n20985), .Z(n20987) );
  AND U22646 ( .A(n20988), .B(n20987), .Z(n21006) );
  XNOR U22647 ( .A(n21007), .B(n21006), .Z(n21008) );
  NANDN U22648 ( .A(n20990), .B(n20989), .Z(n20994) );
  NAND U22649 ( .A(n20992), .B(n20991), .Z(n20993) );
  NAND U22650 ( .A(n20994), .B(n20993), .Z(n21009) );
  XNOR U22651 ( .A(n21008), .B(n21009), .Z(n21000) );
  XNOR U22652 ( .A(n21001), .B(n21000), .Z(n21002) );
  XNOR U22653 ( .A(n21003), .B(n21002), .Z(n21032) );
  XNOR U22654 ( .A(sreg[1473]), .B(n21032), .Z(n21034) );
  NANDN U22655 ( .A(sreg[1472]), .B(n20995), .Z(n20999) );
  NAND U22656 ( .A(n20997), .B(n20996), .Z(n20998) );
  NAND U22657 ( .A(n20999), .B(n20998), .Z(n21033) );
  XNOR U22658 ( .A(n21034), .B(n21033), .Z(c[1473]) );
  NANDN U22659 ( .A(n21001), .B(n21000), .Z(n21005) );
  NANDN U22660 ( .A(n21003), .B(n21002), .Z(n21004) );
  AND U22661 ( .A(n21005), .B(n21004), .Z(n21040) );
  NANDN U22662 ( .A(n21007), .B(n21006), .Z(n21011) );
  NANDN U22663 ( .A(n21009), .B(n21008), .Z(n21010) );
  AND U22664 ( .A(n21011), .B(n21010), .Z(n21038) );
  NAND U22665 ( .A(n42143), .B(n21012), .Z(n21014) );
  XNOR U22666 ( .A(a[452]), .B(n4136), .Z(n21049) );
  NAND U22667 ( .A(n42144), .B(n21049), .Z(n21013) );
  AND U22668 ( .A(n21014), .B(n21013), .Z(n21064) );
  XOR U22669 ( .A(a[456]), .B(n42012), .Z(n21052) );
  XNOR U22670 ( .A(n21064), .B(n21063), .Z(n21066) );
  AND U22671 ( .A(a[458]), .B(b[0]), .Z(n21016) );
  XNOR U22672 ( .A(n21016), .B(n4071), .Z(n21018) );
  NANDN U22673 ( .A(b[0]), .B(a[457]), .Z(n21017) );
  NAND U22674 ( .A(n21018), .B(n21017), .Z(n21060) );
  XOR U22675 ( .A(a[454]), .B(n42085), .Z(n21053) );
  AND U22676 ( .A(a[450]), .B(b[7]), .Z(n21057) );
  XNOR U22677 ( .A(n21058), .B(n21057), .Z(n21059) );
  XNOR U22678 ( .A(n21060), .B(n21059), .Z(n21065) );
  XOR U22679 ( .A(n21066), .B(n21065), .Z(n21044) );
  NANDN U22680 ( .A(n21021), .B(n21020), .Z(n21025) );
  NANDN U22681 ( .A(n21023), .B(n21022), .Z(n21024) );
  AND U22682 ( .A(n21025), .B(n21024), .Z(n21043) );
  XNOR U22683 ( .A(n21044), .B(n21043), .Z(n21045) );
  NANDN U22684 ( .A(n21027), .B(n21026), .Z(n21031) );
  NAND U22685 ( .A(n21029), .B(n21028), .Z(n21030) );
  NAND U22686 ( .A(n21031), .B(n21030), .Z(n21046) );
  XNOR U22687 ( .A(n21045), .B(n21046), .Z(n21037) );
  XNOR U22688 ( .A(n21038), .B(n21037), .Z(n21039) );
  XNOR U22689 ( .A(n21040), .B(n21039), .Z(n21069) );
  XNOR U22690 ( .A(sreg[1474]), .B(n21069), .Z(n21071) );
  NANDN U22691 ( .A(sreg[1473]), .B(n21032), .Z(n21036) );
  NAND U22692 ( .A(n21034), .B(n21033), .Z(n21035) );
  NAND U22693 ( .A(n21036), .B(n21035), .Z(n21070) );
  XNOR U22694 ( .A(n21071), .B(n21070), .Z(c[1474]) );
  NANDN U22695 ( .A(n21038), .B(n21037), .Z(n21042) );
  NANDN U22696 ( .A(n21040), .B(n21039), .Z(n21041) );
  AND U22697 ( .A(n21042), .B(n21041), .Z(n21077) );
  NANDN U22698 ( .A(n21044), .B(n21043), .Z(n21048) );
  NANDN U22699 ( .A(n21046), .B(n21045), .Z(n21047) );
  AND U22700 ( .A(n21048), .B(n21047), .Z(n21075) );
  NAND U22701 ( .A(n42143), .B(n21049), .Z(n21051) );
  XNOR U22702 ( .A(a[453]), .B(n4136), .Z(n21086) );
  NAND U22703 ( .A(n42144), .B(n21086), .Z(n21050) );
  AND U22704 ( .A(n21051), .B(n21050), .Z(n21101) );
  XOR U22705 ( .A(a[457]), .B(n42012), .Z(n21089) );
  XNOR U22706 ( .A(n21101), .B(n21100), .Z(n21103) );
  XOR U22707 ( .A(a[455]), .B(n42085), .Z(n21093) );
  AND U22708 ( .A(a[451]), .B(b[7]), .Z(n21094) );
  XNOR U22709 ( .A(n21095), .B(n21094), .Z(n21096) );
  AND U22710 ( .A(a[459]), .B(b[0]), .Z(n21054) );
  XNOR U22711 ( .A(n21054), .B(n4071), .Z(n21056) );
  NANDN U22712 ( .A(b[0]), .B(a[458]), .Z(n21055) );
  NAND U22713 ( .A(n21056), .B(n21055), .Z(n21097) );
  XNOR U22714 ( .A(n21096), .B(n21097), .Z(n21102) );
  XOR U22715 ( .A(n21103), .B(n21102), .Z(n21081) );
  NANDN U22716 ( .A(n21058), .B(n21057), .Z(n21062) );
  NANDN U22717 ( .A(n21060), .B(n21059), .Z(n21061) );
  AND U22718 ( .A(n21062), .B(n21061), .Z(n21080) );
  XNOR U22719 ( .A(n21081), .B(n21080), .Z(n21082) );
  NANDN U22720 ( .A(n21064), .B(n21063), .Z(n21068) );
  NAND U22721 ( .A(n21066), .B(n21065), .Z(n21067) );
  NAND U22722 ( .A(n21068), .B(n21067), .Z(n21083) );
  XNOR U22723 ( .A(n21082), .B(n21083), .Z(n21074) );
  XNOR U22724 ( .A(n21075), .B(n21074), .Z(n21076) );
  XNOR U22725 ( .A(n21077), .B(n21076), .Z(n21106) );
  XNOR U22726 ( .A(sreg[1475]), .B(n21106), .Z(n21108) );
  NANDN U22727 ( .A(sreg[1474]), .B(n21069), .Z(n21073) );
  NAND U22728 ( .A(n21071), .B(n21070), .Z(n21072) );
  NAND U22729 ( .A(n21073), .B(n21072), .Z(n21107) );
  XNOR U22730 ( .A(n21108), .B(n21107), .Z(c[1475]) );
  NANDN U22731 ( .A(n21075), .B(n21074), .Z(n21079) );
  NANDN U22732 ( .A(n21077), .B(n21076), .Z(n21078) );
  AND U22733 ( .A(n21079), .B(n21078), .Z(n21114) );
  NANDN U22734 ( .A(n21081), .B(n21080), .Z(n21085) );
  NANDN U22735 ( .A(n21083), .B(n21082), .Z(n21084) );
  AND U22736 ( .A(n21085), .B(n21084), .Z(n21112) );
  NAND U22737 ( .A(n42143), .B(n21086), .Z(n21088) );
  XNOR U22738 ( .A(a[454]), .B(n4136), .Z(n21123) );
  NAND U22739 ( .A(n42144), .B(n21123), .Z(n21087) );
  AND U22740 ( .A(n21088), .B(n21087), .Z(n21138) );
  XOR U22741 ( .A(a[458]), .B(n42012), .Z(n21126) );
  XNOR U22742 ( .A(n21138), .B(n21137), .Z(n21140) );
  AND U22743 ( .A(a[460]), .B(b[0]), .Z(n21090) );
  XNOR U22744 ( .A(n21090), .B(n4071), .Z(n21092) );
  NANDN U22745 ( .A(b[0]), .B(a[459]), .Z(n21091) );
  NAND U22746 ( .A(n21092), .B(n21091), .Z(n21134) );
  XOR U22747 ( .A(a[456]), .B(n42085), .Z(n21130) );
  AND U22748 ( .A(a[452]), .B(b[7]), .Z(n21131) );
  XNOR U22749 ( .A(n21132), .B(n21131), .Z(n21133) );
  XNOR U22750 ( .A(n21134), .B(n21133), .Z(n21139) );
  XOR U22751 ( .A(n21140), .B(n21139), .Z(n21118) );
  NANDN U22752 ( .A(n21095), .B(n21094), .Z(n21099) );
  NANDN U22753 ( .A(n21097), .B(n21096), .Z(n21098) );
  AND U22754 ( .A(n21099), .B(n21098), .Z(n21117) );
  XNOR U22755 ( .A(n21118), .B(n21117), .Z(n21119) );
  NANDN U22756 ( .A(n21101), .B(n21100), .Z(n21105) );
  NAND U22757 ( .A(n21103), .B(n21102), .Z(n21104) );
  NAND U22758 ( .A(n21105), .B(n21104), .Z(n21120) );
  XNOR U22759 ( .A(n21119), .B(n21120), .Z(n21111) );
  XNOR U22760 ( .A(n21112), .B(n21111), .Z(n21113) );
  XNOR U22761 ( .A(n21114), .B(n21113), .Z(n21143) );
  XNOR U22762 ( .A(sreg[1476]), .B(n21143), .Z(n21145) );
  NANDN U22763 ( .A(sreg[1475]), .B(n21106), .Z(n21110) );
  NAND U22764 ( .A(n21108), .B(n21107), .Z(n21109) );
  NAND U22765 ( .A(n21110), .B(n21109), .Z(n21144) );
  XNOR U22766 ( .A(n21145), .B(n21144), .Z(c[1476]) );
  NANDN U22767 ( .A(n21112), .B(n21111), .Z(n21116) );
  NANDN U22768 ( .A(n21114), .B(n21113), .Z(n21115) );
  AND U22769 ( .A(n21116), .B(n21115), .Z(n21151) );
  NANDN U22770 ( .A(n21118), .B(n21117), .Z(n21122) );
  NANDN U22771 ( .A(n21120), .B(n21119), .Z(n21121) );
  AND U22772 ( .A(n21122), .B(n21121), .Z(n21149) );
  NAND U22773 ( .A(n42143), .B(n21123), .Z(n21125) );
  XNOR U22774 ( .A(a[455]), .B(n4136), .Z(n21160) );
  NAND U22775 ( .A(n42144), .B(n21160), .Z(n21124) );
  AND U22776 ( .A(n21125), .B(n21124), .Z(n21175) );
  XOR U22777 ( .A(a[459]), .B(n42012), .Z(n21163) );
  XNOR U22778 ( .A(n21175), .B(n21174), .Z(n21177) );
  AND U22779 ( .A(a[461]), .B(b[0]), .Z(n21127) );
  XNOR U22780 ( .A(n21127), .B(n4071), .Z(n21129) );
  NANDN U22781 ( .A(b[0]), .B(a[460]), .Z(n21128) );
  NAND U22782 ( .A(n21129), .B(n21128), .Z(n21171) );
  XOR U22783 ( .A(a[457]), .B(n42085), .Z(n21167) );
  AND U22784 ( .A(a[453]), .B(b[7]), .Z(n21168) );
  XNOR U22785 ( .A(n21169), .B(n21168), .Z(n21170) );
  XNOR U22786 ( .A(n21171), .B(n21170), .Z(n21176) );
  XOR U22787 ( .A(n21177), .B(n21176), .Z(n21155) );
  NANDN U22788 ( .A(n21132), .B(n21131), .Z(n21136) );
  NANDN U22789 ( .A(n21134), .B(n21133), .Z(n21135) );
  AND U22790 ( .A(n21136), .B(n21135), .Z(n21154) );
  XNOR U22791 ( .A(n21155), .B(n21154), .Z(n21156) );
  NANDN U22792 ( .A(n21138), .B(n21137), .Z(n21142) );
  NAND U22793 ( .A(n21140), .B(n21139), .Z(n21141) );
  NAND U22794 ( .A(n21142), .B(n21141), .Z(n21157) );
  XNOR U22795 ( .A(n21156), .B(n21157), .Z(n21148) );
  XNOR U22796 ( .A(n21149), .B(n21148), .Z(n21150) );
  XNOR U22797 ( .A(n21151), .B(n21150), .Z(n21180) );
  XNOR U22798 ( .A(sreg[1477]), .B(n21180), .Z(n21182) );
  NANDN U22799 ( .A(sreg[1476]), .B(n21143), .Z(n21147) );
  NAND U22800 ( .A(n21145), .B(n21144), .Z(n21146) );
  NAND U22801 ( .A(n21147), .B(n21146), .Z(n21181) );
  XNOR U22802 ( .A(n21182), .B(n21181), .Z(c[1477]) );
  NANDN U22803 ( .A(n21149), .B(n21148), .Z(n21153) );
  NANDN U22804 ( .A(n21151), .B(n21150), .Z(n21152) );
  AND U22805 ( .A(n21153), .B(n21152), .Z(n21188) );
  NANDN U22806 ( .A(n21155), .B(n21154), .Z(n21159) );
  NANDN U22807 ( .A(n21157), .B(n21156), .Z(n21158) );
  AND U22808 ( .A(n21159), .B(n21158), .Z(n21186) );
  NAND U22809 ( .A(n42143), .B(n21160), .Z(n21162) );
  XNOR U22810 ( .A(a[456]), .B(n4137), .Z(n21197) );
  NAND U22811 ( .A(n42144), .B(n21197), .Z(n21161) );
  AND U22812 ( .A(n21162), .B(n21161), .Z(n21212) );
  XOR U22813 ( .A(a[460]), .B(n42012), .Z(n21200) );
  XNOR U22814 ( .A(n21212), .B(n21211), .Z(n21214) );
  AND U22815 ( .A(a[462]), .B(b[0]), .Z(n21164) );
  XNOR U22816 ( .A(n21164), .B(n4071), .Z(n21166) );
  NANDN U22817 ( .A(b[0]), .B(a[461]), .Z(n21165) );
  NAND U22818 ( .A(n21166), .B(n21165), .Z(n21208) );
  XOR U22819 ( .A(a[458]), .B(n42085), .Z(n21201) );
  AND U22820 ( .A(a[454]), .B(b[7]), .Z(n21205) );
  XNOR U22821 ( .A(n21206), .B(n21205), .Z(n21207) );
  XNOR U22822 ( .A(n21208), .B(n21207), .Z(n21213) );
  XOR U22823 ( .A(n21214), .B(n21213), .Z(n21192) );
  NANDN U22824 ( .A(n21169), .B(n21168), .Z(n21173) );
  NANDN U22825 ( .A(n21171), .B(n21170), .Z(n21172) );
  AND U22826 ( .A(n21173), .B(n21172), .Z(n21191) );
  XNOR U22827 ( .A(n21192), .B(n21191), .Z(n21193) );
  NANDN U22828 ( .A(n21175), .B(n21174), .Z(n21179) );
  NAND U22829 ( .A(n21177), .B(n21176), .Z(n21178) );
  NAND U22830 ( .A(n21179), .B(n21178), .Z(n21194) );
  XNOR U22831 ( .A(n21193), .B(n21194), .Z(n21185) );
  XNOR U22832 ( .A(n21186), .B(n21185), .Z(n21187) );
  XNOR U22833 ( .A(n21188), .B(n21187), .Z(n21217) );
  XNOR U22834 ( .A(sreg[1478]), .B(n21217), .Z(n21219) );
  NANDN U22835 ( .A(sreg[1477]), .B(n21180), .Z(n21184) );
  NAND U22836 ( .A(n21182), .B(n21181), .Z(n21183) );
  NAND U22837 ( .A(n21184), .B(n21183), .Z(n21218) );
  XNOR U22838 ( .A(n21219), .B(n21218), .Z(c[1478]) );
  NANDN U22839 ( .A(n21186), .B(n21185), .Z(n21190) );
  NANDN U22840 ( .A(n21188), .B(n21187), .Z(n21189) );
  AND U22841 ( .A(n21190), .B(n21189), .Z(n21225) );
  NANDN U22842 ( .A(n21192), .B(n21191), .Z(n21196) );
  NANDN U22843 ( .A(n21194), .B(n21193), .Z(n21195) );
  AND U22844 ( .A(n21196), .B(n21195), .Z(n21223) );
  NAND U22845 ( .A(n42143), .B(n21197), .Z(n21199) );
  XNOR U22846 ( .A(a[457]), .B(n4137), .Z(n21234) );
  NAND U22847 ( .A(n42144), .B(n21234), .Z(n21198) );
  AND U22848 ( .A(n21199), .B(n21198), .Z(n21249) );
  XOR U22849 ( .A(a[461]), .B(n42012), .Z(n21237) );
  XNOR U22850 ( .A(n21249), .B(n21248), .Z(n21251) );
  XOR U22851 ( .A(a[459]), .B(n42085), .Z(n21238) );
  AND U22852 ( .A(a[455]), .B(b[7]), .Z(n21242) );
  XNOR U22853 ( .A(n21243), .B(n21242), .Z(n21244) );
  AND U22854 ( .A(a[463]), .B(b[0]), .Z(n21202) );
  XNOR U22855 ( .A(n21202), .B(n4071), .Z(n21204) );
  NANDN U22856 ( .A(b[0]), .B(a[462]), .Z(n21203) );
  NAND U22857 ( .A(n21204), .B(n21203), .Z(n21245) );
  XNOR U22858 ( .A(n21244), .B(n21245), .Z(n21250) );
  XOR U22859 ( .A(n21251), .B(n21250), .Z(n21229) );
  NANDN U22860 ( .A(n21206), .B(n21205), .Z(n21210) );
  NANDN U22861 ( .A(n21208), .B(n21207), .Z(n21209) );
  AND U22862 ( .A(n21210), .B(n21209), .Z(n21228) );
  XNOR U22863 ( .A(n21229), .B(n21228), .Z(n21230) );
  NANDN U22864 ( .A(n21212), .B(n21211), .Z(n21216) );
  NAND U22865 ( .A(n21214), .B(n21213), .Z(n21215) );
  NAND U22866 ( .A(n21216), .B(n21215), .Z(n21231) );
  XNOR U22867 ( .A(n21230), .B(n21231), .Z(n21222) );
  XNOR U22868 ( .A(n21223), .B(n21222), .Z(n21224) );
  XNOR U22869 ( .A(n21225), .B(n21224), .Z(n21254) );
  XNOR U22870 ( .A(sreg[1479]), .B(n21254), .Z(n21256) );
  NANDN U22871 ( .A(sreg[1478]), .B(n21217), .Z(n21221) );
  NAND U22872 ( .A(n21219), .B(n21218), .Z(n21220) );
  NAND U22873 ( .A(n21221), .B(n21220), .Z(n21255) );
  XNOR U22874 ( .A(n21256), .B(n21255), .Z(c[1479]) );
  NANDN U22875 ( .A(n21223), .B(n21222), .Z(n21227) );
  NANDN U22876 ( .A(n21225), .B(n21224), .Z(n21226) );
  AND U22877 ( .A(n21227), .B(n21226), .Z(n21262) );
  NANDN U22878 ( .A(n21229), .B(n21228), .Z(n21233) );
  NANDN U22879 ( .A(n21231), .B(n21230), .Z(n21232) );
  AND U22880 ( .A(n21233), .B(n21232), .Z(n21260) );
  NAND U22881 ( .A(n42143), .B(n21234), .Z(n21236) );
  XNOR U22882 ( .A(a[458]), .B(n4137), .Z(n21271) );
  NAND U22883 ( .A(n42144), .B(n21271), .Z(n21235) );
  AND U22884 ( .A(n21236), .B(n21235), .Z(n21286) );
  XOR U22885 ( .A(a[462]), .B(n42012), .Z(n21274) );
  XNOR U22886 ( .A(n21286), .B(n21285), .Z(n21288) );
  XOR U22887 ( .A(a[460]), .B(n42085), .Z(n21278) );
  AND U22888 ( .A(a[456]), .B(b[7]), .Z(n21279) );
  XNOR U22889 ( .A(n21280), .B(n21279), .Z(n21281) );
  AND U22890 ( .A(a[464]), .B(b[0]), .Z(n21239) );
  XNOR U22891 ( .A(n21239), .B(n4071), .Z(n21241) );
  NANDN U22892 ( .A(b[0]), .B(a[463]), .Z(n21240) );
  NAND U22893 ( .A(n21241), .B(n21240), .Z(n21282) );
  XNOR U22894 ( .A(n21281), .B(n21282), .Z(n21287) );
  XOR U22895 ( .A(n21288), .B(n21287), .Z(n21266) );
  NANDN U22896 ( .A(n21243), .B(n21242), .Z(n21247) );
  NANDN U22897 ( .A(n21245), .B(n21244), .Z(n21246) );
  AND U22898 ( .A(n21247), .B(n21246), .Z(n21265) );
  XNOR U22899 ( .A(n21266), .B(n21265), .Z(n21267) );
  NANDN U22900 ( .A(n21249), .B(n21248), .Z(n21253) );
  NAND U22901 ( .A(n21251), .B(n21250), .Z(n21252) );
  NAND U22902 ( .A(n21253), .B(n21252), .Z(n21268) );
  XNOR U22903 ( .A(n21267), .B(n21268), .Z(n21259) );
  XNOR U22904 ( .A(n21260), .B(n21259), .Z(n21261) );
  XNOR U22905 ( .A(n21262), .B(n21261), .Z(n21291) );
  XNOR U22906 ( .A(sreg[1480]), .B(n21291), .Z(n21293) );
  NANDN U22907 ( .A(sreg[1479]), .B(n21254), .Z(n21258) );
  NAND U22908 ( .A(n21256), .B(n21255), .Z(n21257) );
  NAND U22909 ( .A(n21258), .B(n21257), .Z(n21292) );
  XNOR U22910 ( .A(n21293), .B(n21292), .Z(c[1480]) );
  NANDN U22911 ( .A(n21260), .B(n21259), .Z(n21264) );
  NANDN U22912 ( .A(n21262), .B(n21261), .Z(n21263) );
  AND U22913 ( .A(n21264), .B(n21263), .Z(n21299) );
  NANDN U22914 ( .A(n21266), .B(n21265), .Z(n21270) );
  NANDN U22915 ( .A(n21268), .B(n21267), .Z(n21269) );
  AND U22916 ( .A(n21270), .B(n21269), .Z(n21297) );
  NAND U22917 ( .A(n42143), .B(n21271), .Z(n21273) );
  XNOR U22918 ( .A(a[459]), .B(n4137), .Z(n21308) );
  NAND U22919 ( .A(n42144), .B(n21308), .Z(n21272) );
  AND U22920 ( .A(n21273), .B(n21272), .Z(n21323) );
  XOR U22921 ( .A(a[463]), .B(n42012), .Z(n21311) );
  XNOR U22922 ( .A(n21323), .B(n21322), .Z(n21325) );
  AND U22923 ( .A(a[465]), .B(b[0]), .Z(n21275) );
  XNOR U22924 ( .A(n21275), .B(n4071), .Z(n21277) );
  NANDN U22925 ( .A(b[0]), .B(a[464]), .Z(n21276) );
  NAND U22926 ( .A(n21277), .B(n21276), .Z(n21319) );
  XOR U22927 ( .A(a[461]), .B(n42085), .Z(n21312) );
  AND U22928 ( .A(a[457]), .B(b[7]), .Z(n21316) );
  XNOR U22929 ( .A(n21317), .B(n21316), .Z(n21318) );
  XNOR U22930 ( .A(n21319), .B(n21318), .Z(n21324) );
  XOR U22931 ( .A(n21325), .B(n21324), .Z(n21303) );
  NANDN U22932 ( .A(n21280), .B(n21279), .Z(n21284) );
  NANDN U22933 ( .A(n21282), .B(n21281), .Z(n21283) );
  AND U22934 ( .A(n21284), .B(n21283), .Z(n21302) );
  XNOR U22935 ( .A(n21303), .B(n21302), .Z(n21304) );
  NANDN U22936 ( .A(n21286), .B(n21285), .Z(n21290) );
  NAND U22937 ( .A(n21288), .B(n21287), .Z(n21289) );
  NAND U22938 ( .A(n21290), .B(n21289), .Z(n21305) );
  XNOR U22939 ( .A(n21304), .B(n21305), .Z(n21296) );
  XNOR U22940 ( .A(n21297), .B(n21296), .Z(n21298) );
  XNOR U22941 ( .A(n21299), .B(n21298), .Z(n21328) );
  XNOR U22942 ( .A(sreg[1481]), .B(n21328), .Z(n21330) );
  NANDN U22943 ( .A(sreg[1480]), .B(n21291), .Z(n21295) );
  NAND U22944 ( .A(n21293), .B(n21292), .Z(n21294) );
  NAND U22945 ( .A(n21295), .B(n21294), .Z(n21329) );
  XNOR U22946 ( .A(n21330), .B(n21329), .Z(c[1481]) );
  NANDN U22947 ( .A(n21297), .B(n21296), .Z(n21301) );
  NANDN U22948 ( .A(n21299), .B(n21298), .Z(n21300) );
  AND U22949 ( .A(n21301), .B(n21300), .Z(n21336) );
  NANDN U22950 ( .A(n21303), .B(n21302), .Z(n21307) );
  NANDN U22951 ( .A(n21305), .B(n21304), .Z(n21306) );
  AND U22952 ( .A(n21307), .B(n21306), .Z(n21334) );
  NAND U22953 ( .A(n42143), .B(n21308), .Z(n21310) );
  XNOR U22954 ( .A(a[460]), .B(n4137), .Z(n21345) );
  NAND U22955 ( .A(n42144), .B(n21345), .Z(n21309) );
  AND U22956 ( .A(n21310), .B(n21309), .Z(n21360) );
  XOR U22957 ( .A(a[464]), .B(n42012), .Z(n21348) );
  XNOR U22958 ( .A(n21360), .B(n21359), .Z(n21362) );
  XOR U22959 ( .A(a[462]), .B(n42085), .Z(n21352) );
  AND U22960 ( .A(a[458]), .B(b[7]), .Z(n21353) );
  XNOR U22961 ( .A(n21354), .B(n21353), .Z(n21355) );
  AND U22962 ( .A(a[466]), .B(b[0]), .Z(n21313) );
  XNOR U22963 ( .A(n21313), .B(n4071), .Z(n21315) );
  NANDN U22964 ( .A(b[0]), .B(a[465]), .Z(n21314) );
  NAND U22965 ( .A(n21315), .B(n21314), .Z(n21356) );
  XNOR U22966 ( .A(n21355), .B(n21356), .Z(n21361) );
  XOR U22967 ( .A(n21362), .B(n21361), .Z(n21340) );
  NANDN U22968 ( .A(n21317), .B(n21316), .Z(n21321) );
  NANDN U22969 ( .A(n21319), .B(n21318), .Z(n21320) );
  AND U22970 ( .A(n21321), .B(n21320), .Z(n21339) );
  XNOR U22971 ( .A(n21340), .B(n21339), .Z(n21341) );
  NANDN U22972 ( .A(n21323), .B(n21322), .Z(n21327) );
  NAND U22973 ( .A(n21325), .B(n21324), .Z(n21326) );
  NAND U22974 ( .A(n21327), .B(n21326), .Z(n21342) );
  XNOR U22975 ( .A(n21341), .B(n21342), .Z(n21333) );
  XNOR U22976 ( .A(n21334), .B(n21333), .Z(n21335) );
  XNOR U22977 ( .A(n21336), .B(n21335), .Z(n21365) );
  XNOR U22978 ( .A(sreg[1482]), .B(n21365), .Z(n21367) );
  NANDN U22979 ( .A(sreg[1481]), .B(n21328), .Z(n21332) );
  NAND U22980 ( .A(n21330), .B(n21329), .Z(n21331) );
  NAND U22981 ( .A(n21332), .B(n21331), .Z(n21366) );
  XNOR U22982 ( .A(n21367), .B(n21366), .Z(c[1482]) );
  NANDN U22983 ( .A(n21334), .B(n21333), .Z(n21338) );
  NANDN U22984 ( .A(n21336), .B(n21335), .Z(n21337) );
  AND U22985 ( .A(n21338), .B(n21337), .Z(n21373) );
  NANDN U22986 ( .A(n21340), .B(n21339), .Z(n21344) );
  NANDN U22987 ( .A(n21342), .B(n21341), .Z(n21343) );
  AND U22988 ( .A(n21344), .B(n21343), .Z(n21371) );
  NAND U22989 ( .A(n42143), .B(n21345), .Z(n21347) );
  XNOR U22990 ( .A(a[461]), .B(n4137), .Z(n21382) );
  NAND U22991 ( .A(n42144), .B(n21382), .Z(n21346) );
  AND U22992 ( .A(n21347), .B(n21346), .Z(n21397) );
  XOR U22993 ( .A(a[465]), .B(n42012), .Z(n21385) );
  XNOR U22994 ( .A(n21397), .B(n21396), .Z(n21399) );
  AND U22995 ( .A(a[467]), .B(b[0]), .Z(n21349) );
  XNOR U22996 ( .A(n21349), .B(n4071), .Z(n21351) );
  NANDN U22997 ( .A(b[0]), .B(a[466]), .Z(n21350) );
  NAND U22998 ( .A(n21351), .B(n21350), .Z(n21393) );
  XOR U22999 ( .A(a[463]), .B(n42085), .Z(n21389) );
  AND U23000 ( .A(a[459]), .B(b[7]), .Z(n21390) );
  XNOR U23001 ( .A(n21391), .B(n21390), .Z(n21392) );
  XNOR U23002 ( .A(n21393), .B(n21392), .Z(n21398) );
  XOR U23003 ( .A(n21399), .B(n21398), .Z(n21377) );
  NANDN U23004 ( .A(n21354), .B(n21353), .Z(n21358) );
  NANDN U23005 ( .A(n21356), .B(n21355), .Z(n21357) );
  AND U23006 ( .A(n21358), .B(n21357), .Z(n21376) );
  XNOR U23007 ( .A(n21377), .B(n21376), .Z(n21378) );
  NANDN U23008 ( .A(n21360), .B(n21359), .Z(n21364) );
  NAND U23009 ( .A(n21362), .B(n21361), .Z(n21363) );
  NAND U23010 ( .A(n21364), .B(n21363), .Z(n21379) );
  XNOR U23011 ( .A(n21378), .B(n21379), .Z(n21370) );
  XNOR U23012 ( .A(n21371), .B(n21370), .Z(n21372) );
  XNOR U23013 ( .A(n21373), .B(n21372), .Z(n21402) );
  XNOR U23014 ( .A(sreg[1483]), .B(n21402), .Z(n21404) );
  NANDN U23015 ( .A(sreg[1482]), .B(n21365), .Z(n21369) );
  NAND U23016 ( .A(n21367), .B(n21366), .Z(n21368) );
  NAND U23017 ( .A(n21369), .B(n21368), .Z(n21403) );
  XNOR U23018 ( .A(n21404), .B(n21403), .Z(c[1483]) );
  NANDN U23019 ( .A(n21371), .B(n21370), .Z(n21375) );
  NANDN U23020 ( .A(n21373), .B(n21372), .Z(n21374) );
  AND U23021 ( .A(n21375), .B(n21374), .Z(n21410) );
  NANDN U23022 ( .A(n21377), .B(n21376), .Z(n21381) );
  NANDN U23023 ( .A(n21379), .B(n21378), .Z(n21380) );
  AND U23024 ( .A(n21381), .B(n21380), .Z(n21408) );
  NAND U23025 ( .A(n42143), .B(n21382), .Z(n21384) );
  XNOR U23026 ( .A(a[462]), .B(n4137), .Z(n21419) );
  NAND U23027 ( .A(n42144), .B(n21419), .Z(n21383) );
  AND U23028 ( .A(n21384), .B(n21383), .Z(n21434) );
  XOR U23029 ( .A(a[466]), .B(n42012), .Z(n21422) );
  XNOR U23030 ( .A(n21434), .B(n21433), .Z(n21436) );
  AND U23031 ( .A(a[468]), .B(b[0]), .Z(n21386) );
  XNOR U23032 ( .A(n21386), .B(n4071), .Z(n21388) );
  NANDN U23033 ( .A(b[0]), .B(a[467]), .Z(n21387) );
  NAND U23034 ( .A(n21388), .B(n21387), .Z(n21430) );
  XOR U23035 ( .A(a[464]), .B(n42085), .Z(n21423) );
  AND U23036 ( .A(a[460]), .B(b[7]), .Z(n21427) );
  XNOR U23037 ( .A(n21428), .B(n21427), .Z(n21429) );
  XNOR U23038 ( .A(n21430), .B(n21429), .Z(n21435) );
  XOR U23039 ( .A(n21436), .B(n21435), .Z(n21414) );
  NANDN U23040 ( .A(n21391), .B(n21390), .Z(n21395) );
  NANDN U23041 ( .A(n21393), .B(n21392), .Z(n21394) );
  AND U23042 ( .A(n21395), .B(n21394), .Z(n21413) );
  XNOR U23043 ( .A(n21414), .B(n21413), .Z(n21415) );
  NANDN U23044 ( .A(n21397), .B(n21396), .Z(n21401) );
  NAND U23045 ( .A(n21399), .B(n21398), .Z(n21400) );
  NAND U23046 ( .A(n21401), .B(n21400), .Z(n21416) );
  XNOR U23047 ( .A(n21415), .B(n21416), .Z(n21407) );
  XNOR U23048 ( .A(n21408), .B(n21407), .Z(n21409) );
  XNOR U23049 ( .A(n21410), .B(n21409), .Z(n21439) );
  XNOR U23050 ( .A(sreg[1484]), .B(n21439), .Z(n21441) );
  NANDN U23051 ( .A(sreg[1483]), .B(n21402), .Z(n21406) );
  NAND U23052 ( .A(n21404), .B(n21403), .Z(n21405) );
  NAND U23053 ( .A(n21406), .B(n21405), .Z(n21440) );
  XNOR U23054 ( .A(n21441), .B(n21440), .Z(c[1484]) );
  NANDN U23055 ( .A(n21408), .B(n21407), .Z(n21412) );
  NANDN U23056 ( .A(n21410), .B(n21409), .Z(n21411) );
  AND U23057 ( .A(n21412), .B(n21411), .Z(n21447) );
  NANDN U23058 ( .A(n21414), .B(n21413), .Z(n21418) );
  NANDN U23059 ( .A(n21416), .B(n21415), .Z(n21417) );
  AND U23060 ( .A(n21418), .B(n21417), .Z(n21445) );
  NAND U23061 ( .A(n42143), .B(n21419), .Z(n21421) );
  XNOR U23062 ( .A(a[463]), .B(n4138), .Z(n21456) );
  NAND U23063 ( .A(n42144), .B(n21456), .Z(n21420) );
  AND U23064 ( .A(n21421), .B(n21420), .Z(n21471) );
  XOR U23065 ( .A(a[467]), .B(n42012), .Z(n21459) );
  XNOR U23066 ( .A(n21471), .B(n21470), .Z(n21473) );
  XOR U23067 ( .A(a[465]), .B(n42085), .Z(n21463) );
  AND U23068 ( .A(a[461]), .B(b[7]), .Z(n21464) );
  XNOR U23069 ( .A(n21465), .B(n21464), .Z(n21466) );
  AND U23070 ( .A(a[469]), .B(b[0]), .Z(n21424) );
  XNOR U23071 ( .A(n21424), .B(n4071), .Z(n21426) );
  NANDN U23072 ( .A(b[0]), .B(a[468]), .Z(n21425) );
  NAND U23073 ( .A(n21426), .B(n21425), .Z(n21467) );
  XNOR U23074 ( .A(n21466), .B(n21467), .Z(n21472) );
  XOR U23075 ( .A(n21473), .B(n21472), .Z(n21451) );
  NANDN U23076 ( .A(n21428), .B(n21427), .Z(n21432) );
  NANDN U23077 ( .A(n21430), .B(n21429), .Z(n21431) );
  AND U23078 ( .A(n21432), .B(n21431), .Z(n21450) );
  XNOR U23079 ( .A(n21451), .B(n21450), .Z(n21452) );
  NANDN U23080 ( .A(n21434), .B(n21433), .Z(n21438) );
  NAND U23081 ( .A(n21436), .B(n21435), .Z(n21437) );
  NAND U23082 ( .A(n21438), .B(n21437), .Z(n21453) );
  XNOR U23083 ( .A(n21452), .B(n21453), .Z(n21444) );
  XNOR U23084 ( .A(n21445), .B(n21444), .Z(n21446) );
  XNOR U23085 ( .A(n21447), .B(n21446), .Z(n21476) );
  XNOR U23086 ( .A(sreg[1485]), .B(n21476), .Z(n21478) );
  NANDN U23087 ( .A(sreg[1484]), .B(n21439), .Z(n21443) );
  NAND U23088 ( .A(n21441), .B(n21440), .Z(n21442) );
  NAND U23089 ( .A(n21443), .B(n21442), .Z(n21477) );
  XNOR U23090 ( .A(n21478), .B(n21477), .Z(c[1485]) );
  NANDN U23091 ( .A(n21445), .B(n21444), .Z(n21449) );
  NANDN U23092 ( .A(n21447), .B(n21446), .Z(n21448) );
  AND U23093 ( .A(n21449), .B(n21448), .Z(n21484) );
  NANDN U23094 ( .A(n21451), .B(n21450), .Z(n21455) );
  NANDN U23095 ( .A(n21453), .B(n21452), .Z(n21454) );
  AND U23096 ( .A(n21455), .B(n21454), .Z(n21482) );
  NAND U23097 ( .A(n42143), .B(n21456), .Z(n21458) );
  XNOR U23098 ( .A(a[464]), .B(n4138), .Z(n21493) );
  NAND U23099 ( .A(n42144), .B(n21493), .Z(n21457) );
  AND U23100 ( .A(n21458), .B(n21457), .Z(n21508) );
  XOR U23101 ( .A(a[468]), .B(n42012), .Z(n21496) );
  XNOR U23102 ( .A(n21508), .B(n21507), .Z(n21510) );
  AND U23103 ( .A(a[470]), .B(b[0]), .Z(n21460) );
  XNOR U23104 ( .A(n21460), .B(n4071), .Z(n21462) );
  NANDN U23105 ( .A(b[0]), .B(a[469]), .Z(n21461) );
  NAND U23106 ( .A(n21462), .B(n21461), .Z(n21504) );
  XOR U23107 ( .A(a[466]), .B(n42085), .Z(n21500) );
  AND U23108 ( .A(a[462]), .B(b[7]), .Z(n21501) );
  XNOR U23109 ( .A(n21502), .B(n21501), .Z(n21503) );
  XNOR U23110 ( .A(n21504), .B(n21503), .Z(n21509) );
  XOR U23111 ( .A(n21510), .B(n21509), .Z(n21488) );
  NANDN U23112 ( .A(n21465), .B(n21464), .Z(n21469) );
  NANDN U23113 ( .A(n21467), .B(n21466), .Z(n21468) );
  AND U23114 ( .A(n21469), .B(n21468), .Z(n21487) );
  XNOR U23115 ( .A(n21488), .B(n21487), .Z(n21489) );
  NANDN U23116 ( .A(n21471), .B(n21470), .Z(n21475) );
  NAND U23117 ( .A(n21473), .B(n21472), .Z(n21474) );
  NAND U23118 ( .A(n21475), .B(n21474), .Z(n21490) );
  XNOR U23119 ( .A(n21489), .B(n21490), .Z(n21481) );
  XNOR U23120 ( .A(n21482), .B(n21481), .Z(n21483) );
  XNOR U23121 ( .A(n21484), .B(n21483), .Z(n21513) );
  XNOR U23122 ( .A(sreg[1486]), .B(n21513), .Z(n21515) );
  NANDN U23123 ( .A(sreg[1485]), .B(n21476), .Z(n21480) );
  NAND U23124 ( .A(n21478), .B(n21477), .Z(n21479) );
  NAND U23125 ( .A(n21480), .B(n21479), .Z(n21514) );
  XNOR U23126 ( .A(n21515), .B(n21514), .Z(c[1486]) );
  NANDN U23127 ( .A(n21482), .B(n21481), .Z(n21486) );
  NANDN U23128 ( .A(n21484), .B(n21483), .Z(n21485) );
  AND U23129 ( .A(n21486), .B(n21485), .Z(n21521) );
  NANDN U23130 ( .A(n21488), .B(n21487), .Z(n21492) );
  NANDN U23131 ( .A(n21490), .B(n21489), .Z(n21491) );
  AND U23132 ( .A(n21492), .B(n21491), .Z(n21519) );
  NAND U23133 ( .A(n42143), .B(n21493), .Z(n21495) );
  XNOR U23134 ( .A(a[465]), .B(n4138), .Z(n21530) );
  NAND U23135 ( .A(n42144), .B(n21530), .Z(n21494) );
  AND U23136 ( .A(n21495), .B(n21494), .Z(n21545) );
  XOR U23137 ( .A(a[469]), .B(n42012), .Z(n21533) );
  XNOR U23138 ( .A(n21545), .B(n21544), .Z(n21547) );
  AND U23139 ( .A(a[471]), .B(b[0]), .Z(n21497) );
  XNOR U23140 ( .A(n21497), .B(n4071), .Z(n21499) );
  NANDN U23141 ( .A(b[0]), .B(a[470]), .Z(n21498) );
  NAND U23142 ( .A(n21499), .B(n21498), .Z(n21541) );
  XOR U23143 ( .A(a[467]), .B(n42085), .Z(n21537) );
  AND U23144 ( .A(a[463]), .B(b[7]), .Z(n21538) );
  XNOR U23145 ( .A(n21539), .B(n21538), .Z(n21540) );
  XNOR U23146 ( .A(n21541), .B(n21540), .Z(n21546) );
  XOR U23147 ( .A(n21547), .B(n21546), .Z(n21525) );
  NANDN U23148 ( .A(n21502), .B(n21501), .Z(n21506) );
  NANDN U23149 ( .A(n21504), .B(n21503), .Z(n21505) );
  AND U23150 ( .A(n21506), .B(n21505), .Z(n21524) );
  XNOR U23151 ( .A(n21525), .B(n21524), .Z(n21526) );
  NANDN U23152 ( .A(n21508), .B(n21507), .Z(n21512) );
  NAND U23153 ( .A(n21510), .B(n21509), .Z(n21511) );
  NAND U23154 ( .A(n21512), .B(n21511), .Z(n21527) );
  XNOR U23155 ( .A(n21526), .B(n21527), .Z(n21518) );
  XNOR U23156 ( .A(n21519), .B(n21518), .Z(n21520) );
  XNOR U23157 ( .A(n21521), .B(n21520), .Z(n21550) );
  XNOR U23158 ( .A(sreg[1487]), .B(n21550), .Z(n21552) );
  NANDN U23159 ( .A(sreg[1486]), .B(n21513), .Z(n21517) );
  NAND U23160 ( .A(n21515), .B(n21514), .Z(n21516) );
  NAND U23161 ( .A(n21517), .B(n21516), .Z(n21551) );
  XNOR U23162 ( .A(n21552), .B(n21551), .Z(c[1487]) );
  NANDN U23163 ( .A(n21519), .B(n21518), .Z(n21523) );
  NANDN U23164 ( .A(n21521), .B(n21520), .Z(n21522) );
  AND U23165 ( .A(n21523), .B(n21522), .Z(n21558) );
  NANDN U23166 ( .A(n21525), .B(n21524), .Z(n21529) );
  NANDN U23167 ( .A(n21527), .B(n21526), .Z(n21528) );
  AND U23168 ( .A(n21529), .B(n21528), .Z(n21556) );
  NAND U23169 ( .A(n42143), .B(n21530), .Z(n21532) );
  XNOR U23170 ( .A(a[466]), .B(n4138), .Z(n21567) );
  NAND U23171 ( .A(n42144), .B(n21567), .Z(n21531) );
  AND U23172 ( .A(n21532), .B(n21531), .Z(n21582) );
  XOR U23173 ( .A(a[470]), .B(n42012), .Z(n21570) );
  XNOR U23174 ( .A(n21582), .B(n21581), .Z(n21584) );
  AND U23175 ( .A(a[472]), .B(b[0]), .Z(n21534) );
  XNOR U23176 ( .A(n21534), .B(n4071), .Z(n21536) );
  NANDN U23177 ( .A(b[0]), .B(a[471]), .Z(n21535) );
  NAND U23178 ( .A(n21536), .B(n21535), .Z(n21578) );
  XOR U23179 ( .A(a[468]), .B(n42085), .Z(n21571) );
  AND U23180 ( .A(a[464]), .B(b[7]), .Z(n21575) );
  XNOR U23181 ( .A(n21576), .B(n21575), .Z(n21577) );
  XNOR U23182 ( .A(n21578), .B(n21577), .Z(n21583) );
  XOR U23183 ( .A(n21584), .B(n21583), .Z(n21562) );
  NANDN U23184 ( .A(n21539), .B(n21538), .Z(n21543) );
  NANDN U23185 ( .A(n21541), .B(n21540), .Z(n21542) );
  AND U23186 ( .A(n21543), .B(n21542), .Z(n21561) );
  XNOR U23187 ( .A(n21562), .B(n21561), .Z(n21563) );
  NANDN U23188 ( .A(n21545), .B(n21544), .Z(n21549) );
  NAND U23189 ( .A(n21547), .B(n21546), .Z(n21548) );
  NAND U23190 ( .A(n21549), .B(n21548), .Z(n21564) );
  XNOR U23191 ( .A(n21563), .B(n21564), .Z(n21555) );
  XNOR U23192 ( .A(n21556), .B(n21555), .Z(n21557) );
  XNOR U23193 ( .A(n21558), .B(n21557), .Z(n21587) );
  XNOR U23194 ( .A(sreg[1488]), .B(n21587), .Z(n21589) );
  NANDN U23195 ( .A(sreg[1487]), .B(n21550), .Z(n21554) );
  NAND U23196 ( .A(n21552), .B(n21551), .Z(n21553) );
  NAND U23197 ( .A(n21554), .B(n21553), .Z(n21588) );
  XNOR U23198 ( .A(n21589), .B(n21588), .Z(c[1488]) );
  NANDN U23199 ( .A(n21556), .B(n21555), .Z(n21560) );
  NANDN U23200 ( .A(n21558), .B(n21557), .Z(n21559) );
  AND U23201 ( .A(n21560), .B(n21559), .Z(n21595) );
  NANDN U23202 ( .A(n21562), .B(n21561), .Z(n21566) );
  NANDN U23203 ( .A(n21564), .B(n21563), .Z(n21565) );
  AND U23204 ( .A(n21566), .B(n21565), .Z(n21593) );
  NAND U23205 ( .A(n42143), .B(n21567), .Z(n21569) );
  XNOR U23206 ( .A(a[467]), .B(n4138), .Z(n21604) );
  NAND U23207 ( .A(n42144), .B(n21604), .Z(n21568) );
  AND U23208 ( .A(n21569), .B(n21568), .Z(n21619) );
  XOR U23209 ( .A(a[471]), .B(n42012), .Z(n21607) );
  XNOR U23210 ( .A(n21619), .B(n21618), .Z(n21621) );
  XOR U23211 ( .A(a[469]), .B(n42085), .Z(n21611) );
  AND U23212 ( .A(a[465]), .B(b[7]), .Z(n21612) );
  XNOR U23213 ( .A(n21613), .B(n21612), .Z(n21614) );
  AND U23214 ( .A(a[473]), .B(b[0]), .Z(n21572) );
  XNOR U23215 ( .A(n21572), .B(n4071), .Z(n21574) );
  NANDN U23216 ( .A(b[0]), .B(a[472]), .Z(n21573) );
  NAND U23217 ( .A(n21574), .B(n21573), .Z(n21615) );
  XNOR U23218 ( .A(n21614), .B(n21615), .Z(n21620) );
  XOR U23219 ( .A(n21621), .B(n21620), .Z(n21599) );
  NANDN U23220 ( .A(n21576), .B(n21575), .Z(n21580) );
  NANDN U23221 ( .A(n21578), .B(n21577), .Z(n21579) );
  AND U23222 ( .A(n21580), .B(n21579), .Z(n21598) );
  XNOR U23223 ( .A(n21599), .B(n21598), .Z(n21600) );
  NANDN U23224 ( .A(n21582), .B(n21581), .Z(n21586) );
  NAND U23225 ( .A(n21584), .B(n21583), .Z(n21585) );
  NAND U23226 ( .A(n21586), .B(n21585), .Z(n21601) );
  XNOR U23227 ( .A(n21600), .B(n21601), .Z(n21592) );
  XNOR U23228 ( .A(n21593), .B(n21592), .Z(n21594) );
  XNOR U23229 ( .A(n21595), .B(n21594), .Z(n21624) );
  XNOR U23230 ( .A(sreg[1489]), .B(n21624), .Z(n21626) );
  NANDN U23231 ( .A(sreg[1488]), .B(n21587), .Z(n21591) );
  NAND U23232 ( .A(n21589), .B(n21588), .Z(n21590) );
  NAND U23233 ( .A(n21591), .B(n21590), .Z(n21625) );
  XNOR U23234 ( .A(n21626), .B(n21625), .Z(c[1489]) );
  NANDN U23235 ( .A(n21593), .B(n21592), .Z(n21597) );
  NANDN U23236 ( .A(n21595), .B(n21594), .Z(n21596) );
  AND U23237 ( .A(n21597), .B(n21596), .Z(n21632) );
  NANDN U23238 ( .A(n21599), .B(n21598), .Z(n21603) );
  NANDN U23239 ( .A(n21601), .B(n21600), .Z(n21602) );
  AND U23240 ( .A(n21603), .B(n21602), .Z(n21630) );
  NAND U23241 ( .A(n42143), .B(n21604), .Z(n21606) );
  XNOR U23242 ( .A(a[468]), .B(n4138), .Z(n21641) );
  NAND U23243 ( .A(n42144), .B(n21641), .Z(n21605) );
  AND U23244 ( .A(n21606), .B(n21605), .Z(n21656) );
  XOR U23245 ( .A(a[472]), .B(n42012), .Z(n21644) );
  XNOR U23246 ( .A(n21656), .B(n21655), .Z(n21658) );
  AND U23247 ( .A(a[474]), .B(b[0]), .Z(n21608) );
  XNOR U23248 ( .A(n21608), .B(n4071), .Z(n21610) );
  NANDN U23249 ( .A(b[0]), .B(a[473]), .Z(n21609) );
  NAND U23250 ( .A(n21610), .B(n21609), .Z(n21652) );
  XOR U23251 ( .A(a[470]), .B(n42085), .Z(n21645) );
  AND U23252 ( .A(a[466]), .B(b[7]), .Z(n21649) );
  XNOR U23253 ( .A(n21650), .B(n21649), .Z(n21651) );
  XNOR U23254 ( .A(n21652), .B(n21651), .Z(n21657) );
  XOR U23255 ( .A(n21658), .B(n21657), .Z(n21636) );
  NANDN U23256 ( .A(n21613), .B(n21612), .Z(n21617) );
  NANDN U23257 ( .A(n21615), .B(n21614), .Z(n21616) );
  AND U23258 ( .A(n21617), .B(n21616), .Z(n21635) );
  XNOR U23259 ( .A(n21636), .B(n21635), .Z(n21637) );
  NANDN U23260 ( .A(n21619), .B(n21618), .Z(n21623) );
  NAND U23261 ( .A(n21621), .B(n21620), .Z(n21622) );
  NAND U23262 ( .A(n21623), .B(n21622), .Z(n21638) );
  XNOR U23263 ( .A(n21637), .B(n21638), .Z(n21629) );
  XNOR U23264 ( .A(n21630), .B(n21629), .Z(n21631) );
  XNOR U23265 ( .A(n21632), .B(n21631), .Z(n21661) );
  XNOR U23266 ( .A(sreg[1490]), .B(n21661), .Z(n21663) );
  NANDN U23267 ( .A(sreg[1489]), .B(n21624), .Z(n21628) );
  NAND U23268 ( .A(n21626), .B(n21625), .Z(n21627) );
  NAND U23269 ( .A(n21628), .B(n21627), .Z(n21662) );
  XNOR U23270 ( .A(n21663), .B(n21662), .Z(c[1490]) );
  NANDN U23271 ( .A(n21630), .B(n21629), .Z(n21634) );
  NANDN U23272 ( .A(n21632), .B(n21631), .Z(n21633) );
  AND U23273 ( .A(n21634), .B(n21633), .Z(n21669) );
  NANDN U23274 ( .A(n21636), .B(n21635), .Z(n21640) );
  NANDN U23275 ( .A(n21638), .B(n21637), .Z(n21639) );
  AND U23276 ( .A(n21640), .B(n21639), .Z(n21667) );
  NAND U23277 ( .A(n42143), .B(n21641), .Z(n21643) );
  XNOR U23278 ( .A(a[469]), .B(n4138), .Z(n21678) );
  NAND U23279 ( .A(n42144), .B(n21678), .Z(n21642) );
  AND U23280 ( .A(n21643), .B(n21642), .Z(n21693) );
  XOR U23281 ( .A(a[473]), .B(n42012), .Z(n21681) );
  XNOR U23282 ( .A(n21693), .B(n21692), .Z(n21695) );
  XOR U23283 ( .A(a[471]), .B(n42085), .Z(n21685) );
  AND U23284 ( .A(a[467]), .B(b[7]), .Z(n21686) );
  XNOR U23285 ( .A(n21687), .B(n21686), .Z(n21688) );
  AND U23286 ( .A(a[475]), .B(b[0]), .Z(n21646) );
  XNOR U23287 ( .A(n21646), .B(n4071), .Z(n21648) );
  NANDN U23288 ( .A(b[0]), .B(a[474]), .Z(n21647) );
  NAND U23289 ( .A(n21648), .B(n21647), .Z(n21689) );
  XNOR U23290 ( .A(n21688), .B(n21689), .Z(n21694) );
  XOR U23291 ( .A(n21695), .B(n21694), .Z(n21673) );
  NANDN U23292 ( .A(n21650), .B(n21649), .Z(n21654) );
  NANDN U23293 ( .A(n21652), .B(n21651), .Z(n21653) );
  AND U23294 ( .A(n21654), .B(n21653), .Z(n21672) );
  XNOR U23295 ( .A(n21673), .B(n21672), .Z(n21674) );
  NANDN U23296 ( .A(n21656), .B(n21655), .Z(n21660) );
  NAND U23297 ( .A(n21658), .B(n21657), .Z(n21659) );
  NAND U23298 ( .A(n21660), .B(n21659), .Z(n21675) );
  XNOR U23299 ( .A(n21674), .B(n21675), .Z(n21666) );
  XNOR U23300 ( .A(n21667), .B(n21666), .Z(n21668) );
  XNOR U23301 ( .A(n21669), .B(n21668), .Z(n21698) );
  XNOR U23302 ( .A(sreg[1491]), .B(n21698), .Z(n21700) );
  NANDN U23303 ( .A(sreg[1490]), .B(n21661), .Z(n21665) );
  NAND U23304 ( .A(n21663), .B(n21662), .Z(n21664) );
  NAND U23305 ( .A(n21665), .B(n21664), .Z(n21699) );
  XNOR U23306 ( .A(n21700), .B(n21699), .Z(c[1491]) );
  NANDN U23307 ( .A(n21667), .B(n21666), .Z(n21671) );
  NANDN U23308 ( .A(n21669), .B(n21668), .Z(n21670) );
  AND U23309 ( .A(n21671), .B(n21670), .Z(n21706) );
  NANDN U23310 ( .A(n21673), .B(n21672), .Z(n21677) );
  NANDN U23311 ( .A(n21675), .B(n21674), .Z(n21676) );
  AND U23312 ( .A(n21677), .B(n21676), .Z(n21704) );
  NAND U23313 ( .A(n42143), .B(n21678), .Z(n21680) );
  XNOR U23314 ( .A(a[470]), .B(n4139), .Z(n21715) );
  NAND U23315 ( .A(n42144), .B(n21715), .Z(n21679) );
  AND U23316 ( .A(n21680), .B(n21679), .Z(n21730) );
  XOR U23317 ( .A(a[474]), .B(n42012), .Z(n21718) );
  XNOR U23318 ( .A(n21730), .B(n21729), .Z(n21732) );
  AND U23319 ( .A(a[476]), .B(b[0]), .Z(n21682) );
  XNOR U23320 ( .A(n21682), .B(n4071), .Z(n21684) );
  NANDN U23321 ( .A(b[0]), .B(a[475]), .Z(n21683) );
  NAND U23322 ( .A(n21684), .B(n21683), .Z(n21726) );
  XOR U23323 ( .A(a[472]), .B(n42085), .Z(n21722) );
  AND U23324 ( .A(a[468]), .B(b[7]), .Z(n21723) );
  XNOR U23325 ( .A(n21724), .B(n21723), .Z(n21725) );
  XNOR U23326 ( .A(n21726), .B(n21725), .Z(n21731) );
  XOR U23327 ( .A(n21732), .B(n21731), .Z(n21710) );
  NANDN U23328 ( .A(n21687), .B(n21686), .Z(n21691) );
  NANDN U23329 ( .A(n21689), .B(n21688), .Z(n21690) );
  AND U23330 ( .A(n21691), .B(n21690), .Z(n21709) );
  XNOR U23331 ( .A(n21710), .B(n21709), .Z(n21711) );
  NANDN U23332 ( .A(n21693), .B(n21692), .Z(n21697) );
  NAND U23333 ( .A(n21695), .B(n21694), .Z(n21696) );
  NAND U23334 ( .A(n21697), .B(n21696), .Z(n21712) );
  XNOR U23335 ( .A(n21711), .B(n21712), .Z(n21703) );
  XNOR U23336 ( .A(n21704), .B(n21703), .Z(n21705) );
  XNOR U23337 ( .A(n21706), .B(n21705), .Z(n21735) );
  XNOR U23338 ( .A(sreg[1492]), .B(n21735), .Z(n21737) );
  NANDN U23339 ( .A(sreg[1491]), .B(n21698), .Z(n21702) );
  NAND U23340 ( .A(n21700), .B(n21699), .Z(n21701) );
  NAND U23341 ( .A(n21702), .B(n21701), .Z(n21736) );
  XNOR U23342 ( .A(n21737), .B(n21736), .Z(c[1492]) );
  NANDN U23343 ( .A(n21704), .B(n21703), .Z(n21708) );
  NANDN U23344 ( .A(n21706), .B(n21705), .Z(n21707) );
  AND U23345 ( .A(n21708), .B(n21707), .Z(n21743) );
  NANDN U23346 ( .A(n21710), .B(n21709), .Z(n21714) );
  NANDN U23347 ( .A(n21712), .B(n21711), .Z(n21713) );
  AND U23348 ( .A(n21714), .B(n21713), .Z(n21741) );
  NAND U23349 ( .A(n42143), .B(n21715), .Z(n21717) );
  XNOR U23350 ( .A(a[471]), .B(n4139), .Z(n21752) );
  NAND U23351 ( .A(n42144), .B(n21752), .Z(n21716) );
  AND U23352 ( .A(n21717), .B(n21716), .Z(n21767) );
  XOR U23353 ( .A(a[475]), .B(n42012), .Z(n21755) );
  XNOR U23354 ( .A(n21767), .B(n21766), .Z(n21769) );
  AND U23355 ( .A(a[477]), .B(b[0]), .Z(n21719) );
  XNOR U23356 ( .A(n21719), .B(n4071), .Z(n21721) );
  NANDN U23357 ( .A(b[0]), .B(a[476]), .Z(n21720) );
  NAND U23358 ( .A(n21721), .B(n21720), .Z(n21763) );
  XOR U23359 ( .A(a[473]), .B(n42085), .Z(n21759) );
  AND U23360 ( .A(a[469]), .B(b[7]), .Z(n21760) );
  XNOR U23361 ( .A(n21761), .B(n21760), .Z(n21762) );
  XNOR U23362 ( .A(n21763), .B(n21762), .Z(n21768) );
  XOR U23363 ( .A(n21769), .B(n21768), .Z(n21747) );
  NANDN U23364 ( .A(n21724), .B(n21723), .Z(n21728) );
  NANDN U23365 ( .A(n21726), .B(n21725), .Z(n21727) );
  AND U23366 ( .A(n21728), .B(n21727), .Z(n21746) );
  XNOR U23367 ( .A(n21747), .B(n21746), .Z(n21748) );
  NANDN U23368 ( .A(n21730), .B(n21729), .Z(n21734) );
  NAND U23369 ( .A(n21732), .B(n21731), .Z(n21733) );
  NAND U23370 ( .A(n21734), .B(n21733), .Z(n21749) );
  XNOR U23371 ( .A(n21748), .B(n21749), .Z(n21740) );
  XNOR U23372 ( .A(n21741), .B(n21740), .Z(n21742) );
  XNOR U23373 ( .A(n21743), .B(n21742), .Z(n21772) );
  XNOR U23374 ( .A(sreg[1493]), .B(n21772), .Z(n21774) );
  NANDN U23375 ( .A(sreg[1492]), .B(n21735), .Z(n21739) );
  NAND U23376 ( .A(n21737), .B(n21736), .Z(n21738) );
  NAND U23377 ( .A(n21739), .B(n21738), .Z(n21773) );
  XNOR U23378 ( .A(n21774), .B(n21773), .Z(c[1493]) );
  NANDN U23379 ( .A(n21741), .B(n21740), .Z(n21745) );
  NANDN U23380 ( .A(n21743), .B(n21742), .Z(n21744) );
  AND U23381 ( .A(n21745), .B(n21744), .Z(n21780) );
  NANDN U23382 ( .A(n21747), .B(n21746), .Z(n21751) );
  NANDN U23383 ( .A(n21749), .B(n21748), .Z(n21750) );
  AND U23384 ( .A(n21751), .B(n21750), .Z(n21778) );
  NAND U23385 ( .A(n42143), .B(n21752), .Z(n21754) );
  XNOR U23386 ( .A(a[472]), .B(n4139), .Z(n21789) );
  NAND U23387 ( .A(n42144), .B(n21789), .Z(n21753) );
  AND U23388 ( .A(n21754), .B(n21753), .Z(n21804) );
  XOR U23389 ( .A(a[476]), .B(n42012), .Z(n21792) );
  XNOR U23390 ( .A(n21804), .B(n21803), .Z(n21806) );
  AND U23391 ( .A(a[478]), .B(b[0]), .Z(n21756) );
  XNOR U23392 ( .A(n21756), .B(n4071), .Z(n21758) );
  NANDN U23393 ( .A(b[0]), .B(a[477]), .Z(n21757) );
  NAND U23394 ( .A(n21758), .B(n21757), .Z(n21800) );
  XOR U23395 ( .A(a[474]), .B(n42085), .Z(n21793) );
  AND U23396 ( .A(a[470]), .B(b[7]), .Z(n21797) );
  XNOR U23397 ( .A(n21798), .B(n21797), .Z(n21799) );
  XNOR U23398 ( .A(n21800), .B(n21799), .Z(n21805) );
  XOR U23399 ( .A(n21806), .B(n21805), .Z(n21784) );
  NANDN U23400 ( .A(n21761), .B(n21760), .Z(n21765) );
  NANDN U23401 ( .A(n21763), .B(n21762), .Z(n21764) );
  AND U23402 ( .A(n21765), .B(n21764), .Z(n21783) );
  XNOR U23403 ( .A(n21784), .B(n21783), .Z(n21785) );
  NANDN U23404 ( .A(n21767), .B(n21766), .Z(n21771) );
  NAND U23405 ( .A(n21769), .B(n21768), .Z(n21770) );
  NAND U23406 ( .A(n21771), .B(n21770), .Z(n21786) );
  XNOR U23407 ( .A(n21785), .B(n21786), .Z(n21777) );
  XNOR U23408 ( .A(n21778), .B(n21777), .Z(n21779) );
  XNOR U23409 ( .A(n21780), .B(n21779), .Z(n21809) );
  XNOR U23410 ( .A(sreg[1494]), .B(n21809), .Z(n21811) );
  NANDN U23411 ( .A(sreg[1493]), .B(n21772), .Z(n21776) );
  NAND U23412 ( .A(n21774), .B(n21773), .Z(n21775) );
  NAND U23413 ( .A(n21776), .B(n21775), .Z(n21810) );
  XNOR U23414 ( .A(n21811), .B(n21810), .Z(c[1494]) );
  NANDN U23415 ( .A(n21778), .B(n21777), .Z(n21782) );
  NANDN U23416 ( .A(n21780), .B(n21779), .Z(n21781) );
  AND U23417 ( .A(n21782), .B(n21781), .Z(n21817) );
  NANDN U23418 ( .A(n21784), .B(n21783), .Z(n21788) );
  NANDN U23419 ( .A(n21786), .B(n21785), .Z(n21787) );
  AND U23420 ( .A(n21788), .B(n21787), .Z(n21815) );
  NAND U23421 ( .A(n42143), .B(n21789), .Z(n21791) );
  XNOR U23422 ( .A(a[473]), .B(n4139), .Z(n21826) );
  NAND U23423 ( .A(n42144), .B(n21826), .Z(n21790) );
  AND U23424 ( .A(n21791), .B(n21790), .Z(n21841) );
  XOR U23425 ( .A(a[477]), .B(n42012), .Z(n21829) );
  XNOR U23426 ( .A(n21841), .B(n21840), .Z(n21843) );
  XOR U23427 ( .A(a[475]), .B(n42085), .Z(n21833) );
  AND U23428 ( .A(a[471]), .B(b[7]), .Z(n21834) );
  XNOR U23429 ( .A(n21835), .B(n21834), .Z(n21836) );
  AND U23430 ( .A(a[479]), .B(b[0]), .Z(n21794) );
  XNOR U23431 ( .A(n21794), .B(n4071), .Z(n21796) );
  NANDN U23432 ( .A(b[0]), .B(a[478]), .Z(n21795) );
  NAND U23433 ( .A(n21796), .B(n21795), .Z(n21837) );
  XNOR U23434 ( .A(n21836), .B(n21837), .Z(n21842) );
  XOR U23435 ( .A(n21843), .B(n21842), .Z(n21821) );
  NANDN U23436 ( .A(n21798), .B(n21797), .Z(n21802) );
  NANDN U23437 ( .A(n21800), .B(n21799), .Z(n21801) );
  AND U23438 ( .A(n21802), .B(n21801), .Z(n21820) );
  XNOR U23439 ( .A(n21821), .B(n21820), .Z(n21822) );
  NANDN U23440 ( .A(n21804), .B(n21803), .Z(n21808) );
  NAND U23441 ( .A(n21806), .B(n21805), .Z(n21807) );
  NAND U23442 ( .A(n21808), .B(n21807), .Z(n21823) );
  XNOR U23443 ( .A(n21822), .B(n21823), .Z(n21814) );
  XNOR U23444 ( .A(n21815), .B(n21814), .Z(n21816) );
  XNOR U23445 ( .A(n21817), .B(n21816), .Z(n21846) );
  XNOR U23446 ( .A(sreg[1495]), .B(n21846), .Z(n21848) );
  NANDN U23447 ( .A(sreg[1494]), .B(n21809), .Z(n21813) );
  NAND U23448 ( .A(n21811), .B(n21810), .Z(n21812) );
  NAND U23449 ( .A(n21813), .B(n21812), .Z(n21847) );
  XNOR U23450 ( .A(n21848), .B(n21847), .Z(c[1495]) );
  NANDN U23451 ( .A(n21815), .B(n21814), .Z(n21819) );
  NANDN U23452 ( .A(n21817), .B(n21816), .Z(n21818) );
  AND U23453 ( .A(n21819), .B(n21818), .Z(n21854) );
  NANDN U23454 ( .A(n21821), .B(n21820), .Z(n21825) );
  NANDN U23455 ( .A(n21823), .B(n21822), .Z(n21824) );
  AND U23456 ( .A(n21825), .B(n21824), .Z(n21852) );
  NAND U23457 ( .A(n42143), .B(n21826), .Z(n21828) );
  XNOR U23458 ( .A(a[474]), .B(n4139), .Z(n21863) );
  NAND U23459 ( .A(n42144), .B(n21863), .Z(n21827) );
  AND U23460 ( .A(n21828), .B(n21827), .Z(n21878) );
  XOR U23461 ( .A(a[478]), .B(n42012), .Z(n21866) );
  XNOR U23462 ( .A(n21878), .B(n21877), .Z(n21880) );
  AND U23463 ( .A(a[480]), .B(b[0]), .Z(n21830) );
  XNOR U23464 ( .A(n21830), .B(n4071), .Z(n21832) );
  NANDN U23465 ( .A(b[0]), .B(a[479]), .Z(n21831) );
  NAND U23466 ( .A(n21832), .B(n21831), .Z(n21874) );
  XOR U23467 ( .A(a[476]), .B(n42085), .Z(n21870) );
  AND U23468 ( .A(a[472]), .B(b[7]), .Z(n21871) );
  XNOR U23469 ( .A(n21872), .B(n21871), .Z(n21873) );
  XNOR U23470 ( .A(n21874), .B(n21873), .Z(n21879) );
  XOR U23471 ( .A(n21880), .B(n21879), .Z(n21858) );
  NANDN U23472 ( .A(n21835), .B(n21834), .Z(n21839) );
  NANDN U23473 ( .A(n21837), .B(n21836), .Z(n21838) );
  AND U23474 ( .A(n21839), .B(n21838), .Z(n21857) );
  XNOR U23475 ( .A(n21858), .B(n21857), .Z(n21859) );
  NANDN U23476 ( .A(n21841), .B(n21840), .Z(n21845) );
  NAND U23477 ( .A(n21843), .B(n21842), .Z(n21844) );
  NAND U23478 ( .A(n21845), .B(n21844), .Z(n21860) );
  XNOR U23479 ( .A(n21859), .B(n21860), .Z(n21851) );
  XNOR U23480 ( .A(n21852), .B(n21851), .Z(n21853) );
  XNOR U23481 ( .A(n21854), .B(n21853), .Z(n21883) );
  XNOR U23482 ( .A(sreg[1496]), .B(n21883), .Z(n21885) );
  NANDN U23483 ( .A(sreg[1495]), .B(n21846), .Z(n21850) );
  NAND U23484 ( .A(n21848), .B(n21847), .Z(n21849) );
  NAND U23485 ( .A(n21850), .B(n21849), .Z(n21884) );
  XNOR U23486 ( .A(n21885), .B(n21884), .Z(c[1496]) );
  NANDN U23487 ( .A(n21852), .B(n21851), .Z(n21856) );
  NANDN U23488 ( .A(n21854), .B(n21853), .Z(n21855) );
  AND U23489 ( .A(n21856), .B(n21855), .Z(n21891) );
  NANDN U23490 ( .A(n21858), .B(n21857), .Z(n21862) );
  NANDN U23491 ( .A(n21860), .B(n21859), .Z(n21861) );
  AND U23492 ( .A(n21862), .B(n21861), .Z(n21889) );
  NAND U23493 ( .A(n42143), .B(n21863), .Z(n21865) );
  XNOR U23494 ( .A(a[475]), .B(n4139), .Z(n21900) );
  NAND U23495 ( .A(n42144), .B(n21900), .Z(n21864) );
  AND U23496 ( .A(n21865), .B(n21864), .Z(n21915) );
  XOR U23497 ( .A(a[479]), .B(n42012), .Z(n21903) );
  XNOR U23498 ( .A(n21915), .B(n21914), .Z(n21917) );
  AND U23499 ( .A(a[481]), .B(b[0]), .Z(n21867) );
  XNOR U23500 ( .A(n21867), .B(n4071), .Z(n21869) );
  NANDN U23501 ( .A(b[0]), .B(a[480]), .Z(n21868) );
  NAND U23502 ( .A(n21869), .B(n21868), .Z(n21911) );
  XOR U23503 ( .A(a[477]), .B(n42085), .Z(n21907) );
  AND U23504 ( .A(a[473]), .B(b[7]), .Z(n21908) );
  XNOR U23505 ( .A(n21909), .B(n21908), .Z(n21910) );
  XNOR U23506 ( .A(n21911), .B(n21910), .Z(n21916) );
  XOR U23507 ( .A(n21917), .B(n21916), .Z(n21895) );
  NANDN U23508 ( .A(n21872), .B(n21871), .Z(n21876) );
  NANDN U23509 ( .A(n21874), .B(n21873), .Z(n21875) );
  AND U23510 ( .A(n21876), .B(n21875), .Z(n21894) );
  XNOR U23511 ( .A(n21895), .B(n21894), .Z(n21896) );
  NANDN U23512 ( .A(n21878), .B(n21877), .Z(n21882) );
  NAND U23513 ( .A(n21880), .B(n21879), .Z(n21881) );
  NAND U23514 ( .A(n21882), .B(n21881), .Z(n21897) );
  XNOR U23515 ( .A(n21896), .B(n21897), .Z(n21888) );
  XNOR U23516 ( .A(n21889), .B(n21888), .Z(n21890) );
  XNOR U23517 ( .A(n21891), .B(n21890), .Z(n21920) );
  XNOR U23518 ( .A(sreg[1497]), .B(n21920), .Z(n21922) );
  NANDN U23519 ( .A(sreg[1496]), .B(n21883), .Z(n21887) );
  NAND U23520 ( .A(n21885), .B(n21884), .Z(n21886) );
  NAND U23521 ( .A(n21887), .B(n21886), .Z(n21921) );
  XNOR U23522 ( .A(n21922), .B(n21921), .Z(c[1497]) );
  NANDN U23523 ( .A(n21889), .B(n21888), .Z(n21893) );
  NANDN U23524 ( .A(n21891), .B(n21890), .Z(n21892) );
  AND U23525 ( .A(n21893), .B(n21892), .Z(n21928) );
  NANDN U23526 ( .A(n21895), .B(n21894), .Z(n21899) );
  NANDN U23527 ( .A(n21897), .B(n21896), .Z(n21898) );
  AND U23528 ( .A(n21899), .B(n21898), .Z(n21926) );
  NAND U23529 ( .A(n42143), .B(n21900), .Z(n21902) );
  XNOR U23530 ( .A(a[476]), .B(n4139), .Z(n21937) );
  NAND U23531 ( .A(n42144), .B(n21937), .Z(n21901) );
  AND U23532 ( .A(n21902), .B(n21901), .Z(n21952) );
  XOR U23533 ( .A(a[480]), .B(n42012), .Z(n21940) );
  XNOR U23534 ( .A(n21952), .B(n21951), .Z(n21954) );
  AND U23535 ( .A(a[482]), .B(b[0]), .Z(n21904) );
  XNOR U23536 ( .A(n21904), .B(n4071), .Z(n21906) );
  NANDN U23537 ( .A(b[0]), .B(a[481]), .Z(n21905) );
  NAND U23538 ( .A(n21906), .B(n21905), .Z(n21948) );
  XOR U23539 ( .A(a[478]), .B(n42085), .Z(n21941) );
  AND U23540 ( .A(a[474]), .B(b[7]), .Z(n21945) );
  XNOR U23541 ( .A(n21946), .B(n21945), .Z(n21947) );
  XNOR U23542 ( .A(n21948), .B(n21947), .Z(n21953) );
  XOR U23543 ( .A(n21954), .B(n21953), .Z(n21932) );
  NANDN U23544 ( .A(n21909), .B(n21908), .Z(n21913) );
  NANDN U23545 ( .A(n21911), .B(n21910), .Z(n21912) );
  AND U23546 ( .A(n21913), .B(n21912), .Z(n21931) );
  XNOR U23547 ( .A(n21932), .B(n21931), .Z(n21933) );
  NANDN U23548 ( .A(n21915), .B(n21914), .Z(n21919) );
  NAND U23549 ( .A(n21917), .B(n21916), .Z(n21918) );
  NAND U23550 ( .A(n21919), .B(n21918), .Z(n21934) );
  XNOR U23551 ( .A(n21933), .B(n21934), .Z(n21925) );
  XNOR U23552 ( .A(n21926), .B(n21925), .Z(n21927) );
  XNOR U23553 ( .A(n21928), .B(n21927), .Z(n21957) );
  XNOR U23554 ( .A(sreg[1498]), .B(n21957), .Z(n21959) );
  NANDN U23555 ( .A(sreg[1497]), .B(n21920), .Z(n21924) );
  NAND U23556 ( .A(n21922), .B(n21921), .Z(n21923) );
  NAND U23557 ( .A(n21924), .B(n21923), .Z(n21958) );
  XNOR U23558 ( .A(n21959), .B(n21958), .Z(c[1498]) );
  NANDN U23559 ( .A(n21926), .B(n21925), .Z(n21930) );
  NANDN U23560 ( .A(n21928), .B(n21927), .Z(n21929) );
  AND U23561 ( .A(n21930), .B(n21929), .Z(n21965) );
  NANDN U23562 ( .A(n21932), .B(n21931), .Z(n21936) );
  NANDN U23563 ( .A(n21934), .B(n21933), .Z(n21935) );
  AND U23564 ( .A(n21936), .B(n21935), .Z(n21963) );
  NAND U23565 ( .A(n42143), .B(n21937), .Z(n21939) );
  XNOR U23566 ( .A(a[477]), .B(n4140), .Z(n21974) );
  NAND U23567 ( .A(n42144), .B(n21974), .Z(n21938) );
  AND U23568 ( .A(n21939), .B(n21938), .Z(n21989) );
  XOR U23569 ( .A(a[481]), .B(n42012), .Z(n21977) );
  XNOR U23570 ( .A(n21989), .B(n21988), .Z(n21991) );
  XOR U23571 ( .A(a[479]), .B(n42085), .Z(n21981) );
  AND U23572 ( .A(a[475]), .B(b[7]), .Z(n21982) );
  XNOR U23573 ( .A(n21983), .B(n21982), .Z(n21984) );
  AND U23574 ( .A(a[483]), .B(b[0]), .Z(n21942) );
  XNOR U23575 ( .A(n21942), .B(n4071), .Z(n21944) );
  NANDN U23576 ( .A(b[0]), .B(a[482]), .Z(n21943) );
  NAND U23577 ( .A(n21944), .B(n21943), .Z(n21985) );
  XNOR U23578 ( .A(n21984), .B(n21985), .Z(n21990) );
  XOR U23579 ( .A(n21991), .B(n21990), .Z(n21969) );
  NANDN U23580 ( .A(n21946), .B(n21945), .Z(n21950) );
  NANDN U23581 ( .A(n21948), .B(n21947), .Z(n21949) );
  AND U23582 ( .A(n21950), .B(n21949), .Z(n21968) );
  XNOR U23583 ( .A(n21969), .B(n21968), .Z(n21970) );
  NANDN U23584 ( .A(n21952), .B(n21951), .Z(n21956) );
  NAND U23585 ( .A(n21954), .B(n21953), .Z(n21955) );
  NAND U23586 ( .A(n21956), .B(n21955), .Z(n21971) );
  XNOR U23587 ( .A(n21970), .B(n21971), .Z(n21962) );
  XNOR U23588 ( .A(n21963), .B(n21962), .Z(n21964) );
  XNOR U23589 ( .A(n21965), .B(n21964), .Z(n21994) );
  XNOR U23590 ( .A(sreg[1499]), .B(n21994), .Z(n21996) );
  NANDN U23591 ( .A(sreg[1498]), .B(n21957), .Z(n21961) );
  NAND U23592 ( .A(n21959), .B(n21958), .Z(n21960) );
  NAND U23593 ( .A(n21961), .B(n21960), .Z(n21995) );
  XNOR U23594 ( .A(n21996), .B(n21995), .Z(c[1499]) );
  NANDN U23595 ( .A(n21963), .B(n21962), .Z(n21967) );
  NANDN U23596 ( .A(n21965), .B(n21964), .Z(n21966) );
  AND U23597 ( .A(n21967), .B(n21966), .Z(n22002) );
  NANDN U23598 ( .A(n21969), .B(n21968), .Z(n21973) );
  NANDN U23599 ( .A(n21971), .B(n21970), .Z(n21972) );
  AND U23600 ( .A(n21973), .B(n21972), .Z(n22000) );
  NAND U23601 ( .A(n42143), .B(n21974), .Z(n21976) );
  XNOR U23602 ( .A(a[478]), .B(n4140), .Z(n22011) );
  NAND U23603 ( .A(n42144), .B(n22011), .Z(n21975) );
  AND U23604 ( .A(n21976), .B(n21975), .Z(n22026) );
  XOR U23605 ( .A(a[482]), .B(n42012), .Z(n22014) );
  XNOR U23606 ( .A(n22026), .B(n22025), .Z(n22028) );
  AND U23607 ( .A(a[484]), .B(b[0]), .Z(n21978) );
  XNOR U23608 ( .A(n21978), .B(n4071), .Z(n21980) );
  NANDN U23609 ( .A(b[0]), .B(a[483]), .Z(n21979) );
  NAND U23610 ( .A(n21980), .B(n21979), .Z(n22022) );
  XOR U23611 ( .A(a[480]), .B(n42085), .Z(n22018) );
  AND U23612 ( .A(a[476]), .B(b[7]), .Z(n22019) );
  XNOR U23613 ( .A(n22020), .B(n22019), .Z(n22021) );
  XNOR U23614 ( .A(n22022), .B(n22021), .Z(n22027) );
  XOR U23615 ( .A(n22028), .B(n22027), .Z(n22006) );
  NANDN U23616 ( .A(n21983), .B(n21982), .Z(n21987) );
  NANDN U23617 ( .A(n21985), .B(n21984), .Z(n21986) );
  AND U23618 ( .A(n21987), .B(n21986), .Z(n22005) );
  XNOR U23619 ( .A(n22006), .B(n22005), .Z(n22007) );
  NANDN U23620 ( .A(n21989), .B(n21988), .Z(n21993) );
  NAND U23621 ( .A(n21991), .B(n21990), .Z(n21992) );
  NAND U23622 ( .A(n21993), .B(n21992), .Z(n22008) );
  XNOR U23623 ( .A(n22007), .B(n22008), .Z(n21999) );
  XNOR U23624 ( .A(n22000), .B(n21999), .Z(n22001) );
  XNOR U23625 ( .A(n22002), .B(n22001), .Z(n22031) );
  XNOR U23626 ( .A(sreg[1500]), .B(n22031), .Z(n22033) );
  NANDN U23627 ( .A(sreg[1499]), .B(n21994), .Z(n21998) );
  NAND U23628 ( .A(n21996), .B(n21995), .Z(n21997) );
  NAND U23629 ( .A(n21998), .B(n21997), .Z(n22032) );
  XNOR U23630 ( .A(n22033), .B(n22032), .Z(c[1500]) );
  NANDN U23631 ( .A(n22000), .B(n21999), .Z(n22004) );
  NANDN U23632 ( .A(n22002), .B(n22001), .Z(n22003) );
  AND U23633 ( .A(n22004), .B(n22003), .Z(n22039) );
  NANDN U23634 ( .A(n22006), .B(n22005), .Z(n22010) );
  NANDN U23635 ( .A(n22008), .B(n22007), .Z(n22009) );
  AND U23636 ( .A(n22010), .B(n22009), .Z(n22037) );
  NAND U23637 ( .A(n42143), .B(n22011), .Z(n22013) );
  XNOR U23638 ( .A(a[479]), .B(n4140), .Z(n22048) );
  NAND U23639 ( .A(n42144), .B(n22048), .Z(n22012) );
  AND U23640 ( .A(n22013), .B(n22012), .Z(n22063) );
  XOR U23641 ( .A(a[483]), .B(n42012), .Z(n22051) );
  XNOR U23642 ( .A(n22063), .B(n22062), .Z(n22065) );
  AND U23643 ( .A(a[485]), .B(b[0]), .Z(n22015) );
  XNOR U23644 ( .A(n22015), .B(n4071), .Z(n22017) );
  NANDN U23645 ( .A(b[0]), .B(a[484]), .Z(n22016) );
  NAND U23646 ( .A(n22017), .B(n22016), .Z(n22059) );
  XOR U23647 ( .A(a[481]), .B(n42085), .Z(n22052) );
  AND U23648 ( .A(a[477]), .B(b[7]), .Z(n22056) );
  XNOR U23649 ( .A(n22057), .B(n22056), .Z(n22058) );
  XNOR U23650 ( .A(n22059), .B(n22058), .Z(n22064) );
  XOR U23651 ( .A(n22065), .B(n22064), .Z(n22043) );
  NANDN U23652 ( .A(n22020), .B(n22019), .Z(n22024) );
  NANDN U23653 ( .A(n22022), .B(n22021), .Z(n22023) );
  AND U23654 ( .A(n22024), .B(n22023), .Z(n22042) );
  XNOR U23655 ( .A(n22043), .B(n22042), .Z(n22044) );
  NANDN U23656 ( .A(n22026), .B(n22025), .Z(n22030) );
  NAND U23657 ( .A(n22028), .B(n22027), .Z(n22029) );
  NAND U23658 ( .A(n22030), .B(n22029), .Z(n22045) );
  XNOR U23659 ( .A(n22044), .B(n22045), .Z(n22036) );
  XNOR U23660 ( .A(n22037), .B(n22036), .Z(n22038) );
  XNOR U23661 ( .A(n22039), .B(n22038), .Z(n22068) );
  XNOR U23662 ( .A(sreg[1501]), .B(n22068), .Z(n22070) );
  NANDN U23663 ( .A(sreg[1500]), .B(n22031), .Z(n22035) );
  NAND U23664 ( .A(n22033), .B(n22032), .Z(n22034) );
  NAND U23665 ( .A(n22035), .B(n22034), .Z(n22069) );
  XNOR U23666 ( .A(n22070), .B(n22069), .Z(c[1501]) );
  NANDN U23667 ( .A(n22037), .B(n22036), .Z(n22041) );
  NANDN U23668 ( .A(n22039), .B(n22038), .Z(n22040) );
  AND U23669 ( .A(n22041), .B(n22040), .Z(n22076) );
  NANDN U23670 ( .A(n22043), .B(n22042), .Z(n22047) );
  NANDN U23671 ( .A(n22045), .B(n22044), .Z(n22046) );
  AND U23672 ( .A(n22047), .B(n22046), .Z(n22074) );
  NAND U23673 ( .A(n42143), .B(n22048), .Z(n22050) );
  XNOR U23674 ( .A(a[480]), .B(n4140), .Z(n22085) );
  NAND U23675 ( .A(n42144), .B(n22085), .Z(n22049) );
  AND U23676 ( .A(n22050), .B(n22049), .Z(n22100) );
  XOR U23677 ( .A(a[484]), .B(n42012), .Z(n22088) );
  XNOR U23678 ( .A(n22100), .B(n22099), .Z(n22102) );
  XOR U23679 ( .A(a[482]), .B(n42085), .Z(n22092) );
  AND U23680 ( .A(a[478]), .B(b[7]), .Z(n22093) );
  XNOR U23681 ( .A(n22094), .B(n22093), .Z(n22095) );
  AND U23682 ( .A(a[486]), .B(b[0]), .Z(n22053) );
  XNOR U23683 ( .A(n22053), .B(n4071), .Z(n22055) );
  NANDN U23684 ( .A(b[0]), .B(a[485]), .Z(n22054) );
  NAND U23685 ( .A(n22055), .B(n22054), .Z(n22096) );
  XNOR U23686 ( .A(n22095), .B(n22096), .Z(n22101) );
  XOR U23687 ( .A(n22102), .B(n22101), .Z(n22080) );
  NANDN U23688 ( .A(n22057), .B(n22056), .Z(n22061) );
  NANDN U23689 ( .A(n22059), .B(n22058), .Z(n22060) );
  AND U23690 ( .A(n22061), .B(n22060), .Z(n22079) );
  XNOR U23691 ( .A(n22080), .B(n22079), .Z(n22081) );
  NANDN U23692 ( .A(n22063), .B(n22062), .Z(n22067) );
  NAND U23693 ( .A(n22065), .B(n22064), .Z(n22066) );
  NAND U23694 ( .A(n22067), .B(n22066), .Z(n22082) );
  XNOR U23695 ( .A(n22081), .B(n22082), .Z(n22073) );
  XNOR U23696 ( .A(n22074), .B(n22073), .Z(n22075) );
  XNOR U23697 ( .A(n22076), .B(n22075), .Z(n22105) );
  XNOR U23698 ( .A(sreg[1502]), .B(n22105), .Z(n22107) );
  NANDN U23699 ( .A(sreg[1501]), .B(n22068), .Z(n22072) );
  NAND U23700 ( .A(n22070), .B(n22069), .Z(n22071) );
  NAND U23701 ( .A(n22072), .B(n22071), .Z(n22106) );
  XNOR U23702 ( .A(n22107), .B(n22106), .Z(c[1502]) );
  NANDN U23703 ( .A(n22074), .B(n22073), .Z(n22078) );
  NANDN U23704 ( .A(n22076), .B(n22075), .Z(n22077) );
  AND U23705 ( .A(n22078), .B(n22077), .Z(n22113) );
  NANDN U23706 ( .A(n22080), .B(n22079), .Z(n22084) );
  NANDN U23707 ( .A(n22082), .B(n22081), .Z(n22083) );
  AND U23708 ( .A(n22084), .B(n22083), .Z(n22111) );
  NAND U23709 ( .A(n42143), .B(n22085), .Z(n22087) );
  XNOR U23710 ( .A(a[481]), .B(n4140), .Z(n22122) );
  NAND U23711 ( .A(n42144), .B(n22122), .Z(n22086) );
  AND U23712 ( .A(n22087), .B(n22086), .Z(n22137) );
  XOR U23713 ( .A(a[485]), .B(n42012), .Z(n22125) );
  XNOR U23714 ( .A(n22137), .B(n22136), .Z(n22139) );
  AND U23715 ( .A(a[487]), .B(b[0]), .Z(n22089) );
  XNOR U23716 ( .A(n22089), .B(n4071), .Z(n22091) );
  NANDN U23717 ( .A(b[0]), .B(a[486]), .Z(n22090) );
  NAND U23718 ( .A(n22091), .B(n22090), .Z(n22133) );
  XOR U23719 ( .A(a[483]), .B(n42085), .Z(n22126) );
  AND U23720 ( .A(a[479]), .B(b[7]), .Z(n22130) );
  XNOR U23721 ( .A(n22131), .B(n22130), .Z(n22132) );
  XNOR U23722 ( .A(n22133), .B(n22132), .Z(n22138) );
  XOR U23723 ( .A(n22139), .B(n22138), .Z(n22117) );
  NANDN U23724 ( .A(n22094), .B(n22093), .Z(n22098) );
  NANDN U23725 ( .A(n22096), .B(n22095), .Z(n22097) );
  AND U23726 ( .A(n22098), .B(n22097), .Z(n22116) );
  XNOR U23727 ( .A(n22117), .B(n22116), .Z(n22118) );
  NANDN U23728 ( .A(n22100), .B(n22099), .Z(n22104) );
  NAND U23729 ( .A(n22102), .B(n22101), .Z(n22103) );
  NAND U23730 ( .A(n22104), .B(n22103), .Z(n22119) );
  XNOR U23731 ( .A(n22118), .B(n22119), .Z(n22110) );
  XNOR U23732 ( .A(n22111), .B(n22110), .Z(n22112) );
  XNOR U23733 ( .A(n22113), .B(n22112), .Z(n22142) );
  XNOR U23734 ( .A(sreg[1503]), .B(n22142), .Z(n22144) );
  NANDN U23735 ( .A(sreg[1502]), .B(n22105), .Z(n22109) );
  NAND U23736 ( .A(n22107), .B(n22106), .Z(n22108) );
  NAND U23737 ( .A(n22109), .B(n22108), .Z(n22143) );
  XNOR U23738 ( .A(n22144), .B(n22143), .Z(c[1503]) );
  NANDN U23739 ( .A(n22111), .B(n22110), .Z(n22115) );
  NANDN U23740 ( .A(n22113), .B(n22112), .Z(n22114) );
  AND U23741 ( .A(n22115), .B(n22114), .Z(n22150) );
  NANDN U23742 ( .A(n22117), .B(n22116), .Z(n22121) );
  NANDN U23743 ( .A(n22119), .B(n22118), .Z(n22120) );
  AND U23744 ( .A(n22121), .B(n22120), .Z(n22148) );
  NAND U23745 ( .A(n42143), .B(n22122), .Z(n22124) );
  XNOR U23746 ( .A(a[482]), .B(n4140), .Z(n22159) );
  NAND U23747 ( .A(n42144), .B(n22159), .Z(n22123) );
  AND U23748 ( .A(n22124), .B(n22123), .Z(n22174) );
  XOR U23749 ( .A(a[486]), .B(n42012), .Z(n22162) );
  XNOR U23750 ( .A(n22174), .B(n22173), .Z(n22176) );
  XOR U23751 ( .A(a[484]), .B(n42085), .Z(n22166) );
  AND U23752 ( .A(a[480]), .B(b[7]), .Z(n22167) );
  XNOR U23753 ( .A(n22168), .B(n22167), .Z(n22169) );
  AND U23754 ( .A(a[488]), .B(b[0]), .Z(n22127) );
  XNOR U23755 ( .A(n22127), .B(n4071), .Z(n22129) );
  NANDN U23756 ( .A(b[0]), .B(a[487]), .Z(n22128) );
  NAND U23757 ( .A(n22129), .B(n22128), .Z(n22170) );
  XNOR U23758 ( .A(n22169), .B(n22170), .Z(n22175) );
  XOR U23759 ( .A(n22176), .B(n22175), .Z(n22154) );
  NANDN U23760 ( .A(n22131), .B(n22130), .Z(n22135) );
  NANDN U23761 ( .A(n22133), .B(n22132), .Z(n22134) );
  AND U23762 ( .A(n22135), .B(n22134), .Z(n22153) );
  XNOR U23763 ( .A(n22154), .B(n22153), .Z(n22155) );
  NANDN U23764 ( .A(n22137), .B(n22136), .Z(n22141) );
  NAND U23765 ( .A(n22139), .B(n22138), .Z(n22140) );
  NAND U23766 ( .A(n22141), .B(n22140), .Z(n22156) );
  XNOR U23767 ( .A(n22155), .B(n22156), .Z(n22147) );
  XNOR U23768 ( .A(n22148), .B(n22147), .Z(n22149) );
  XNOR U23769 ( .A(n22150), .B(n22149), .Z(n22179) );
  XNOR U23770 ( .A(sreg[1504]), .B(n22179), .Z(n22181) );
  NANDN U23771 ( .A(sreg[1503]), .B(n22142), .Z(n22146) );
  NAND U23772 ( .A(n22144), .B(n22143), .Z(n22145) );
  NAND U23773 ( .A(n22146), .B(n22145), .Z(n22180) );
  XNOR U23774 ( .A(n22181), .B(n22180), .Z(c[1504]) );
  NANDN U23775 ( .A(n22148), .B(n22147), .Z(n22152) );
  NANDN U23776 ( .A(n22150), .B(n22149), .Z(n22151) );
  AND U23777 ( .A(n22152), .B(n22151), .Z(n22187) );
  NANDN U23778 ( .A(n22154), .B(n22153), .Z(n22158) );
  NANDN U23779 ( .A(n22156), .B(n22155), .Z(n22157) );
  AND U23780 ( .A(n22158), .B(n22157), .Z(n22185) );
  NAND U23781 ( .A(n42143), .B(n22159), .Z(n22161) );
  XNOR U23782 ( .A(a[483]), .B(n4140), .Z(n22196) );
  NAND U23783 ( .A(n42144), .B(n22196), .Z(n22160) );
  AND U23784 ( .A(n22161), .B(n22160), .Z(n22211) );
  XOR U23785 ( .A(a[487]), .B(n42012), .Z(n22199) );
  XNOR U23786 ( .A(n22211), .B(n22210), .Z(n22213) );
  AND U23787 ( .A(a[489]), .B(b[0]), .Z(n22163) );
  XNOR U23788 ( .A(n22163), .B(n4071), .Z(n22165) );
  NANDN U23789 ( .A(b[0]), .B(a[488]), .Z(n22164) );
  NAND U23790 ( .A(n22165), .B(n22164), .Z(n22207) );
  XOR U23791 ( .A(a[485]), .B(n42085), .Z(n22203) );
  AND U23792 ( .A(a[481]), .B(b[7]), .Z(n22204) );
  XNOR U23793 ( .A(n22205), .B(n22204), .Z(n22206) );
  XNOR U23794 ( .A(n22207), .B(n22206), .Z(n22212) );
  XOR U23795 ( .A(n22213), .B(n22212), .Z(n22191) );
  NANDN U23796 ( .A(n22168), .B(n22167), .Z(n22172) );
  NANDN U23797 ( .A(n22170), .B(n22169), .Z(n22171) );
  AND U23798 ( .A(n22172), .B(n22171), .Z(n22190) );
  XNOR U23799 ( .A(n22191), .B(n22190), .Z(n22192) );
  NANDN U23800 ( .A(n22174), .B(n22173), .Z(n22178) );
  NAND U23801 ( .A(n22176), .B(n22175), .Z(n22177) );
  NAND U23802 ( .A(n22178), .B(n22177), .Z(n22193) );
  XNOR U23803 ( .A(n22192), .B(n22193), .Z(n22184) );
  XNOR U23804 ( .A(n22185), .B(n22184), .Z(n22186) );
  XNOR U23805 ( .A(n22187), .B(n22186), .Z(n22216) );
  XNOR U23806 ( .A(sreg[1505]), .B(n22216), .Z(n22218) );
  NANDN U23807 ( .A(sreg[1504]), .B(n22179), .Z(n22183) );
  NAND U23808 ( .A(n22181), .B(n22180), .Z(n22182) );
  NAND U23809 ( .A(n22183), .B(n22182), .Z(n22217) );
  XNOR U23810 ( .A(n22218), .B(n22217), .Z(c[1505]) );
  NANDN U23811 ( .A(n22185), .B(n22184), .Z(n22189) );
  NANDN U23812 ( .A(n22187), .B(n22186), .Z(n22188) );
  AND U23813 ( .A(n22189), .B(n22188), .Z(n22224) );
  NANDN U23814 ( .A(n22191), .B(n22190), .Z(n22195) );
  NANDN U23815 ( .A(n22193), .B(n22192), .Z(n22194) );
  AND U23816 ( .A(n22195), .B(n22194), .Z(n22222) );
  NAND U23817 ( .A(n42143), .B(n22196), .Z(n22198) );
  XNOR U23818 ( .A(a[484]), .B(n4141), .Z(n22233) );
  NAND U23819 ( .A(n42144), .B(n22233), .Z(n22197) );
  AND U23820 ( .A(n22198), .B(n22197), .Z(n22248) );
  XOR U23821 ( .A(a[488]), .B(n42012), .Z(n22236) );
  XNOR U23822 ( .A(n22248), .B(n22247), .Z(n22250) );
  AND U23823 ( .A(a[490]), .B(b[0]), .Z(n22200) );
  XNOR U23824 ( .A(n22200), .B(n4071), .Z(n22202) );
  NANDN U23825 ( .A(b[0]), .B(a[489]), .Z(n22201) );
  NAND U23826 ( .A(n22202), .B(n22201), .Z(n22244) );
  XOR U23827 ( .A(a[486]), .B(n42085), .Z(n22237) );
  AND U23828 ( .A(a[482]), .B(b[7]), .Z(n22241) );
  XNOR U23829 ( .A(n22242), .B(n22241), .Z(n22243) );
  XNOR U23830 ( .A(n22244), .B(n22243), .Z(n22249) );
  XOR U23831 ( .A(n22250), .B(n22249), .Z(n22228) );
  NANDN U23832 ( .A(n22205), .B(n22204), .Z(n22209) );
  NANDN U23833 ( .A(n22207), .B(n22206), .Z(n22208) );
  AND U23834 ( .A(n22209), .B(n22208), .Z(n22227) );
  XNOR U23835 ( .A(n22228), .B(n22227), .Z(n22229) );
  NANDN U23836 ( .A(n22211), .B(n22210), .Z(n22215) );
  NAND U23837 ( .A(n22213), .B(n22212), .Z(n22214) );
  NAND U23838 ( .A(n22215), .B(n22214), .Z(n22230) );
  XNOR U23839 ( .A(n22229), .B(n22230), .Z(n22221) );
  XNOR U23840 ( .A(n22222), .B(n22221), .Z(n22223) );
  XNOR U23841 ( .A(n22224), .B(n22223), .Z(n22253) );
  XNOR U23842 ( .A(sreg[1506]), .B(n22253), .Z(n22255) );
  NANDN U23843 ( .A(sreg[1505]), .B(n22216), .Z(n22220) );
  NAND U23844 ( .A(n22218), .B(n22217), .Z(n22219) );
  NAND U23845 ( .A(n22220), .B(n22219), .Z(n22254) );
  XNOR U23846 ( .A(n22255), .B(n22254), .Z(c[1506]) );
  NANDN U23847 ( .A(n22222), .B(n22221), .Z(n22226) );
  NANDN U23848 ( .A(n22224), .B(n22223), .Z(n22225) );
  AND U23849 ( .A(n22226), .B(n22225), .Z(n22261) );
  NANDN U23850 ( .A(n22228), .B(n22227), .Z(n22232) );
  NANDN U23851 ( .A(n22230), .B(n22229), .Z(n22231) );
  AND U23852 ( .A(n22232), .B(n22231), .Z(n22259) );
  NAND U23853 ( .A(n42143), .B(n22233), .Z(n22235) );
  XNOR U23854 ( .A(a[485]), .B(n4141), .Z(n22270) );
  NAND U23855 ( .A(n42144), .B(n22270), .Z(n22234) );
  AND U23856 ( .A(n22235), .B(n22234), .Z(n22285) );
  XOR U23857 ( .A(a[489]), .B(n42012), .Z(n22273) );
  XNOR U23858 ( .A(n22285), .B(n22284), .Z(n22287) );
  XOR U23859 ( .A(a[487]), .B(n42085), .Z(n22277) );
  AND U23860 ( .A(a[483]), .B(b[7]), .Z(n22278) );
  XNOR U23861 ( .A(n22279), .B(n22278), .Z(n22280) );
  AND U23862 ( .A(a[491]), .B(b[0]), .Z(n22238) );
  XNOR U23863 ( .A(n22238), .B(n4071), .Z(n22240) );
  NANDN U23864 ( .A(b[0]), .B(a[490]), .Z(n22239) );
  NAND U23865 ( .A(n22240), .B(n22239), .Z(n22281) );
  XNOR U23866 ( .A(n22280), .B(n22281), .Z(n22286) );
  XOR U23867 ( .A(n22287), .B(n22286), .Z(n22265) );
  NANDN U23868 ( .A(n22242), .B(n22241), .Z(n22246) );
  NANDN U23869 ( .A(n22244), .B(n22243), .Z(n22245) );
  AND U23870 ( .A(n22246), .B(n22245), .Z(n22264) );
  XNOR U23871 ( .A(n22265), .B(n22264), .Z(n22266) );
  NANDN U23872 ( .A(n22248), .B(n22247), .Z(n22252) );
  NAND U23873 ( .A(n22250), .B(n22249), .Z(n22251) );
  NAND U23874 ( .A(n22252), .B(n22251), .Z(n22267) );
  XNOR U23875 ( .A(n22266), .B(n22267), .Z(n22258) );
  XNOR U23876 ( .A(n22259), .B(n22258), .Z(n22260) );
  XNOR U23877 ( .A(n22261), .B(n22260), .Z(n22290) );
  XNOR U23878 ( .A(sreg[1507]), .B(n22290), .Z(n22292) );
  NANDN U23879 ( .A(sreg[1506]), .B(n22253), .Z(n22257) );
  NAND U23880 ( .A(n22255), .B(n22254), .Z(n22256) );
  NAND U23881 ( .A(n22257), .B(n22256), .Z(n22291) );
  XNOR U23882 ( .A(n22292), .B(n22291), .Z(c[1507]) );
  NANDN U23883 ( .A(n22259), .B(n22258), .Z(n22263) );
  NANDN U23884 ( .A(n22261), .B(n22260), .Z(n22262) );
  AND U23885 ( .A(n22263), .B(n22262), .Z(n22298) );
  NANDN U23886 ( .A(n22265), .B(n22264), .Z(n22269) );
  NANDN U23887 ( .A(n22267), .B(n22266), .Z(n22268) );
  AND U23888 ( .A(n22269), .B(n22268), .Z(n22296) );
  NAND U23889 ( .A(n42143), .B(n22270), .Z(n22272) );
  XNOR U23890 ( .A(a[486]), .B(n4141), .Z(n22307) );
  NAND U23891 ( .A(n42144), .B(n22307), .Z(n22271) );
  AND U23892 ( .A(n22272), .B(n22271), .Z(n22322) );
  XOR U23893 ( .A(a[490]), .B(n42012), .Z(n22310) );
  XNOR U23894 ( .A(n22322), .B(n22321), .Z(n22324) );
  AND U23895 ( .A(a[492]), .B(b[0]), .Z(n22274) );
  XNOR U23896 ( .A(n22274), .B(n4071), .Z(n22276) );
  NANDN U23897 ( .A(b[0]), .B(a[491]), .Z(n22275) );
  NAND U23898 ( .A(n22276), .B(n22275), .Z(n22318) );
  XOR U23899 ( .A(a[488]), .B(n42085), .Z(n22314) );
  AND U23900 ( .A(a[484]), .B(b[7]), .Z(n22315) );
  XNOR U23901 ( .A(n22316), .B(n22315), .Z(n22317) );
  XNOR U23902 ( .A(n22318), .B(n22317), .Z(n22323) );
  XOR U23903 ( .A(n22324), .B(n22323), .Z(n22302) );
  NANDN U23904 ( .A(n22279), .B(n22278), .Z(n22283) );
  NANDN U23905 ( .A(n22281), .B(n22280), .Z(n22282) );
  AND U23906 ( .A(n22283), .B(n22282), .Z(n22301) );
  XNOR U23907 ( .A(n22302), .B(n22301), .Z(n22303) );
  NANDN U23908 ( .A(n22285), .B(n22284), .Z(n22289) );
  NAND U23909 ( .A(n22287), .B(n22286), .Z(n22288) );
  NAND U23910 ( .A(n22289), .B(n22288), .Z(n22304) );
  XNOR U23911 ( .A(n22303), .B(n22304), .Z(n22295) );
  XNOR U23912 ( .A(n22296), .B(n22295), .Z(n22297) );
  XNOR U23913 ( .A(n22298), .B(n22297), .Z(n22327) );
  XNOR U23914 ( .A(sreg[1508]), .B(n22327), .Z(n22329) );
  NANDN U23915 ( .A(sreg[1507]), .B(n22290), .Z(n22294) );
  NAND U23916 ( .A(n22292), .B(n22291), .Z(n22293) );
  NAND U23917 ( .A(n22294), .B(n22293), .Z(n22328) );
  XNOR U23918 ( .A(n22329), .B(n22328), .Z(c[1508]) );
  NANDN U23919 ( .A(n22296), .B(n22295), .Z(n22300) );
  NANDN U23920 ( .A(n22298), .B(n22297), .Z(n22299) );
  AND U23921 ( .A(n22300), .B(n22299), .Z(n22335) );
  NANDN U23922 ( .A(n22302), .B(n22301), .Z(n22306) );
  NANDN U23923 ( .A(n22304), .B(n22303), .Z(n22305) );
  AND U23924 ( .A(n22306), .B(n22305), .Z(n22333) );
  NAND U23925 ( .A(n42143), .B(n22307), .Z(n22309) );
  XNOR U23926 ( .A(a[487]), .B(n4141), .Z(n22344) );
  NAND U23927 ( .A(n42144), .B(n22344), .Z(n22308) );
  AND U23928 ( .A(n22309), .B(n22308), .Z(n22359) );
  XOR U23929 ( .A(a[491]), .B(n42012), .Z(n22347) );
  XNOR U23930 ( .A(n22359), .B(n22358), .Z(n22361) );
  AND U23931 ( .A(a[493]), .B(b[0]), .Z(n22311) );
  XNOR U23932 ( .A(n22311), .B(n4071), .Z(n22313) );
  NANDN U23933 ( .A(b[0]), .B(a[492]), .Z(n22312) );
  NAND U23934 ( .A(n22313), .B(n22312), .Z(n22355) );
  XOR U23935 ( .A(a[489]), .B(n42085), .Z(n22351) );
  AND U23936 ( .A(a[485]), .B(b[7]), .Z(n22352) );
  XNOR U23937 ( .A(n22353), .B(n22352), .Z(n22354) );
  XNOR U23938 ( .A(n22355), .B(n22354), .Z(n22360) );
  XOR U23939 ( .A(n22361), .B(n22360), .Z(n22339) );
  NANDN U23940 ( .A(n22316), .B(n22315), .Z(n22320) );
  NANDN U23941 ( .A(n22318), .B(n22317), .Z(n22319) );
  AND U23942 ( .A(n22320), .B(n22319), .Z(n22338) );
  XNOR U23943 ( .A(n22339), .B(n22338), .Z(n22340) );
  NANDN U23944 ( .A(n22322), .B(n22321), .Z(n22326) );
  NAND U23945 ( .A(n22324), .B(n22323), .Z(n22325) );
  NAND U23946 ( .A(n22326), .B(n22325), .Z(n22341) );
  XNOR U23947 ( .A(n22340), .B(n22341), .Z(n22332) );
  XNOR U23948 ( .A(n22333), .B(n22332), .Z(n22334) );
  XNOR U23949 ( .A(n22335), .B(n22334), .Z(n22364) );
  XNOR U23950 ( .A(sreg[1509]), .B(n22364), .Z(n22366) );
  NANDN U23951 ( .A(sreg[1508]), .B(n22327), .Z(n22331) );
  NAND U23952 ( .A(n22329), .B(n22328), .Z(n22330) );
  NAND U23953 ( .A(n22331), .B(n22330), .Z(n22365) );
  XNOR U23954 ( .A(n22366), .B(n22365), .Z(c[1509]) );
  NANDN U23955 ( .A(n22333), .B(n22332), .Z(n22337) );
  NANDN U23956 ( .A(n22335), .B(n22334), .Z(n22336) );
  AND U23957 ( .A(n22337), .B(n22336), .Z(n22372) );
  NANDN U23958 ( .A(n22339), .B(n22338), .Z(n22343) );
  NANDN U23959 ( .A(n22341), .B(n22340), .Z(n22342) );
  AND U23960 ( .A(n22343), .B(n22342), .Z(n22370) );
  NAND U23961 ( .A(n42143), .B(n22344), .Z(n22346) );
  XNOR U23962 ( .A(a[488]), .B(n4141), .Z(n22381) );
  NAND U23963 ( .A(n42144), .B(n22381), .Z(n22345) );
  AND U23964 ( .A(n22346), .B(n22345), .Z(n22396) );
  XOR U23965 ( .A(a[492]), .B(n42012), .Z(n22384) );
  XNOR U23966 ( .A(n22396), .B(n22395), .Z(n22398) );
  AND U23967 ( .A(a[494]), .B(b[0]), .Z(n22348) );
  XNOR U23968 ( .A(n22348), .B(n4071), .Z(n22350) );
  NANDN U23969 ( .A(b[0]), .B(a[493]), .Z(n22349) );
  NAND U23970 ( .A(n22350), .B(n22349), .Z(n22392) );
  XOR U23971 ( .A(a[490]), .B(n42085), .Z(n22388) );
  AND U23972 ( .A(a[486]), .B(b[7]), .Z(n22389) );
  XNOR U23973 ( .A(n22390), .B(n22389), .Z(n22391) );
  XNOR U23974 ( .A(n22392), .B(n22391), .Z(n22397) );
  XOR U23975 ( .A(n22398), .B(n22397), .Z(n22376) );
  NANDN U23976 ( .A(n22353), .B(n22352), .Z(n22357) );
  NANDN U23977 ( .A(n22355), .B(n22354), .Z(n22356) );
  AND U23978 ( .A(n22357), .B(n22356), .Z(n22375) );
  XNOR U23979 ( .A(n22376), .B(n22375), .Z(n22377) );
  NANDN U23980 ( .A(n22359), .B(n22358), .Z(n22363) );
  NAND U23981 ( .A(n22361), .B(n22360), .Z(n22362) );
  NAND U23982 ( .A(n22363), .B(n22362), .Z(n22378) );
  XNOR U23983 ( .A(n22377), .B(n22378), .Z(n22369) );
  XNOR U23984 ( .A(n22370), .B(n22369), .Z(n22371) );
  XNOR U23985 ( .A(n22372), .B(n22371), .Z(n22401) );
  XNOR U23986 ( .A(sreg[1510]), .B(n22401), .Z(n22403) );
  NANDN U23987 ( .A(sreg[1509]), .B(n22364), .Z(n22368) );
  NAND U23988 ( .A(n22366), .B(n22365), .Z(n22367) );
  NAND U23989 ( .A(n22368), .B(n22367), .Z(n22402) );
  XNOR U23990 ( .A(n22403), .B(n22402), .Z(c[1510]) );
  NANDN U23991 ( .A(n22370), .B(n22369), .Z(n22374) );
  NANDN U23992 ( .A(n22372), .B(n22371), .Z(n22373) );
  AND U23993 ( .A(n22374), .B(n22373), .Z(n22409) );
  NANDN U23994 ( .A(n22376), .B(n22375), .Z(n22380) );
  NANDN U23995 ( .A(n22378), .B(n22377), .Z(n22379) );
  AND U23996 ( .A(n22380), .B(n22379), .Z(n22407) );
  NAND U23997 ( .A(n42143), .B(n22381), .Z(n22383) );
  XNOR U23998 ( .A(a[489]), .B(n4141), .Z(n22418) );
  NAND U23999 ( .A(n42144), .B(n22418), .Z(n22382) );
  AND U24000 ( .A(n22383), .B(n22382), .Z(n22433) );
  XOR U24001 ( .A(a[493]), .B(n42012), .Z(n22421) );
  XNOR U24002 ( .A(n22433), .B(n22432), .Z(n22435) );
  AND U24003 ( .A(a[495]), .B(b[0]), .Z(n22385) );
  XNOR U24004 ( .A(n22385), .B(n4071), .Z(n22387) );
  NANDN U24005 ( .A(b[0]), .B(a[494]), .Z(n22386) );
  NAND U24006 ( .A(n22387), .B(n22386), .Z(n22429) );
  XOR U24007 ( .A(a[491]), .B(n42085), .Z(n22425) );
  AND U24008 ( .A(a[487]), .B(b[7]), .Z(n22426) );
  XNOR U24009 ( .A(n22427), .B(n22426), .Z(n22428) );
  XNOR U24010 ( .A(n22429), .B(n22428), .Z(n22434) );
  XOR U24011 ( .A(n22435), .B(n22434), .Z(n22413) );
  NANDN U24012 ( .A(n22390), .B(n22389), .Z(n22394) );
  NANDN U24013 ( .A(n22392), .B(n22391), .Z(n22393) );
  AND U24014 ( .A(n22394), .B(n22393), .Z(n22412) );
  XNOR U24015 ( .A(n22413), .B(n22412), .Z(n22414) );
  NANDN U24016 ( .A(n22396), .B(n22395), .Z(n22400) );
  NAND U24017 ( .A(n22398), .B(n22397), .Z(n22399) );
  NAND U24018 ( .A(n22400), .B(n22399), .Z(n22415) );
  XNOR U24019 ( .A(n22414), .B(n22415), .Z(n22406) );
  XNOR U24020 ( .A(n22407), .B(n22406), .Z(n22408) );
  XNOR U24021 ( .A(n22409), .B(n22408), .Z(n22438) );
  XNOR U24022 ( .A(sreg[1511]), .B(n22438), .Z(n22440) );
  NANDN U24023 ( .A(sreg[1510]), .B(n22401), .Z(n22405) );
  NAND U24024 ( .A(n22403), .B(n22402), .Z(n22404) );
  NAND U24025 ( .A(n22405), .B(n22404), .Z(n22439) );
  XNOR U24026 ( .A(n22440), .B(n22439), .Z(c[1511]) );
  NANDN U24027 ( .A(n22407), .B(n22406), .Z(n22411) );
  NANDN U24028 ( .A(n22409), .B(n22408), .Z(n22410) );
  AND U24029 ( .A(n22411), .B(n22410), .Z(n22446) );
  NANDN U24030 ( .A(n22413), .B(n22412), .Z(n22417) );
  NANDN U24031 ( .A(n22415), .B(n22414), .Z(n22416) );
  AND U24032 ( .A(n22417), .B(n22416), .Z(n22444) );
  NAND U24033 ( .A(n42143), .B(n22418), .Z(n22420) );
  XNOR U24034 ( .A(a[490]), .B(n4141), .Z(n22455) );
  NAND U24035 ( .A(n42144), .B(n22455), .Z(n22419) );
  AND U24036 ( .A(n22420), .B(n22419), .Z(n22470) );
  XOR U24037 ( .A(a[494]), .B(n42012), .Z(n22458) );
  XNOR U24038 ( .A(n22470), .B(n22469), .Z(n22472) );
  AND U24039 ( .A(a[496]), .B(b[0]), .Z(n22422) );
  XNOR U24040 ( .A(n22422), .B(n4071), .Z(n22424) );
  NANDN U24041 ( .A(b[0]), .B(a[495]), .Z(n22423) );
  NAND U24042 ( .A(n22424), .B(n22423), .Z(n22466) );
  XOR U24043 ( .A(a[492]), .B(n42085), .Z(n22462) );
  AND U24044 ( .A(a[488]), .B(b[7]), .Z(n22463) );
  XNOR U24045 ( .A(n22464), .B(n22463), .Z(n22465) );
  XNOR U24046 ( .A(n22466), .B(n22465), .Z(n22471) );
  XOR U24047 ( .A(n22472), .B(n22471), .Z(n22450) );
  NANDN U24048 ( .A(n22427), .B(n22426), .Z(n22431) );
  NANDN U24049 ( .A(n22429), .B(n22428), .Z(n22430) );
  AND U24050 ( .A(n22431), .B(n22430), .Z(n22449) );
  XNOR U24051 ( .A(n22450), .B(n22449), .Z(n22451) );
  NANDN U24052 ( .A(n22433), .B(n22432), .Z(n22437) );
  NAND U24053 ( .A(n22435), .B(n22434), .Z(n22436) );
  NAND U24054 ( .A(n22437), .B(n22436), .Z(n22452) );
  XNOR U24055 ( .A(n22451), .B(n22452), .Z(n22443) );
  XNOR U24056 ( .A(n22444), .B(n22443), .Z(n22445) );
  XNOR U24057 ( .A(n22446), .B(n22445), .Z(n22475) );
  XNOR U24058 ( .A(sreg[1512]), .B(n22475), .Z(n22477) );
  NANDN U24059 ( .A(sreg[1511]), .B(n22438), .Z(n22442) );
  NAND U24060 ( .A(n22440), .B(n22439), .Z(n22441) );
  NAND U24061 ( .A(n22442), .B(n22441), .Z(n22476) );
  XNOR U24062 ( .A(n22477), .B(n22476), .Z(c[1512]) );
  NANDN U24063 ( .A(n22444), .B(n22443), .Z(n22448) );
  NANDN U24064 ( .A(n22446), .B(n22445), .Z(n22447) );
  AND U24065 ( .A(n22448), .B(n22447), .Z(n22483) );
  NANDN U24066 ( .A(n22450), .B(n22449), .Z(n22454) );
  NANDN U24067 ( .A(n22452), .B(n22451), .Z(n22453) );
  AND U24068 ( .A(n22454), .B(n22453), .Z(n22481) );
  NAND U24069 ( .A(n42143), .B(n22455), .Z(n22457) );
  XNOR U24070 ( .A(a[491]), .B(n4142), .Z(n22492) );
  NAND U24071 ( .A(n42144), .B(n22492), .Z(n22456) );
  AND U24072 ( .A(n22457), .B(n22456), .Z(n22507) );
  XOR U24073 ( .A(a[495]), .B(n42012), .Z(n22495) );
  XNOR U24074 ( .A(n22507), .B(n22506), .Z(n22509) );
  AND U24075 ( .A(a[497]), .B(b[0]), .Z(n22459) );
  XNOR U24076 ( .A(n22459), .B(n4071), .Z(n22461) );
  NANDN U24077 ( .A(b[0]), .B(a[496]), .Z(n22460) );
  NAND U24078 ( .A(n22461), .B(n22460), .Z(n22503) );
  XOR U24079 ( .A(a[493]), .B(n42085), .Z(n22496) );
  AND U24080 ( .A(a[489]), .B(b[7]), .Z(n22500) );
  XNOR U24081 ( .A(n22501), .B(n22500), .Z(n22502) );
  XNOR U24082 ( .A(n22503), .B(n22502), .Z(n22508) );
  XOR U24083 ( .A(n22509), .B(n22508), .Z(n22487) );
  NANDN U24084 ( .A(n22464), .B(n22463), .Z(n22468) );
  NANDN U24085 ( .A(n22466), .B(n22465), .Z(n22467) );
  AND U24086 ( .A(n22468), .B(n22467), .Z(n22486) );
  XNOR U24087 ( .A(n22487), .B(n22486), .Z(n22488) );
  NANDN U24088 ( .A(n22470), .B(n22469), .Z(n22474) );
  NAND U24089 ( .A(n22472), .B(n22471), .Z(n22473) );
  NAND U24090 ( .A(n22474), .B(n22473), .Z(n22489) );
  XNOR U24091 ( .A(n22488), .B(n22489), .Z(n22480) );
  XNOR U24092 ( .A(n22481), .B(n22480), .Z(n22482) );
  XNOR U24093 ( .A(n22483), .B(n22482), .Z(n22512) );
  XNOR U24094 ( .A(sreg[1513]), .B(n22512), .Z(n22514) );
  NANDN U24095 ( .A(sreg[1512]), .B(n22475), .Z(n22479) );
  NAND U24096 ( .A(n22477), .B(n22476), .Z(n22478) );
  NAND U24097 ( .A(n22479), .B(n22478), .Z(n22513) );
  XNOR U24098 ( .A(n22514), .B(n22513), .Z(c[1513]) );
  NANDN U24099 ( .A(n22481), .B(n22480), .Z(n22485) );
  NANDN U24100 ( .A(n22483), .B(n22482), .Z(n22484) );
  AND U24101 ( .A(n22485), .B(n22484), .Z(n22520) );
  NANDN U24102 ( .A(n22487), .B(n22486), .Z(n22491) );
  NANDN U24103 ( .A(n22489), .B(n22488), .Z(n22490) );
  AND U24104 ( .A(n22491), .B(n22490), .Z(n22518) );
  NAND U24105 ( .A(n42143), .B(n22492), .Z(n22494) );
  XNOR U24106 ( .A(a[492]), .B(n4142), .Z(n22529) );
  NAND U24107 ( .A(n42144), .B(n22529), .Z(n22493) );
  AND U24108 ( .A(n22494), .B(n22493), .Z(n22544) );
  XOR U24109 ( .A(a[496]), .B(n42012), .Z(n22532) );
  XNOR U24110 ( .A(n22544), .B(n22543), .Z(n22546) );
  XOR U24111 ( .A(a[494]), .B(n42085), .Z(n22536) );
  AND U24112 ( .A(a[490]), .B(b[7]), .Z(n22537) );
  XNOR U24113 ( .A(n22538), .B(n22537), .Z(n22539) );
  AND U24114 ( .A(a[498]), .B(b[0]), .Z(n22497) );
  XNOR U24115 ( .A(n22497), .B(n4071), .Z(n22499) );
  NANDN U24116 ( .A(b[0]), .B(a[497]), .Z(n22498) );
  NAND U24117 ( .A(n22499), .B(n22498), .Z(n22540) );
  XNOR U24118 ( .A(n22539), .B(n22540), .Z(n22545) );
  XOR U24119 ( .A(n22546), .B(n22545), .Z(n22524) );
  NANDN U24120 ( .A(n22501), .B(n22500), .Z(n22505) );
  NANDN U24121 ( .A(n22503), .B(n22502), .Z(n22504) );
  AND U24122 ( .A(n22505), .B(n22504), .Z(n22523) );
  XNOR U24123 ( .A(n22524), .B(n22523), .Z(n22525) );
  NANDN U24124 ( .A(n22507), .B(n22506), .Z(n22511) );
  NAND U24125 ( .A(n22509), .B(n22508), .Z(n22510) );
  NAND U24126 ( .A(n22511), .B(n22510), .Z(n22526) );
  XNOR U24127 ( .A(n22525), .B(n22526), .Z(n22517) );
  XNOR U24128 ( .A(n22518), .B(n22517), .Z(n22519) );
  XNOR U24129 ( .A(n22520), .B(n22519), .Z(n22549) );
  XNOR U24130 ( .A(sreg[1514]), .B(n22549), .Z(n22551) );
  NANDN U24131 ( .A(sreg[1513]), .B(n22512), .Z(n22516) );
  NAND U24132 ( .A(n22514), .B(n22513), .Z(n22515) );
  NAND U24133 ( .A(n22516), .B(n22515), .Z(n22550) );
  XNOR U24134 ( .A(n22551), .B(n22550), .Z(c[1514]) );
  NANDN U24135 ( .A(n22518), .B(n22517), .Z(n22522) );
  NANDN U24136 ( .A(n22520), .B(n22519), .Z(n22521) );
  AND U24137 ( .A(n22522), .B(n22521), .Z(n22557) );
  NANDN U24138 ( .A(n22524), .B(n22523), .Z(n22528) );
  NANDN U24139 ( .A(n22526), .B(n22525), .Z(n22527) );
  AND U24140 ( .A(n22528), .B(n22527), .Z(n22555) );
  NAND U24141 ( .A(n42143), .B(n22529), .Z(n22531) );
  XNOR U24142 ( .A(a[493]), .B(n4142), .Z(n22566) );
  NAND U24143 ( .A(n42144), .B(n22566), .Z(n22530) );
  AND U24144 ( .A(n22531), .B(n22530), .Z(n22581) );
  XOR U24145 ( .A(a[497]), .B(n42012), .Z(n22569) );
  XNOR U24146 ( .A(n22581), .B(n22580), .Z(n22583) );
  AND U24147 ( .A(b[0]), .B(a[499]), .Z(n22533) );
  XOR U24148 ( .A(b[1]), .B(n22533), .Z(n22535) );
  NANDN U24149 ( .A(b[0]), .B(a[498]), .Z(n22534) );
  AND U24150 ( .A(n22535), .B(n22534), .Z(n22576) );
  XOR U24151 ( .A(a[495]), .B(n42085), .Z(n22573) );
  AND U24152 ( .A(a[491]), .B(b[7]), .Z(n22574) );
  XOR U24153 ( .A(n22575), .B(n22574), .Z(n22577) );
  XNOR U24154 ( .A(n22576), .B(n22577), .Z(n22582) );
  XOR U24155 ( .A(n22583), .B(n22582), .Z(n22561) );
  NANDN U24156 ( .A(n22538), .B(n22537), .Z(n22542) );
  NANDN U24157 ( .A(n22540), .B(n22539), .Z(n22541) );
  AND U24158 ( .A(n22542), .B(n22541), .Z(n22560) );
  XNOR U24159 ( .A(n22561), .B(n22560), .Z(n22562) );
  NANDN U24160 ( .A(n22544), .B(n22543), .Z(n22548) );
  NAND U24161 ( .A(n22546), .B(n22545), .Z(n22547) );
  NAND U24162 ( .A(n22548), .B(n22547), .Z(n22563) );
  XNOR U24163 ( .A(n22562), .B(n22563), .Z(n22554) );
  XNOR U24164 ( .A(n22555), .B(n22554), .Z(n22556) );
  XNOR U24165 ( .A(n22557), .B(n22556), .Z(n22586) );
  XNOR U24166 ( .A(sreg[1515]), .B(n22586), .Z(n22588) );
  NANDN U24167 ( .A(sreg[1514]), .B(n22549), .Z(n22553) );
  NAND U24168 ( .A(n22551), .B(n22550), .Z(n22552) );
  NAND U24169 ( .A(n22553), .B(n22552), .Z(n22587) );
  XNOR U24170 ( .A(n22588), .B(n22587), .Z(c[1515]) );
  NANDN U24171 ( .A(n22555), .B(n22554), .Z(n22559) );
  NANDN U24172 ( .A(n22557), .B(n22556), .Z(n22558) );
  AND U24173 ( .A(n22559), .B(n22558), .Z(n22594) );
  NANDN U24174 ( .A(n22561), .B(n22560), .Z(n22565) );
  NANDN U24175 ( .A(n22563), .B(n22562), .Z(n22564) );
  AND U24176 ( .A(n22565), .B(n22564), .Z(n22592) );
  NAND U24177 ( .A(n42143), .B(n22566), .Z(n22568) );
  XNOR U24178 ( .A(a[494]), .B(n4142), .Z(n22603) );
  NAND U24179 ( .A(n42144), .B(n22603), .Z(n22567) );
  AND U24180 ( .A(n22568), .B(n22567), .Z(n22618) );
  XOR U24181 ( .A(a[498]), .B(n42012), .Z(n22606) );
  XNOR U24182 ( .A(n22618), .B(n22617), .Z(n22620) );
  AND U24183 ( .A(a[500]), .B(b[0]), .Z(n22570) );
  XNOR U24184 ( .A(n22570), .B(n4071), .Z(n22572) );
  NANDN U24185 ( .A(b[0]), .B(a[499]), .Z(n22571) );
  NAND U24186 ( .A(n22572), .B(n22571), .Z(n22614) );
  XOR U24187 ( .A(a[496]), .B(n42085), .Z(n22610) );
  AND U24188 ( .A(a[492]), .B(b[7]), .Z(n22611) );
  XNOR U24189 ( .A(n22612), .B(n22611), .Z(n22613) );
  XNOR U24190 ( .A(n22614), .B(n22613), .Z(n22619) );
  XOR U24191 ( .A(n22620), .B(n22619), .Z(n22598) );
  NANDN U24192 ( .A(n22575), .B(n22574), .Z(n22579) );
  NANDN U24193 ( .A(n22577), .B(n22576), .Z(n22578) );
  AND U24194 ( .A(n22579), .B(n22578), .Z(n22597) );
  XNOR U24195 ( .A(n22598), .B(n22597), .Z(n22599) );
  NANDN U24196 ( .A(n22581), .B(n22580), .Z(n22585) );
  NAND U24197 ( .A(n22583), .B(n22582), .Z(n22584) );
  NAND U24198 ( .A(n22585), .B(n22584), .Z(n22600) );
  XNOR U24199 ( .A(n22599), .B(n22600), .Z(n22591) );
  XNOR U24200 ( .A(n22592), .B(n22591), .Z(n22593) );
  XNOR U24201 ( .A(n22594), .B(n22593), .Z(n22623) );
  XNOR U24202 ( .A(sreg[1516]), .B(n22623), .Z(n22625) );
  NANDN U24203 ( .A(sreg[1515]), .B(n22586), .Z(n22590) );
  NAND U24204 ( .A(n22588), .B(n22587), .Z(n22589) );
  NAND U24205 ( .A(n22590), .B(n22589), .Z(n22624) );
  XNOR U24206 ( .A(n22625), .B(n22624), .Z(c[1516]) );
  NANDN U24207 ( .A(n22592), .B(n22591), .Z(n22596) );
  NANDN U24208 ( .A(n22594), .B(n22593), .Z(n22595) );
  AND U24209 ( .A(n22596), .B(n22595), .Z(n22631) );
  NANDN U24210 ( .A(n22598), .B(n22597), .Z(n22602) );
  NANDN U24211 ( .A(n22600), .B(n22599), .Z(n22601) );
  AND U24212 ( .A(n22602), .B(n22601), .Z(n22629) );
  NAND U24213 ( .A(n42143), .B(n22603), .Z(n22605) );
  XNOR U24214 ( .A(a[495]), .B(n4142), .Z(n22640) );
  NAND U24215 ( .A(n42144), .B(n22640), .Z(n22604) );
  AND U24216 ( .A(n22605), .B(n22604), .Z(n22655) );
  XOR U24217 ( .A(a[499]), .B(n42012), .Z(n22643) );
  XNOR U24218 ( .A(n22655), .B(n22654), .Z(n22657) );
  AND U24219 ( .A(a[501]), .B(b[0]), .Z(n22607) );
  XNOR U24220 ( .A(n22607), .B(n4071), .Z(n22609) );
  NANDN U24221 ( .A(b[0]), .B(a[500]), .Z(n22608) );
  NAND U24222 ( .A(n22609), .B(n22608), .Z(n22651) );
  XOR U24223 ( .A(a[497]), .B(n42085), .Z(n22647) );
  AND U24224 ( .A(a[493]), .B(b[7]), .Z(n22648) );
  XNOR U24225 ( .A(n22649), .B(n22648), .Z(n22650) );
  XNOR U24226 ( .A(n22651), .B(n22650), .Z(n22656) );
  XOR U24227 ( .A(n22657), .B(n22656), .Z(n22635) );
  NANDN U24228 ( .A(n22612), .B(n22611), .Z(n22616) );
  NANDN U24229 ( .A(n22614), .B(n22613), .Z(n22615) );
  AND U24230 ( .A(n22616), .B(n22615), .Z(n22634) );
  XNOR U24231 ( .A(n22635), .B(n22634), .Z(n22636) );
  NANDN U24232 ( .A(n22618), .B(n22617), .Z(n22622) );
  NAND U24233 ( .A(n22620), .B(n22619), .Z(n22621) );
  NAND U24234 ( .A(n22622), .B(n22621), .Z(n22637) );
  XNOR U24235 ( .A(n22636), .B(n22637), .Z(n22628) );
  XNOR U24236 ( .A(n22629), .B(n22628), .Z(n22630) );
  XNOR U24237 ( .A(n22631), .B(n22630), .Z(n22660) );
  XNOR U24238 ( .A(sreg[1517]), .B(n22660), .Z(n22662) );
  NANDN U24239 ( .A(sreg[1516]), .B(n22623), .Z(n22627) );
  NAND U24240 ( .A(n22625), .B(n22624), .Z(n22626) );
  NAND U24241 ( .A(n22627), .B(n22626), .Z(n22661) );
  XNOR U24242 ( .A(n22662), .B(n22661), .Z(c[1517]) );
  NANDN U24243 ( .A(n22629), .B(n22628), .Z(n22633) );
  NANDN U24244 ( .A(n22631), .B(n22630), .Z(n22632) );
  AND U24245 ( .A(n22633), .B(n22632), .Z(n22668) );
  NANDN U24246 ( .A(n22635), .B(n22634), .Z(n22639) );
  NANDN U24247 ( .A(n22637), .B(n22636), .Z(n22638) );
  AND U24248 ( .A(n22639), .B(n22638), .Z(n22666) );
  NAND U24249 ( .A(n42143), .B(n22640), .Z(n22642) );
  XNOR U24250 ( .A(a[496]), .B(n4142), .Z(n22677) );
  NAND U24251 ( .A(n42144), .B(n22677), .Z(n22641) );
  AND U24252 ( .A(n22642), .B(n22641), .Z(n22692) );
  XOR U24253 ( .A(a[500]), .B(n42012), .Z(n22680) );
  XNOR U24254 ( .A(n22692), .B(n22691), .Z(n22694) );
  AND U24255 ( .A(a[502]), .B(b[0]), .Z(n22644) );
  XNOR U24256 ( .A(n22644), .B(n4071), .Z(n22646) );
  NANDN U24257 ( .A(b[0]), .B(a[501]), .Z(n22645) );
  NAND U24258 ( .A(n22646), .B(n22645), .Z(n22688) );
  XOR U24259 ( .A(a[498]), .B(n42085), .Z(n22684) );
  AND U24260 ( .A(a[494]), .B(b[7]), .Z(n22685) );
  XNOR U24261 ( .A(n22686), .B(n22685), .Z(n22687) );
  XNOR U24262 ( .A(n22688), .B(n22687), .Z(n22693) );
  XOR U24263 ( .A(n22694), .B(n22693), .Z(n22672) );
  NANDN U24264 ( .A(n22649), .B(n22648), .Z(n22653) );
  NANDN U24265 ( .A(n22651), .B(n22650), .Z(n22652) );
  AND U24266 ( .A(n22653), .B(n22652), .Z(n22671) );
  XNOR U24267 ( .A(n22672), .B(n22671), .Z(n22673) );
  NANDN U24268 ( .A(n22655), .B(n22654), .Z(n22659) );
  NAND U24269 ( .A(n22657), .B(n22656), .Z(n22658) );
  NAND U24270 ( .A(n22659), .B(n22658), .Z(n22674) );
  XNOR U24271 ( .A(n22673), .B(n22674), .Z(n22665) );
  XNOR U24272 ( .A(n22666), .B(n22665), .Z(n22667) );
  XNOR U24273 ( .A(n22668), .B(n22667), .Z(n22697) );
  XNOR U24274 ( .A(sreg[1518]), .B(n22697), .Z(n22699) );
  NANDN U24275 ( .A(sreg[1517]), .B(n22660), .Z(n22664) );
  NAND U24276 ( .A(n22662), .B(n22661), .Z(n22663) );
  NAND U24277 ( .A(n22664), .B(n22663), .Z(n22698) );
  XNOR U24278 ( .A(n22699), .B(n22698), .Z(c[1518]) );
  NANDN U24279 ( .A(n22666), .B(n22665), .Z(n22670) );
  NANDN U24280 ( .A(n22668), .B(n22667), .Z(n22669) );
  AND U24281 ( .A(n22670), .B(n22669), .Z(n22705) );
  NANDN U24282 ( .A(n22672), .B(n22671), .Z(n22676) );
  NANDN U24283 ( .A(n22674), .B(n22673), .Z(n22675) );
  AND U24284 ( .A(n22676), .B(n22675), .Z(n22703) );
  NAND U24285 ( .A(n42143), .B(n22677), .Z(n22679) );
  XNOR U24286 ( .A(a[497]), .B(n4142), .Z(n22714) );
  NAND U24287 ( .A(n42144), .B(n22714), .Z(n22678) );
  AND U24288 ( .A(n22679), .B(n22678), .Z(n22729) );
  XOR U24289 ( .A(a[501]), .B(n42012), .Z(n22717) );
  XNOR U24290 ( .A(n22729), .B(n22728), .Z(n22731) );
  AND U24291 ( .A(a[503]), .B(b[0]), .Z(n22681) );
  XNOR U24292 ( .A(n22681), .B(n4071), .Z(n22683) );
  NANDN U24293 ( .A(b[0]), .B(a[502]), .Z(n22682) );
  NAND U24294 ( .A(n22683), .B(n22682), .Z(n22725) );
  XOR U24295 ( .A(a[499]), .B(n42085), .Z(n22718) );
  AND U24296 ( .A(a[495]), .B(b[7]), .Z(n22722) );
  XNOR U24297 ( .A(n22723), .B(n22722), .Z(n22724) );
  XNOR U24298 ( .A(n22725), .B(n22724), .Z(n22730) );
  XOR U24299 ( .A(n22731), .B(n22730), .Z(n22709) );
  NANDN U24300 ( .A(n22686), .B(n22685), .Z(n22690) );
  NANDN U24301 ( .A(n22688), .B(n22687), .Z(n22689) );
  AND U24302 ( .A(n22690), .B(n22689), .Z(n22708) );
  XNOR U24303 ( .A(n22709), .B(n22708), .Z(n22710) );
  NANDN U24304 ( .A(n22692), .B(n22691), .Z(n22696) );
  NAND U24305 ( .A(n22694), .B(n22693), .Z(n22695) );
  NAND U24306 ( .A(n22696), .B(n22695), .Z(n22711) );
  XNOR U24307 ( .A(n22710), .B(n22711), .Z(n22702) );
  XNOR U24308 ( .A(n22703), .B(n22702), .Z(n22704) );
  XNOR U24309 ( .A(n22705), .B(n22704), .Z(n22734) );
  XNOR U24310 ( .A(sreg[1519]), .B(n22734), .Z(n22736) );
  NANDN U24311 ( .A(sreg[1518]), .B(n22697), .Z(n22701) );
  NAND U24312 ( .A(n22699), .B(n22698), .Z(n22700) );
  NAND U24313 ( .A(n22701), .B(n22700), .Z(n22735) );
  XNOR U24314 ( .A(n22736), .B(n22735), .Z(c[1519]) );
  NANDN U24315 ( .A(n22703), .B(n22702), .Z(n22707) );
  NANDN U24316 ( .A(n22705), .B(n22704), .Z(n22706) );
  AND U24317 ( .A(n22707), .B(n22706), .Z(n22746) );
  NANDN U24318 ( .A(n22709), .B(n22708), .Z(n22713) );
  NANDN U24319 ( .A(n22711), .B(n22710), .Z(n22712) );
  AND U24320 ( .A(n22713), .B(n22712), .Z(n22745) );
  NAND U24321 ( .A(n42143), .B(n22714), .Z(n22716) );
  XNOR U24322 ( .A(a[498]), .B(n4143), .Z(n22756) );
  NAND U24323 ( .A(n42144), .B(n22756), .Z(n22715) );
  AND U24324 ( .A(n22716), .B(n22715), .Z(n22771) );
  XOR U24325 ( .A(a[502]), .B(n42012), .Z(n22759) );
  XNOR U24326 ( .A(n22771), .B(n22770), .Z(n22773) );
  XOR U24327 ( .A(a[500]), .B(n42085), .Z(n22763) );
  AND U24328 ( .A(a[496]), .B(b[7]), .Z(n22764) );
  XNOR U24329 ( .A(n22765), .B(n22764), .Z(n22766) );
  AND U24330 ( .A(a[504]), .B(b[0]), .Z(n22719) );
  XNOR U24331 ( .A(n22719), .B(n4071), .Z(n22721) );
  NANDN U24332 ( .A(b[0]), .B(a[503]), .Z(n22720) );
  NAND U24333 ( .A(n22721), .B(n22720), .Z(n22767) );
  XNOR U24334 ( .A(n22766), .B(n22767), .Z(n22772) );
  XOR U24335 ( .A(n22773), .B(n22772), .Z(n22751) );
  NANDN U24336 ( .A(n22723), .B(n22722), .Z(n22727) );
  NANDN U24337 ( .A(n22725), .B(n22724), .Z(n22726) );
  AND U24338 ( .A(n22727), .B(n22726), .Z(n22750) );
  XNOR U24339 ( .A(n22751), .B(n22750), .Z(n22752) );
  NANDN U24340 ( .A(n22729), .B(n22728), .Z(n22733) );
  NAND U24341 ( .A(n22731), .B(n22730), .Z(n22732) );
  NAND U24342 ( .A(n22733), .B(n22732), .Z(n22753) );
  XNOR U24343 ( .A(n22752), .B(n22753), .Z(n22744) );
  XOR U24344 ( .A(n22745), .B(n22744), .Z(n22747) );
  XOR U24345 ( .A(n22746), .B(n22747), .Z(n22739) );
  XNOR U24346 ( .A(n22739), .B(sreg[1520]), .Z(n22741) );
  NANDN U24347 ( .A(sreg[1519]), .B(n22734), .Z(n22738) );
  NAND U24348 ( .A(n22736), .B(n22735), .Z(n22737) );
  AND U24349 ( .A(n22738), .B(n22737), .Z(n22740) );
  XOR U24350 ( .A(n22741), .B(n22740), .Z(c[1520]) );
  NANDN U24351 ( .A(n22739), .B(sreg[1520]), .Z(n22743) );
  NAND U24352 ( .A(n22741), .B(n22740), .Z(n22742) );
  AND U24353 ( .A(n22743), .B(n22742), .Z(n22810) );
  NANDN U24354 ( .A(n22745), .B(n22744), .Z(n22749) );
  OR U24355 ( .A(n22747), .B(n22746), .Z(n22748) );
  AND U24356 ( .A(n22749), .B(n22748), .Z(n22779) );
  NANDN U24357 ( .A(n22751), .B(n22750), .Z(n22755) );
  NANDN U24358 ( .A(n22753), .B(n22752), .Z(n22754) );
  AND U24359 ( .A(n22755), .B(n22754), .Z(n22777) );
  NAND U24360 ( .A(n42143), .B(n22756), .Z(n22758) );
  XNOR U24361 ( .A(a[499]), .B(n4143), .Z(n22788) );
  NAND U24362 ( .A(n42144), .B(n22788), .Z(n22757) );
  AND U24363 ( .A(n22758), .B(n22757), .Z(n22803) );
  XOR U24364 ( .A(a[503]), .B(n42012), .Z(n22791) );
  XNOR U24365 ( .A(n22803), .B(n22802), .Z(n22805) );
  AND U24366 ( .A(a[505]), .B(b[0]), .Z(n22760) );
  XNOR U24367 ( .A(n22760), .B(n4071), .Z(n22762) );
  NANDN U24368 ( .A(b[0]), .B(a[504]), .Z(n22761) );
  NAND U24369 ( .A(n22762), .B(n22761), .Z(n22799) );
  XOR U24370 ( .A(a[501]), .B(n42085), .Z(n22792) );
  AND U24371 ( .A(a[497]), .B(b[7]), .Z(n22796) );
  XNOR U24372 ( .A(n22797), .B(n22796), .Z(n22798) );
  XNOR U24373 ( .A(n22799), .B(n22798), .Z(n22804) );
  XOR U24374 ( .A(n22805), .B(n22804), .Z(n22783) );
  NANDN U24375 ( .A(n22765), .B(n22764), .Z(n22769) );
  NANDN U24376 ( .A(n22767), .B(n22766), .Z(n22768) );
  AND U24377 ( .A(n22769), .B(n22768), .Z(n22782) );
  XNOR U24378 ( .A(n22783), .B(n22782), .Z(n22784) );
  NANDN U24379 ( .A(n22771), .B(n22770), .Z(n22775) );
  NAND U24380 ( .A(n22773), .B(n22772), .Z(n22774) );
  NAND U24381 ( .A(n22775), .B(n22774), .Z(n22785) );
  XNOR U24382 ( .A(n22784), .B(n22785), .Z(n22776) );
  XNOR U24383 ( .A(n22777), .B(n22776), .Z(n22778) );
  XNOR U24384 ( .A(n22779), .B(n22778), .Z(n22808) );
  XNOR U24385 ( .A(sreg[1521]), .B(n22808), .Z(n22809) );
  XNOR U24386 ( .A(n22810), .B(n22809), .Z(c[1521]) );
  NANDN U24387 ( .A(n22777), .B(n22776), .Z(n22781) );
  NANDN U24388 ( .A(n22779), .B(n22778), .Z(n22780) );
  AND U24389 ( .A(n22781), .B(n22780), .Z(n22816) );
  NANDN U24390 ( .A(n22783), .B(n22782), .Z(n22787) );
  NANDN U24391 ( .A(n22785), .B(n22784), .Z(n22786) );
  AND U24392 ( .A(n22787), .B(n22786), .Z(n22814) );
  NAND U24393 ( .A(n42143), .B(n22788), .Z(n22790) );
  XNOR U24394 ( .A(a[500]), .B(n4143), .Z(n22825) );
  NAND U24395 ( .A(n42144), .B(n22825), .Z(n22789) );
  AND U24396 ( .A(n22790), .B(n22789), .Z(n22840) );
  XOR U24397 ( .A(a[504]), .B(n42012), .Z(n22828) );
  XNOR U24398 ( .A(n22840), .B(n22839), .Z(n22842) );
  XOR U24399 ( .A(a[502]), .B(n42085), .Z(n22829) );
  AND U24400 ( .A(a[498]), .B(b[7]), .Z(n22833) );
  XNOR U24401 ( .A(n22834), .B(n22833), .Z(n22835) );
  AND U24402 ( .A(a[506]), .B(b[0]), .Z(n22793) );
  XNOR U24403 ( .A(n22793), .B(n4071), .Z(n22795) );
  NANDN U24404 ( .A(b[0]), .B(a[505]), .Z(n22794) );
  NAND U24405 ( .A(n22795), .B(n22794), .Z(n22836) );
  XNOR U24406 ( .A(n22835), .B(n22836), .Z(n22841) );
  XOR U24407 ( .A(n22842), .B(n22841), .Z(n22820) );
  NANDN U24408 ( .A(n22797), .B(n22796), .Z(n22801) );
  NANDN U24409 ( .A(n22799), .B(n22798), .Z(n22800) );
  AND U24410 ( .A(n22801), .B(n22800), .Z(n22819) );
  XNOR U24411 ( .A(n22820), .B(n22819), .Z(n22821) );
  NANDN U24412 ( .A(n22803), .B(n22802), .Z(n22807) );
  NAND U24413 ( .A(n22805), .B(n22804), .Z(n22806) );
  NAND U24414 ( .A(n22807), .B(n22806), .Z(n22822) );
  XNOR U24415 ( .A(n22821), .B(n22822), .Z(n22813) );
  XNOR U24416 ( .A(n22814), .B(n22813), .Z(n22815) );
  XNOR U24417 ( .A(n22816), .B(n22815), .Z(n22845) );
  XNOR U24418 ( .A(sreg[1522]), .B(n22845), .Z(n22847) );
  NANDN U24419 ( .A(sreg[1521]), .B(n22808), .Z(n22812) );
  NAND U24420 ( .A(n22810), .B(n22809), .Z(n22811) );
  NAND U24421 ( .A(n22812), .B(n22811), .Z(n22846) );
  XNOR U24422 ( .A(n22847), .B(n22846), .Z(c[1522]) );
  NANDN U24423 ( .A(n22814), .B(n22813), .Z(n22818) );
  NANDN U24424 ( .A(n22816), .B(n22815), .Z(n22817) );
  AND U24425 ( .A(n22818), .B(n22817), .Z(n22853) );
  NANDN U24426 ( .A(n22820), .B(n22819), .Z(n22824) );
  NANDN U24427 ( .A(n22822), .B(n22821), .Z(n22823) );
  AND U24428 ( .A(n22824), .B(n22823), .Z(n22851) );
  NAND U24429 ( .A(n42143), .B(n22825), .Z(n22827) );
  XNOR U24430 ( .A(a[501]), .B(n4143), .Z(n22862) );
  NAND U24431 ( .A(n42144), .B(n22862), .Z(n22826) );
  AND U24432 ( .A(n22827), .B(n22826), .Z(n22877) );
  XOR U24433 ( .A(a[505]), .B(n42012), .Z(n22865) );
  XNOR U24434 ( .A(n22877), .B(n22876), .Z(n22879) );
  XOR U24435 ( .A(a[503]), .B(n42085), .Z(n22869) );
  AND U24436 ( .A(a[499]), .B(b[7]), .Z(n22870) );
  XNOR U24437 ( .A(n22871), .B(n22870), .Z(n22872) );
  AND U24438 ( .A(a[507]), .B(b[0]), .Z(n22830) );
  XNOR U24439 ( .A(n22830), .B(n4071), .Z(n22832) );
  NANDN U24440 ( .A(b[0]), .B(a[506]), .Z(n22831) );
  NAND U24441 ( .A(n22832), .B(n22831), .Z(n22873) );
  XNOR U24442 ( .A(n22872), .B(n22873), .Z(n22878) );
  XOR U24443 ( .A(n22879), .B(n22878), .Z(n22857) );
  NANDN U24444 ( .A(n22834), .B(n22833), .Z(n22838) );
  NANDN U24445 ( .A(n22836), .B(n22835), .Z(n22837) );
  AND U24446 ( .A(n22838), .B(n22837), .Z(n22856) );
  XNOR U24447 ( .A(n22857), .B(n22856), .Z(n22858) );
  NANDN U24448 ( .A(n22840), .B(n22839), .Z(n22844) );
  NAND U24449 ( .A(n22842), .B(n22841), .Z(n22843) );
  NAND U24450 ( .A(n22844), .B(n22843), .Z(n22859) );
  XNOR U24451 ( .A(n22858), .B(n22859), .Z(n22850) );
  XNOR U24452 ( .A(n22851), .B(n22850), .Z(n22852) );
  XNOR U24453 ( .A(n22853), .B(n22852), .Z(n22882) );
  XNOR U24454 ( .A(sreg[1523]), .B(n22882), .Z(n22884) );
  NANDN U24455 ( .A(sreg[1522]), .B(n22845), .Z(n22849) );
  NAND U24456 ( .A(n22847), .B(n22846), .Z(n22848) );
  NAND U24457 ( .A(n22849), .B(n22848), .Z(n22883) );
  XNOR U24458 ( .A(n22884), .B(n22883), .Z(c[1523]) );
  NANDN U24459 ( .A(n22851), .B(n22850), .Z(n22855) );
  NANDN U24460 ( .A(n22853), .B(n22852), .Z(n22854) );
  AND U24461 ( .A(n22855), .B(n22854), .Z(n22890) );
  NANDN U24462 ( .A(n22857), .B(n22856), .Z(n22861) );
  NANDN U24463 ( .A(n22859), .B(n22858), .Z(n22860) );
  AND U24464 ( .A(n22861), .B(n22860), .Z(n22888) );
  NAND U24465 ( .A(n42143), .B(n22862), .Z(n22864) );
  XNOR U24466 ( .A(a[502]), .B(n4143), .Z(n22899) );
  NAND U24467 ( .A(n42144), .B(n22899), .Z(n22863) );
  AND U24468 ( .A(n22864), .B(n22863), .Z(n22914) );
  XOR U24469 ( .A(a[506]), .B(n42012), .Z(n22902) );
  XNOR U24470 ( .A(n22914), .B(n22913), .Z(n22916) );
  AND U24471 ( .A(a[508]), .B(b[0]), .Z(n22866) );
  XNOR U24472 ( .A(n22866), .B(n4071), .Z(n22868) );
  NANDN U24473 ( .A(b[0]), .B(a[507]), .Z(n22867) );
  NAND U24474 ( .A(n22868), .B(n22867), .Z(n22910) );
  XOR U24475 ( .A(a[504]), .B(n42085), .Z(n22903) );
  AND U24476 ( .A(a[500]), .B(b[7]), .Z(n22907) );
  XNOR U24477 ( .A(n22908), .B(n22907), .Z(n22909) );
  XNOR U24478 ( .A(n22910), .B(n22909), .Z(n22915) );
  XOR U24479 ( .A(n22916), .B(n22915), .Z(n22894) );
  NANDN U24480 ( .A(n22871), .B(n22870), .Z(n22875) );
  NANDN U24481 ( .A(n22873), .B(n22872), .Z(n22874) );
  AND U24482 ( .A(n22875), .B(n22874), .Z(n22893) );
  XNOR U24483 ( .A(n22894), .B(n22893), .Z(n22895) );
  NANDN U24484 ( .A(n22877), .B(n22876), .Z(n22881) );
  NAND U24485 ( .A(n22879), .B(n22878), .Z(n22880) );
  NAND U24486 ( .A(n22881), .B(n22880), .Z(n22896) );
  XNOR U24487 ( .A(n22895), .B(n22896), .Z(n22887) );
  XNOR U24488 ( .A(n22888), .B(n22887), .Z(n22889) );
  XNOR U24489 ( .A(n22890), .B(n22889), .Z(n22919) );
  XNOR U24490 ( .A(sreg[1524]), .B(n22919), .Z(n22921) );
  NANDN U24491 ( .A(sreg[1523]), .B(n22882), .Z(n22886) );
  NAND U24492 ( .A(n22884), .B(n22883), .Z(n22885) );
  NAND U24493 ( .A(n22886), .B(n22885), .Z(n22920) );
  XNOR U24494 ( .A(n22921), .B(n22920), .Z(c[1524]) );
  NANDN U24495 ( .A(n22888), .B(n22887), .Z(n22892) );
  NANDN U24496 ( .A(n22890), .B(n22889), .Z(n22891) );
  AND U24497 ( .A(n22892), .B(n22891), .Z(n22927) );
  NANDN U24498 ( .A(n22894), .B(n22893), .Z(n22898) );
  NANDN U24499 ( .A(n22896), .B(n22895), .Z(n22897) );
  AND U24500 ( .A(n22898), .B(n22897), .Z(n22925) );
  NAND U24501 ( .A(n42143), .B(n22899), .Z(n22901) );
  XNOR U24502 ( .A(a[503]), .B(n4143), .Z(n22936) );
  NAND U24503 ( .A(n42144), .B(n22936), .Z(n22900) );
  AND U24504 ( .A(n22901), .B(n22900), .Z(n22951) );
  XOR U24505 ( .A(a[507]), .B(n42012), .Z(n22939) );
  XNOR U24506 ( .A(n22951), .B(n22950), .Z(n22953) );
  XOR U24507 ( .A(a[505]), .B(n42085), .Z(n22943) );
  AND U24508 ( .A(a[501]), .B(b[7]), .Z(n22944) );
  XNOR U24509 ( .A(n22945), .B(n22944), .Z(n22946) );
  AND U24510 ( .A(a[509]), .B(b[0]), .Z(n22904) );
  XNOR U24511 ( .A(n22904), .B(n4071), .Z(n22906) );
  NANDN U24512 ( .A(b[0]), .B(a[508]), .Z(n22905) );
  NAND U24513 ( .A(n22906), .B(n22905), .Z(n22947) );
  XNOR U24514 ( .A(n22946), .B(n22947), .Z(n22952) );
  XOR U24515 ( .A(n22953), .B(n22952), .Z(n22931) );
  NANDN U24516 ( .A(n22908), .B(n22907), .Z(n22912) );
  NANDN U24517 ( .A(n22910), .B(n22909), .Z(n22911) );
  AND U24518 ( .A(n22912), .B(n22911), .Z(n22930) );
  XNOR U24519 ( .A(n22931), .B(n22930), .Z(n22932) );
  NANDN U24520 ( .A(n22914), .B(n22913), .Z(n22918) );
  NAND U24521 ( .A(n22916), .B(n22915), .Z(n22917) );
  NAND U24522 ( .A(n22918), .B(n22917), .Z(n22933) );
  XNOR U24523 ( .A(n22932), .B(n22933), .Z(n22924) );
  XNOR U24524 ( .A(n22925), .B(n22924), .Z(n22926) );
  XNOR U24525 ( .A(n22927), .B(n22926), .Z(n22956) );
  XNOR U24526 ( .A(sreg[1525]), .B(n22956), .Z(n22958) );
  NANDN U24527 ( .A(sreg[1524]), .B(n22919), .Z(n22923) );
  NAND U24528 ( .A(n22921), .B(n22920), .Z(n22922) );
  NAND U24529 ( .A(n22923), .B(n22922), .Z(n22957) );
  XNOR U24530 ( .A(n22958), .B(n22957), .Z(c[1525]) );
  NANDN U24531 ( .A(n22925), .B(n22924), .Z(n22929) );
  NANDN U24532 ( .A(n22927), .B(n22926), .Z(n22928) );
  AND U24533 ( .A(n22929), .B(n22928), .Z(n22964) );
  NANDN U24534 ( .A(n22931), .B(n22930), .Z(n22935) );
  NANDN U24535 ( .A(n22933), .B(n22932), .Z(n22934) );
  AND U24536 ( .A(n22935), .B(n22934), .Z(n22962) );
  NAND U24537 ( .A(n42143), .B(n22936), .Z(n22938) );
  XNOR U24538 ( .A(a[504]), .B(n4143), .Z(n22973) );
  NAND U24539 ( .A(n42144), .B(n22973), .Z(n22937) );
  AND U24540 ( .A(n22938), .B(n22937), .Z(n22988) );
  XOR U24541 ( .A(a[508]), .B(n42012), .Z(n22976) );
  XNOR U24542 ( .A(n22988), .B(n22987), .Z(n22990) );
  AND U24543 ( .A(a[510]), .B(b[0]), .Z(n22940) );
  XNOR U24544 ( .A(n22940), .B(n4071), .Z(n22942) );
  NANDN U24545 ( .A(b[0]), .B(a[509]), .Z(n22941) );
  NAND U24546 ( .A(n22942), .B(n22941), .Z(n22984) );
  XOR U24547 ( .A(a[506]), .B(n42085), .Z(n22980) );
  AND U24548 ( .A(a[502]), .B(b[7]), .Z(n22981) );
  XNOR U24549 ( .A(n22982), .B(n22981), .Z(n22983) );
  XNOR U24550 ( .A(n22984), .B(n22983), .Z(n22989) );
  XOR U24551 ( .A(n22990), .B(n22989), .Z(n22968) );
  NANDN U24552 ( .A(n22945), .B(n22944), .Z(n22949) );
  NANDN U24553 ( .A(n22947), .B(n22946), .Z(n22948) );
  AND U24554 ( .A(n22949), .B(n22948), .Z(n22967) );
  XNOR U24555 ( .A(n22968), .B(n22967), .Z(n22969) );
  NANDN U24556 ( .A(n22951), .B(n22950), .Z(n22955) );
  NAND U24557 ( .A(n22953), .B(n22952), .Z(n22954) );
  NAND U24558 ( .A(n22955), .B(n22954), .Z(n22970) );
  XNOR U24559 ( .A(n22969), .B(n22970), .Z(n22961) );
  XNOR U24560 ( .A(n22962), .B(n22961), .Z(n22963) );
  XNOR U24561 ( .A(n22964), .B(n22963), .Z(n22993) );
  XNOR U24562 ( .A(sreg[1526]), .B(n22993), .Z(n22995) );
  NANDN U24563 ( .A(sreg[1525]), .B(n22956), .Z(n22960) );
  NAND U24564 ( .A(n22958), .B(n22957), .Z(n22959) );
  NAND U24565 ( .A(n22960), .B(n22959), .Z(n22994) );
  XNOR U24566 ( .A(n22995), .B(n22994), .Z(c[1526]) );
  NANDN U24567 ( .A(n22962), .B(n22961), .Z(n22966) );
  NANDN U24568 ( .A(n22964), .B(n22963), .Z(n22965) );
  AND U24569 ( .A(n22966), .B(n22965), .Z(n23001) );
  NANDN U24570 ( .A(n22968), .B(n22967), .Z(n22972) );
  NANDN U24571 ( .A(n22970), .B(n22969), .Z(n22971) );
  AND U24572 ( .A(n22972), .B(n22971), .Z(n22999) );
  NAND U24573 ( .A(n42143), .B(n22973), .Z(n22975) );
  XNOR U24574 ( .A(a[505]), .B(n4144), .Z(n23010) );
  NAND U24575 ( .A(n42144), .B(n23010), .Z(n22974) );
  AND U24576 ( .A(n22975), .B(n22974), .Z(n23025) );
  XOR U24577 ( .A(a[509]), .B(n42012), .Z(n23013) );
  XNOR U24578 ( .A(n23025), .B(n23024), .Z(n23027) );
  AND U24579 ( .A(a[511]), .B(b[0]), .Z(n22977) );
  XNOR U24580 ( .A(n22977), .B(n4071), .Z(n22979) );
  NANDN U24581 ( .A(b[0]), .B(a[510]), .Z(n22978) );
  NAND U24582 ( .A(n22979), .B(n22978), .Z(n23021) );
  XOR U24583 ( .A(a[507]), .B(n42085), .Z(n23017) );
  AND U24584 ( .A(a[503]), .B(b[7]), .Z(n23018) );
  XNOR U24585 ( .A(n23019), .B(n23018), .Z(n23020) );
  XNOR U24586 ( .A(n23021), .B(n23020), .Z(n23026) );
  XOR U24587 ( .A(n23027), .B(n23026), .Z(n23005) );
  NANDN U24588 ( .A(n22982), .B(n22981), .Z(n22986) );
  NANDN U24589 ( .A(n22984), .B(n22983), .Z(n22985) );
  AND U24590 ( .A(n22986), .B(n22985), .Z(n23004) );
  XNOR U24591 ( .A(n23005), .B(n23004), .Z(n23006) );
  NANDN U24592 ( .A(n22988), .B(n22987), .Z(n22992) );
  NAND U24593 ( .A(n22990), .B(n22989), .Z(n22991) );
  NAND U24594 ( .A(n22992), .B(n22991), .Z(n23007) );
  XNOR U24595 ( .A(n23006), .B(n23007), .Z(n22998) );
  XNOR U24596 ( .A(n22999), .B(n22998), .Z(n23000) );
  XNOR U24597 ( .A(n23001), .B(n23000), .Z(n23030) );
  XNOR U24598 ( .A(sreg[1527]), .B(n23030), .Z(n23032) );
  NANDN U24599 ( .A(sreg[1526]), .B(n22993), .Z(n22997) );
  NAND U24600 ( .A(n22995), .B(n22994), .Z(n22996) );
  NAND U24601 ( .A(n22997), .B(n22996), .Z(n23031) );
  XNOR U24602 ( .A(n23032), .B(n23031), .Z(c[1527]) );
  NANDN U24603 ( .A(n22999), .B(n22998), .Z(n23003) );
  NANDN U24604 ( .A(n23001), .B(n23000), .Z(n23002) );
  AND U24605 ( .A(n23003), .B(n23002), .Z(n23038) );
  NANDN U24606 ( .A(n23005), .B(n23004), .Z(n23009) );
  NANDN U24607 ( .A(n23007), .B(n23006), .Z(n23008) );
  AND U24608 ( .A(n23009), .B(n23008), .Z(n23036) );
  NAND U24609 ( .A(n42143), .B(n23010), .Z(n23012) );
  XNOR U24610 ( .A(a[506]), .B(n4144), .Z(n23047) );
  NAND U24611 ( .A(n42144), .B(n23047), .Z(n23011) );
  AND U24612 ( .A(n23012), .B(n23011), .Z(n23062) );
  XOR U24613 ( .A(a[510]), .B(n42012), .Z(n23050) );
  XNOR U24614 ( .A(n23062), .B(n23061), .Z(n23064) );
  AND U24615 ( .A(a[512]), .B(b[0]), .Z(n23014) );
  XNOR U24616 ( .A(n23014), .B(n4071), .Z(n23016) );
  NANDN U24617 ( .A(b[0]), .B(a[511]), .Z(n23015) );
  NAND U24618 ( .A(n23016), .B(n23015), .Z(n23058) );
  XOR U24619 ( .A(a[508]), .B(n42085), .Z(n23054) );
  AND U24620 ( .A(a[504]), .B(b[7]), .Z(n23055) );
  XNOR U24621 ( .A(n23056), .B(n23055), .Z(n23057) );
  XNOR U24622 ( .A(n23058), .B(n23057), .Z(n23063) );
  XOR U24623 ( .A(n23064), .B(n23063), .Z(n23042) );
  NANDN U24624 ( .A(n23019), .B(n23018), .Z(n23023) );
  NANDN U24625 ( .A(n23021), .B(n23020), .Z(n23022) );
  AND U24626 ( .A(n23023), .B(n23022), .Z(n23041) );
  XNOR U24627 ( .A(n23042), .B(n23041), .Z(n23043) );
  NANDN U24628 ( .A(n23025), .B(n23024), .Z(n23029) );
  NAND U24629 ( .A(n23027), .B(n23026), .Z(n23028) );
  NAND U24630 ( .A(n23029), .B(n23028), .Z(n23044) );
  XNOR U24631 ( .A(n23043), .B(n23044), .Z(n23035) );
  XNOR U24632 ( .A(n23036), .B(n23035), .Z(n23037) );
  XNOR U24633 ( .A(n23038), .B(n23037), .Z(n23067) );
  XNOR U24634 ( .A(sreg[1528]), .B(n23067), .Z(n23069) );
  NANDN U24635 ( .A(sreg[1527]), .B(n23030), .Z(n23034) );
  NAND U24636 ( .A(n23032), .B(n23031), .Z(n23033) );
  NAND U24637 ( .A(n23034), .B(n23033), .Z(n23068) );
  XNOR U24638 ( .A(n23069), .B(n23068), .Z(c[1528]) );
  NANDN U24639 ( .A(n23036), .B(n23035), .Z(n23040) );
  NANDN U24640 ( .A(n23038), .B(n23037), .Z(n23039) );
  AND U24641 ( .A(n23040), .B(n23039), .Z(n23075) );
  NANDN U24642 ( .A(n23042), .B(n23041), .Z(n23046) );
  NANDN U24643 ( .A(n23044), .B(n23043), .Z(n23045) );
  AND U24644 ( .A(n23046), .B(n23045), .Z(n23073) );
  NAND U24645 ( .A(n42143), .B(n23047), .Z(n23049) );
  XNOR U24646 ( .A(a[507]), .B(n4144), .Z(n23084) );
  NAND U24647 ( .A(n42144), .B(n23084), .Z(n23048) );
  AND U24648 ( .A(n23049), .B(n23048), .Z(n23099) );
  XOR U24649 ( .A(a[511]), .B(n42012), .Z(n23087) );
  XNOR U24650 ( .A(n23099), .B(n23098), .Z(n23101) );
  AND U24651 ( .A(a[513]), .B(b[0]), .Z(n23051) );
  XNOR U24652 ( .A(n23051), .B(n4071), .Z(n23053) );
  NANDN U24653 ( .A(b[0]), .B(a[512]), .Z(n23052) );
  NAND U24654 ( .A(n23053), .B(n23052), .Z(n23095) );
  XOR U24655 ( .A(a[509]), .B(n42085), .Z(n23088) );
  AND U24656 ( .A(a[505]), .B(b[7]), .Z(n23092) );
  XNOR U24657 ( .A(n23093), .B(n23092), .Z(n23094) );
  XNOR U24658 ( .A(n23095), .B(n23094), .Z(n23100) );
  XOR U24659 ( .A(n23101), .B(n23100), .Z(n23079) );
  NANDN U24660 ( .A(n23056), .B(n23055), .Z(n23060) );
  NANDN U24661 ( .A(n23058), .B(n23057), .Z(n23059) );
  AND U24662 ( .A(n23060), .B(n23059), .Z(n23078) );
  XNOR U24663 ( .A(n23079), .B(n23078), .Z(n23080) );
  NANDN U24664 ( .A(n23062), .B(n23061), .Z(n23066) );
  NAND U24665 ( .A(n23064), .B(n23063), .Z(n23065) );
  NAND U24666 ( .A(n23066), .B(n23065), .Z(n23081) );
  XNOR U24667 ( .A(n23080), .B(n23081), .Z(n23072) );
  XNOR U24668 ( .A(n23073), .B(n23072), .Z(n23074) );
  XNOR U24669 ( .A(n23075), .B(n23074), .Z(n23104) );
  XNOR U24670 ( .A(sreg[1529]), .B(n23104), .Z(n23106) );
  NANDN U24671 ( .A(sreg[1528]), .B(n23067), .Z(n23071) );
  NAND U24672 ( .A(n23069), .B(n23068), .Z(n23070) );
  NAND U24673 ( .A(n23071), .B(n23070), .Z(n23105) );
  XNOR U24674 ( .A(n23106), .B(n23105), .Z(c[1529]) );
  NANDN U24675 ( .A(n23073), .B(n23072), .Z(n23077) );
  NANDN U24676 ( .A(n23075), .B(n23074), .Z(n23076) );
  AND U24677 ( .A(n23077), .B(n23076), .Z(n23112) );
  NANDN U24678 ( .A(n23079), .B(n23078), .Z(n23083) );
  NANDN U24679 ( .A(n23081), .B(n23080), .Z(n23082) );
  AND U24680 ( .A(n23083), .B(n23082), .Z(n23110) );
  NAND U24681 ( .A(n42143), .B(n23084), .Z(n23086) );
  XNOR U24682 ( .A(a[508]), .B(n4144), .Z(n23121) );
  NAND U24683 ( .A(n42144), .B(n23121), .Z(n23085) );
  AND U24684 ( .A(n23086), .B(n23085), .Z(n23136) );
  XOR U24685 ( .A(a[512]), .B(n42012), .Z(n23124) );
  XNOR U24686 ( .A(n23136), .B(n23135), .Z(n23138) );
  XOR U24687 ( .A(a[510]), .B(n42085), .Z(n23128) );
  AND U24688 ( .A(a[506]), .B(b[7]), .Z(n23129) );
  XNOR U24689 ( .A(n23130), .B(n23129), .Z(n23131) );
  AND U24690 ( .A(a[514]), .B(b[0]), .Z(n23089) );
  XNOR U24691 ( .A(n23089), .B(n4071), .Z(n23091) );
  NANDN U24692 ( .A(b[0]), .B(a[513]), .Z(n23090) );
  NAND U24693 ( .A(n23091), .B(n23090), .Z(n23132) );
  XNOR U24694 ( .A(n23131), .B(n23132), .Z(n23137) );
  XOR U24695 ( .A(n23138), .B(n23137), .Z(n23116) );
  NANDN U24696 ( .A(n23093), .B(n23092), .Z(n23097) );
  NANDN U24697 ( .A(n23095), .B(n23094), .Z(n23096) );
  AND U24698 ( .A(n23097), .B(n23096), .Z(n23115) );
  XNOR U24699 ( .A(n23116), .B(n23115), .Z(n23117) );
  NANDN U24700 ( .A(n23099), .B(n23098), .Z(n23103) );
  NAND U24701 ( .A(n23101), .B(n23100), .Z(n23102) );
  NAND U24702 ( .A(n23103), .B(n23102), .Z(n23118) );
  XNOR U24703 ( .A(n23117), .B(n23118), .Z(n23109) );
  XNOR U24704 ( .A(n23110), .B(n23109), .Z(n23111) );
  XNOR U24705 ( .A(n23112), .B(n23111), .Z(n23141) );
  XNOR U24706 ( .A(sreg[1530]), .B(n23141), .Z(n23143) );
  NANDN U24707 ( .A(sreg[1529]), .B(n23104), .Z(n23108) );
  NAND U24708 ( .A(n23106), .B(n23105), .Z(n23107) );
  NAND U24709 ( .A(n23108), .B(n23107), .Z(n23142) );
  XNOR U24710 ( .A(n23143), .B(n23142), .Z(c[1530]) );
  NANDN U24711 ( .A(n23110), .B(n23109), .Z(n23114) );
  NANDN U24712 ( .A(n23112), .B(n23111), .Z(n23113) );
  AND U24713 ( .A(n23114), .B(n23113), .Z(n23149) );
  NANDN U24714 ( .A(n23116), .B(n23115), .Z(n23120) );
  NANDN U24715 ( .A(n23118), .B(n23117), .Z(n23119) );
  AND U24716 ( .A(n23120), .B(n23119), .Z(n23147) );
  NAND U24717 ( .A(n42143), .B(n23121), .Z(n23123) );
  XNOR U24718 ( .A(a[509]), .B(n4144), .Z(n23158) );
  NAND U24719 ( .A(n42144), .B(n23158), .Z(n23122) );
  AND U24720 ( .A(n23123), .B(n23122), .Z(n23173) );
  XOR U24721 ( .A(a[513]), .B(n42012), .Z(n23161) );
  XNOR U24722 ( .A(n23173), .B(n23172), .Z(n23175) );
  AND U24723 ( .A(a[515]), .B(b[0]), .Z(n23125) );
  XNOR U24724 ( .A(n23125), .B(n4071), .Z(n23127) );
  NANDN U24725 ( .A(b[0]), .B(a[514]), .Z(n23126) );
  NAND U24726 ( .A(n23127), .B(n23126), .Z(n23169) );
  XOR U24727 ( .A(a[511]), .B(n42085), .Z(n23165) );
  AND U24728 ( .A(a[507]), .B(b[7]), .Z(n23166) );
  XNOR U24729 ( .A(n23167), .B(n23166), .Z(n23168) );
  XNOR U24730 ( .A(n23169), .B(n23168), .Z(n23174) );
  XOR U24731 ( .A(n23175), .B(n23174), .Z(n23153) );
  NANDN U24732 ( .A(n23130), .B(n23129), .Z(n23134) );
  NANDN U24733 ( .A(n23132), .B(n23131), .Z(n23133) );
  AND U24734 ( .A(n23134), .B(n23133), .Z(n23152) );
  XNOR U24735 ( .A(n23153), .B(n23152), .Z(n23154) );
  NANDN U24736 ( .A(n23136), .B(n23135), .Z(n23140) );
  NAND U24737 ( .A(n23138), .B(n23137), .Z(n23139) );
  NAND U24738 ( .A(n23140), .B(n23139), .Z(n23155) );
  XNOR U24739 ( .A(n23154), .B(n23155), .Z(n23146) );
  XNOR U24740 ( .A(n23147), .B(n23146), .Z(n23148) );
  XNOR U24741 ( .A(n23149), .B(n23148), .Z(n23178) );
  XNOR U24742 ( .A(sreg[1531]), .B(n23178), .Z(n23180) );
  NANDN U24743 ( .A(sreg[1530]), .B(n23141), .Z(n23145) );
  NAND U24744 ( .A(n23143), .B(n23142), .Z(n23144) );
  NAND U24745 ( .A(n23145), .B(n23144), .Z(n23179) );
  XNOR U24746 ( .A(n23180), .B(n23179), .Z(c[1531]) );
  NANDN U24747 ( .A(n23147), .B(n23146), .Z(n23151) );
  NANDN U24748 ( .A(n23149), .B(n23148), .Z(n23150) );
  AND U24749 ( .A(n23151), .B(n23150), .Z(n23186) );
  NANDN U24750 ( .A(n23153), .B(n23152), .Z(n23157) );
  NANDN U24751 ( .A(n23155), .B(n23154), .Z(n23156) );
  AND U24752 ( .A(n23157), .B(n23156), .Z(n23184) );
  NAND U24753 ( .A(n42143), .B(n23158), .Z(n23160) );
  XNOR U24754 ( .A(a[510]), .B(n4144), .Z(n23195) );
  NAND U24755 ( .A(n42144), .B(n23195), .Z(n23159) );
  AND U24756 ( .A(n23160), .B(n23159), .Z(n23210) );
  XOR U24757 ( .A(a[514]), .B(n42012), .Z(n23198) );
  XNOR U24758 ( .A(n23210), .B(n23209), .Z(n23212) );
  AND U24759 ( .A(a[516]), .B(b[0]), .Z(n23162) );
  XNOR U24760 ( .A(n23162), .B(n4071), .Z(n23164) );
  NANDN U24761 ( .A(b[0]), .B(a[515]), .Z(n23163) );
  NAND U24762 ( .A(n23164), .B(n23163), .Z(n23206) );
  XOR U24763 ( .A(a[512]), .B(n42085), .Z(n23199) );
  AND U24764 ( .A(a[508]), .B(b[7]), .Z(n23203) );
  XNOR U24765 ( .A(n23204), .B(n23203), .Z(n23205) );
  XNOR U24766 ( .A(n23206), .B(n23205), .Z(n23211) );
  XOR U24767 ( .A(n23212), .B(n23211), .Z(n23190) );
  NANDN U24768 ( .A(n23167), .B(n23166), .Z(n23171) );
  NANDN U24769 ( .A(n23169), .B(n23168), .Z(n23170) );
  AND U24770 ( .A(n23171), .B(n23170), .Z(n23189) );
  XNOR U24771 ( .A(n23190), .B(n23189), .Z(n23191) );
  NANDN U24772 ( .A(n23173), .B(n23172), .Z(n23177) );
  NAND U24773 ( .A(n23175), .B(n23174), .Z(n23176) );
  NAND U24774 ( .A(n23177), .B(n23176), .Z(n23192) );
  XNOR U24775 ( .A(n23191), .B(n23192), .Z(n23183) );
  XNOR U24776 ( .A(n23184), .B(n23183), .Z(n23185) );
  XNOR U24777 ( .A(n23186), .B(n23185), .Z(n23215) );
  XNOR U24778 ( .A(sreg[1532]), .B(n23215), .Z(n23217) );
  NANDN U24779 ( .A(sreg[1531]), .B(n23178), .Z(n23182) );
  NAND U24780 ( .A(n23180), .B(n23179), .Z(n23181) );
  NAND U24781 ( .A(n23182), .B(n23181), .Z(n23216) );
  XNOR U24782 ( .A(n23217), .B(n23216), .Z(c[1532]) );
  NANDN U24783 ( .A(n23184), .B(n23183), .Z(n23188) );
  NANDN U24784 ( .A(n23186), .B(n23185), .Z(n23187) );
  AND U24785 ( .A(n23188), .B(n23187), .Z(n23223) );
  NANDN U24786 ( .A(n23190), .B(n23189), .Z(n23194) );
  NANDN U24787 ( .A(n23192), .B(n23191), .Z(n23193) );
  AND U24788 ( .A(n23194), .B(n23193), .Z(n23221) );
  NAND U24789 ( .A(n42143), .B(n23195), .Z(n23197) );
  XNOR U24790 ( .A(a[511]), .B(n4144), .Z(n23232) );
  NAND U24791 ( .A(n42144), .B(n23232), .Z(n23196) );
  AND U24792 ( .A(n23197), .B(n23196), .Z(n23247) );
  XOR U24793 ( .A(a[515]), .B(n42012), .Z(n23235) );
  XNOR U24794 ( .A(n23247), .B(n23246), .Z(n23249) );
  XOR U24795 ( .A(a[513]), .B(n42085), .Z(n23239) );
  AND U24796 ( .A(a[509]), .B(b[7]), .Z(n23240) );
  XNOR U24797 ( .A(n23241), .B(n23240), .Z(n23242) );
  AND U24798 ( .A(a[517]), .B(b[0]), .Z(n23200) );
  XNOR U24799 ( .A(n23200), .B(n4071), .Z(n23202) );
  NANDN U24800 ( .A(b[0]), .B(a[516]), .Z(n23201) );
  NAND U24801 ( .A(n23202), .B(n23201), .Z(n23243) );
  XNOR U24802 ( .A(n23242), .B(n23243), .Z(n23248) );
  XOR U24803 ( .A(n23249), .B(n23248), .Z(n23227) );
  NANDN U24804 ( .A(n23204), .B(n23203), .Z(n23208) );
  NANDN U24805 ( .A(n23206), .B(n23205), .Z(n23207) );
  AND U24806 ( .A(n23208), .B(n23207), .Z(n23226) );
  XNOR U24807 ( .A(n23227), .B(n23226), .Z(n23228) );
  NANDN U24808 ( .A(n23210), .B(n23209), .Z(n23214) );
  NAND U24809 ( .A(n23212), .B(n23211), .Z(n23213) );
  NAND U24810 ( .A(n23214), .B(n23213), .Z(n23229) );
  XNOR U24811 ( .A(n23228), .B(n23229), .Z(n23220) );
  XNOR U24812 ( .A(n23221), .B(n23220), .Z(n23222) );
  XNOR U24813 ( .A(n23223), .B(n23222), .Z(n23252) );
  XNOR U24814 ( .A(sreg[1533]), .B(n23252), .Z(n23254) );
  NANDN U24815 ( .A(sreg[1532]), .B(n23215), .Z(n23219) );
  NAND U24816 ( .A(n23217), .B(n23216), .Z(n23218) );
  NAND U24817 ( .A(n23219), .B(n23218), .Z(n23253) );
  XNOR U24818 ( .A(n23254), .B(n23253), .Z(c[1533]) );
  NANDN U24819 ( .A(n23221), .B(n23220), .Z(n23225) );
  NANDN U24820 ( .A(n23223), .B(n23222), .Z(n23224) );
  AND U24821 ( .A(n23225), .B(n23224), .Z(n23260) );
  NANDN U24822 ( .A(n23227), .B(n23226), .Z(n23231) );
  NANDN U24823 ( .A(n23229), .B(n23228), .Z(n23230) );
  AND U24824 ( .A(n23231), .B(n23230), .Z(n23258) );
  NAND U24825 ( .A(n42143), .B(n23232), .Z(n23234) );
  XNOR U24826 ( .A(a[512]), .B(n4145), .Z(n23269) );
  NAND U24827 ( .A(n42144), .B(n23269), .Z(n23233) );
  AND U24828 ( .A(n23234), .B(n23233), .Z(n23284) );
  XOR U24829 ( .A(a[516]), .B(n42012), .Z(n23272) );
  XNOR U24830 ( .A(n23284), .B(n23283), .Z(n23286) );
  AND U24831 ( .A(a[518]), .B(b[0]), .Z(n23236) );
  XNOR U24832 ( .A(n23236), .B(n4071), .Z(n23238) );
  NANDN U24833 ( .A(b[0]), .B(a[517]), .Z(n23237) );
  NAND U24834 ( .A(n23238), .B(n23237), .Z(n23280) );
  XOR U24835 ( .A(a[514]), .B(n42085), .Z(n23273) );
  AND U24836 ( .A(a[510]), .B(b[7]), .Z(n23277) );
  XNOR U24837 ( .A(n23278), .B(n23277), .Z(n23279) );
  XNOR U24838 ( .A(n23280), .B(n23279), .Z(n23285) );
  XOR U24839 ( .A(n23286), .B(n23285), .Z(n23264) );
  NANDN U24840 ( .A(n23241), .B(n23240), .Z(n23245) );
  NANDN U24841 ( .A(n23243), .B(n23242), .Z(n23244) );
  AND U24842 ( .A(n23245), .B(n23244), .Z(n23263) );
  XNOR U24843 ( .A(n23264), .B(n23263), .Z(n23265) );
  NANDN U24844 ( .A(n23247), .B(n23246), .Z(n23251) );
  NAND U24845 ( .A(n23249), .B(n23248), .Z(n23250) );
  NAND U24846 ( .A(n23251), .B(n23250), .Z(n23266) );
  XNOR U24847 ( .A(n23265), .B(n23266), .Z(n23257) );
  XNOR U24848 ( .A(n23258), .B(n23257), .Z(n23259) );
  XNOR U24849 ( .A(n23260), .B(n23259), .Z(n23289) );
  XNOR U24850 ( .A(sreg[1534]), .B(n23289), .Z(n23291) );
  NANDN U24851 ( .A(sreg[1533]), .B(n23252), .Z(n23256) );
  NAND U24852 ( .A(n23254), .B(n23253), .Z(n23255) );
  NAND U24853 ( .A(n23256), .B(n23255), .Z(n23290) );
  XNOR U24854 ( .A(n23291), .B(n23290), .Z(c[1534]) );
  NANDN U24855 ( .A(n23258), .B(n23257), .Z(n23262) );
  NANDN U24856 ( .A(n23260), .B(n23259), .Z(n23261) );
  AND U24857 ( .A(n23262), .B(n23261), .Z(n23297) );
  NANDN U24858 ( .A(n23264), .B(n23263), .Z(n23268) );
  NANDN U24859 ( .A(n23266), .B(n23265), .Z(n23267) );
  AND U24860 ( .A(n23268), .B(n23267), .Z(n23295) );
  NAND U24861 ( .A(n42143), .B(n23269), .Z(n23271) );
  XNOR U24862 ( .A(a[513]), .B(n4145), .Z(n23306) );
  NAND U24863 ( .A(n42144), .B(n23306), .Z(n23270) );
  AND U24864 ( .A(n23271), .B(n23270), .Z(n23321) );
  XOR U24865 ( .A(a[517]), .B(n42012), .Z(n23309) );
  XNOR U24866 ( .A(n23321), .B(n23320), .Z(n23323) );
  XOR U24867 ( .A(a[515]), .B(n42085), .Z(n23313) );
  AND U24868 ( .A(a[511]), .B(b[7]), .Z(n23314) );
  XNOR U24869 ( .A(n23315), .B(n23314), .Z(n23316) );
  AND U24870 ( .A(a[519]), .B(b[0]), .Z(n23274) );
  XNOR U24871 ( .A(n23274), .B(n4071), .Z(n23276) );
  NANDN U24872 ( .A(b[0]), .B(a[518]), .Z(n23275) );
  NAND U24873 ( .A(n23276), .B(n23275), .Z(n23317) );
  XNOR U24874 ( .A(n23316), .B(n23317), .Z(n23322) );
  XOR U24875 ( .A(n23323), .B(n23322), .Z(n23301) );
  NANDN U24876 ( .A(n23278), .B(n23277), .Z(n23282) );
  NANDN U24877 ( .A(n23280), .B(n23279), .Z(n23281) );
  AND U24878 ( .A(n23282), .B(n23281), .Z(n23300) );
  XNOR U24879 ( .A(n23301), .B(n23300), .Z(n23302) );
  NANDN U24880 ( .A(n23284), .B(n23283), .Z(n23288) );
  NAND U24881 ( .A(n23286), .B(n23285), .Z(n23287) );
  NAND U24882 ( .A(n23288), .B(n23287), .Z(n23303) );
  XNOR U24883 ( .A(n23302), .B(n23303), .Z(n23294) );
  XNOR U24884 ( .A(n23295), .B(n23294), .Z(n23296) );
  XNOR U24885 ( .A(n23297), .B(n23296), .Z(n23326) );
  XNOR U24886 ( .A(sreg[1535]), .B(n23326), .Z(n23328) );
  NANDN U24887 ( .A(sreg[1534]), .B(n23289), .Z(n23293) );
  NAND U24888 ( .A(n23291), .B(n23290), .Z(n23292) );
  NAND U24889 ( .A(n23293), .B(n23292), .Z(n23327) );
  XNOR U24890 ( .A(n23328), .B(n23327), .Z(c[1535]) );
  NANDN U24891 ( .A(n23295), .B(n23294), .Z(n23299) );
  NANDN U24892 ( .A(n23297), .B(n23296), .Z(n23298) );
  AND U24893 ( .A(n23299), .B(n23298), .Z(n23334) );
  NANDN U24894 ( .A(n23301), .B(n23300), .Z(n23305) );
  NANDN U24895 ( .A(n23303), .B(n23302), .Z(n23304) );
  AND U24896 ( .A(n23305), .B(n23304), .Z(n23332) );
  NAND U24897 ( .A(n42143), .B(n23306), .Z(n23308) );
  XNOR U24898 ( .A(a[514]), .B(n4145), .Z(n23343) );
  NAND U24899 ( .A(n42144), .B(n23343), .Z(n23307) );
  AND U24900 ( .A(n23308), .B(n23307), .Z(n23358) );
  XOR U24901 ( .A(a[518]), .B(n42012), .Z(n23346) );
  XNOR U24902 ( .A(n23358), .B(n23357), .Z(n23360) );
  AND U24903 ( .A(a[520]), .B(b[0]), .Z(n23310) );
  XNOR U24904 ( .A(n23310), .B(n4071), .Z(n23312) );
  NANDN U24905 ( .A(b[0]), .B(a[519]), .Z(n23311) );
  NAND U24906 ( .A(n23312), .B(n23311), .Z(n23354) );
  XOR U24907 ( .A(a[516]), .B(n42085), .Z(n23350) );
  AND U24908 ( .A(a[512]), .B(b[7]), .Z(n23351) );
  XNOR U24909 ( .A(n23352), .B(n23351), .Z(n23353) );
  XNOR U24910 ( .A(n23354), .B(n23353), .Z(n23359) );
  XOR U24911 ( .A(n23360), .B(n23359), .Z(n23338) );
  NANDN U24912 ( .A(n23315), .B(n23314), .Z(n23319) );
  NANDN U24913 ( .A(n23317), .B(n23316), .Z(n23318) );
  AND U24914 ( .A(n23319), .B(n23318), .Z(n23337) );
  XNOR U24915 ( .A(n23338), .B(n23337), .Z(n23339) );
  NANDN U24916 ( .A(n23321), .B(n23320), .Z(n23325) );
  NAND U24917 ( .A(n23323), .B(n23322), .Z(n23324) );
  NAND U24918 ( .A(n23325), .B(n23324), .Z(n23340) );
  XNOR U24919 ( .A(n23339), .B(n23340), .Z(n23331) );
  XNOR U24920 ( .A(n23332), .B(n23331), .Z(n23333) );
  XNOR U24921 ( .A(n23334), .B(n23333), .Z(n23363) );
  XNOR U24922 ( .A(sreg[1536]), .B(n23363), .Z(n23365) );
  NANDN U24923 ( .A(sreg[1535]), .B(n23326), .Z(n23330) );
  NAND U24924 ( .A(n23328), .B(n23327), .Z(n23329) );
  NAND U24925 ( .A(n23330), .B(n23329), .Z(n23364) );
  XNOR U24926 ( .A(n23365), .B(n23364), .Z(c[1536]) );
  NANDN U24927 ( .A(n23332), .B(n23331), .Z(n23336) );
  NANDN U24928 ( .A(n23334), .B(n23333), .Z(n23335) );
  AND U24929 ( .A(n23336), .B(n23335), .Z(n23371) );
  NANDN U24930 ( .A(n23338), .B(n23337), .Z(n23342) );
  NANDN U24931 ( .A(n23340), .B(n23339), .Z(n23341) );
  AND U24932 ( .A(n23342), .B(n23341), .Z(n23369) );
  NAND U24933 ( .A(n42143), .B(n23343), .Z(n23345) );
  XNOR U24934 ( .A(a[515]), .B(n4145), .Z(n23380) );
  NAND U24935 ( .A(n42144), .B(n23380), .Z(n23344) );
  AND U24936 ( .A(n23345), .B(n23344), .Z(n23395) );
  XOR U24937 ( .A(a[519]), .B(n42012), .Z(n23383) );
  XNOR U24938 ( .A(n23395), .B(n23394), .Z(n23397) );
  AND U24939 ( .A(a[521]), .B(b[0]), .Z(n23347) );
  XNOR U24940 ( .A(n23347), .B(n4071), .Z(n23349) );
  NANDN U24941 ( .A(b[0]), .B(a[520]), .Z(n23348) );
  NAND U24942 ( .A(n23349), .B(n23348), .Z(n23391) );
  XOR U24943 ( .A(a[517]), .B(n42085), .Z(n23384) );
  AND U24944 ( .A(a[513]), .B(b[7]), .Z(n23388) );
  XNOR U24945 ( .A(n23389), .B(n23388), .Z(n23390) );
  XNOR U24946 ( .A(n23391), .B(n23390), .Z(n23396) );
  XOR U24947 ( .A(n23397), .B(n23396), .Z(n23375) );
  NANDN U24948 ( .A(n23352), .B(n23351), .Z(n23356) );
  NANDN U24949 ( .A(n23354), .B(n23353), .Z(n23355) );
  AND U24950 ( .A(n23356), .B(n23355), .Z(n23374) );
  XNOR U24951 ( .A(n23375), .B(n23374), .Z(n23376) );
  NANDN U24952 ( .A(n23358), .B(n23357), .Z(n23362) );
  NAND U24953 ( .A(n23360), .B(n23359), .Z(n23361) );
  NAND U24954 ( .A(n23362), .B(n23361), .Z(n23377) );
  XNOR U24955 ( .A(n23376), .B(n23377), .Z(n23368) );
  XNOR U24956 ( .A(n23369), .B(n23368), .Z(n23370) );
  XNOR U24957 ( .A(n23371), .B(n23370), .Z(n23400) );
  XNOR U24958 ( .A(sreg[1537]), .B(n23400), .Z(n23402) );
  NANDN U24959 ( .A(sreg[1536]), .B(n23363), .Z(n23367) );
  NAND U24960 ( .A(n23365), .B(n23364), .Z(n23366) );
  NAND U24961 ( .A(n23367), .B(n23366), .Z(n23401) );
  XNOR U24962 ( .A(n23402), .B(n23401), .Z(c[1537]) );
  NANDN U24963 ( .A(n23369), .B(n23368), .Z(n23373) );
  NANDN U24964 ( .A(n23371), .B(n23370), .Z(n23372) );
  AND U24965 ( .A(n23373), .B(n23372), .Z(n23408) );
  NANDN U24966 ( .A(n23375), .B(n23374), .Z(n23379) );
  NANDN U24967 ( .A(n23377), .B(n23376), .Z(n23378) );
  AND U24968 ( .A(n23379), .B(n23378), .Z(n23406) );
  NAND U24969 ( .A(n42143), .B(n23380), .Z(n23382) );
  XNOR U24970 ( .A(a[516]), .B(n4145), .Z(n23417) );
  NAND U24971 ( .A(n42144), .B(n23417), .Z(n23381) );
  AND U24972 ( .A(n23382), .B(n23381), .Z(n23432) );
  XOR U24973 ( .A(a[520]), .B(n42012), .Z(n23420) );
  XNOR U24974 ( .A(n23432), .B(n23431), .Z(n23434) );
  XOR U24975 ( .A(a[518]), .B(n42085), .Z(n23421) );
  AND U24976 ( .A(a[514]), .B(b[7]), .Z(n23425) );
  XNOR U24977 ( .A(n23426), .B(n23425), .Z(n23427) );
  AND U24978 ( .A(a[522]), .B(b[0]), .Z(n23385) );
  XNOR U24979 ( .A(n23385), .B(n4071), .Z(n23387) );
  NANDN U24980 ( .A(b[0]), .B(a[521]), .Z(n23386) );
  NAND U24981 ( .A(n23387), .B(n23386), .Z(n23428) );
  XNOR U24982 ( .A(n23427), .B(n23428), .Z(n23433) );
  XOR U24983 ( .A(n23434), .B(n23433), .Z(n23412) );
  NANDN U24984 ( .A(n23389), .B(n23388), .Z(n23393) );
  NANDN U24985 ( .A(n23391), .B(n23390), .Z(n23392) );
  AND U24986 ( .A(n23393), .B(n23392), .Z(n23411) );
  XNOR U24987 ( .A(n23412), .B(n23411), .Z(n23413) );
  NANDN U24988 ( .A(n23395), .B(n23394), .Z(n23399) );
  NAND U24989 ( .A(n23397), .B(n23396), .Z(n23398) );
  NAND U24990 ( .A(n23399), .B(n23398), .Z(n23414) );
  XNOR U24991 ( .A(n23413), .B(n23414), .Z(n23405) );
  XNOR U24992 ( .A(n23406), .B(n23405), .Z(n23407) );
  XNOR U24993 ( .A(n23408), .B(n23407), .Z(n23437) );
  XNOR U24994 ( .A(sreg[1538]), .B(n23437), .Z(n23439) );
  NANDN U24995 ( .A(sreg[1537]), .B(n23400), .Z(n23404) );
  NAND U24996 ( .A(n23402), .B(n23401), .Z(n23403) );
  NAND U24997 ( .A(n23404), .B(n23403), .Z(n23438) );
  XNOR U24998 ( .A(n23439), .B(n23438), .Z(c[1538]) );
  NANDN U24999 ( .A(n23406), .B(n23405), .Z(n23410) );
  NANDN U25000 ( .A(n23408), .B(n23407), .Z(n23409) );
  AND U25001 ( .A(n23410), .B(n23409), .Z(n23445) );
  NANDN U25002 ( .A(n23412), .B(n23411), .Z(n23416) );
  NANDN U25003 ( .A(n23414), .B(n23413), .Z(n23415) );
  AND U25004 ( .A(n23416), .B(n23415), .Z(n23443) );
  NAND U25005 ( .A(n42143), .B(n23417), .Z(n23419) );
  XNOR U25006 ( .A(a[517]), .B(n4145), .Z(n23454) );
  NAND U25007 ( .A(n42144), .B(n23454), .Z(n23418) );
  AND U25008 ( .A(n23419), .B(n23418), .Z(n23469) );
  XOR U25009 ( .A(a[521]), .B(n42012), .Z(n23457) );
  XNOR U25010 ( .A(n23469), .B(n23468), .Z(n23471) );
  XOR U25011 ( .A(a[519]), .B(n42085), .Z(n23458) );
  AND U25012 ( .A(a[515]), .B(b[7]), .Z(n23462) );
  XNOR U25013 ( .A(n23463), .B(n23462), .Z(n23464) );
  AND U25014 ( .A(a[523]), .B(b[0]), .Z(n23422) );
  XNOR U25015 ( .A(n23422), .B(n4071), .Z(n23424) );
  NANDN U25016 ( .A(b[0]), .B(a[522]), .Z(n23423) );
  NAND U25017 ( .A(n23424), .B(n23423), .Z(n23465) );
  XNOR U25018 ( .A(n23464), .B(n23465), .Z(n23470) );
  XOR U25019 ( .A(n23471), .B(n23470), .Z(n23449) );
  NANDN U25020 ( .A(n23426), .B(n23425), .Z(n23430) );
  NANDN U25021 ( .A(n23428), .B(n23427), .Z(n23429) );
  AND U25022 ( .A(n23430), .B(n23429), .Z(n23448) );
  XNOR U25023 ( .A(n23449), .B(n23448), .Z(n23450) );
  NANDN U25024 ( .A(n23432), .B(n23431), .Z(n23436) );
  NAND U25025 ( .A(n23434), .B(n23433), .Z(n23435) );
  NAND U25026 ( .A(n23436), .B(n23435), .Z(n23451) );
  XNOR U25027 ( .A(n23450), .B(n23451), .Z(n23442) );
  XNOR U25028 ( .A(n23443), .B(n23442), .Z(n23444) );
  XNOR U25029 ( .A(n23445), .B(n23444), .Z(n23474) );
  XNOR U25030 ( .A(sreg[1539]), .B(n23474), .Z(n23476) );
  NANDN U25031 ( .A(sreg[1538]), .B(n23437), .Z(n23441) );
  NAND U25032 ( .A(n23439), .B(n23438), .Z(n23440) );
  NAND U25033 ( .A(n23441), .B(n23440), .Z(n23475) );
  XNOR U25034 ( .A(n23476), .B(n23475), .Z(c[1539]) );
  NANDN U25035 ( .A(n23443), .B(n23442), .Z(n23447) );
  NANDN U25036 ( .A(n23445), .B(n23444), .Z(n23446) );
  AND U25037 ( .A(n23447), .B(n23446), .Z(n23482) );
  NANDN U25038 ( .A(n23449), .B(n23448), .Z(n23453) );
  NANDN U25039 ( .A(n23451), .B(n23450), .Z(n23452) );
  AND U25040 ( .A(n23453), .B(n23452), .Z(n23480) );
  NAND U25041 ( .A(n42143), .B(n23454), .Z(n23456) );
  XNOR U25042 ( .A(a[518]), .B(n4145), .Z(n23491) );
  NAND U25043 ( .A(n42144), .B(n23491), .Z(n23455) );
  AND U25044 ( .A(n23456), .B(n23455), .Z(n23506) );
  XOR U25045 ( .A(a[522]), .B(n42012), .Z(n23494) );
  XNOR U25046 ( .A(n23506), .B(n23505), .Z(n23508) );
  XOR U25047 ( .A(a[520]), .B(n42085), .Z(n23498) );
  AND U25048 ( .A(a[516]), .B(b[7]), .Z(n23499) );
  XNOR U25049 ( .A(n23500), .B(n23499), .Z(n23501) );
  AND U25050 ( .A(a[524]), .B(b[0]), .Z(n23459) );
  XNOR U25051 ( .A(n23459), .B(n4071), .Z(n23461) );
  NANDN U25052 ( .A(b[0]), .B(a[523]), .Z(n23460) );
  NAND U25053 ( .A(n23461), .B(n23460), .Z(n23502) );
  XNOR U25054 ( .A(n23501), .B(n23502), .Z(n23507) );
  XOR U25055 ( .A(n23508), .B(n23507), .Z(n23486) );
  NANDN U25056 ( .A(n23463), .B(n23462), .Z(n23467) );
  NANDN U25057 ( .A(n23465), .B(n23464), .Z(n23466) );
  AND U25058 ( .A(n23467), .B(n23466), .Z(n23485) );
  XNOR U25059 ( .A(n23486), .B(n23485), .Z(n23487) );
  NANDN U25060 ( .A(n23469), .B(n23468), .Z(n23473) );
  NAND U25061 ( .A(n23471), .B(n23470), .Z(n23472) );
  NAND U25062 ( .A(n23473), .B(n23472), .Z(n23488) );
  XNOR U25063 ( .A(n23487), .B(n23488), .Z(n23479) );
  XNOR U25064 ( .A(n23480), .B(n23479), .Z(n23481) );
  XNOR U25065 ( .A(n23482), .B(n23481), .Z(n23511) );
  XNOR U25066 ( .A(sreg[1540]), .B(n23511), .Z(n23513) );
  NANDN U25067 ( .A(sreg[1539]), .B(n23474), .Z(n23478) );
  NAND U25068 ( .A(n23476), .B(n23475), .Z(n23477) );
  NAND U25069 ( .A(n23478), .B(n23477), .Z(n23512) );
  XNOR U25070 ( .A(n23513), .B(n23512), .Z(c[1540]) );
  NANDN U25071 ( .A(n23480), .B(n23479), .Z(n23484) );
  NANDN U25072 ( .A(n23482), .B(n23481), .Z(n23483) );
  AND U25073 ( .A(n23484), .B(n23483), .Z(n23519) );
  NANDN U25074 ( .A(n23486), .B(n23485), .Z(n23490) );
  NANDN U25075 ( .A(n23488), .B(n23487), .Z(n23489) );
  AND U25076 ( .A(n23490), .B(n23489), .Z(n23517) );
  NAND U25077 ( .A(n42143), .B(n23491), .Z(n23493) );
  XNOR U25078 ( .A(a[519]), .B(n4146), .Z(n23528) );
  NAND U25079 ( .A(n42144), .B(n23528), .Z(n23492) );
  AND U25080 ( .A(n23493), .B(n23492), .Z(n23543) );
  XOR U25081 ( .A(a[523]), .B(n42012), .Z(n23531) );
  XNOR U25082 ( .A(n23543), .B(n23542), .Z(n23545) );
  AND U25083 ( .A(a[525]), .B(b[0]), .Z(n23495) );
  XNOR U25084 ( .A(n23495), .B(n4071), .Z(n23497) );
  NANDN U25085 ( .A(b[0]), .B(a[524]), .Z(n23496) );
  NAND U25086 ( .A(n23497), .B(n23496), .Z(n23539) );
  XOR U25087 ( .A(a[521]), .B(n42085), .Z(n23535) );
  AND U25088 ( .A(a[517]), .B(b[7]), .Z(n23536) );
  XNOR U25089 ( .A(n23537), .B(n23536), .Z(n23538) );
  XNOR U25090 ( .A(n23539), .B(n23538), .Z(n23544) );
  XOR U25091 ( .A(n23545), .B(n23544), .Z(n23523) );
  NANDN U25092 ( .A(n23500), .B(n23499), .Z(n23504) );
  NANDN U25093 ( .A(n23502), .B(n23501), .Z(n23503) );
  AND U25094 ( .A(n23504), .B(n23503), .Z(n23522) );
  XNOR U25095 ( .A(n23523), .B(n23522), .Z(n23524) );
  NANDN U25096 ( .A(n23506), .B(n23505), .Z(n23510) );
  NAND U25097 ( .A(n23508), .B(n23507), .Z(n23509) );
  NAND U25098 ( .A(n23510), .B(n23509), .Z(n23525) );
  XNOR U25099 ( .A(n23524), .B(n23525), .Z(n23516) );
  XNOR U25100 ( .A(n23517), .B(n23516), .Z(n23518) );
  XNOR U25101 ( .A(n23519), .B(n23518), .Z(n23548) );
  XNOR U25102 ( .A(sreg[1541]), .B(n23548), .Z(n23550) );
  NANDN U25103 ( .A(sreg[1540]), .B(n23511), .Z(n23515) );
  NAND U25104 ( .A(n23513), .B(n23512), .Z(n23514) );
  NAND U25105 ( .A(n23515), .B(n23514), .Z(n23549) );
  XNOR U25106 ( .A(n23550), .B(n23549), .Z(c[1541]) );
  NANDN U25107 ( .A(n23517), .B(n23516), .Z(n23521) );
  NANDN U25108 ( .A(n23519), .B(n23518), .Z(n23520) );
  AND U25109 ( .A(n23521), .B(n23520), .Z(n23556) );
  NANDN U25110 ( .A(n23523), .B(n23522), .Z(n23527) );
  NANDN U25111 ( .A(n23525), .B(n23524), .Z(n23526) );
  AND U25112 ( .A(n23527), .B(n23526), .Z(n23554) );
  NAND U25113 ( .A(n42143), .B(n23528), .Z(n23530) );
  XNOR U25114 ( .A(a[520]), .B(n4146), .Z(n23565) );
  NAND U25115 ( .A(n42144), .B(n23565), .Z(n23529) );
  AND U25116 ( .A(n23530), .B(n23529), .Z(n23580) );
  XOR U25117 ( .A(a[524]), .B(n42012), .Z(n23568) );
  XNOR U25118 ( .A(n23580), .B(n23579), .Z(n23582) );
  AND U25119 ( .A(a[526]), .B(b[0]), .Z(n23532) );
  XNOR U25120 ( .A(n23532), .B(n4071), .Z(n23534) );
  NANDN U25121 ( .A(b[0]), .B(a[525]), .Z(n23533) );
  NAND U25122 ( .A(n23534), .B(n23533), .Z(n23576) );
  XOR U25123 ( .A(a[522]), .B(n42085), .Z(n23572) );
  AND U25124 ( .A(a[518]), .B(b[7]), .Z(n23573) );
  XNOR U25125 ( .A(n23574), .B(n23573), .Z(n23575) );
  XNOR U25126 ( .A(n23576), .B(n23575), .Z(n23581) );
  XOR U25127 ( .A(n23582), .B(n23581), .Z(n23560) );
  NANDN U25128 ( .A(n23537), .B(n23536), .Z(n23541) );
  NANDN U25129 ( .A(n23539), .B(n23538), .Z(n23540) );
  AND U25130 ( .A(n23541), .B(n23540), .Z(n23559) );
  XNOR U25131 ( .A(n23560), .B(n23559), .Z(n23561) );
  NANDN U25132 ( .A(n23543), .B(n23542), .Z(n23547) );
  NAND U25133 ( .A(n23545), .B(n23544), .Z(n23546) );
  NAND U25134 ( .A(n23547), .B(n23546), .Z(n23562) );
  XNOR U25135 ( .A(n23561), .B(n23562), .Z(n23553) );
  XNOR U25136 ( .A(n23554), .B(n23553), .Z(n23555) );
  XNOR U25137 ( .A(n23556), .B(n23555), .Z(n23585) );
  XNOR U25138 ( .A(sreg[1542]), .B(n23585), .Z(n23587) );
  NANDN U25139 ( .A(sreg[1541]), .B(n23548), .Z(n23552) );
  NAND U25140 ( .A(n23550), .B(n23549), .Z(n23551) );
  NAND U25141 ( .A(n23552), .B(n23551), .Z(n23586) );
  XNOR U25142 ( .A(n23587), .B(n23586), .Z(c[1542]) );
  NANDN U25143 ( .A(n23554), .B(n23553), .Z(n23558) );
  NANDN U25144 ( .A(n23556), .B(n23555), .Z(n23557) );
  AND U25145 ( .A(n23558), .B(n23557), .Z(n23593) );
  NANDN U25146 ( .A(n23560), .B(n23559), .Z(n23564) );
  NANDN U25147 ( .A(n23562), .B(n23561), .Z(n23563) );
  AND U25148 ( .A(n23564), .B(n23563), .Z(n23591) );
  NAND U25149 ( .A(n42143), .B(n23565), .Z(n23567) );
  XNOR U25150 ( .A(a[521]), .B(n4146), .Z(n23602) );
  NAND U25151 ( .A(n42144), .B(n23602), .Z(n23566) );
  AND U25152 ( .A(n23567), .B(n23566), .Z(n23617) );
  XOR U25153 ( .A(a[525]), .B(n42012), .Z(n23605) );
  XNOR U25154 ( .A(n23617), .B(n23616), .Z(n23619) );
  AND U25155 ( .A(a[527]), .B(b[0]), .Z(n23569) );
  XNOR U25156 ( .A(n23569), .B(n4071), .Z(n23571) );
  NANDN U25157 ( .A(b[0]), .B(a[526]), .Z(n23570) );
  NAND U25158 ( .A(n23571), .B(n23570), .Z(n23613) );
  XOR U25159 ( .A(a[523]), .B(n42085), .Z(n23606) );
  AND U25160 ( .A(a[519]), .B(b[7]), .Z(n23610) );
  XNOR U25161 ( .A(n23611), .B(n23610), .Z(n23612) );
  XNOR U25162 ( .A(n23613), .B(n23612), .Z(n23618) );
  XOR U25163 ( .A(n23619), .B(n23618), .Z(n23597) );
  NANDN U25164 ( .A(n23574), .B(n23573), .Z(n23578) );
  NANDN U25165 ( .A(n23576), .B(n23575), .Z(n23577) );
  AND U25166 ( .A(n23578), .B(n23577), .Z(n23596) );
  XNOR U25167 ( .A(n23597), .B(n23596), .Z(n23598) );
  NANDN U25168 ( .A(n23580), .B(n23579), .Z(n23584) );
  NAND U25169 ( .A(n23582), .B(n23581), .Z(n23583) );
  NAND U25170 ( .A(n23584), .B(n23583), .Z(n23599) );
  XNOR U25171 ( .A(n23598), .B(n23599), .Z(n23590) );
  XNOR U25172 ( .A(n23591), .B(n23590), .Z(n23592) );
  XNOR U25173 ( .A(n23593), .B(n23592), .Z(n23622) );
  XNOR U25174 ( .A(sreg[1543]), .B(n23622), .Z(n23624) );
  NANDN U25175 ( .A(sreg[1542]), .B(n23585), .Z(n23589) );
  NAND U25176 ( .A(n23587), .B(n23586), .Z(n23588) );
  NAND U25177 ( .A(n23589), .B(n23588), .Z(n23623) );
  XNOR U25178 ( .A(n23624), .B(n23623), .Z(c[1543]) );
  NANDN U25179 ( .A(n23591), .B(n23590), .Z(n23595) );
  NANDN U25180 ( .A(n23593), .B(n23592), .Z(n23594) );
  AND U25181 ( .A(n23595), .B(n23594), .Z(n23630) );
  NANDN U25182 ( .A(n23597), .B(n23596), .Z(n23601) );
  NANDN U25183 ( .A(n23599), .B(n23598), .Z(n23600) );
  AND U25184 ( .A(n23601), .B(n23600), .Z(n23628) );
  NAND U25185 ( .A(n42143), .B(n23602), .Z(n23604) );
  XNOR U25186 ( .A(a[522]), .B(n4146), .Z(n23639) );
  NAND U25187 ( .A(n42144), .B(n23639), .Z(n23603) );
  AND U25188 ( .A(n23604), .B(n23603), .Z(n23654) );
  XOR U25189 ( .A(a[526]), .B(n42012), .Z(n23642) );
  XNOR U25190 ( .A(n23654), .B(n23653), .Z(n23656) );
  XOR U25191 ( .A(a[524]), .B(n42085), .Z(n23646) );
  AND U25192 ( .A(a[520]), .B(b[7]), .Z(n23647) );
  XNOR U25193 ( .A(n23648), .B(n23647), .Z(n23649) );
  AND U25194 ( .A(a[528]), .B(b[0]), .Z(n23607) );
  XNOR U25195 ( .A(n23607), .B(n4071), .Z(n23609) );
  NANDN U25196 ( .A(b[0]), .B(a[527]), .Z(n23608) );
  NAND U25197 ( .A(n23609), .B(n23608), .Z(n23650) );
  XNOR U25198 ( .A(n23649), .B(n23650), .Z(n23655) );
  XOR U25199 ( .A(n23656), .B(n23655), .Z(n23634) );
  NANDN U25200 ( .A(n23611), .B(n23610), .Z(n23615) );
  NANDN U25201 ( .A(n23613), .B(n23612), .Z(n23614) );
  AND U25202 ( .A(n23615), .B(n23614), .Z(n23633) );
  XNOR U25203 ( .A(n23634), .B(n23633), .Z(n23635) );
  NANDN U25204 ( .A(n23617), .B(n23616), .Z(n23621) );
  NAND U25205 ( .A(n23619), .B(n23618), .Z(n23620) );
  NAND U25206 ( .A(n23621), .B(n23620), .Z(n23636) );
  XNOR U25207 ( .A(n23635), .B(n23636), .Z(n23627) );
  XNOR U25208 ( .A(n23628), .B(n23627), .Z(n23629) );
  XNOR U25209 ( .A(n23630), .B(n23629), .Z(n23659) );
  XNOR U25210 ( .A(sreg[1544]), .B(n23659), .Z(n23661) );
  NANDN U25211 ( .A(sreg[1543]), .B(n23622), .Z(n23626) );
  NAND U25212 ( .A(n23624), .B(n23623), .Z(n23625) );
  NAND U25213 ( .A(n23626), .B(n23625), .Z(n23660) );
  XNOR U25214 ( .A(n23661), .B(n23660), .Z(c[1544]) );
  NANDN U25215 ( .A(n23628), .B(n23627), .Z(n23632) );
  NANDN U25216 ( .A(n23630), .B(n23629), .Z(n23631) );
  AND U25217 ( .A(n23632), .B(n23631), .Z(n23667) );
  NANDN U25218 ( .A(n23634), .B(n23633), .Z(n23638) );
  NANDN U25219 ( .A(n23636), .B(n23635), .Z(n23637) );
  AND U25220 ( .A(n23638), .B(n23637), .Z(n23665) );
  NAND U25221 ( .A(n42143), .B(n23639), .Z(n23641) );
  XNOR U25222 ( .A(a[523]), .B(n4146), .Z(n23676) );
  NAND U25223 ( .A(n42144), .B(n23676), .Z(n23640) );
  AND U25224 ( .A(n23641), .B(n23640), .Z(n23691) );
  XOR U25225 ( .A(a[527]), .B(n42012), .Z(n23679) );
  XNOR U25226 ( .A(n23691), .B(n23690), .Z(n23693) );
  AND U25227 ( .A(a[529]), .B(b[0]), .Z(n23643) );
  XNOR U25228 ( .A(n23643), .B(n4071), .Z(n23645) );
  NANDN U25229 ( .A(b[0]), .B(a[528]), .Z(n23644) );
  NAND U25230 ( .A(n23645), .B(n23644), .Z(n23687) );
  XOR U25231 ( .A(a[525]), .B(n42085), .Z(n23683) );
  AND U25232 ( .A(a[521]), .B(b[7]), .Z(n23684) );
  XNOR U25233 ( .A(n23685), .B(n23684), .Z(n23686) );
  XNOR U25234 ( .A(n23687), .B(n23686), .Z(n23692) );
  XOR U25235 ( .A(n23693), .B(n23692), .Z(n23671) );
  NANDN U25236 ( .A(n23648), .B(n23647), .Z(n23652) );
  NANDN U25237 ( .A(n23650), .B(n23649), .Z(n23651) );
  AND U25238 ( .A(n23652), .B(n23651), .Z(n23670) );
  XNOR U25239 ( .A(n23671), .B(n23670), .Z(n23672) );
  NANDN U25240 ( .A(n23654), .B(n23653), .Z(n23658) );
  NAND U25241 ( .A(n23656), .B(n23655), .Z(n23657) );
  NAND U25242 ( .A(n23658), .B(n23657), .Z(n23673) );
  XNOR U25243 ( .A(n23672), .B(n23673), .Z(n23664) );
  XNOR U25244 ( .A(n23665), .B(n23664), .Z(n23666) );
  XNOR U25245 ( .A(n23667), .B(n23666), .Z(n23696) );
  XNOR U25246 ( .A(sreg[1545]), .B(n23696), .Z(n23698) );
  NANDN U25247 ( .A(sreg[1544]), .B(n23659), .Z(n23663) );
  NAND U25248 ( .A(n23661), .B(n23660), .Z(n23662) );
  NAND U25249 ( .A(n23663), .B(n23662), .Z(n23697) );
  XNOR U25250 ( .A(n23698), .B(n23697), .Z(c[1545]) );
  NANDN U25251 ( .A(n23665), .B(n23664), .Z(n23669) );
  NANDN U25252 ( .A(n23667), .B(n23666), .Z(n23668) );
  AND U25253 ( .A(n23669), .B(n23668), .Z(n23704) );
  NANDN U25254 ( .A(n23671), .B(n23670), .Z(n23675) );
  NANDN U25255 ( .A(n23673), .B(n23672), .Z(n23674) );
  AND U25256 ( .A(n23675), .B(n23674), .Z(n23702) );
  NAND U25257 ( .A(n42143), .B(n23676), .Z(n23678) );
  XNOR U25258 ( .A(a[524]), .B(n4146), .Z(n23713) );
  NAND U25259 ( .A(n42144), .B(n23713), .Z(n23677) );
  AND U25260 ( .A(n23678), .B(n23677), .Z(n23728) );
  XOR U25261 ( .A(a[528]), .B(n42012), .Z(n23716) );
  XNOR U25262 ( .A(n23728), .B(n23727), .Z(n23730) );
  AND U25263 ( .A(a[530]), .B(b[0]), .Z(n23680) );
  XNOR U25264 ( .A(n23680), .B(n4071), .Z(n23682) );
  NANDN U25265 ( .A(b[0]), .B(a[529]), .Z(n23681) );
  NAND U25266 ( .A(n23682), .B(n23681), .Z(n23724) );
  XOR U25267 ( .A(a[526]), .B(n42085), .Z(n23717) );
  AND U25268 ( .A(a[522]), .B(b[7]), .Z(n23721) );
  XNOR U25269 ( .A(n23722), .B(n23721), .Z(n23723) );
  XNOR U25270 ( .A(n23724), .B(n23723), .Z(n23729) );
  XOR U25271 ( .A(n23730), .B(n23729), .Z(n23708) );
  NANDN U25272 ( .A(n23685), .B(n23684), .Z(n23689) );
  NANDN U25273 ( .A(n23687), .B(n23686), .Z(n23688) );
  AND U25274 ( .A(n23689), .B(n23688), .Z(n23707) );
  XNOR U25275 ( .A(n23708), .B(n23707), .Z(n23709) );
  NANDN U25276 ( .A(n23691), .B(n23690), .Z(n23695) );
  NAND U25277 ( .A(n23693), .B(n23692), .Z(n23694) );
  NAND U25278 ( .A(n23695), .B(n23694), .Z(n23710) );
  XNOR U25279 ( .A(n23709), .B(n23710), .Z(n23701) );
  XNOR U25280 ( .A(n23702), .B(n23701), .Z(n23703) );
  XNOR U25281 ( .A(n23704), .B(n23703), .Z(n23733) );
  XNOR U25282 ( .A(sreg[1546]), .B(n23733), .Z(n23735) );
  NANDN U25283 ( .A(sreg[1545]), .B(n23696), .Z(n23700) );
  NAND U25284 ( .A(n23698), .B(n23697), .Z(n23699) );
  NAND U25285 ( .A(n23700), .B(n23699), .Z(n23734) );
  XNOR U25286 ( .A(n23735), .B(n23734), .Z(c[1546]) );
  NANDN U25287 ( .A(n23702), .B(n23701), .Z(n23706) );
  NANDN U25288 ( .A(n23704), .B(n23703), .Z(n23705) );
  AND U25289 ( .A(n23706), .B(n23705), .Z(n23741) );
  NANDN U25290 ( .A(n23708), .B(n23707), .Z(n23712) );
  NANDN U25291 ( .A(n23710), .B(n23709), .Z(n23711) );
  AND U25292 ( .A(n23712), .B(n23711), .Z(n23739) );
  NAND U25293 ( .A(n42143), .B(n23713), .Z(n23715) );
  XNOR U25294 ( .A(a[525]), .B(n4146), .Z(n23750) );
  NAND U25295 ( .A(n42144), .B(n23750), .Z(n23714) );
  AND U25296 ( .A(n23715), .B(n23714), .Z(n23765) );
  XOR U25297 ( .A(a[529]), .B(n42012), .Z(n23753) );
  XNOR U25298 ( .A(n23765), .B(n23764), .Z(n23767) );
  XOR U25299 ( .A(a[527]), .B(n42085), .Z(n23757) );
  AND U25300 ( .A(a[523]), .B(b[7]), .Z(n23758) );
  XNOR U25301 ( .A(n23759), .B(n23758), .Z(n23760) );
  AND U25302 ( .A(a[531]), .B(b[0]), .Z(n23718) );
  XNOR U25303 ( .A(n23718), .B(n4071), .Z(n23720) );
  NANDN U25304 ( .A(b[0]), .B(a[530]), .Z(n23719) );
  NAND U25305 ( .A(n23720), .B(n23719), .Z(n23761) );
  XNOR U25306 ( .A(n23760), .B(n23761), .Z(n23766) );
  XOR U25307 ( .A(n23767), .B(n23766), .Z(n23745) );
  NANDN U25308 ( .A(n23722), .B(n23721), .Z(n23726) );
  NANDN U25309 ( .A(n23724), .B(n23723), .Z(n23725) );
  AND U25310 ( .A(n23726), .B(n23725), .Z(n23744) );
  XNOR U25311 ( .A(n23745), .B(n23744), .Z(n23746) );
  NANDN U25312 ( .A(n23728), .B(n23727), .Z(n23732) );
  NAND U25313 ( .A(n23730), .B(n23729), .Z(n23731) );
  NAND U25314 ( .A(n23732), .B(n23731), .Z(n23747) );
  XNOR U25315 ( .A(n23746), .B(n23747), .Z(n23738) );
  XNOR U25316 ( .A(n23739), .B(n23738), .Z(n23740) );
  XNOR U25317 ( .A(n23741), .B(n23740), .Z(n23770) );
  XNOR U25318 ( .A(sreg[1547]), .B(n23770), .Z(n23772) );
  NANDN U25319 ( .A(sreg[1546]), .B(n23733), .Z(n23737) );
  NAND U25320 ( .A(n23735), .B(n23734), .Z(n23736) );
  NAND U25321 ( .A(n23737), .B(n23736), .Z(n23771) );
  XNOR U25322 ( .A(n23772), .B(n23771), .Z(c[1547]) );
  NANDN U25323 ( .A(n23739), .B(n23738), .Z(n23743) );
  NANDN U25324 ( .A(n23741), .B(n23740), .Z(n23742) );
  AND U25325 ( .A(n23743), .B(n23742), .Z(n23778) );
  NANDN U25326 ( .A(n23745), .B(n23744), .Z(n23749) );
  NANDN U25327 ( .A(n23747), .B(n23746), .Z(n23748) );
  AND U25328 ( .A(n23749), .B(n23748), .Z(n23776) );
  NAND U25329 ( .A(n42143), .B(n23750), .Z(n23752) );
  XNOR U25330 ( .A(a[526]), .B(n4147), .Z(n23787) );
  NAND U25331 ( .A(n42144), .B(n23787), .Z(n23751) );
  AND U25332 ( .A(n23752), .B(n23751), .Z(n23802) );
  XOR U25333 ( .A(a[530]), .B(n42012), .Z(n23790) );
  XNOR U25334 ( .A(n23802), .B(n23801), .Z(n23804) );
  AND U25335 ( .A(a[532]), .B(b[0]), .Z(n23754) );
  XNOR U25336 ( .A(n23754), .B(n4071), .Z(n23756) );
  NANDN U25337 ( .A(b[0]), .B(a[531]), .Z(n23755) );
  NAND U25338 ( .A(n23756), .B(n23755), .Z(n23798) );
  XOR U25339 ( .A(a[528]), .B(n42085), .Z(n23794) );
  AND U25340 ( .A(a[524]), .B(b[7]), .Z(n23795) );
  XNOR U25341 ( .A(n23796), .B(n23795), .Z(n23797) );
  XNOR U25342 ( .A(n23798), .B(n23797), .Z(n23803) );
  XOR U25343 ( .A(n23804), .B(n23803), .Z(n23782) );
  NANDN U25344 ( .A(n23759), .B(n23758), .Z(n23763) );
  NANDN U25345 ( .A(n23761), .B(n23760), .Z(n23762) );
  AND U25346 ( .A(n23763), .B(n23762), .Z(n23781) );
  XNOR U25347 ( .A(n23782), .B(n23781), .Z(n23783) );
  NANDN U25348 ( .A(n23765), .B(n23764), .Z(n23769) );
  NAND U25349 ( .A(n23767), .B(n23766), .Z(n23768) );
  NAND U25350 ( .A(n23769), .B(n23768), .Z(n23784) );
  XNOR U25351 ( .A(n23783), .B(n23784), .Z(n23775) );
  XNOR U25352 ( .A(n23776), .B(n23775), .Z(n23777) );
  XNOR U25353 ( .A(n23778), .B(n23777), .Z(n23807) );
  XNOR U25354 ( .A(sreg[1548]), .B(n23807), .Z(n23809) );
  NANDN U25355 ( .A(sreg[1547]), .B(n23770), .Z(n23774) );
  NAND U25356 ( .A(n23772), .B(n23771), .Z(n23773) );
  NAND U25357 ( .A(n23774), .B(n23773), .Z(n23808) );
  XNOR U25358 ( .A(n23809), .B(n23808), .Z(c[1548]) );
  NANDN U25359 ( .A(n23776), .B(n23775), .Z(n23780) );
  NANDN U25360 ( .A(n23778), .B(n23777), .Z(n23779) );
  AND U25361 ( .A(n23780), .B(n23779), .Z(n23815) );
  NANDN U25362 ( .A(n23782), .B(n23781), .Z(n23786) );
  NANDN U25363 ( .A(n23784), .B(n23783), .Z(n23785) );
  AND U25364 ( .A(n23786), .B(n23785), .Z(n23813) );
  NAND U25365 ( .A(n42143), .B(n23787), .Z(n23789) );
  XNOR U25366 ( .A(a[527]), .B(n4147), .Z(n23824) );
  NAND U25367 ( .A(n42144), .B(n23824), .Z(n23788) );
  AND U25368 ( .A(n23789), .B(n23788), .Z(n23839) );
  XOR U25369 ( .A(a[531]), .B(n42012), .Z(n23827) );
  XNOR U25370 ( .A(n23839), .B(n23838), .Z(n23841) );
  AND U25371 ( .A(a[533]), .B(b[0]), .Z(n23791) );
  XNOR U25372 ( .A(n23791), .B(n4071), .Z(n23793) );
  NANDN U25373 ( .A(b[0]), .B(a[532]), .Z(n23792) );
  NAND U25374 ( .A(n23793), .B(n23792), .Z(n23835) );
  XOR U25375 ( .A(a[529]), .B(n42085), .Z(n23828) );
  AND U25376 ( .A(a[525]), .B(b[7]), .Z(n23832) );
  XNOR U25377 ( .A(n23833), .B(n23832), .Z(n23834) );
  XNOR U25378 ( .A(n23835), .B(n23834), .Z(n23840) );
  XOR U25379 ( .A(n23841), .B(n23840), .Z(n23819) );
  NANDN U25380 ( .A(n23796), .B(n23795), .Z(n23800) );
  NANDN U25381 ( .A(n23798), .B(n23797), .Z(n23799) );
  AND U25382 ( .A(n23800), .B(n23799), .Z(n23818) );
  XNOR U25383 ( .A(n23819), .B(n23818), .Z(n23820) );
  NANDN U25384 ( .A(n23802), .B(n23801), .Z(n23806) );
  NAND U25385 ( .A(n23804), .B(n23803), .Z(n23805) );
  NAND U25386 ( .A(n23806), .B(n23805), .Z(n23821) );
  XNOR U25387 ( .A(n23820), .B(n23821), .Z(n23812) );
  XNOR U25388 ( .A(n23813), .B(n23812), .Z(n23814) );
  XNOR U25389 ( .A(n23815), .B(n23814), .Z(n23844) );
  XNOR U25390 ( .A(sreg[1549]), .B(n23844), .Z(n23846) );
  NANDN U25391 ( .A(sreg[1548]), .B(n23807), .Z(n23811) );
  NAND U25392 ( .A(n23809), .B(n23808), .Z(n23810) );
  NAND U25393 ( .A(n23811), .B(n23810), .Z(n23845) );
  XNOR U25394 ( .A(n23846), .B(n23845), .Z(c[1549]) );
  NANDN U25395 ( .A(n23813), .B(n23812), .Z(n23817) );
  NANDN U25396 ( .A(n23815), .B(n23814), .Z(n23816) );
  AND U25397 ( .A(n23817), .B(n23816), .Z(n23852) );
  NANDN U25398 ( .A(n23819), .B(n23818), .Z(n23823) );
  NANDN U25399 ( .A(n23821), .B(n23820), .Z(n23822) );
  AND U25400 ( .A(n23823), .B(n23822), .Z(n23850) );
  NAND U25401 ( .A(n42143), .B(n23824), .Z(n23826) );
  XNOR U25402 ( .A(a[528]), .B(n4147), .Z(n23861) );
  NAND U25403 ( .A(n42144), .B(n23861), .Z(n23825) );
  AND U25404 ( .A(n23826), .B(n23825), .Z(n23876) );
  XOR U25405 ( .A(a[532]), .B(n42012), .Z(n23864) );
  XNOR U25406 ( .A(n23876), .B(n23875), .Z(n23878) );
  XOR U25407 ( .A(a[530]), .B(n42085), .Z(n23868) );
  AND U25408 ( .A(a[526]), .B(b[7]), .Z(n23869) );
  XNOR U25409 ( .A(n23870), .B(n23869), .Z(n23871) );
  AND U25410 ( .A(a[534]), .B(b[0]), .Z(n23829) );
  XNOR U25411 ( .A(n23829), .B(n4071), .Z(n23831) );
  NANDN U25412 ( .A(b[0]), .B(a[533]), .Z(n23830) );
  NAND U25413 ( .A(n23831), .B(n23830), .Z(n23872) );
  XNOR U25414 ( .A(n23871), .B(n23872), .Z(n23877) );
  XOR U25415 ( .A(n23878), .B(n23877), .Z(n23856) );
  NANDN U25416 ( .A(n23833), .B(n23832), .Z(n23837) );
  NANDN U25417 ( .A(n23835), .B(n23834), .Z(n23836) );
  AND U25418 ( .A(n23837), .B(n23836), .Z(n23855) );
  XNOR U25419 ( .A(n23856), .B(n23855), .Z(n23857) );
  NANDN U25420 ( .A(n23839), .B(n23838), .Z(n23843) );
  NAND U25421 ( .A(n23841), .B(n23840), .Z(n23842) );
  NAND U25422 ( .A(n23843), .B(n23842), .Z(n23858) );
  XNOR U25423 ( .A(n23857), .B(n23858), .Z(n23849) );
  XNOR U25424 ( .A(n23850), .B(n23849), .Z(n23851) );
  XNOR U25425 ( .A(n23852), .B(n23851), .Z(n23881) );
  XNOR U25426 ( .A(sreg[1550]), .B(n23881), .Z(n23883) );
  NANDN U25427 ( .A(sreg[1549]), .B(n23844), .Z(n23848) );
  NAND U25428 ( .A(n23846), .B(n23845), .Z(n23847) );
  NAND U25429 ( .A(n23848), .B(n23847), .Z(n23882) );
  XNOR U25430 ( .A(n23883), .B(n23882), .Z(c[1550]) );
  NANDN U25431 ( .A(n23850), .B(n23849), .Z(n23854) );
  NANDN U25432 ( .A(n23852), .B(n23851), .Z(n23853) );
  AND U25433 ( .A(n23854), .B(n23853), .Z(n23889) );
  NANDN U25434 ( .A(n23856), .B(n23855), .Z(n23860) );
  NANDN U25435 ( .A(n23858), .B(n23857), .Z(n23859) );
  AND U25436 ( .A(n23860), .B(n23859), .Z(n23887) );
  NAND U25437 ( .A(n42143), .B(n23861), .Z(n23863) );
  XNOR U25438 ( .A(a[529]), .B(n4147), .Z(n23898) );
  NAND U25439 ( .A(n42144), .B(n23898), .Z(n23862) );
  AND U25440 ( .A(n23863), .B(n23862), .Z(n23913) );
  XOR U25441 ( .A(a[533]), .B(n42012), .Z(n23901) );
  XNOR U25442 ( .A(n23913), .B(n23912), .Z(n23915) );
  AND U25443 ( .A(a[535]), .B(b[0]), .Z(n23865) );
  XNOR U25444 ( .A(n23865), .B(n4071), .Z(n23867) );
  NANDN U25445 ( .A(b[0]), .B(a[534]), .Z(n23866) );
  NAND U25446 ( .A(n23867), .B(n23866), .Z(n23909) );
  XOR U25447 ( .A(a[531]), .B(n42085), .Z(n23905) );
  AND U25448 ( .A(a[527]), .B(b[7]), .Z(n23906) );
  XNOR U25449 ( .A(n23907), .B(n23906), .Z(n23908) );
  XNOR U25450 ( .A(n23909), .B(n23908), .Z(n23914) );
  XOR U25451 ( .A(n23915), .B(n23914), .Z(n23893) );
  NANDN U25452 ( .A(n23870), .B(n23869), .Z(n23874) );
  NANDN U25453 ( .A(n23872), .B(n23871), .Z(n23873) );
  AND U25454 ( .A(n23874), .B(n23873), .Z(n23892) );
  XNOR U25455 ( .A(n23893), .B(n23892), .Z(n23894) );
  NANDN U25456 ( .A(n23876), .B(n23875), .Z(n23880) );
  NAND U25457 ( .A(n23878), .B(n23877), .Z(n23879) );
  NAND U25458 ( .A(n23880), .B(n23879), .Z(n23895) );
  XNOR U25459 ( .A(n23894), .B(n23895), .Z(n23886) );
  XNOR U25460 ( .A(n23887), .B(n23886), .Z(n23888) );
  XNOR U25461 ( .A(n23889), .B(n23888), .Z(n23918) );
  XNOR U25462 ( .A(sreg[1551]), .B(n23918), .Z(n23920) );
  NANDN U25463 ( .A(sreg[1550]), .B(n23881), .Z(n23885) );
  NAND U25464 ( .A(n23883), .B(n23882), .Z(n23884) );
  NAND U25465 ( .A(n23885), .B(n23884), .Z(n23919) );
  XNOR U25466 ( .A(n23920), .B(n23919), .Z(c[1551]) );
  NANDN U25467 ( .A(n23887), .B(n23886), .Z(n23891) );
  NANDN U25468 ( .A(n23889), .B(n23888), .Z(n23890) );
  AND U25469 ( .A(n23891), .B(n23890), .Z(n23926) );
  NANDN U25470 ( .A(n23893), .B(n23892), .Z(n23897) );
  NANDN U25471 ( .A(n23895), .B(n23894), .Z(n23896) );
  AND U25472 ( .A(n23897), .B(n23896), .Z(n23924) );
  NAND U25473 ( .A(n42143), .B(n23898), .Z(n23900) );
  XNOR U25474 ( .A(a[530]), .B(n4147), .Z(n23935) );
  NAND U25475 ( .A(n42144), .B(n23935), .Z(n23899) );
  AND U25476 ( .A(n23900), .B(n23899), .Z(n23950) );
  XOR U25477 ( .A(a[534]), .B(n42012), .Z(n23938) );
  XNOR U25478 ( .A(n23950), .B(n23949), .Z(n23952) );
  AND U25479 ( .A(a[536]), .B(b[0]), .Z(n23902) );
  XNOR U25480 ( .A(n23902), .B(n4071), .Z(n23904) );
  NANDN U25481 ( .A(b[0]), .B(a[535]), .Z(n23903) );
  NAND U25482 ( .A(n23904), .B(n23903), .Z(n23946) );
  XOR U25483 ( .A(a[532]), .B(n42085), .Z(n23939) );
  AND U25484 ( .A(a[528]), .B(b[7]), .Z(n23943) );
  XNOR U25485 ( .A(n23944), .B(n23943), .Z(n23945) );
  XNOR U25486 ( .A(n23946), .B(n23945), .Z(n23951) );
  XOR U25487 ( .A(n23952), .B(n23951), .Z(n23930) );
  NANDN U25488 ( .A(n23907), .B(n23906), .Z(n23911) );
  NANDN U25489 ( .A(n23909), .B(n23908), .Z(n23910) );
  AND U25490 ( .A(n23911), .B(n23910), .Z(n23929) );
  XNOR U25491 ( .A(n23930), .B(n23929), .Z(n23931) );
  NANDN U25492 ( .A(n23913), .B(n23912), .Z(n23917) );
  NAND U25493 ( .A(n23915), .B(n23914), .Z(n23916) );
  NAND U25494 ( .A(n23917), .B(n23916), .Z(n23932) );
  XNOR U25495 ( .A(n23931), .B(n23932), .Z(n23923) );
  XNOR U25496 ( .A(n23924), .B(n23923), .Z(n23925) );
  XNOR U25497 ( .A(n23926), .B(n23925), .Z(n23955) );
  XNOR U25498 ( .A(sreg[1552]), .B(n23955), .Z(n23957) );
  NANDN U25499 ( .A(sreg[1551]), .B(n23918), .Z(n23922) );
  NAND U25500 ( .A(n23920), .B(n23919), .Z(n23921) );
  NAND U25501 ( .A(n23922), .B(n23921), .Z(n23956) );
  XNOR U25502 ( .A(n23957), .B(n23956), .Z(c[1552]) );
  NANDN U25503 ( .A(n23924), .B(n23923), .Z(n23928) );
  NANDN U25504 ( .A(n23926), .B(n23925), .Z(n23927) );
  AND U25505 ( .A(n23928), .B(n23927), .Z(n23963) );
  NANDN U25506 ( .A(n23930), .B(n23929), .Z(n23934) );
  NANDN U25507 ( .A(n23932), .B(n23931), .Z(n23933) );
  AND U25508 ( .A(n23934), .B(n23933), .Z(n23961) );
  NAND U25509 ( .A(n42143), .B(n23935), .Z(n23937) );
  XNOR U25510 ( .A(a[531]), .B(n4147), .Z(n23972) );
  NAND U25511 ( .A(n42144), .B(n23972), .Z(n23936) );
  AND U25512 ( .A(n23937), .B(n23936), .Z(n23987) );
  XOR U25513 ( .A(a[535]), .B(n42012), .Z(n23975) );
  XNOR U25514 ( .A(n23987), .B(n23986), .Z(n23989) );
  XOR U25515 ( .A(a[533]), .B(n42085), .Z(n23979) );
  AND U25516 ( .A(a[529]), .B(b[7]), .Z(n23980) );
  XNOR U25517 ( .A(n23981), .B(n23980), .Z(n23982) );
  AND U25518 ( .A(a[537]), .B(b[0]), .Z(n23940) );
  XNOR U25519 ( .A(n23940), .B(n4071), .Z(n23942) );
  NANDN U25520 ( .A(b[0]), .B(a[536]), .Z(n23941) );
  NAND U25521 ( .A(n23942), .B(n23941), .Z(n23983) );
  XNOR U25522 ( .A(n23982), .B(n23983), .Z(n23988) );
  XOR U25523 ( .A(n23989), .B(n23988), .Z(n23967) );
  NANDN U25524 ( .A(n23944), .B(n23943), .Z(n23948) );
  NANDN U25525 ( .A(n23946), .B(n23945), .Z(n23947) );
  AND U25526 ( .A(n23948), .B(n23947), .Z(n23966) );
  XNOR U25527 ( .A(n23967), .B(n23966), .Z(n23968) );
  NANDN U25528 ( .A(n23950), .B(n23949), .Z(n23954) );
  NAND U25529 ( .A(n23952), .B(n23951), .Z(n23953) );
  NAND U25530 ( .A(n23954), .B(n23953), .Z(n23969) );
  XNOR U25531 ( .A(n23968), .B(n23969), .Z(n23960) );
  XNOR U25532 ( .A(n23961), .B(n23960), .Z(n23962) );
  XNOR U25533 ( .A(n23963), .B(n23962), .Z(n23992) );
  XNOR U25534 ( .A(sreg[1553]), .B(n23992), .Z(n23994) );
  NANDN U25535 ( .A(sreg[1552]), .B(n23955), .Z(n23959) );
  NAND U25536 ( .A(n23957), .B(n23956), .Z(n23958) );
  NAND U25537 ( .A(n23959), .B(n23958), .Z(n23993) );
  XNOR U25538 ( .A(n23994), .B(n23993), .Z(c[1553]) );
  NANDN U25539 ( .A(n23961), .B(n23960), .Z(n23965) );
  NANDN U25540 ( .A(n23963), .B(n23962), .Z(n23964) );
  AND U25541 ( .A(n23965), .B(n23964), .Z(n24000) );
  NANDN U25542 ( .A(n23967), .B(n23966), .Z(n23971) );
  NANDN U25543 ( .A(n23969), .B(n23968), .Z(n23970) );
  AND U25544 ( .A(n23971), .B(n23970), .Z(n23998) );
  NAND U25545 ( .A(n42143), .B(n23972), .Z(n23974) );
  XNOR U25546 ( .A(a[532]), .B(n4147), .Z(n24009) );
  NAND U25547 ( .A(n42144), .B(n24009), .Z(n23973) );
  AND U25548 ( .A(n23974), .B(n23973), .Z(n24024) );
  XOR U25549 ( .A(a[536]), .B(n42012), .Z(n24012) );
  XNOR U25550 ( .A(n24024), .B(n24023), .Z(n24026) );
  AND U25551 ( .A(a[538]), .B(b[0]), .Z(n23976) );
  XNOR U25552 ( .A(n23976), .B(n4071), .Z(n23978) );
  NANDN U25553 ( .A(b[0]), .B(a[537]), .Z(n23977) );
  NAND U25554 ( .A(n23978), .B(n23977), .Z(n24020) );
  XOR U25555 ( .A(a[534]), .B(n42085), .Z(n24016) );
  AND U25556 ( .A(a[530]), .B(b[7]), .Z(n24017) );
  XNOR U25557 ( .A(n24018), .B(n24017), .Z(n24019) );
  XNOR U25558 ( .A(n24020), .B(n24019), .Z(n24025) );
  XOR U25559 ( .A(n24026), .B(n24025), .Z(n24004) );
  NANDN U25560 ( .A(n23981), .B(n23980), .Z(n23985) );
  NANDN U25561 ( .A(n23983), .B(n23982), .Z(n23984) );
  AND U25562 ( .A(n23985), .B(n23984), .Z(n24003) );
  XNOR U25563 ( .A(n24004), .B(n24003), .Z(n24005) );
  NANDN U25564 ( .A(n23987), .B(n23986), .Z(n23991) );
  NAND U25565 ( .A(n23989), .B(n23988), .Z(n23990) );
  NAND U25566 ( .A(n23991), .B(n23990), .Z(n24006) );
  XNOR U25567 ( .A(n24005), .B(n24006), .Z(n23997) );
  XNOR U25568 ( .A(n23998), .B(n23997), .Z(n23999) );
  XNOR U25569 ( .A(n24000), .B(n23999), .Z(n24029) );
  XNOR U25570 ( .A(sreg[1554]), .B(n24029), .Z(n24031) );
  NANDN U25571 ( .A(sreg[1553]), .B(n23992), .Z(n23996) );
  NAND U25572 ( .A(n23994), .B(n23993), .Z(n23995) );
  NAND U25573 ( .A(n23996), .B(n23995), .Z(n24030) );
  XNOR U25574 ( .A(n24031), .B(n24030), .Z(c[1554]) );
  NANDN U25575 ( .A(n23998), .B(n23997), .Z(n24002) );
  NANDN U25576 ( .A(n24000), .B(n23999), .Z(n24001) );
  AND U25577 ( .A(n24002), .B(n24001), .Z(n24037) );
  NANDN U25578 ( .A(n24004), .B(n24003), .Z(n24008) );
  NANDN U25579 ( .A(n24006), .B(n24005), .Z(n24007) );
  AND U25580 ( .A(n24008), .B(n24007), .Z(n24035) );
  NAND U25581 ( .A(n42143), .B(n24009), .Z(n24011) );
  XNOR U25582 ( .A(a[533]), .B(n4148), .Z(n24046) );
  NAND U25583 ( .A(n42144), .B(n24046), .Z(n24010) );
  AND U25584 ( .A(n24011), .B(n24010), .Z(n24061) );
  XOR U25585 ( .A(a[537]), .B(n42012), .Z(n24049) );
  XNOR U25586 ( .A(n24061), .B(n24060), .Z(n24063) );
  AND U25587 ( .A(a[539]), .B(b[0]), .Z(n24013) );
  XNOR U25588 ( .A(n24013), .B(n4071), .Z(n24015) );
  NANDN U25589 ( .A(b[0]), .B(a[538]), .Z(n24014) );
  NAND U25590 ( .A(n24015), .B(n24014), .Z(n24057) );
  XOR U25591 ( .A(a[535]), .B(n42085), .Z(n24053) );
  AND U25592 ( .A(a[531]), .B(b[7]), .Z(n24054) );
  XNOR U25593 ( .A(n24055), .B(n24054), .Z(n24056) );
  XNOR U25594 ( .A(n24057), .B(n24056), .Z(n24062) );
  XOR U25595 ( .A(n24063), .B(n24062), .Z(n24041) );
  NANDN U25596 ( .A(n24018), .B(n24017), .Z(n24022) );
  NANDN U25597 ( .A(n24020), .B(n24019), .Z(n24021) );
  AND U25598 ( .A(n24022), .B(n24021), .Z(n24040) );
  XNOR U25599 ( .A(n24041), .B(n24040), .Z(n24042) );
  NANDN U25600 ( .A(n24024), .B(n24023), .Z(n24028) );
  NAND U25601 ( .A(n24026), .B(n24025), .Z(n24027) );
  NAND U25602 ( .A(n24028), .B(n24027), .Z(n24043) );
  XNOR U25603 ( .A(n24042), .B(n24043), .Z(n24034) );
  XNOR U25604 ( .A(n24035), .B(n24034), .Z(n24036) );
  XNOR U25605 ( .A(n24037), .B(n24036), .Z(n24066) );
  XNOR U25606 ( .A(sreg[1555]), .B(n24066), .Z(n24068) );
  NANDN U25607 ( .A(sreg[1554]), .B(n24029), .Z(n24033) );
  NAND U25608 ( .A(n24031), .B(n24030), .Z(n24032) );
  NAND U25609 ( .A(n24033), .B(n24032), .Z(n24067) );
  XNOR U25610 ( .A(n24068), .B(n24067), .Z(c[1555]) );
  NANDN U25611 ( .A(n24035), .B(n24034), .Z(n24039) );
  NANDN U25612 ( .A(n24037), .B(n24036), .Z(n24038) );
  AND U25613 ( .A(n24039), .B(n24038), .Z(n24074) );
  NANDN U25614 ( .A(n24041), .B(n24040), .Z(n24045) );
  NANDN U25615 ( .A(n24043), .B(n24042), .Z(n24044) );
  AND U25616 ( .A(n24045), .B(n24044), .Z(n24072) );
  NAND U25617 ( .A(n42143), .B(n24046), .Z(n24048) );
  XNOR U25618 ( .A(a[534]), .B(n4148), .Z(n24083) );
  NAND U25619 ( .A(n42144), .B(n24083), .Z(n24047) );
  AND U25620 ( .A(n24048), .B(n24047), .Z(n24098) );
  XOR U25621 ( .A(a[538]), .B(n42012), .Z(n24086) );
  XNOR U25622 ( .A(n24098), .B(n24097), .Z(n24100) );
  AND U25623 ( .A(a[540]), .B(b[0]), .Z(n24050) );
  XNOR U25624 ( .A(n24050), .B(n4071), .Z(n24052) );
  NANDN U25625 ( .A(b[0]), .B(a[539]), .Z(n24051) );
  NAND U25626 ( .A(n24052), .B(n24051), .Z(n24094) );
  XOR U25627 ( .A(a[536]), .B(n42085), .Z(n24087) );
  AND U25628 ( .A(a[532]), .B(b[7]), .Z(n24091) );
  XNOR U25629 ( .A(n24092), .B(n24091), .Z(n24093) );
  XNOR U25630 ( .A(n24094), .B(n24093), .Z(n24099) );
  XOR U25631 ( .A(n24100), .B(n24099), .Z(n24078) );
  NANDN U25632 ( .A(n24055), .B(n24054), .Z(n24059) );
  NANDN U25633 ( .A(n24057), .B(n24056), .Z(n24058) );
  AND U25634 ( .A(n24059), .B(n24058), .Z(n24077) );
  XNOR U25635 ( .A(n24078), .B(n24077), .Z(n24079) );
  NANDN U25636 ( .A(n24061), .B(n24060), .Z(n24065) );
  NAND U25637 ( .A(n24063), .B(n24062), .Z(n24064) );
  NAND U25638 ( .A(n24065), .B(n24064), .Z(n24080) );
  XNOR U25639 ( .A(n24079), .B(n24080), .Z(n24071) );
  XNOR U25640 ( .A(n24072), .B(n24071), .Z(n24073) );
  XNOR U25641 ( .A(n24074), .B(n24073), .Z(n24103) );
  XNOR U25642 ( .A(sreg[1556]), .B(n24103), .Z(n24105) );
  NANDN U25643 ( .A(sreg[1555]), .B(n24066), .Z(n24070) );
  NAND U25644 ( .A(n24068), .B(n24067), .Z(n24069) );
  NAND U25645 ( .A(n24070), .B(n24069), .Z(n24104) );
  XNOR U25646 ( .A(n24105), .B(n24104), .Z(c[1556]) );
  NANDN U25647 ( .A(n24072), .B(n24071), .Z(n24076) );
  NANDN U25648 ( .A(n24074), .B(n24073), .Z(n24075) );
  AND U25649 ( .A(n24076), .B(n24075), .Z(n24111) );
  NANDN U25650 ( .A(n24078), .B(n24077), .Z(n24082) );
  NANDN U25651 ( .A(n24080), .B(n24079), .Z(n24081) );
  AND U25652 ( .A(n24082), .B(n24081), .Z(n24109) );
  NAND U25653 ( .A(n42143), .B(n24083), .Z(n24085) );
  XNOR U25654 ( .A(a[535]), .B(n4148), .Z(n24120) );
  NAND U25655 ( .A(n42144), .B(n24120), .Z(n24084) );
  AND U25656 ( .A(n24085), .B(n24084), .Z(n24135) );
  XOR U25657 ( .A(a[539]), .B(n42012), .Z(n24123) );
  XNOR U25658 ( .A(n24135), .B(n24134), .Z(n24137) );
  XOR U25659 ( .A(a[537]), .B(n42085), .Z(n24124) );
  AND U25660 ( .A(a[533]), .B(b[7]), .Z(n24128) );
  XNOR U25661 ( .A(n24129), .B(n24128), .Z(n24130) );
  AND U25662 ( .A(a[541]), .B(b[0]), .Z(n24088) );
  XNOR U25663 ( .A(n24088), .B(n4071), .Z(n24090) );
  NANDN U25664 ( .A(b[0]), .B(a[540]), .Z(n24089) );
  NAND U25665 ( .A(n24090), .B(n24089), .Z(n24131) );
  XNOR U25666 ( .A(n24130), .B(n24131), .Z(n24136) );
  XOR U25667 ( .A(n24137), .B(n24136), .Z(n24115) );
  NANDN U25668 ( .A(n24092), .B(n24091), .Z(n24096) );
  NANDN U25669 ( .A(n24094), .B(n24093), .Z(n24095) );
  AND U25670 ( .A(n24096), .B(n24095), .Z(n24114) );
  XNOR U25671 ( .A(n24115), .B(n24114), .Z(n24116) );
  NANDN U25672 ( .A(n24098), .B(n24097), .Z(n24102) );
  NAND U25673 ( .A(n24100), .B(n24099), .Z(n24101) );
  NAND U25674 ( .A(n24102), .B(n24101), .Z(n24117) );
  XNOR U25675 ( .A(n24116), .B(n24117), .Z(n24108) );
  XNOR U25676 ( .A(n24109), .B(n24108), .Z(n24110) );
  XNOR U25677 ( .A(n24111), .B(n24110), .Z(n24140) );
  XNOR U25678 ( .A(sreg[1557]), .B(n24140), .Z(n24142) );
  NANDN U25679 ( .A(sreg[1556]), .B(n24103), .Z(n24107) );
  NAND U25680 ( .A(n24105), .B(n24104), .Z(n24106) );
  NAND U25681 ( .A(n24107), .B(n24106), .Z(n24141) );
  XNOR U25682 ( .A(n24142), .B(n24141), .Z(c[1557]) );
  NANDN U25683 ( .A(n24109), .B(n24108), .Z(n24113) );
  NANDN U25684 ( .A(n24111), .B(n24110), .Z(n24112) );
  AND U25685 ( .A(n24113), .B(n24112), .Z(n24148) );
  NANDN U25686 ( .A(n24115), .B(n24114), .Z(n24119) );
  NANDN U25687 ( .A(n24117), .B(n24116), .Z(n24118) );
  AND U25688 ( .A(n24119), .B(n24118), .Z(n24146) );
  NAND U25689 ( .A(n42143), .B(n24120), .Z(n24122) );
  XNOR U25690 ( .A(a[536]), .B(n4148), .Z(n24157) );
  NAND U25691 ( .A(n42144), .B(n24157), .Z(n24121) );
  AND U25692 ( .A(n24122), .B(n24121), .Z(n24172) );
  XOR U25693 ( .A(a[540]), .B(n42012), .Z(n24160) );
  XNOR U25694 ( .A(n24172), .B(n24171), .Z(n24174) );
  XOR U25695 ( .A(a[538]), .B(n42085), .Z(n24164) );
  AND U25696 ( .A(a[534]), .B(b[7]), .Z(n24165) );
  XNOR U25697 ( .A(n24166), .B(n24165), .Z(n24167) );
  AND U25698 ( .A(a[542]), .B(b[0]), .Z(n24125) );
  XNOR U25699 ( .A(n24125), .B(n4071), .Z(n24127) );
  NANDN U25700 ( .A(b[0]), .B(a[541]), .Z(n24126) );
  NAND U25701 ( .A(n24127), .B(n24126), .Z(n24168) );
  XNOR U25702 ( .A(n24167), .B(n24168), .Z(n24173) );
  XOR U25703 ( .A(n24174), .B(n24173), .Z(n24152) );
  NANDN U25704 ( .A(n24129), .B(n24128), .Z(n24133) );
  NANDN U25705 ( .A(n24131), .B(n24130), .Z(n24132) );
  AND U25706 ( .A(n24133), .B(n24132), .Z(n24151) );
  XNOR U25707 ( .A(n24152), .B(n24151), .Z(n24153) );
  NANDN U25708 ( .A(n24135), .B(n24134), .Z(n24139) );
  NAND U25709 ( .A(n24137), .B(n24136), .Z(n24138) );
  NAND U25710 ( .A(n24139), .B(n24138), .Z(n24154) );
  XNOR U25711 ( .A(n24153), .B(n24154), .Z(n24145) );
  XNOR U25712 ( .A(n24146), .B(n24145), .Z(n24147) );
  XNOR U25713 ( .A(n24148), .B(n24147), .Z(n24177) );
  XNOR U25714 ( .A(sreg[1558]), .B(n24177), .Z(n24179) );
  NANDN U25715 ( .A(sreg[1557]), .B(n24140), .Z(n24144) );
  NAND U25716 ( .A(n24142), .B(n24141), .Z(n24143) );
  NAND U25717 ( .A(n24144), .B(n24143), .Z(n24178) );
  XNOR U25718 ( .A(n24179), .B(n24178), .Z(c[1558]) );
  NANDN U25719 ( .A(n24146), .B(n24145), .Z(n24150) );
  NANDN U25720 ( .A(n24148), .B(n24147), .Z(n24149) );
  AND U25721 ( .A(n24150), .B(n24149), .Z(n24185) );
  NANDN U25722 ( .A(n24152), .B(n24151), .Z(n24156) );
  NANDN U25723 ( .A(n24154), .B(n24153), .Z(n24155) );
  AND U25724 ( .A(n24156), .B(n24155), .Z(n24183) );
  NAND U25725 ( .A(n42143), .B(n24157), .Z(n24159) );
  XNOR U25726 ( .A(a[537]), .B(n4148), .Z(n24194) );
  NAND U25727 ( .A(n42144), .B(n24194), .Z(n24158) );
  AND U25728 ( .A(n24159), .B(n24158), .Z(n24209) );
  XOR U25729 ( .A(a[541]), .B(n42012), .Z(n24197) );
  XNOR U25730 ( .A(n24209), .B(n24208), .Z(n24211) );
  AND U25731 ( .A(a[543]), .B(b[0]), .Z(n24161) );
  XNOR U25732 ( .A(n24161), .B(n4071), .Z(n24163) );
  NANDN U25733 ( .A(b[0]), .B(a[542]), .Z(n24162) );
  NAND U25734 ( .A(n24163), .B(n24162), .Z(n24205) );
  XOR U25735 ( .A(a[539]), .B(n42085), .Z(n24201) );
  AND U25736 ( .A(a[535]), .B(b[7]), .Z(n24202) );
  XNOR U25737 ( .A(n24203), .B(n24202), .Z(n24204) );
  XNOR U25738 ( .A(n24205), .B(n24204), .Z(n24210) );
  XOR U25739 ( .A(n24211), .B(n24210), .Z(n24189) );
  NANDN U25740 ( .A(n24166), .B(n24165), .Z(n24170) );
  NANDN U25741 ( .A(n24168), .B(n24167), .Z(n24169) );
  AND U25742 ( .A(n24170), .B(n24169), .Z(n24188) );
  XNOR U25743 ( .A(n24189), .B(n24188), .Z(n24190) );
  NANDN U25744 ( .A(n24172), .B(n24171), .Z(n24176) );
  NAND U25745 ( .A(n24174), .B(n24173), .Z(n24175) );
  NAND U25746 ( .A(n24176), .B(n24175), .Z(n24191) );
  XNOR U25747 ( .A(n24190), .B(n24191), .Z(n24182) );
  XNOR U25748 ( .A(n24183), .B(n24182), .Z(n24184) );
  XNOR U25749 ( .A(n24185), .B(n24184), .Z(n24214) );
  XNOR U25750 ( .A(sreg[1559]), .B(n24214), .Z(n24216) );
  NANDN U25751 ( .A(sreg[1558]), .B(n24177), .Z(n24181) );
  NAND U25752 ( .A(n24179), .B(n24178), .Z(n24180) );
  NAND U25753 ( .A(n24181), .B(n24180), .Z(n24215) );
  XNOR U25754 ( .A(n24216), .B(n24215), .Z(c[1559]) );
  NANDN U25755 ( .A(n24183), .B(n24182), .Z(n24187) );
  NANDN U25756 ( .A(n24185), .B(n24184), .Z(n24186) );
  AND U25757 ( .A(n24187), .B(n24186), .Z(n24222) );
  NANDN U25758 ( .A(n24189), .B(n24188), .Z(n24193) );
  NANDN U25759 ( .A(n24191), .B(n24190), .Z(n24192) );
  AND U25760 ( .A(n24193), .B(n24192), .Z(n24220) );
  NAND U25761 ( .A(n42143), .B(n24194), .Z(n24196) );
  XNOR U25762 ( .A(a[538]), .B(n4148), .Z(n24231) );
  NAND U25763 ( .A(n42144), .B(n24231), .Z(n24195) );
  AND U25764 ( .A(n24196), .B(n24195), .Z(n24246) );
  XOR U25765 ( .A(a[542]), .B(n42012), .Z(n24234) );
  XNOR U25766 ( .A(n24246), .B(n24245), .Z(n24248) );
  AND U25767 ( .A(a[544]), .B(b[0]), .Z(n24198) );
  XNOR U25768 ( .A(n24198), .B(n4071), .Z(n24200) );
  NANDN U25769 ( .A(b[0]), .B(a[543]), .Z(n24199) );
  NAND U25770 ( .A(n24200), .B(n24199), .Z(n24242) );
  XOR U25771 ( .A(a[540]), .B(n42085), .Z(n24238) );
  AND U25772 ( .A(a[536]), .B(b[7]), .Z(n24239) );
  XNOR U25773 ( .A(n24240), .B(n24239), .Z(n24241) );
  XNOR U25774 ( .A(n24242), .B(n24241), .Z(n24247) );
  XOR U25775 ( .A(n24248), .B(n24247), .Z(n24226) );
  NANDN U25776 ( .A(n24203), .B(n24202), .Z(n24207) );
  NANDN U25777 ( .A(n24205), .B(n24204), .Z(n24206) );
  AND U25778 ( .A(n24207), .B(n24206), .Z(n24225) );
  XNOR U25779 ( .A(n24226), .B(n24225), .Z(n24227) );
  NANDN U25780 ( .A(n24209), .B(n24208), .Z(n24213) );
  NAND U25781 ( .A(n24211), .B(n24210), .Z(n24212) );
  NAND U25782 ( .A(n24213), .B(n24212), .Z(n24228) );
  XNOR U25783 ( .A(n24227), .B(n24228), .Z(n24219) );
  XNOR U25784 ( .A(n24220), .B(n24219), .Z(n24221) );
  XNOR U25785 ( .A(n24222), .B(n24221), .Z(n24251) );
  XNOR U25786 ( .A(sreg[1560]), .B(n24251), .Z(n24253) );
  NANDN U25787 ( .A(sreg[1559]), .B(n24214), .Z(n24218) );
  NAND U25788 ( .A(n24216), .B(n24215), .Z(n24217) );
  NAND U25789 ( .A(n24218), .B(n24217), .Z(n24252) );
  XNOR U25790 ( .A(n24253), .B(n24252), .Z(c[1560]) );
  NANDN U25791 ( .A(n24220), .B(n24219), .Z(n24224) );
  NANDN U25792 ( .A(n24222), .B(n24221), .Z(n24223) );
  AND U25793 ( .A(n24224), .B(n24223), .Z(n24259) );
  NANDN U25794 ( .A(n24226), .B(n24225), .Z(n24230) );
  NANDN U25795 ( .A(n24228), .B(n24227), .Z(n24229) );
  AND U25796 ( .A(n24230), .B(n24229), .Z(n24257) );
  NAND U25797 ( .A(n42143), .B(n24231), .Z(n24233) );
  XNOR U25798 ( .A(a[539]), .B(n4148), .Z(n24268) );
  NAND U25799 ( .A(n42144), .B(n24268), .Z(n24232) );
  AND U25800 ( .A(n24233), .B(n24232), .Z(n24283) );
  XOR U25801 ( .A(a[543]), .B(n42012), .Z(n24271) );
  XNOR U25802 ( .A(n24283), .B(n24282), .Z(n24285) );
  AND U25803 ( .A(a[545]), .B(b[0]), .Z(n24235) );
  XNOR U25804 ( .A(n24235), .B(n4071), .Z(n24237) );
  NANDN U25805 ( .A(b[0]), .B(a[544]), .Z(n24236) );
  NAND U25806 ( .A(n24237), .B(n24236), .Z(n24279) );
  XOR U25807 ( .A(a[541]), .B(n42085), .Z(n24275) );
  AND U25808 ( .A(a[537]), .B(b[7]), .Z(n24276) );
  XNOR U25809 ( .A(n24277), .B(n24276), .Z(n24278) );
  XNOR U25810 ( .A(n24279), .B(n24278), .Z(n24284) );
  XOR U25811 ( .A(n24285), .B(n24284), .Z(n24263) );
  NANDN U25812 ( .A(n24240), .B(n24239), .Z(n24244) );
  NANDN U25813 ( .A(n24242), .B(n24241), .Z(n24243) );
  AND U25814 ( .A(n24244), .B(n24243), .Z(n24262) );
  XNOR U25815 ( .A(n24263), .B(n24262), .Z(n24264) );
  NANDN U25816 ( .A(n24246), .B(n24245), .Z(n24250) );
  NAND U25817 ( .A(n24248), .B(n24247), .Z(n24249) );
  NAND U25818 ( .A(n24250), .B(n24249), .Z(n24265) );
  XNOR U25819 ( .A(n24264), .B(n24265), .Z(n24256) );
  XNOR U25820 ( .A(n24257), .B(n24256), .Z(n24258) );
  XNOR U25821 ( .A(n24259), .B(n24258), .Z(n24288) );
  XNOR U25822 ( .A(sreg[1561]), .B(n24288), .Z(n24290) );
  NANDN U25823 ( .A(sreg[1560]), .B(n24251), .Z(n24255) );
  NAND U25824 ( .A(n24253), .B(n24252), .Z(n24254) );
  NAND U25825 ( .A(n24255), .B(n24254), .Z(n24289) );
  XNOR U25826 ( .A(n24290), .B(n24289), .Z(c[1561]) );
  NANDN U25827 ( .A(n24257), .B(n24256), .Z(n24261) );
  NANDN U25828 ( .A(n24259), .B(n24258), .Z(n24260) );
  AND U25829 ( .A(n24261), .B(n24260), .Z(n24296) );
  NANDN U25830 ( .A(n24263), .B(n24262), .Z(n24267) );
  NANDN U25831 ( .A(n24265), .B(n24264), .Z(n24266) );
  AND U25832 ( .A(n24267), .B(n24266), .Z(n24294) );
  NAND U25833 ( .A(n42143), .B(n24268), .Z(n24270) );
  XNOR U25834 ( .A(a[540]), .B(n4149), .Z(n24305) );
  NAND U25835 ( .A(n42144), .B(n24305), .Z(n24269) );
  AND U25836 ( .A(n24270), .B(n24269), .Z(n24320) );
  XOR U25837 ( .A(a[544]), .B(n42012), .Z(n24308) );
  XNOR U25838 ( .A(n24320), .B(n24319), .Z(n24322) );
  AND U25839 ( .A(a[546]), .B(b[0]), .Z(n24272) );
  XNOR U25840 ( .A(n24272), .B(n4071), .Z(n24274) );
  NANDN U25841 ( .A(b[0]), .B(a[545]), .Z(n24273) );
  NAND U25842 ( .A(n24274), .B(n24273), .Z(n24316) );
  XOR U25843 ( .A(a[542]), .B(n42085), .Z(n24312) );
  AND U25844 ( .A(a[538]), .B(b[7]), .Z(n24313) );
  XNOR U25845 ( .A(n24314), .B(n24313), .Z(n24315) );
  XNOR U25846 ( .A(n24316), .B(n24315), .Z(n24321) );
  XOR U25847 ( .A(n24322), .B(n24321), .Z(n24300) );
  NANDN U25848 ( .A(n24277), .B(n24276), .Z(n24281) );
  NANDN U25849 ( .A(n24279), .B(n24278), .Z(n24280) );
  AND U25850 ( .A(n24281), .B(n24280), .Z(n24299) );
  XNOR U25851 ( .A(n24300), .B(n24299), .Z(n24301) );
  NANDN U25852 ( .A(n24283), .B(n24282), .Z(n24287) );
  NAND U25853 ( .A(n24285), .B(n24284), .Z(n24286) );
  NAND U25854 ( .A(n24287), .B(n24286), .Z(n24302) );
  XNOR U25855 ( .A(n24301), .B(n24302), .Z(n24293) );
  XNOR U25856 ( .A(n24294), .B(n24293), .Z(n24295) );
  XNOR U25857 ( .A(n24296), .B(n24295), .Z(n24325) );
  XNOR U25858 ( .A(sreg[1562]), .B(n24325), .Z(n24327) );
  NANDN U25859 ( .A(sreg[1561]), .B(n24288), .Z(n24292) );
  NAND U25860 ( .A(n24290), .B(n24289), .Z(n24291) );
  NAND U25861 ( .A(n24292), .B(n24291), .Z(n24326) );
  XNOR U25862 ( .A(n24327), .B(n24326), .Z(c[1562]) );
  NANDN U25863 ( .A(n24294), .B(n24293), .Z(n24298) );
  NANDN U25864 ( .A(n24296), .B(n24295), .Z(n24297) );
  AND U25865 ( .A(n24298), .B(n24297), .Z(n24333) );
  NANDN U25866 ( .A(n24300), .B(n24299), .Z(n24304) );
  NANDN U25867 ( .A(n24302), .B(n24301), .Z(n24303) );
  AND U25868 ( .A(n24304), .B(n24303), .Z(n24331) );
  NAND U25869 ( .A(n42143), .B(n24305), .Z(n24307) );
  XNOR U25870 ( .A(a[541]), .B(n4149), .Z(n24342) );
  NAND U25871 ( .A(n42144), .B(n24342), .Z(n24306) );
  AND U25872 ( .A(n24307), .B(n24306), .Z(n24357) );
  XOR U25873 ( .A(a[545]), .B(n42012), .Z(n24345) );
  XNOR U25874 ( .A(n24357), .B(n24356), .Z(n24359) );
  AND U25875 ( .A(a[547]), .B(b[0]), .Z(n24309) );
  XNOR U25876 ( .A(n24309), .B(n4071), .Z(n24311) );
  NANDN U25877 ( .A(b[0]), .B(a[546]), .Z(n24310) );
  NAND U25878 ( .A(n24311), .B(n24310), .Z(n24353) );
  XOR U25879 ( .A(a[543]), .B(n42085), .Z(n24349) );
  AND U25880 ( .A(a[539]), .B(b[7]), .Z(n24350) );
  XNOR U25881 ( .A(n24351), .B(n24350), .Z(n24352) );
  XNOR U25882 ( .A(n24353), .B(n24352), .Z(n24358) );
  XOR U25883 ( .A(n24359), .B(n24358), .Z(n24337) );
  NANDN U25884 ( .A(n24314), .B(n24313), .Z(n24318) );
  NANDN U25885 ( .A(n24316), .B(n24315), .Z(n24317) );
  AND U25886 ( .A(n24318), .B(n24317), .Z(n24336) );
  XNOR U25887 ( .A(n24337), .B(n24336), .Z(n24338) );
  NANDN U25888 ( .A(n24320), .B(n24319), .Z(n24324) );
  NAND U25889 ( .A(n24322), .B(n24321), .Z(n24323) );
  NAND U25890 ( .A(n24324), .B(n24323), .Z(n24339) );
  XNOR U25891 ( .A(n24338), .B(n24339), .Z(n24330) );
  XNOR U25892 ( .A(n24331), .B(n24330), .Z(n24332) );
  XNOR U25893 ( .A(n24333), .B(n24332), .Z(n24362) );
  XNOR U25894 ( .A(sreg[1563]), .B(n24362), .Z(n24364) );
  NANDN U25895 ( .A(sreg[1562]), .B(n24325), .Z(n24329) );
  NAND U25896 ( .A(n24327), .B(n24326), .Z(n24328) );
  NAND U25897 ( .A(n24329), .B(n24328), .Z(n24363) );
  XNOR U25898 ( .A(n24364), .B(n24363), .Z(c[1563]) );
  NANDN U25899 ( .A(n24331), .B(n24330), .Z(n24335) );
  NANDN U25900 ( .A(n24333), .B(n24332), .Z(n24334) );
  AND U25901 ( .A(n24335), .B(n24334), .Z(n24370) );
  NANDN U25902 ( .A(n24337), .B(n24336), .Z(n24341) );
  NANDN U25903 ( .A(n24339), .B(n24338), .Z(n24340) );
  AND U25904 ( .A(n24341), .B(n24340), .Z(n24368) );
  NAND U25905 ( .A(n42143), .B(n24342), .Z(n24344) );
  XNOR U25906 ( .A(a[542]), .B(n4149), .Z(n24379) );
  NAND U25907 ( .A(n42144), .B(n24379), .Z(n24343) );
  AND U25908 ( .A(n24344), .B(n24343), .Z(n24394) );
  XOR U25909 ( .A(a[546]), .B(n42012), .Z(n24382) );
  XNOR U25910 ( .A(n24394), .B(n24393), .Z(n24396) );
  AND U25911 ( .A(a[548]), .B(b[0]), .Z(n24346) );
  XNOR U25912 ( .A(n24346), .B(n4071), .Z(n24348) );
  NANDN U25913 ( .A(b[0]), .B(a[547]), .Z(n24347) );
  NAND U25914 ( .A(n24348), .B(n24347), .Z(n24390) );
  XOR U25915 ( .A(a[544]), .B(n42085), .Z(n24386) );
  AND U25916 ( .A(a[540]), .B(b[7]), .Z(n24387) );
  XNOR U25917 ( .A(n24388), .B(n24387), .Z(n24389) );
  XNOR U25918 ( .A(n24390), .B(n24389), .Z(n24395) );
  XOR U25919 ( .A(n24396), .B(n24395), .Z(n24374) );
  NANDN U25920 ( .A(n24351), .B(n24350), .Z(n24355) );
  NANDN U25921 ( .A(n24353), .B(n24352), .Z(n24354) );
  AND U25922 ( .A(n24355), .B(n24354), .Z(n24373) );
  XNOR U25923 ( .A(n24374), .B(n24373), .Z(n24375) );
  NANDN U25924 ( .A(n24357), .B(n24356), .Z(n24361) );
  NAND U25925 ( .A(n24359), .B(n24358), .Z(n24360) );
  NAND U25926 ( .A(n24361), .B(n24360), .Z(n24376) );
  XNOR U25927 ( .A(n24375), .B(n24376), .Z(n24367) );
  XNOR U25928 ( .A(n24368), .B(n24367), .Z(n24369) );
  XNOR U25929 ( .A(n24370), .B(n24369), .Z(n24399) );
  XNOR U25930 ( .A(sreg[1564]), .B(n24399), .Z(n24401) );
  NANDN U25931 ( .A(sreg[1563]), .B(n24362), .Z(n24366) );
  NAND U25932 ( .A(n24364), .B(n24363), .Z(n24365) );
  NAND U25933 ( .A(n24366), .B(n24365), .Z(n24400) );
  XNOR U25934 ( .A(n24401), .B(n24400), .Z(c[1564]) );
  NANDN U25935 ( .A(n24368), .B(n24367), .Z(n24372) );
  NANDN U25936 ( .A(n24370), .B(n24369), .Z(n24371) );
  AND U25937 ( .A(n24372), .B(n24371), .Z(n24407) );
  NANDN U25938 ( .A(n24374), .B(n24373), .Z(n24378) );
  NANDN U25939 ( .A(n24376), .B(n24375), .Z(n24377) );
  AND U25940 ( .A(n24378), .B(n24377), .Z(n24405) );
  NAND U25941 ( .A(n42143), .B(n24379), .Z(n24381) );
  XNOR U25942 ( .A(a[543]), .B(n4149), .Z(n24416) );
  NAND U25943 ( .A(n42144), .B(n24416), .Z(n24380) );
  AND U25944 ( .A(n24381), .B(n24380), .Z(n24431) );
  XOR U25945 ( .A(a[547]), .B(n42012), .Z(n24419) );
  XNOR U25946 ( .A(n24431), .B(n24430), .Z(n24433) );
  AND U25947 ( .A(a[549]), .B(b[0]), .Z(n24383) );
  XNOR U25948 ( .A(n24383), .B(n4071), .Z(n24385) );
  NANDN U25949 ( .A(b[0]), .B(a[548]), .Z(n24384) );
  NAND U25950 ( .A(n24385), .B(n24384), .Z(n24427) );
  XOR U25951 ( .A(a[545]), .B(n42085), .Z(n24423) );
  AND U25952 ( .A(a[541]), .B(b[7]), .Z(n24424) );
  XNOR U25953 ( .A(n24425), .B(n24424), .Z(n24426) );
  XNOR U25954 ( .A(n24427), .B(n24426), .Z(n24432) );
  XOR U25955 ( .A(n24433), .B(n24432), .Z(n24411) );
  NANDN U25956 ( .A(n24388), .B(n24387), .Z(n24392) );
  NANDN U25957 ( .A(n24390), .B(n24389), .Z(n24391) );
  AND U25958 ( .A(n24392), .B(n24391), .Z(n24410) );
  XNOR U25959 ( .A(n24411), .B(n24410), .Z(n24412) );
  NANDN U25960 ( .A(n24394), .B(n24393), .Z(n24398) );
  NAND U25961 ( .A(n24396), .B(n24395), .Z(n24397) );
  NAND U25962 ( .A(n24398), .B(n24397), .Z(n24413) );
  XNOR U25963 ( .A(n24412), .B(n24413), .Z(n24404) );
  XNOR U25964 ( .A(n24405), .B(n24404), .Z(n24406) );
  XNOR U25965 ( .A(n24407), .B(n24406), .Z(n24436) );
  XNOR U25966 ( .A(sreg[1565]), .B(n24436), .Z(n24438) );
  NANDN U25967 ( .A(sreg[1564]), .B(n24399), .Z(n24403) );
  NAND U25968 ( .A(n24401), .B(n24400), .Z(n24402) );
  NAND U25969 ( .A(n24403), .B(n24402), .Z(n24437) );
  XNOR U25970 ( .A(n24438), .B(n24437), .Z(c[1565]) );
  NANDN U25971 ( .A(n24405), .B(n24404), .Z(n24409) );
  NANDN U25972 ( .A(n24407), .B(n24406), .Z(n24408) );
  AND U25973 ( .A(n24409), .B(n24408), .Z(n24444) );
  NANDN U25974 ( .A(n24411), .B(n24410), .Z(n24415) );
  NANDN U25975 ( .A(n24413), .B(n24412), .Z(n24414) );
  AND U25976 ( .A(n24415), .B(n24414), .Z(n24442) );
  NAND U25977 ( .A(n42143), .B(n24416), .Z(n24418) );
  XNOR U25978 ( .A(a[544]), .B(n4149), .Z(n24453) );
  NAND U25979 ( .A(n42144), .B(n24453), .Z(n24417) );
  AND U25980 ( .A(n24418), .B(n24417), .Z(n24468) );
  XOR U25981 ( .A(a[548]), .B(n42012), .Z(n24456) );
  XNOR U25982 ( .A(n24468), .B(n24467), .Z(n24470) );
  AND U25983 ( .A(a[550]), .B(b[0]), .Z(n24420) );
  XNOR U25984 ( .A(n24420), .B(n4071), .Z(n24422) );
  NANDN U25985 ( .A(b[0]), .B(a[549]), .Z(n24421) );
  NAND U25986 ( .A(n24422), .B(n24421), .Z(n24464) );
  XOR U25987 ( .A(a[546]), .B(n42085), .Z(n24460) );
  AND U25988 ( .A(a[542]), .B(b[7]), .Z(n24461) );
  XNOR U25989 ( .A(n24462), .B(n24461), .Z(n24463) );
  XNOR U25990 ( .A(n24464), .B(n24463), .Z(n24469) );
  XOR U25991 ( .A(n24470), .B(n24469), .Z(n24448) );
  NANDN U25992 ( .A(n24425), .B(n24424), .Z(n24429) );
  NANDN U25993 ( .A(n24427), .B(n24426), .Z(n24428) );
  AND U25994 ( .A(n24429), .B(n24428), .Z(n24447) );
  XNOR U25995 ( .A(n24448), .B(n24447), .Z(n24449) );
  NANDN U25996 ( .A(n24431), .B(n24430), .Z(n24435) );
  NAND U25997 ( .A(n24433), .B(n24432), .Z(n24434) );
  NAND U25998 ( .A(n24435), .B(n24434), .Z(n24450) );
  XNOR U25999 ( .A(n24449), .B(n24450), .Z(n24441) );
  XNOR U26000 ( .A(n24442), .B(n24441), .Z(n24443) );
  XNOR U26001 ( .A(n24444), .B(n24443), .Z(n24473) );
  XNOR U26002 ( .A(sreg[1566]), .B(n24473), .Z(n24475) );
  NANDN U26003 ( .A(sreg[1565]), .B(n24436), .Z(n24440) );
  NAND U26004 ( .A(n24438), .B(n24437), .Z(n24439) );
  NAND U26005 ( .A(n24440), .B(n24439), .Z(n24474) );
  XNOR U26006 ( .A(n24475), .B(n24474), .Z(c[1566]) );
  NANDN U26007 ( .A(n24442), .B(n24441), .Z(n24446) );
  NANDN U26008 ( .A(n24444), .B(n24443), .Z(n24445) );
  AND U26009 ( .A(n24446), .B(n24445), .Z(n24481) );
  NANDN U26010 ( .A(n24448), .B(n24447), .Z(n24452) );
  NANDN U26011 ( .A(n24450), .B(n24449), .Z(n24451) );
  AND U26012 ( .A(n24452), .B(n24451), .Z(n24479) );
  NAND U26013 ( .A(n42143), .B(n24453), .Z(n24455) );
  XNOR U26014 ( .A(a[545]), .B(n4149), .Z(n24490) );
  NAND U26015 ( .A(n42144), .B(n24490), .Z(n24454) );
  AND U26016 ( .A(n24455), .B(n24454), .Z(n24505) );
  XOR U26017 ( .A(a[549]), .B(n42012), .Z(n24493) );
  XNOR U26018 ( .A(n24505), .B(n24504), .Z(n24507) );
  AND U26019 ( .A(a[551]), .B(b[0]), .Z(n24457) );
  XNOR U26020 ( .A(n24457), .B(n4071), .Z(n24459) );
  NANDN U26021 ( .A(b[0]), .B(a[550]), .Z(n24458) );
  NAND U26022 ( .A(n24459), .B(n24458), .Z(n24501) );
  XOR U26023 ( .A(a[547]), .B(n42085), .Z(n24497) );
  AND U26024 ( .A(a[543]), .B(b[7]), .Z(n24498) );
  XNOR U26025 ( .A(n24499), .B(n24498), .Z(n24500) );
  XNOR U26026 ( .A(n24501), .B(n24500), .Z(n24506) );
  XOR U26027 ( .A(n24507), .B(n24506), .Z(n24485) );
  NANDN U26028 ( .A(n24462), .B(n24461), .Z(n24466) );
  NANDN U26029 ( .A(n24464), .B(n24463), .Z(n24465) );
  AND U26030 ( .A(n24466), .B(n24465), .Z(n24484) );
  XNOR U26031 ( .A(n24485), .B(n24484), .Z(n24486) );
  NANDN U26032 ( .A(n24468), .B(n24467), .Z(n24472) );
  NAND U26033 ( .A(n24470), .B(n24469), .Z(n24471) );
  NAND U26034 ( .A(n24472), .B(n24471), .Z(n24487) );
  XNOR U26035 ( .A(n24486), .B(n24487), .Z(n24478) );
  XNOR U26036 ( .A(n24479), .B(n24478), .Z(n24480) );
  XNOR U26037 ( .A(n24481), .B(n24480), .Z(n24510) );
  XNOR U26038 ( .A(sreg[1567]), .B(n24510), .Z(n24512) );
  NANDN U26039 ( .A(sreg[1566]), .B(n24473), .Z(n24477) );
  NAND U26040 ( .A(n24475), .B(n24474), .Z(n24476) );
  NAND U26041 ( .A(n24477), .B(n24476), .Z(n24511) );
  XNOR U26042 ( .A(n24512), .B(n24511), .Z(c[1567]) );
  NANDN U26043 ( .A(n24479), .B(n24478), .Z(n24483) );
  NANDN U26044 ( .A(n24481), .B(n24480), .Z(n24482) );
  AND U26045 ( .A(n24483), .B(n24482), .Z(n24518) );
  NANDN U26046 ( .A(n24485), .B(n24484), .Z(n24489) );
  NANDN U26047 ( .A(n24487), .B(n24486), .Z(n24488) );
  AND U26048 ( .A(n24489), .B(n24488), .Z(n24516) );
  NAND U26049 ( .A(n42143), .B(n24490), .Z(n24492) );
  XNOR U26050 ( .A(a[546]), .B(n4149), .Z(n24527) );
  NAND U26051 ( .A(n42144), .B(n24527), .Z(n24491) );
  AND U26052 ( .A(n24492), .B(n24491), .Z(n24542) );
  XOR U26053 ( .A(a[550]), .B(n42012), .Z(n24530) );
  XNOR U26054 ( .A(n24542), .B(n24541), .Z(n24544) );
  AND U26055 ( .A(a[552]), .B(b[0]), .Z(n24494) );
  XNOR U26056 ( .A(n24494), .B(n4071), .Z(n24496) );
  NANDN U26057 ( .A(b[0]), .B(a[551]), .Z(n24495) );
  NAND U26058 ( .A(n24496), .B(n24495), .Z(n24538) );
  XOR U26059 ( .A(a[548]), .B(n42085), .Z(n24531) );
  AND U26060 ( .A(a[544]), .B(b[7]), .Z(n24535) );
  XNOR U26061 ( .A(n24536), .B(n24535), .Z(n24537) );
  XNOR U26062 ( .A(n24538), .B(n24537), .Z(n24543) );
  XOR U26063 ( .A(n24544), .B(n24543), .Z(n24522) );
  NANDN U26064 ( .A(n24499), .B(n24498), .Z(n24503) );
  NANDN U26065 ( .A(n24501), .B(n24500), .Z(n24502) );
  AND U26066 ( .A(n24503), .B(n24502), .Z(n24521) );
  XNOR U26067 ( .A(n24522), .B(n24521), .Z(n24523) );
  NANDN U26068 ( .A(n24505), .B(n24504), .Z(n24509) );
  NAND U26069 ( .A(n24507), .B(n24506), .Z(n24508) );
  NAND U26070 ( .A(n24509), .B(n24508), .Z(n24524) );
  XNOR U26071 ( .A(n24523), .B(n24524), .Z(n24515) );
  XNOR U26072 ( .A(n24516), .B(n24515), .Z(n24517) );
  XNOR U26073 ( .A(n24518), .B(n24517), .Z(n24547) );
  XNOR U26074 ( .A(sreg[1568]), .B(n24547), .Z(n24549) );
  NANDN U26075 ( .A(sreg[1567]), .B(n24510), .Z(n24514) );
  NAND U26076 ( .A(n24512), .B(n24511), .Z(n24513) );
  NAND U26077 ( .A(n24514), .B(n24513), .Z(n24548) );
  XNOR U26078 ( .A(n24549), .B(n24548), .Z(c[1568]) );
  NANDN U26079 ( .A(n24516), .B(n24515), .Z(n24520) );
  NANDN U26080 ( .A(n24518), .B(n24517), .Z(n24519) );
  AND U26081 ( .A(n24520), .B(n24519), .Z(n24555) );
  NANDN U26082 ( .A(n24522), .B(n24521), .Z(n24526) );
  NANDN U26083 ( .A(n24524), .B(n24523), .Z(n24525) );
  AND U26084 ( .A(n24526), .B(n24525), .Z(n24553) );
  NAND U26085 ( .A(n42143), .B(n24527), .Z(n24529) );
  XNOR U26086 ( .A(a[547]), .B(n4150), .Z(n24564) );
  NAND U26087 ( .A(n42144), .B(n24564), .Z(n24528) );
  AND U26088 ( .A(n24529), .B(n24528), .Z(n24579) );
  XOR U26089 ( .A(a[551]), .B(n42012), .Z(n24567) );
  XNOR U26090 ( .A(n24579), .B(n24578), .Z(n24581) );
  XOR U26091 ( .A(a[549]), .B(n42085), .Z(n24571) );
  AND U26092 ( .A(a[545]), .B(b[7]), .Z(n24572) );
  XNOR U26093 ( .A(n24573), .B(n24572), .Z(n24574) );
  AND U26094 ( .A(a[553]), .B(b[0]), .Z(n24532) );
  XNOR U26095 ( .A(n24532), .B(n4071), .Z(n24534) );
  NANDN U26096 ( .A(b[0]), .B(a[552]), .Z(n24533) );
  NAND U26097 ( .A(n24534), .B(n24533), .Z(n24575) );
  XNOR U26098 ( .A(n24574), .B(n24575), .Z(n24580) );
  XOR U26099 ( .A(n24581), .B(n24580), .Z(n24559) );
  NANDN U26100 ( .A(n24536), .B(n24535), .Z(n24540) );
  NANDN U26101 ( .A(n24538), .B(n24537), .Z(n24539) );
  AND U26102 ( .A(n24540), .B(n24539), .Z(n24558) );
  XNOR U26103 ( .A(n24559), .B(n24558), .Z(n24560) );
  NANDN U26104 ( .A(n24542), .B(n24541), .Z(n24546) );
  NAND U26105 ( .A(n24544), .B(n24543), .Z(n24545) );
  NAND U26106 ( .A(n24546), .B(n24545), .Z(n24561) );
  XNOR U26107 ( .A(n24560), .B(n24561), .Z(n24552) );
  XNOR U26108 ( .A(n24553), .B(n24552), .Z(n24554) );
  XNOR U26109 ( .A(n24555), .B(n24554), .Z(n24584) );
  XNOR U26110 ( .A(sreg[1569]), .B(n24584), .Z(n24586) );
  NANDN U26111 ( .A(sreg[1568]), .B(n24547), .Z(n24551) );
  NAND U26112 ( .A(n24549), .B(n24548), .Z(n24550) );
  NAND U26113 ( .A(n24551), .B(n24550), .Z(n24585) );
  XNOR U26114 ( .A(n24586), .B(n24585), .Z(c[1569]) );
  NANDN U26115 ( .A(n24553), .B(n24552), .Z(n24557) );
  NANDN U26116 ( .A(n24555), .B(n24554), .Z(n24556) );
  AND U26117 ( .A(n24557), .B(n24556), .Z(n24592) );
  NANDN U26118 ( .A(n24559), .B(n24558), .Z(n24563) );
  NANDN U26119 ( .A(n24561), .B(n24560), .Z(n24562) );
  AND U26120 ( .A(n24563), .B(n24562), .Z(n24590) );
  NAND U26121 ( .A(n42143), .B(n24564), .Z(n24566) );
  XNOR U26122 ( .A(a[548]), .B(n4150), .Z(n24601) );
  NAND U26123 ( .A(n42144), .B(n24601), .Z(n24565) );
  AND U26124 ( .A(n24566), .B(n24565), .Z(n24616) );
  XOR U26125 ( .A(a[552]), .B(n42012), .Z(n24604) );
  XNOR U26126 ( .A(n24616), .B(n24615), .Z(n24618) );
  AND U26127 ( .A(a[554]), .B(b[0]), .Z(n24568) );
  XNOR U26128 ( .A(n24568), .B(n4071), .Z(n24570) );
  NANDN U26129 ( .A(b[0]), .B(a[553]), .Z(n24569) );
  NAND U26130 ( .A(n24570), .B(n24569), .Z(n24612) );
  XOR U26131 ( .A(a[550]), .B(n42085), .Z(n24605) );
  AND U26132 ( .A(a[546]), .B(b[7]), .Z(n24609) );
  XNOR U26133 ( .A(n24610), .B(n24609), .Z(n24611) );
  XNOR U26134 ( .A(n24612), .B(n24611), .Z(n24617) );
  XOR U26135 ( .A(n24618), .B(n24617), .Z(n24596) );
  NANDN U26136 ( .A(n24573), .B(n24572), .Z(n24577) );
  NANDN U26137 ( .A(n24575), .B(n24574), .Z(n24576) );
  AND U26138 ( .A(n24577), .B(n24576), .Z(n24595) );
  XNOR U26139 ( .A(n24596), .B(n24595), .Z(n24597) );
  NANDN U26140 ( .A(n24579), .B(n24578), .Z(n24583) );
  NAND U26141 ( .A(n24581), .B(n24580), .Z(n24582) );
  NAND U26142 ( .A(n24583), .B(n24582), .Z(n24598) );
  XNOR U26143 ( .A(n24597), .B(n24598), .Z(n24589) );
  XNOR U26144 ( .A(n24590), .B(n24589), .Z(n24591) );
  XNOR U26145 ( .A(n24592), .B(n24591), .Z(n24621) );
  XNOR U26146 ( .A(sreg[1570]), .B(n24621), .Z(n24623) );
  NANDN U26147 ( .A(sreg[1569]), .B(n24584), .Z(n24588) );
  NAND U26148 ( .A(n24586), .B(n24585), .Z(n24587) );
  NAND U26149 ( .A(n24588), .B(n24587), .Z(n24622) );
  XNOR U26150 ( .A(n24623), .B(n24622), .Z(c[1570]) );
  NANDN U26151 ( .A(n24590), .B(n24589), .Z(n24594) );
  NANDN U26152 ( .A(n24592), .B(n24591), .Z(n24593) );
  AND U26153 ( .A(n24594), .B(n24593), .Z(n24629) );
  NANDN U26154 ( .A(n24596), .B(n24595), .Z(n24600) );
  NANDN U26155 ( .A(n24598), .B(n24597), .Z(n24599) );
  AND U26156 ( .A(n24600), .B(n24599), .Z(n24627) );
  NAND U26157 ( .A(n42143), .B(n24601), .Z(n24603) );
  XNOR U26158 ( .A(a[549]), .B(n4150), .Z(n24638) );
  NAND U26159 ( .A(n42144), .B(n24638), .Z(n24602) );
  AND U26160 ( .A(n24603), .B(n24602), .Z(n24653) );
  XOR U26161 ( .A(a[553]), .B(n42012), .Z(n24641) );
  XNOR U26162 ( .A(n24653), .B(n24652), .Z(n24655) );
  XOR U26163 ( .A(a[551]), .B(n42085), .Z(n24645) );
  AND U26164 ( .A(a[547]), .B(b[7]), .Z(n24646) );
  XNOR U26165 ( .A(n24647), .B(n24646), .Z(n24648) );
  AND U26166 ( .A(a[555]), .B(b[0]), .Z(n24606) );
  XNOR U26167 ( .A(n24606), .B(n4071), .Z(n24608) );
  NANDN U26168 ( .A(b[0]), .B(a[554]), .Z(n24607) );
  NAND U26169 ( .A(n24608), .B(n24607), .Z(n24649) );
  XNOR U26170 ( .A(n24648), .B(n24649), .Z(n24654) );
  XOR U26171 ( .A(n24655), .B(n24654), .Z(n24633) );
  NANDN U26172 ( .A(n24610), .B(n24609), .Z(n24614) );
  NANDN U26173 ( .A(n24612), .B(n24611), .Z(n24613) );
  AND U26174 ( .A(n24614), .B(n24613), .Z(n24632) );
  XNOR U26175 ( .A(n24633), .B(n24632), .Z(n24634) );
  NANDN U26176 ( .A(n24616), .B(n24615), .Z(n24620) );
  NAND U26177 ( .A(n24618), .B(n24617), .Z(n24619) );
  NAND U26178 ( .A(n24620), .B(n24619), .Z(n24635) );
  XNOR U26179 ( .A(n24634), .B(n24635), .Z(n24626) );
  XNOR U26180 ( .A(n24627), .B(n24626), .Z(n24628) );
  XNOR U26181 ( .A(n24629), .B(n24628), .Z(n24658) );
  XNOR U26182 ( .A(sreg[1571]), .B(n24658), .Z(n24660) );
  NANDN U26183 ( .A(sreg[1570]), .B(n24621), .Z(n24625) );
  NAND U26184 ( .A(n24623), .B(n24622), .Z(n24624) );
  NAND U26185 ( .A(n24625), .B(n24624), .Z(n24659) );
  XNOR U26186 ( .A(n24660), .B(n24659), .Z(c[1571]) );
  NANDN U26187 ( .A(n24627), .B(n24626), .Z(n24631) );
  NANDN U26188 ( .A(n24629), .B(n24628), .Z(n24630) );
  AND U26189 ( .A(n24631), .B(n24630), .Z(n24666) );
  NANDN U26190 ( .A(n24633), .B(n24632), .Z(n24637) );
  NANDN U26191 ( .A(n24635), .B(n24634), .Z(n24636) );
  AND U26192 ( .A(n24637), .B(n24636), .Z(n24664) );
  NAND U26193 ( .A(n42143), .B(n24638), .Z(n24640) );
  XNOR U26194 ( .A(a[550]), .B(n4150), .Z(n24675) );
  NAND U26195 ( .A(n42144), .B(n24675), .Z(n24639) );
  AND U26196 ( .A(n24640), .B(n24639), .Z(n24690) );
  XOR U26197 ( .A(a[554]), .B(n42012), .Z(n24678) );
  XNOR U26198 ( .A(n24690), .B(n24689), .Z(n24692) );
  AND U26199 ( .A(a[556]), .B(b[0]), .Z(n24642) );
  XNOR U26200 ( .A(n24642), .B(n4071), .Z(n24644) );
  NANDN U26201 ( .A(b[0]), .B(a[555]), .Z(n24643) );
  NAND U26202 ( .A(n24644), .B(n24643), .Z(n24686) );
  XOR U26203 ( .A(a[552]), .B(n42085), .Z(n24682) );
  AND U26204 ( .A(a[548]), .B(b[7]), .Z(n24683) );
  XNOR U26205 ( .A(n24684), .B(n24683), .Z(n24685) );
  XNOR U26206 ( .A(n24686), .B(n24685), .Z(n24691) );
  XOR U26207 ( .A(n24692), .B(n24691), .Z(n24670) );
  NANDN U26208 ( .A(n24647), .B(n24646), .Z(n24651) );
  NANDN U26209 ( .A(n24649), .B(n24648), .Z(n24650) );
  AND U26210 ( .A(n24651), .B(n24650), .Z(n24669) );
  XNOR U26211 ( .A(n24670), .B(n24669), .Z(n24671) );
  NANDN U26212 ( .A(n24653), .B(n24652), .Z(n24657) );
  NAND U26213 ( .A(n24655), .B(n24654), .Z(n24656) );
  NAND U26214 ( .A(n24657), .B(n24656), .Z(n24672) );
  XNOR U26215 ( .A(n24671), .B(n24672), .Z(n24663) );
  XNOR U26216 ( .A(n24664), .B(n24663), .Z(n24665) );
  XNOR U26217 ( .A(n24666), .B(n24665), .Z(n24695) );
  XNOR U26218 ( .A(sreg[1572]), .B(n24695), .Z(n24697) );
  NANDN U26219 ( .A(sreg[1571]), .B(n24658), .Z(n24662) );
  NAND U26220 ( .A(n24660), .B(n24659), .Z(n24661) );
  NAND U26221 ( .A(n24662), .B(n24661), .Z(n24696) );
  XNOR U26222 ( .A(n24697), .B(n24696), .Z(c[1572]) );
  NANDN U26223 ( .A(n24664), .B(n24663), .Z(n24668) );
  NANDN U26224 ( .A(n24666), .B(n24665), .Z(n24667) );
  AND U26225 ( .A(n24668), .B(n24667), .Z(n24703) );
  NANDN U26226 ( .A(n24670), .B(n24669), .Z(n24674) );
  NANDN U26227 ( .A(n24672), .B(n24671), .Z(n24673) );
  AND U26228 ( .A(n24674), .B(n24673), .Z(n24701) );
  NAND U26229 ( .A(n42143), .B(n24675), .Z(n24677) );
  XNOR U26230 ( .A(a[551]), .B(n4150), .Z(n24712) );
  NAND U26231 ( .A(n42144), .B(n24712), .Z(n24676) );
  AND U26232 ( .A(n24677), .B(n24676), .Z(n24727) );
  XOR U26233 ( .A(a[555]), .B(n42012), .Z(n24715) );
  XNOR U26234 ( .A(n24727), .B(n24726), .Z(n24729) );
  AND U26235 ( .A(a[557]), .B(b[0]), .Z(n24679) );
  XNOR U26236 ( .A(n24679), .B(n4071), .Z(n24681) );
  NANDN U26237 ( .A(b[0]), .B(a[556]), .Z(n24680) );
  NAND U26238 ( .A(n24681), .B(n24680), .Z(n24723) );
  XOR U26239 ( .A(a[553]), .B(n42085), .Z(n24716) );
  AND U26240 ( .A(a[549]), .B(b[7]), .Z(n24720) );
  XNOR U26241 ( .A(n24721), .B(n24720), .Z(n24722) );
  XNOR U26242 ( .A(n24723), .B(n24722), .Z(n24728) );
  XOR U26243 ( .A(n24729), .B(n24728), .Z(n24707) );
  NANDN U26244 ( .A(n24684), .B(n24683), .Z(n24688) );
  NANDN U26245 ( .A(n24686), .B(n24685), .Z(n24687) );
  AND U26246 ( .A(n24688), .B(n24687), .Z(n24706) );
  XNOR U26247 ( .A(n24707), .B(n24706), .Z(n24708) );
  NANDN U26248 ( .A(n24690), .B(n24689), .Z(n24694) );
  NAND U26249 ( .A(n24692), .B(n24691), .Z(n24693) );
  NAND U26250 ( .A(n24694), .B(n24693), .Z(n24709) );
  XNOR U26251 ( .A(n24708), .B(n24709), .Z(n24700) );
  XNOR U26252 ( .A(n24701), .B(n24700), .Z(n24702) );
  XNOR U26253 ( .A(n24703), .B(n24702), .Z(n24732) );
  XNOR U26254 ( .A(sreg[1573]), .B(n24732), .Z(n24734) );
  NANDN U26255 ( .A(sreg[1572]), .B(n24695), .Z(n24699) );
  NAND U26256 ( .A(n24697), .B(n24696), .Z(n24698) );
  NAND U26257 ( .A(n24699), .B(n24698), .Z(n24733) );
  XNOR U26258 ( .A(n24734), .B(n24733), .Z(c[1573]) );
  NANDN U26259 ( .A(n24701), .B(n24700), .Z(n24705) );
  NANDN U26260 ( .A(n24703), .B(n24702), .Z(n24704) );
  AND U26261 ( .A(n24705), .B(n24704), .Z(n24740) );
  NANDN U26262 ( .A(n24707), .B(n24706), .Z(n24711) );
  NANDN U26263 ( .A(n24709), .B(n24708), .Z(n24710) );
  AND U26264 ( .A(n24711), .B(n24710), .Z(n24738) );
  NAND U26265 ( .A(n42143), .B(n24712), .Z(n24714) );
  XNOR U26266 ( .A(a[552]), .B(n4150), .Z(n24749) );
  NAND U26267 ( .A(n42144), .B(n24749), .Z(n24713) );
  AND U26268 ( .A(n24714), .B(n24713), .Z(n24764) );
  XOR U26269 ( .A(a[556]), .B(n42012), .Z(n24752) );
  XNOR U26270 ( .A(n24764), .B(n24763), .Z(n24766) );
  XOR U26271 ( .A(a[554]), .B(n42085), .Z(n24756) );
  AND U26272 ( .A(a[550]), .B(b[7]), .Z(n24757) );
  XNOR U26273 ( .A(n24758), .B(n24757), .Z(n24759) );
  AND U26274 ( .A(a[558]), .B(b[0]), .Z(n24717) );
  XNOR U26275 ( .A(n24717), .B(n4071), .Z(n24719) );
  NANDN U26276 ( .A(b[0]), .B(a[557]), .Z(n24718) );
  NAND U26277 ( .A(n24719), .B(n24718), .Z(n24760) );
  XNOR U26278 ( .A(n24759), .B(n24760), .Z(n24765) );
  XOR U26279 ( .A(n24766), .B(n24765), .Z(n24744) );
  NANDN U26280 ( .A(n24721), .B(n24720), .Z(n24725) );
  NANDN U26281 ( .A(n24723), .B(n24722), .Z(n24724) );
  AND U26282 ( .A(n24725), .B(n24724), .Z(n24743) );
  XNOR U26283 ( .A(n24744), .B(n24743), .Z(n24745) );
  NANDN U26284 ( .A(n24727), .B(n24726), .Z(n24731) );
  NAND U26285 ( .A(n24729), .B(n24728), .Z(n24730) );
  NAND U26286 ( .A(n24731), .B(n24730), .Z(n24746) );
  XNOR U26287 ( .A(n24745), .B(n24746), .Z(n24737) );
  XNOR U26288 ( .A(n24738), .B(n24737), .Z(n24739) );
  XNOR U26289 ( .A(n24740), .B(n24739), .Z(n24769) );
  XNOR U26290 ( .A(sreg[1574]), .B(n24769), .Z(n24771) );
  NANDN U26291 ( .A(sreg[1573]), .B(n24732), .Z(n24736) );
  NAND U26292 ( .A(n24734), .B(n24733), .Z(n24735) );
  NAND U26293 ( .A(n24736), .B(n24735), .Z(n24770) );
  XNOR U26294 ( .A(n24771), .B(n24770), .Z(c[1574]) );
  NANDN U26295 ( .A(n24738), .B(n24737), .Z(n24742) );
  NANDN U26296 ( .A(n24740), .B(n24739), .Z(n24741) );
  AND U26297 ( .A(n24742), .B(n24741), .Z(n24777) );
  NANDN U26298 ( .A(n24744), .B(n24743), .Z(n24748) );
  NANDN U26299 ( .A(n24746), .B(n24745), .Z(n24747) );
  AND U26300 ( .A(n24748), .B(n24747), .Z(n24775) );
  NAND U26301 ( .A(n42143), .B(n24749), .Z(n24751) );
  XNOR U26302 ( .A(a[553]), .B(n4150), .Z(n24786) );
  NAND U26303 ( .A(n42144), .B(n24786), .Z(n24750) );
  AND U26304 ( .A(n24751), .B(n24750), .Z(n24801) );
  XOR U26305 ( .A(a[557]), .B(n42012), .Z(n24789) );
  XNOR U26306 ( .A(n24801), .B(n24800), .Z(n24803) );
  AND U26307 ( .A(a[559]), .B(b[0]), .Z(n24753) );
  XNOR U26308 ( .A(n24753), .B(n4071), .Z(n24755) );
  NANDN U26309 ( .A(b[0]), .B(a[558]), .Z(n24754) );
  NAND U26310 ( .A(n24755), .B(n24754), .Z(n24797) );
  XOR U26311 ( .A(a[555]), .B(n42085), .Z(n24790) );
  AND U26312 ( .A(a[551]), .B(b[7]), .Z(n24794) );
  XNOR U26313 ( .A(n24795), .B(n24794), .Z(n24796) );
  XNOR U26314 ( .A(n24797), .B(n24796), .Z(n24802) );
  XOR U26315 ( .A(n24803), .B(n24802), .Z(n24781) );
  NANDN U26316 ( .A(n24758), .B(n24757), .Z(n24762) );
  NANDN U26317 ( .A(n24760), .B(n24759), .Z(n24761) );
  AND U26318 ( .A(n24762), .B(n24761), .Z(n24780) );
  XNOR U26319 ( .A(n24781), .B(n24780), .Z(n24782) );
  NANDN U26320 ( .A(n24764), .B(n24763), .Z(n24768) );
  NAND U26321 ( .A(n24766), .B(n24765), .Z(n24767) );
  NAND U26322 ( .A(n24768), .B(n24767), .Z(n24783) );
  XNOR U26323 ( .A(n24782), .B(n24783), .Z(n24774) );
  XNOR U26324 ( .A(n24775), .B(n24774), .Z(n24776) );
  XNOR U26325 ( .A(n24777), .B(n24776), .Z(n24806) );
  XNOR U26326 ( .A(sreg[1575]), .B(n24806), .Z(n24808) );
  NANDN U26327 ( .A(sreg[1574]), .B(n24769), .Z(n24773) );
  NAND U26328 ( .A(n24771), .B(n24770), .Z(n24772) );
  NAND U26329 ( .A(n24773), .B(n24772), .Z(n24807) );
  XNOR U26330 ( .A(n24808), .B(n24807), .Z(c[1575]) );
  NANDN U26331 ( .A(n24775), .B(n24774), .Z(n24779) );
  NANDN U26332 ( .A(n24777), .B(n24776), .Z(n24778) );
  AND U26333 ( .A(n24779), .B(n24778), .Z(n24814) );
  NANDN U26334 ( .A(n24781), .B(n24780), .Z(n24785) );
  NANDN U26335 ( .A(n24783), .B(n24782), .Z(n24784) );
  AND U26336 ( .A(n24785), .B(n24784), .Z(n24812) );
  NAND U26337 ( .A(n42143), .B(n24786), .Z(n24788) );
  XNOR U26338 ( .A(a[554]), .B(n4151), .Z(n24823) );
  NAND U26339 ( .A(n42144), .B(n24823), .Z(n24787) );
  AND U26340 ( .A(n24788), .B(n24787), .Z(n24838) );
  XOR U26341 ( .A(a[558]), .B(n42012), .Z(n24826) );
  XNOR U26342 ( .A(n24838), .B(n24837), .Z(n24840) );
  XOR U26343 ( .A(a[556]), .B(n42085), .Z(n24830) );
  AND U26344 ( .A(a[552]), .B(b[7]), .Z(n24831) );
  XNOR U26345 ( .A(n24832), .B(n24831), .Z(n24833) );
  AND U26346 ( .A(a[560]), .B(b[0]), .Z(n24791) );
  XNOR U26347 ( .A(n24791), .B(n4071), .Z(n24793) );
  NANDN U26348 ( .A(b[0]), .B(a[559]), .Z(n24792) );
  NAND U26349 ( .A(n24793), .B(n24792), .Z(n24834) );
  XNOR U26350 ( .A(n24833), .B(n24834), .Z(n24839) );
  XOR U26351 ( .A(n24840), .B(n24839), .Z(n24818) );
  NANDN U26352 ( .A(n24795), .B(n24794), .Z(n24799) );
  NANDN U26353 ( .A(n24797), .B(n24796), .Z(n24798) );
  AND U26354 ( .A(n24799), .B(n24798), .Z(n24817) );
  XNOR U26355 ( .A(n24818), .B(n24817), .Z(n24819) );
  NANDN U26356 ( .A(n24801), .B(n24800), .Z(n24805) );
  NAND U26357 ( .A(n24803), .B(n24802), .Z(n24804) );
  NAND U26358 ( .A(n24805), .B(n24804), .Z(n24820) );
  XNOR U26359 ( .A(n24819), .B(n24820), .Z(n24811) );
  XNOR U26360 ( .A(n24812), .B(n24811), .Z(n24813) );
  XNOR U26361 ( .A(n24814), .B(n24813), .Z(n24843) );
  XNOR U26362 ( .A(sreg[1576]), .B(n24843), .Z(n24845) );
  NANDN U26363 ( .A(sreg[1575]), .B(n24806), .Z(n24810) );
  NAND U26364 ( .A(n24808), .B(n24807), .Z(n24809) );
  NAND U26365 ( .A(n24810), .B(n24809), .Z(n24844) );
  XNOR U26366 ( .A(n24845), .B(n24844), .Z(c[1576]) );
  NANDN U26367 ( .A(n24812), .B(n24811), .Z(n24816) );
  NANDN U26368 ( .A(n24814), .B(n24813), .Z(n24815) );
  AND U26369 ( .A(n24816), .B(n24815), .Z(n24851) );
  NANDN U26370 ( .A(n24818), .B(n24817), .Z(n24822) );
  NANDN U26371 ( .A(n24820), .B(n24819), .Z(n24821) );
  AND U26372 ( .A(n24822), .B(n24821), .Z(n24849) );
  NAND U26373 ( .A(n42143), .B(n24823), .Z(n24825) );
  XNOR U26374 ( .A(a[555]), .B(n4151), .Z(n24860) );
  NAND U26375 ( .A(n42144), .B(n24860), .Z(n24824) );
  AND U26376 ( .A(n24825), .B(n24824), .Z(n24875) );
  XOR U26377 ( .A(a[559]), .B(n42012), .Z(n24863) );
  XNOR U26378 ( .A(n24875), .B(n24874), .Z(n24877) );
  AND U26379 ( .A(a[561]), .B(b[0]), .Z(n24827) );
  XNOR U26380 ( .A(n24827), .B(n4071), .Z(n24829) );
  NANDN U26381 ( .A(b[0]), .B(a[560]), .Z(n24828) );
  NAND U26382 ( .A(n24829), .B(n24828), .Z(n24871) );
  XOR U26383 ( .A(a[557]), .B(n42085), .Z(n24867) );
  AND U26384 ( .A(a[553]), .B(b[7]), .Z(n24868) );
  XNOR U26385 ( .A(n24869), .B(n24868), .Z(n24870) );
  XNOR U26386 ( .A(n24871), .B(n24870), .Z(n24876) );
  XOR U26387 ( .A(n24877), .B(n24876), .Z(n24855) );
  NANDN U26388 ( .A(n24832), .B(n24831), .Z(n24836) );
  NANDN U26389 ( .A(n24834), .B(n24833), .Z(n24835) );
  AND U26390 ( .A(n24836), .B(n24835), .Z(n24854) );
  XNOR U26391 ( .A(n24855), .B(n24854), .Z(n24856) );
  NANDN U26392 ( .A(n24838), .B(n24837), .Z(n24842) );
  NAND U26393 ( .A(n24840), .B(n24839), .Z(n24841) );
  NAND U26394 ( .A(n24842), .B(n24841), .Z(n24857) );
  XNOR U26395 ( .A(n24856), .B(n24857), .Z(n24848) );
  XNOR U26396 ( .A(n24849), .B(n24848), .Z(n24850) );
  XNOR U26397 ( .A(n24851), .B(n24850), .Z(n24880) );
  XNOR U26398 ( .A(sreg[1577]), .B(n24880), .Z(n24882) );
  NANDN U26399 ( .A(sreg[1576]), .B(n24843), .Z(n24847) );
  NAND U26400 ( .A(n24845), .B(n24844), .Z(n24846) );
  NAND U26401 ( .A(n24847), .B(n24846), .Z(n24881) );
  XNOR U26402 ( .A(n24882), .B(n24881), .Z(c[1577]) );
  NANDN U26403 ( .A(n24849), .B(n24848), .Z(n24853) );
  NANDN U26404 ( .A(n24851), .B(n24850), .Z(n24852) );
  AND U26405 ( .A(n24853), .B(n24852), .Z(n24888) );
  NANDN U26406 ( .A(n24855), .B(n24854), .Z(n24859) );
  NANDN U26407 ( .A(n24857), .B(n24856), .Z(n24858) );
  AND U26408 ( .A(n24859), .B(n24858), .Z(n24886) );
  NAND U26409 ( .A(n42143), .B(n24860), .Z(n24862) );
  XNOR U26410 ( .A(a[556]), .B(n4151), .Z(n24897) );
  NAND U26411 ( .A(n42144), .B(n24897), .Z(n24861) );
  AND U26412 ( .A(n24862), .B(n24861), .Z(n24912) );
  XOR U26413 ( .A(a[560]), .B(n42012), .Z(n24900) );
  XNOR U26414 ( .A(n24912), .B(n24911), .Z(n24914) );
  AND U26415 ( .A(a[562]), .B(b[0]), .Z(n24864) );
  XNOR U26416 ( .A(n24864), .B(n4071), .Z(n24866) );
  NANDN U26417 ( .A(b[0]), .B(a[561]), .Z(n24865) );
  NAND U26418 ( .A(n24866), .B(n24865), .Z(n24908) );
  XOR U26419 ( .A(a[558]), .B(n42085), .Z(n24901) );
  AND U26420 ( .A(a[554]), .B(b[7]), .Z(n24905) );
  XNOR U26421 ( .A(n24906), .B(n24905), .Z(n24907) );
  XNOR U26422 ( .A(n24908), .B(n24907), .Z(n24913) );
  XOR U26423 ( .A(n24914), .B(n24913), .Z(n24892) );
  NANDN U26424 ( .A(n24869), .B(n24868), .Z(n24873) );
  NANDN U26425 ( .A(n24871), .B(n24870), .Z(n24872) );
  AND U26426 ( .A(n24873), .B(n24872), .Z(n24891) );
  XNOR U26427 ( .A(n24892), .B(n24891), .Z(n24893) );
  NANDN U26428 ( .A(n24875), .B(n24874), .Z(n24879) );
  NAND U26429 ( .A(n24877), .B(n24876), .Z(n24878) );
  NAND U26430 ( .A(n24879), .B(n24878), .Z(n24894) );
  XNOR U26431 ( .A(n24893), .B(n24894), .Z(n24885) );
  XNOR U26432 ( .A(n24886), .B(n24885), .Z(n24887) );
  XNOR U26433 ( .A(n24888), .B(n24887), .Z(n24917) );
  XNOR U26434 ( .A(sreg[1578]), .B(n24917), .Z(n24919) );
  NANDN U26435 ( .A(sreg[1577]), .B(n24880), .Z(n24884) );
  NAND U26436 ( .A(n24882), .B(n24881), .Z(n24883) );
  NAND U26437 ( .A(n24884), .B(n24883), .Z(n24918) );
  XNOR U26438 ( .A(n24919), .B(n24918), .Z(c[1578]) );
  NANDN U26439 ( .A(n24886), .B(n24885), .Z(n24890) );
  NANDN U26440 ( .A(n24888), .B(n24887), .Z(n24889) );
  AND U26441 ( .A(n24890), .B(n24889), .Z(n24925) );
  NANDN U26442 ( .A(n24892), .B(n24891), .Z(n24896) );
  NANDN U26443 ( .A(n24894), .B(n24893), .Z(n24895) );
  AND U26444 ( .A(n24896), .B(n24895), .Z(n24923) );
  NAND U26445 ( .A(n42143), .B(n24897), .Z(n24899) );
  XNOR U26446 ( .A(a[557]), .B(n4151), .Z(n24934) );
  NAND U26447 ( .A(n42144), .B(n24934), .Z(n24898) );
  AND U26448 ( .A(n24899), .B(n24898), .Z(n24949) );
  XOR U26449 ( .A(a[561]), .B(n42012), .Z(n24937) );
  XNOR U26450 ( .A(n24949), .B(n24948), .Z(n24951) );
  XOR U26451 ( .A(a[559]), .B(n42085), .Z(n24941) );
  AND U26452 ( .A(a[555]), .B(b[7]), .Z(n24942) );
  XNOR U26453 ( .A(n24943), .B(n24942), .Z(n24944) );
  AND U26454 ( .A(a[563]), .B(b[0]), .Z(n24902) );
  XNOR U26455 ( .A(n24902), .B(n4071), .Z(n24904) );
  NANDN U26456 ( .A(b[0]), .B(a[562]), .Z(n24903) );
  NAND U26457 ( .A(n24904), .B(n24903), .Z(n24945) );
  XNOR U26458 ( .A(n24944), .B(n24945), .Z(n24950) );
  XOR U26459 ( .A(n24951), .B(n24950), .Z(n24929) );
  NANDN U26460 ( .A(n24906), .B(n24905), .Z(n24910) );
  NANDN U26461 ( .A(n24908), .B(n24907), .Z(n24909) );
  AND U26462 ( .A(n24910), .B(n24909), .Z(n24928) );
  XNOR U26463 ( .A(n24929), .B(n24928), .Z(n24930) );
  NANDN U26464 ( .A(n24912), .B(n24911), .Z(n24916) );
  NAND U26465 ( .A(n24914), .B(n24913), .Z(n24915) );
  NAND U26466 ( .A(n24916), .B(n24915), .Z(n24931) );
  XNOR U26467 ( .A(n24930), .B(n24931), .Z(n24922) );
  XNOR U26468 ( .A(n24923), .B(n24922), .Z(n24924) );
  XNOR U26469 ( .A(n24925), .B(n24924), .Z(n24954) );
  XNOR U26470 ( .A(sreg[1579]), .B(n24954), .Z(n24956) );
  NANDN U26471 ( .A(sreg[1578]), .B(n24917), .Z(n24921) );
  NAND U26472 ( .A(n24919), .B(n24918), .Z(n24920) );
  NAND U26473 ( .A(n24921), .B(n24920), .Z(n24955) );
  XNOR U26474 ( .A(n24956), .B(n24955), .Z(c[1579]) );
  NANDN U26475 ( .A(n24923), .B(n24922), .Z(n24927) );
  NANDN U26476 ( .A(n24925), .B(n24924), .Z(n24926) );
  AND U26477 ( .A(n24927), .B(n24926), .Z(n24962) );
  NANDN U26478 ( .A(n24929), .B(n24928), .Z(n24933) );
  NANDN U26479 ( .A(n24931), .B(n24930), .Z(n24932) );
  AND U26480 ( .A(n24933), .B(n24932), .Z(n24960) );
  NAND U26481 ( .A(n42143), .B(n24934), .Z(n24936) );
  XNOR U26482 ( .A(a[558]), .B(n4151), .Z(n24971) );
  NAND U26483 ( .A(n42144), .B(n24971), .Z(n24935) );
  AND U26484 ( .A(n24936), .B(n24935), .Z(n24986) );
  XOR U26485 ( .A(a[562]), .B(n42012), .Z(n24974) );
  XNOR U26486 ( .A(n24986), .B(n24985), .Z(n24988) );
  AND U26487 ( .A(b[0]), .B(a[564]), .Z(n24938) );
  XOR U26488 ( .A(b[1]), .B(n24938), .Z(n24940) );
  NANDN U26489 ( .A(n29564), .B(a[563]), .Z(n24939) );
  AND U26490 ( .A(n24940), .B(n24939), .Z(n24981) );
  XOR U26491 ( .A(a[560]), .B(n42085), .Z(n24978) );
  AND U26492 ( .A(a[556]), .B(b[7]), .Z(n24979) );
  XOR U26493 ( .A(n24980), .B(n24979), .Z(n24982) );
  XNOR U26494 ( .A(n24981), .B(n24982), .Z(n24987) );
  XOR U26495 ( .A(n24988), .B(n24987), .Z(n24966) );
  NANDN U26496 ( .A(n24943), .B(n24942), .Z(n24947) );
  NANDN U26497 ( .A(n24945), .B(n24944), .Z(n24946) );
  AND U26498 ( .A(n24947), .B(n24946), .Z(n24965) );
  XNOR U26499 ( .A(n24966), .B(n24965), .Z(n24967) );
  NANDN U26500 ( .A(n24949), .B(n24948), .Z(n24953) );
  NAND U26501 ( .A(n24951), .B(n24950), .Z(n24952) );
  NAND U26502 ( .A(n24953), .B(n24952), .Z(n24968) );
  XNOR U26503 ( .A(n24967), .B(n24968), .Z(n24959) );
  XNOR U26504 ( .A(n24960), .B(n24959), .Z(n24961) );
  XNOR U26505 ( .A(n24962), .B(n24961), .Z(n24991) );
  XNOR U26506 ( .A(sreg[1580]), .B(n24991), .Z(n24993) );
  NANDN U26507 ( .A(sreg[1579]), .B(n24954), .Z(n24958) );
  NAND U26508 ( .A(n24956), .B(n24955), .Z(n24957) );
  NAND U26509 ( .A(n24958), .B(n24957), .Z(n24992) );
  XNOR U26510 ( .A(n24993), .B(n24992), .Z(c[1580]) );
  NANDN U26511 ( .A(n24960), .B(n24959), .Z(n24964) );
  NANDN U26512 ( .A(n24962), .B(n24961), .Z(n24963) );
  AND U26513 ( .A(n24964), .B(n24963), .Z(n24999) );
  NANDN U26514 ( .A(n24966), .B(n24965), .Z(n24970) );
  NANDN U26515 ( .A(n24968), .B(n24967), .Z(n24969) );
  AND U26516 ( .A(n24970), .B(n24969), .Z(n24997) );
  NAND U26517 ( .A(n42143), .B(n24971), .Z(n24973) );
  XNOR U26518 ( .A(a[559]), .B(n4151), .Z(n25008) );
  NAND U26519 ( .A(n42144), .B(n25008), .Z(n24972) );
  AND U26520 ( .A(n24973), .B(n24972), .Z(n25023) );
  XOR U26521 ( .A(a[563]), .B(n42012), .Z(n25011) );
  XNOR U26522 ( .A(n25023), .B(n25022), .Z(n25025) );
  AND U26523 ( .A(a[565]), .B(b[0]), .Z(n24975) );
  XNOR U26524 ( .A(n24975), .B(n4071), .Z(n24977) );
  NANDN U26525 ( .A(b[0]), .B(a[564]), .Z(n24976) );
  NAND U26526 ( .A(n24977), .B(n24976), .Z(n25019) );
  XOR U26527 ( .A(a[561]), .B(n42085), .Z(n25015) );
  AND U26528 ( .A(a[557]), .B(b[7]), .Z(n25016) );
  XNOR U26529 ( .A(n25017), .B(n25016), .Z(n25018) );
  XNOR U26530 ( .A(n25019), .B(n25018), .Z(n25024) );
  XOR U26531 ( .A(n25025), .B(n25024), .Z(n25003) );
  NANDN U26532 ( .A(n24980), .B(n24979), .Z(n24984) );
  NANDN U26533 ( .A(n24982), .B(n24981), .Z(n24983) );
  AND U26534 ( .A(n24984), .B(n24983), .Z(n25002) );
  XNOR U26535 ( .A(n25003), .B(n25002), .Z(n25004) );
  NANDN U26536 ( .A(n24986), .B(n24985), .Z(n24990) );
  NAND U26537 ( .A(n24988), .B(n24987), .Z(n24989) );
  NAND U26538 ( .A(n24990), .B(n24989), .Z(n25005) );
  XNOR U26539 ( .A(n25004), .B(n25005), .Z(n24996) );
  XNOR U26540 ( .A(n24997), .B(n24996), .Z(n24998) );
  XNOR U26541 ( .A(n24999), .B(n24998), .Z(n25028) );
  XNOR U26542 ( .A(sreg[1581]), .B(n25028), .Z(n25030) );
  NANDN U26543 ( .A(sreg[1580]), .B(n24991), .Z(n24995) );
  NAND U26544 ( .A(n24993), .B(n24992), .Z(n24994) );
  NAND U26545 ( .A(n24995), .B(n24994), .Z(n25029) );
  XNOR U26546 ( .A(n25030), .B(n25029), .Z(c[1581]) );
  NANDN U26547 ( .A(n24997), .B(n24996), .Z(n25001) );
  NANDN U26548 ( .A(n24999), .B(n24998), .Z(n25000) );
  AND U26549 ( .A(n25001), .B(n25000), .Z(n25036) );
  NANDN U26550 ( .A(n25003), .B(n25002), .Z(n25007) );
  NANDN U26551 ( .A(n25005), .B(n25004), .Z(n25006) );
  AND U26552 ( .A(n25007), .B(n25006), .Z(n25034) );
  NAND U26553 ( .A(n42143), .B(n25008), .Z(n25010) );
  XNOR U26554 ( .A(a[560]), .B(n4151), .Z(n25045) );
  NAND U26555 ( .A(n42144), .B(n25045), .Z(n25009) );
  AND U26556 ( .A(n25010), .B(n25009), .Z(n25060) );
  XOR U26557 ( .A(a[564]), .B(n42012), .Z(n25048) );
  XNOR U26558 ( .A(n25060), .B(n25059), .Z(n25062) );
  AND U26559 ( .A(a[566]), .B(b[0]), .Z(n25012) );
  XNOR U26560 ( .A(n25012), .B(n4071), .Z(n25014) );
  NANDN U26561 ( .A(b[0]), .B(a[565]), .Z(n25013) );
  NAND U26562 ( .A(n25014), .B(n25013), .Z(n25056) );
  XOR U26563 ( .A(a[562]), .B(n42085), .Z(n25052) );
  AND U26564 ( .A(a[558]), .B(b[7]), .Z(n25053) );
  XNOR U26565 ( .A(n25054), .B(n25053), .Z(n25055) );
  XNOR U26566 ( .A(n25056), .B(n25055), .Z(n25061) );
  XOR U26567 ( .A(n25062), .B(n25061), .Z(n25040) );
  NANDN U26568 ( .A(n25017), .B(n25016), .Z(n25021) );
  NANDN U26569 ( .A(n25019), .B(n25018), .Z(n25020) );
  AND U26570 ( .A(n25021), .B(n25020), .Z(n25039) );
  XNOR U26571 ( .A(n25040), .B(n25039), .Z(n25041) );
  NANDN U26572 ( .A(n25023), .B(n25022), .Z(n25027) );
  NAND U26573 ( .A(n25025), .B(n25024), .Z(n25026) );
  NAND U26574 ( .A(n25027), .B(n25026), .Z(n25042) );
  XNOR U26575 ( .A(n25041), .B(n25042), .Z(n25033) );
  XNOR U26576 ( .A(n25034), .B(n25033), .Z(n25035) );
  XNOR U26577 ( .A(n25036), .B(n25035), .Z(n25065) );
  XNOR U26578 ( .A(sreg[1582]), .B(n25065), .Z(n25067) );
  NANDN U26579 ( .A(sreg[1581]), .B(n25028), .Z(n25032) );
  NAND U26580 ( .A(n25030), .B(n25029), .Z(n25031) );
  NAND U26581 ( .A(n25032), .B(n25031), .Z(n25066) );
  XNOR U26582 ( .A(n25067), .B(n25066), .Z(c[1582]) );
  NANDN U26583 ( .A(n25034), .B(n25033), .Z(n25038) );
  NANDN U26584 ( .A(n25036), .B(n25035), .Z(n25037) );
  AND U26585 ( .A(n25038), .B(n25037), .Z(n25073) );
  NANDN U26586 ( .A(n25040), .B(n25039), .Z(n25044) );
  NANDN U26587 ( .A(n25042), .B(n25041), .Z(n25043) );
  AND U26588 ( .A(n25044), .B(n25043), .Z(n25071) );
  NAND U26589 ( .A(n42143), .B(n25045), .Z(n25047) );
  XNOR U26590 ( .A(a[561]), .B(n4152), .Z(n25082) );
  NAND U26591 ( .A(n42144), .B(n25082), .Z(n25046) );
  AND U26592 ( .A(n25047), .B(n25046), .Z(n25097) );
  XOR U26593 ( .A(a[565]), .B(n42012), .Z(n25085) );
  XNOR U26594 ( .A(n25097), .B(n25096), .Z(n25099) );
  AND U26595 ( .A(b[0]), .B(a[567]), .Z(n25049) );
  XOR U26596 ( .A(b[1]), .B(n25049), .Z(n25051) );
  NANDN U26597 ( .A(b[0]), .B(a[566]), .Z(n25050) );
  AND U26598 ( .A(n25051), .B(n25050), .Z(n25092) );
  XOR U26599 ( .A(a[563]), .B(n42085), .Z(n25089) );
  AND U26600 ( .A(a[559]), .B(b[7]), .Z(n25090) );
  XOR U26601 ( .A(n25091), .B(n25090), .Z(n25093) );
  XNOR U26602 ( .A(n25092), .B(n25093), .Z(n25098) );
  XOR U26603 ( .A(n25099), .B(n25098), .Z(n25077) );
  NANDN U26604 ( .A(n25054), .B(n25053), .Z(n25058) );
  NANDN U26605 ( .A(n25056), .B(n25055), .Z(n25057) );
  AND U26606 ( .A(n25058), .B(n25057), .Z(n25076) );
  XNOR U26607 ( .A(n25077), .B(n25076), .Z(n25078) );
  NANDN U26608 ( .A(n25060), .B(n25059), .Z(n25064) );
  NAND U26609 ( .A(n25062), .B(n25061), .Z(n25063) );
  NAND U26610 ( .A(n25064), .B(n25063), .Z(n25079) );
  XNOR U26611 ( .A(n25078), .B(n25079), .Z(n25070) );
  XNOR U26612 ( .A(n25071), .B(n25070), .Z(n25072) );
  XNOR U26613 ( .A(n25073), .B(n25072), .Z(n25102) );
  XNOR U26614 ( .A(sreg[1583]), .B(n25102), .Z(n25104) );
  NANDN U26615 ( .A(sreg[1582]), .B(n25065), .Z(n25069) );
  NAND U26616 ( .A(n25067), .B(n25066), .Z(n25068) );
  NAND U26617 ( .A(n25069), .B(n25068), .Z(n25103) );
  XNOR U26618 ( .A(n25104), .B(n25103), .Z(c[1583]) );
  NANDN U26619 ( .A(n25071), .B(n25070), .Z(n25075) );
  NANDN U26620 ( .A(n25073), .B(n25072), .Z(n25074) );
  AND U26621 ( .A(n25075), .B(n25074), .Z(n25110) );
  NANDN U26622 ( .A(n25077), .B(n25076), .Z(n25081) );
  NANDN U26623 ( .A(n25079), .B(n25078), .Z(n25080) );
  AND U26624 ( .A(n25081), .B(n25080), .Z(n25108) );
  NAND U26625 ( .A(n42143), .B(n25082), .Z(n25084) );
  XNOR U26626 ( .A(a[562]), .B(n4152), .Z(n25119) );
  NAND U26627 ( .A(n42144), .B(n25119), .Z(n25083) );
  AND U26628 ( .A(n25084), .B(n25083), .Z(n25134) );
  XOR U26629 ( .A(a[566]), .B(n42012), .Z(n25122) );
  XNOR U26630 ( .A(n25134), .B(n25133), .Z(n25136) );
  AND U26631 ( .A(a[568]), .B(b[0]), .Z(n25086) );
  XNOR U26632 ( .A(n25086), .B(n4071), .Z(n25088) );
  NANDN U26633 ( .A(b[0]), .B(a[567]), .Z(n25087) );
  NAND U26634 ( .A(n25088), .B(n25087), .Z(n25130) );
  XOR U26635 ( .A(a[564]), .B(n42085), .Z(n25126) );
  AND U26636 ( .A(a[560]), .B(b[7]), .Z(n25127) );
  XNOR U26637 ( .A(n25128), .B(n25127), .Z(n25129) );
  XNOR U26638 ( .A(n25130), .B(n25129), .Z(n25135) );
  XOR U26639 ( .A(n25136), .B(n25135), .Z(n25114) );
  NANDN U26640 ( .A(n25091), .B(n25090), .Z(n25095) );
  NANDN U26641 ( .A(n25093), .B(n25092), .Z(n25094) );
  AND U26642 ( .A(n25095), .B(n25094), .Z(n25113) );
  XNOR U26643 ( .A(n25114), .B(n25113), .Z(n25115) );
  NANDN U26644 ( .A(n25097), .B(n25096), .Z(n25101) );
  NAND U26645 ( .A(n25099), .B(n25098), .Z(n25100) );
  NAND U26646 ( .A(n25101), .B(n25100), .Z(n25116) );
  XNOR U26647 ( .A(n25115), .B(n25116), .Z(n25107) );
  XNOR U26648 ( .A(n25108), .B(n25107), .Z(n25109) );
  XNOR U26649 ( .A(n25110), .B(n25109), .Z(n25139) );
  XNOR U26650 ( .A(sreg[1584]), .B(n25139), .Z(n25141) );
  NANDN U26651 ( .A(sreg[1583]), .B(n25102), .Z(n25106) );
  NAND U26652 ( .A(n25104), .B(n25103), .Z(n25105) );
  NAND U26653 ( .A(n25106), .B(n25105), .Z(n25140) );
  XNOR U26654 ( .A(n25141), .B(n25140), .Z(c[1584]) );
  NANDN U26655 ( .A(n25108), .B(n25107), .Z(n25112) );
  NANDN U26656 ( .A(n25110), .B(n25109), .Z(n25111) );
  AND U26657 ( .A(n25112), .B(n25111), .Z(n25147) );
  NANDN U26658 ( .A(n25114), .B(n25113), .Z(n25118) );
  NANDN U26659 ( .A(n25116), .B(n25115), .Z(n25117) );
  AND U26660 ( .A(n25118), .B(n25117), .Z(n25145) );
  NAND U26661 ( .A(n42143), .B(n25119), .Z(n25121) );
  XNOR U26662 ( .A(a[563]), .B(n4152), .Z(n25156) );
  NAND U26663 ( .A(n42144), .B(n25156), .Z(n25120) );
  AND U26664 ( .A(n25121), .B(n25120), .Z(n25171) );
  XOR U26665 ( .A(a[567]), .B(n42012), .Z(n25159) );
  XNOR U26666 ( .A(n25171), .B(n25170), .Z(n25173) );
  AND U26667 ( .A(a[569]), .B(b[0]), .Z(n25123) );
  XNOR U26668 ( .A(n25123), .B(n4071), .Z(n25125) );
  NANDN U26669 ( .A(b[0]), .B(a[568]), .Z(n25124) );
  NAND U26670 ( .A(n25125), .B(n25124), .Z(n25167) );
  XOR U26671 ( .A(a[565]), .B(n42085), .Z(n25163) );
  AND U26672 ( .A(a[561]), .B(b[7]), .Z(n25164) );
  XNOR U26673 ( .A(n25165), .B(n25164), .Z(n25166) );
  XNOR U26674 ( .A(n25167), .B(n25166), .Z(n25172) );
  XOR U26675 ( .A(n25173), .B(n25172), .Z(n25151) );
  NANDN U26676 ( .A(n25128), .B(n25127), .Z(n25132) );
  NANDN U26677 ( .A(n25130), .B(n25129), .Z(n25131) );
  AND U26678 ( .A(n25132), .B(n25131), .Z(n25150) );
  XNOR U26679 ( .A(n25151), .B(n25150), .Z(n25152) );
  NANDN U26680 ( .A(n25134), .B(n25133), .Z(n25138) );
  NAND U26681 ( .A(n25136), .B(n25135), .Z(n25137) );
  NAND U26682 ( .A(n25138), .B(n25137), .Z(n25153) );
  XNOR U26683 ( .A(n25152), .B(n25153), .Z(n25144) );
  XNOR U26684 ( .A(n25145), .B(n25144), .Z(n25146) );
  XNOR U26685 ( .A(n25147), .B(n25146), .Z(n25176) );
  XNOR U26686 ( .A(sreg[1585]), .B(n25176), .Z(n25178) );
  NANDN U26687 ( .A(sreg[1584]), .B(n25139), .Z(n25143) );
  NAND U26688 ( .A(n25141), .B(n25140), .Z(n25142) );
  NAND U26689 ( .A(n25143), .B(n25142), .Z(n25177) );
  XNOR U26690 ( .A(n25178), .B(n25177), .Z(c[1585]) );
  NANDN U26691 ( .A(n25145), .B(n25144), .Z(n25149) );
  NANDN U26692 ( .A(n25147), .B(n25146), .Z(n25148) );
  AND U26693 ( .A(n25149), .B(n25148), .Z(n25184) );
  NANDN U26694 ( .A(n25151), .B(n25150), .Z(n25155) );
  NANDN U26695 ( .A(n25153), .B(n25152), .Z(n25154) );
  AND U26696 ( .A(n25155), .B(n25154), .Z(n25182) );
  NAND U26697 ( .A(n42143), .B(n25156), .Z(n25158) );
  XNOR U26698 ( .A(a[564]), .B(n4152), .Z(n25193) );
  NAND U26699 ( .A(n42144), .B(n25193), .Z(n25157) );
  AND U26700 ( .A(n25158), .B(n25157), .Z(n25208) );
  XOR U26701 ( .A(a[568]), .B(n42012), .Z(n25196) );
  XNOR U26702 ( .A(n25208), .B(n25207), .Z(n25210) );
  AND U26703 ( .A(a[570]), .B(b[0]), .Z(n25160) );
  XNOR U26704 ( .A(n25160), .B(n4071), .Z(n25162) );
  NANDN U26705 ( .A(b[0]), .B(a[569]), .Z(n25161) );
  NAND U26706 ( .A(n25162), .B(n25161), .Z(n25204) );
  XOR U26707 ( .A(a[566]), .B(n42085), .Z(n25200) );
  AND U26708 ( .A(a[562]), .B(b[7]), .Z(n25201) );
  XNOR U26709 ( .A(n25202), .B(n25201), .Z(n25203) );
  XNOR U26710 ( .A(n25204), .B(n25203), .Z(n25209) );
  XOR U26711 ( .A(n25210), .B(n25209), .Z(n25188) );
  NANDN U26712 ( .A(n25165), .B(n25164), .Z(n25169) );
  NANDN U26713 ( .A(n25167), .B(n25166), .Z(n25168) );
  AND U26714 ( .A(n25169), .B(n25168), .Z(n25187) );
  XNOR U26715 ( .A(n25188), .B(n25187), .Z(n25189) );
  NANDN U26716 ( .A(n25171), .B(n25170), .Z(n25175) );
  NAND U26717 ( .A(n25173), .B(n25172), .Z(n25174) );
  NAND U26718 ( .A(n25175), .B(n25174), .Z(n25190) );
  XNOR U26719 ( .A(n25189), .B(n25190), .Z(n25181) );
  XNOR U26720 ( .A(n25182), .B(n25181), .Z(n25183) );
  XNOR U26721 ( .A(n25184), .B(n25183), .Z(n25213) );
  XNOR U26722 ( .A(sreg[1586]), .B(n25213), .Z(n25215) );
  NANDN U26723 ( .A(sreg[1585]), .B(n25176), .Z(n25180) );
  NAND U26724 ( .A(n25178), .B(n25177), .Z(n25179) );
  NAND U26725 ( .A(n25180), .B(n25179), .Z(n25214) );
  XNOR U26726 ( .A(n25215), .B(n25214), .Z(c[1586]) );
  NANDN U26727 ( .A(n25182), .B(n25181), .Z(n25186) );
  NANDN U26728 ( .A(n25184), .B(n25183), .Z(n25185) );
  AND U26729 ( .A(n25186), .B(n25185), .Z(n25221) );
  NANDN U26730 ( .A(n25188), .B(n25187), .Z(n25192) );
  NANDN U26731 ( .A(n25190), .B(n25189), .Z(n25191) );
  AND U26732 ( .A(n25192), .B(n25191), .Z(n25219) );
  NAND U26733 ( .A(n42143), .B(n25193), .Z(n25195) );
  XNOR U26734 ( .A(a[565]), .B(n4152), .Z(n25230) );
  NAND U26735 ( .A(n42144), .B(n25230), .Z(n25194) );
  AND U26736 ( .A(n25195), .B(n25194), .Z(n25245) );
  XOR U26737 ( .A(a[569]), .B(n42012), .Z(n25233) );
  XNOR U26738 ( .A(n25245), .B(n25244), .Z(n25247) );
  AND U26739 ( .A(a[571]), .B(b[0]), .Z(n25197) );
  XNOR U26740 ( .A(n25197), .B(n4071), .Z(n25199) );
  NANDN U26741 ( .A(b[0]), .B(a[570]), .Z(n25198) );
  NAND U26742 ( .A(n25199), .B(n25198), .Z(n25241) );
  XOR U26743 ( .A(a[567]), .B(n42085), .Z(n25234) );
  AND U26744 ( .A(a[563]), .B(b[7]), .Z(n25238) );
  XNOR U26745 ( .A(n25239), .B(n25238), .Z(n25240) );
  XNOR U26746 ( .A(n25241), .B(n25240), .Z(n25246) );
  XOR U26747 ( .A(n25247), .B(n25246), .Z(n25225) );
  NANDN U26748 ( .A(n25202), .B(n25201), .Z(n25206) );
  NANDN U26749 ( .A(n25204), .B(n25203), .Z(n25205) );
  AND U26750 ( .A(n25206), .B(n25205), .Z(n25224) );
  XNOR U26751 ( .A(n25225), .B(n25224), .Z(n25226) );
  NANDN U26752 ( .A(n25208), .B(n25207), .Z(n25212) );
  NAND U26753 ( .A(n25210), .B(n25209), .Z(n25211) );
  NAND U26754 ( .A(n25212), .B(n25211), .Z(n25227) );
  XNOR U26755 ( .A(n25226), .B(n25227), .Z(n25218) );
  XNOR U26756 ( .A(n25219), .B(n25218), .Z(n25220) );
  XNOR U26757 ( .A(n25221), .B(n25220), .Z(n25250) );
  XNOR U26758 ( .A(sreg[1587]), .B(n25250), .Z(n25252) );
  NANDN U26759 ( .A(sreg[1586]), .B(n25213), .Z(n25217) );
  NAND U26760 ( .A(n25215), .B(n25214), .Z(n25216) );
  NAND U26761 ( .A(n25217), .B(n25216), .Z(n25251) );
  XNOR U26762 ( .A(n25252), .B(n25251), .Z(c[1587]) );
  NANDN U26763 ( .A(n25219), .B(n25218), .Z(n25223) );
  NANDN U26764 ( .A(n25221), .B(n25220), .Z(n25222) );
  AND U26765 ( .A(n25223), .B(n25222), .Z(n25258) );
  NANDN U26766 ( .A(n25225), .B(n25224), .Z(n25229) );
  NANDN U26767 ( .A(n25227), .B(n25226), .Z(n25228) );
  AND U26768 ( .A(n25229), .B(n25228), .Z(n25256) );
  NAND U26769 ( .A(n42143), .B(n25230), .Z(n25232) );
  XNOR U26770 ( .A(a[566]), .B(n4152), .Z(n25267) );
  NAND U26771 ( .A(n42144), .B(n25267), .Z(n25231) );
  AND U26772 ( .A(n25232), .B(n25231), .Z(n25282) );
  XOR U26773 ( .A(a[570]), .B(n42012), .Z(n25270) );
  XNOR U26774 ( .A(n25282), .B(n25281), .Z(n25284) );
  XOR U26775 ( .A(a[568]), .B(n42085), .Z(n25271) );
  AND U26776 ( .A(a[564]), .B(b[7]), .Z(n25275) );
  XNOR U26777 ( .A(n25276), .B(n25275), .Z(n25277) );
  AND U26778 ( .A(a[572]), .B(b[0]), .Z(n25235) );
  XNOR U26779 ( .A(n25235), .B(n4071), .Z(n25237) );
  NANDN U26780 ( .A(b[0]), .B(a[571]), .Z(n25236) );
  NAND U26781 ( .A(n25237), .B(n25236), .Z(n25278) );
  XNOR U26782 ( .A(n25277), .B(n25278), .Z(n25283) );
  XOR U26783 ( .A(n25284), .B(n25283), .Z(n25262) );
  NANDN U26784 ( .A(n25239), .B(n25238), .Z(n25243) );
  NANDN U26785 ( .A(n25241), .B(n25240), .Z(n25242) );
  AND U26786 ( .A(n25243), .B(n25242), .Z(n25261) );
  XNOR U26787 ( .A(n25262), .B(n25261), .Z(n25263) );
  NANDN U26788 ( .A(n25245), .B(n25244), .Z(n25249) );
  NAND U26789 ( .A(n25247), .B(n25246), .Z(n25248) );
  NAND U26790 ( .A(n25249), .B(n25248), .Z(n25264) );
  XNOR U26791 ( .A(n25263), .B(n25264), .Z(n25255) );
  XNOR U26792 ( .A(n25256), .B(n25255), .Z(n25257) );
  XNOR U26793 ( .A(n25258), .B(n25257), .Z(n25287) );
  XNOR U26794 ( .A(sreg[1588]), .B(n25287), .Z(n25289) );
  NANDN U26795 ( .A(sreg[1587]), .B(n25250), .Z(n25254) );
  NAND U26796 ( .A(n25252), .B(n25251), .Z(n25253) );
  NAND U26797 ( .A(n25254), .B(n25253), .Z(n25288) );
  XNOR U26798 ( .A(n25289), .B(n25288), .Z(c[1588]) );
  NANDN U26799 ( .A(n25256), .B(n25255), .Z(n25260) );
  NANDN U26800 ( .A(n25258), .B(n25257), .Z(n25259) );
  AND U26801 ( .A(n25260), .B(n25259), .Z(n25295) );
  NANDN U26802 ( .A(n25262), .B(n25261), .Z(n25266) );
  NANDN U26803 ( .A(n25264), .B(n25263), .Z(n25265) );
  AND U26804 ( .A(n25266), .B(n25265), .Z(n25293) );
  NAND U26805 ( .A(n42143), .B(n25267), .Z(n25269) );
  XNOR U26806 ( .A(a[567]), .B(n4152), .Z(n25304) );
  NAND U26807 ( .A(n42144), .B(n25304), .Z(n25268) );
  AND U26808 ( .A(n25269), .B(n25268), .Z(n25319) );
  XOR U26809 ( .A(a[571]), .B(n42012), .Z(n25307) );
  XNOR U26810 ( .A(n25319), .B(n25318), .Z(n25321) );
  XOR U26811 ( .A(a[569]), .B(n42085), .Z(n25311) );
  AND U26812 ( .A(a[565]), .B(b[7]), .Z(n25312) );
  XNOR U26813 ( .A(n25313), .B(n25312), .Z(n25314) );
  AND U26814 ( .A(a[573]), .B(b[0]), .Z(n25272) );
  XNOR U26815 ( .A(n25272), .B(n4071), .Z(n25274) );
  NANDN U26816 ( .A(b[0]), .B(a[572]), .Z(n25273) );
  NAND U26817 ( .A(n25274), .B(n25273), .Z(n25315) );
  XNOR U26818 ( .A(n25314), .B(n25315), .Z(n25320) );
  XOR U26819 ( .A(n25321), .B(n25320), .Z(n25299) );
  NANDN U26820 ( .A(n25276), .B(n25275), .Z(n25280) );
  NANDN U26821 ( .A(n25278), .B(n25277), .Z(n25279) );
  AND U26822 ( .A(n25280), .B(n25279), .Z(n25298) );
  XNOR U26823 ( .A(n25299), .B(n25298), .Z(n25300) );
  NANDN U26824 ( .A(n25282), .B(n25281), .Z(n25286) );
  NAND U26825 ( .A(n25284), .B(n25283), .Z(n25285) );
  NAND U26826 ( .A(n25286), .B(n25285), .Z(n25301) );
  XNOR U26827 ( .A(n25300), .B(n25301), .Z(n25292) );
  XNOR U26828 ( .A(n25293), .B(n25292), .Z(n25294) );
  XNOR U26829 ( .A(n25295), .B(n25294), .Z(n25324) );
  XNOR U26830 ( .A(sreg[1589]), .B(n25324), .Z(n25326) );
  NANDN U26831 ( .A(sreg[1588]), .B(n25287), .Z(n25291) );
  NAND U26832 ( .A(n25289), .B(n25288), .Z(n25290) );
  NAND U26833 ( .A(n25291), .B(n25290), .Z(n25325) );
  XNOR U26834 ( .A(n25326), .B(n25325), .Z(c[1589]) );
  NANDN U26835 ( .A(n25293), .B(n25292), .Z(n25297) );
  NANDN U26836 ( .A(n25295), .B(n25294), .Z(n25296) );
  AND U26837 ( .A(n25297), .B(n25296), .Z(n25332) );
  NANDN U26838 ( .A(n25299), .B(n25298), .Z(n25303) );
  NANDN U26839 ( .A(n25301), .B(n25300), .Z(n25302) );
  AND U26840 ( .A(n25303), .B(n25302), .Z(n25330) );
  NAND U26841 ( .A(n42143), .B(n25304), .Z(n25306) );
  XNOR U26842 ( .A(a[568]), .B(n4153), .Z(n25341) );
  NAND U26843 ( .A(n42144), .B(n25341), .Z(n25305) );
  AND U26844 ( .A(n25306), .B(n25305), .Z(n25356) );
  XOR U26845 ( .A(a[572]), .B(n42012), .Z(n25344) );
  XNOR U26846 ( .A(n25356), .B(n25355), .Z(n25358) );
  AND U26847 ( .A(a[574]), .B(b[0]), .Z(n25308) );
  XNOR U26848 ( .A(n25308), .B(n4071), .Z(n25310) );
  NANDN U26849 ( .A(b[0]), .B(a[573]), .Z(n25309) );
  NAND U26850 ( .A(n25310), .B(n25309), .Z(n25352) );
  XOR U26851 ( .A(a[570]), .B(n42085), .Z(n25348) );
  AND U26852 ( .A(a[566]), .B(b[7]), .Z(n25349) );
  XNOR U26853 ( .A(n25350), .B(n25349), .Z(n25351) );
  XNOR U26854 ( .A(n25352), .B(n25351), .Z(n25357) );
  XOR U26855 ( .A(n25358), .B(n25357), .Z(n25336) );
  NANDN U26856 ( .A(n25313), .B(n25312), .Z(n25317) );
  NANDN U26857 ( .A(n25315), .B(n25314), .Z(n25316) );
  AND U26858 ( .A(n25317), .B(n25316), .Z(n25335) );
  XNOR U26859 ( .A(n25336), .B(n25335), .Z(n25337) );
  NANDN U26860 ( .A(n25319), .B(n25318), .Z(n25323) );
  NAND U26861 ( .A(n25321), .B(n25320), .Z(n25322) );
  NAND U26862 ( .A(n25323), .B(n25322), .Z(n25338) );
  XNOR U26863 ( .A(n25337), .B(n25338), .Z(n25329) );
  XNOR U26864 ( .A(n25330), .B(n25329), .Z(n25331) );
  XNOR U26865 ( .A(n25332), .B(n25331), .Z(n25361) );
  XNOR U26866 ( .A(sreg[1590]), .B(n25361), .Z(n25363) );
  NANDN U26867 ( .A(sreg[1589]), .B(n25324), .Z(n25328) );
  NAND U26868 ( .A(n25326), .B(n25325), .Z(n25327) );
  NAND U26869 ( .A(n25328), .B(n25327), .Z(n25362) );
  XNOR U26870 ( .A(n25363), .B(n25362), .Z(c[1590]) );
  NANDN U26871 ( .A(n25330), .B(n25329), .Z(n25334) );
  NANDN U26872 ( .A(n25332), .B(n25331), .Z(n25333) );
  AND U26873 ( .A(n25334), .B(n25333), .Z(n25369) );
  NANDN U26874 ( .A(n25336), .B(n25335), .Z(n25340) );
  NANDN U26875 ( .A(n25338), .B(n25337), .Z(n25339) );
  AND U26876 ( .A(n25340), .B(n25339), .Z(n25367) );
  NAND U26877 ( .A(n42143), .B(n25341), .Z(n25343) );
  XNOR U26878 ( .A(a[569]), .B(n4153), .Z(n25378) );
  NAND U26879 ( .A(n42144), .B(n25378), .Z(n25342) );
  AND U26880 ( .A(n25343), .B(n25342), .Z(n25393) );
  XOR U26881 ( .A(a[573]), .B(n42012), .Z(n25381) );
  XNOR U26882 ( .A(n25393), .B(n25392), .Z(n25395) );
  AND U26883 ( .A(a[575]), .B(b[0]), .Z(n25345) );
  XNOR U26884 ( .A(n25345), .B(n4071), .Z(n25347) );
  NANDN U26885 ( .A(b[0]), .B(a[574]), .Z(n25346) );
  NAND U26886 ( .A(n25347), .B(n25346), .Z(n25389) );
  XOR U26887 ( .A(a[571]), .B(n42085), .Z(n25382) );
  AND U26888 ( .A(a[567]), .B(b[7]), .Z(n25386) );
  XNOR U26889 ( .A(n25387), .B(n25386), .Z(n25388) );
  XNOR U26890 ( .A(n25389), .B(n25388), .Z(n25394) );
  XOR U26891 ( .A(n25395), .B(n25394), .Z(n25373) );
  NANDN U26892 ( .A(n25350), .B(n25349), .Z(n25354) );
  NANDN U26893 ( .A(n25352), .B(n25351), .Z(n25353) );
  AND U26894 ( .A(n25354), .B(n25353), .Z(n25372) );
  XNOR U26895 ( .A(n25373), .B(n25372), .Z(n25374) );
  NANDN U26896 ( .A(n25356), .B(n25355), .Z(n25360) );
  NAND U26897 ( .A(n25358), .B(n25357), .Z(n25359) );
  NAND U26898 ( .A(n25360), .B(n25359), .Z(n25375) );
  XNOR U26899 ( .A(n25374), .B(n25375), .Z(n25366) );
  XNOR U26900 ( .A(n25367), .B(n25366), .Z(n25368) );
  XNOR U26901 ( .A(n25369), .B(n25368), .Z(n25398) );
  XNOR U26902 ( .A(sreg[1591]), .B(n25398), .Z(n25400) );
  NANDN U26903 ( .A(sreg[1590]), .B(n25361), .Z(n25365) );
  NAND U26904 ( .A(n25363), .B(n25362), .Z(n25364) );
  NAND U26905 ( .A(n25365), .B(n25364), .Z(n25399) );
  XNOR U26906 ( .A(n25400), .B(n25399), .Z(c[1591]) );
  NANDN U26907 ( .A(n25367), .B(n25366), .Z(n25371) );
  NANDN U26908 ( .A(n25369), .B(n25368), .Z(n25370) );
  AND U26909 ( .A(n25371), .B(n25370), .Z(n25406) );
  NANDN U26910 ( .A(n25373), .B(n25372), .Z(n25377) );
  NANDN U26911 ( .A(n25375), .B(n25374), .Z(n25376) );
  AND U26912 ( .A(n25377), .B(n25376), .Z(n25404) );
  NAND U26913 ( .A(n42143), .B(n25378), .Z(n25380) );
  XNOR U26914 ( .A(a[570]), .B(n4153), .Z(n25415) );
  NAND U26915 ( .A(n42144), .B(n25415), .Z(n25379) );
  AND U26916 ( .A(n25380), .B(n25379), .Z(n25430) );
  XOR U26917 ( .A(a[574]), .B(n42012), .Z(n25418) );
  XNOR U26918 ( .A(n25430), .B(n25429), .Z(n25432) );
  XOR U26919 ( .A(a[572]), .B(n42085), .Z(n25422) );
  AND U26920 ( .A(a[568]), .B(b[7]), .Z(n25423) );
  XNOR U26921 ( .A(n25424), .B(n25423), .Z(n25425) );
  AND U26922 ( .A(a[576]), .B(b[0]), .Z(n25383) );
  XNOR U26923 ( .A(n25383), .B(n4071), .Z(n25385) );
  NANDN U26924 ( .A(b[0]), .B(a[575]), .Z(n25384) );
  NAND U26925 ( .A(n25385), .B(n25384), .Z(n25426) );
  XNOR U26926 ( .A(n25425), .B(n25426), .Z(n25431) );
  XOR U26927 ( .A(n25432), .B(n25431), .Z(n25410) );
  NANDN U26928 ( .A(n25387), .B(n25386), .Z(n25391) );
  NANDN U26929 ( .A(n25389), .B(n25388), .Z(n25390) );
  AND U26930 ( .A(n25391), .B(n25390), .Z(n25409) );
  XNOR U26931 ( .A(n25410), .B(n25409), .Z(n25411) );
  NANDN U26932 ( .A(n25393), .B(n25392), .Z(n25397) );
  NAND U26933 ( .A(n25395), .B(n25394), .Z(n25396) );
  NAND U26934 ( .A(n25397), .B(n25396), .Z(n25412) );
  XNOR U26935 ( .A(n25411), .B(n25412), .Z(n25403) );
  XNOR U26936 ( .A(n25404), .B(n25403), .Z(n25405) );
  XNOR U26937 ( .A(n25406), .B(n25405), .Z(n25435) );
  XNOR U26938 ( .A(sreg[1592]), .B(n25435), .Z(n25437) );
  NANDN U26939 ( .A(sreg[1591]), .B(n25398), .Z(n25402) );
  NAND U26940 ( .A(n25400), .B(n25399), .Z(n25401) );
  NAND U26941 ( .A(n25402), .B(n25401), .Z(n25436) );
  XNOR U26942 ( .A(n25437), .B(n25436), .Z(c[1592]) );
  NANDN U26943 ( .A(n25404), .B(n25403), .Z(n25408) );
  NANDN U26944 ( .A(n25406), .B(n25405), .Z(n25407) );
  AND U26945 ( .A(n25408), .B(n25407), .Z(n25443) );
  NANDN U26946 ( .A(n25410), .B(n25409), .Z(n25414) );
  NANDN U26947 ( .A(n25412), .B(n25411), .Z(n25413) );
  AND U26948 ( .A(n25414), .B(n25413), .Z(n25441) );
  NAND U26949 ( .A(n42143), .B(n25415), .Z(n25417) );
  XNOR U26950 ( .A(a[571]), .B(n4153), .Z(n25452) );
  NAND U26951 ( .A(n42144), .B(n25452), .Z(n25416) );
  AND U26952 ( .A(n25417), .B(n25416), .Z(n25467) );
  XOR U26953 ( .A(a[575]), .B(n42012), .Z(n25455) );
  XNOR U26954 ( .A(n25467), .B(n25466), .Z(n25469) );
  AND U26955 ( .A(a[577]), .B(b[0]), .Z(n25419) );
  XNOR U26956 ( .A(n25419), .B(n4071), .Z(n25421) );
  NANDN U26957 ( .A(b[0]), .B(a[576]), .Z(n25420) );
  NAND U26958 ( .A(n25421), .B(n25420), .Z(n25463) );
  XOR U26959 ( .A(a[573]), .B(n42085), .Z(n25459) );
  AND U26960 ( .A(a[569]), .B(b[7]), .Z(n25460) );
  XNOR U26961 ( .A(n25461), .B(n25460), .Z(n25462) );
  XNOR U26962 ( .A(n25463), .B(n25462), .Z(n25468) );
  XOR U26963 ( .A(n25469), .B(n25468), .Z(n25447) );
  NANDN U26964 ( .A(n25424), .B(n25423), .Z(n25428) );
  NANDN U26965 ( .A(n25426), .B(n25425), .Z(n25427) );
  AND U26966 ( .A(n25428), .B(n25427), .Z(n25446) );
  XNOR U26967 ( .A(n25447), .B(n25446), .Z(n25448) );
  NANDN U26968 ( .A(n25430), .B(n25429), .Z(n25434) );
  NAND U26969 ( .A(n25432), .B(n25431), .Z(n25433) );
  NAND U26970 ( .A(n25434), .B(n25433), .Z(n25449) );
  XNOR U26971 ( .A(n25448), .B(n25449), .Z(n25440) );
  XNOR U26972 ( .A(n25441), .B(n25440), .Z(n25442) );
  XNOR U26973 ( .A(n25443), .B(n25442), .Z(n25472) );
  XNOR U26974 ( .A(sreg[1593]), .B(n25472), .Z(n25474) );
  NANDN U26975 ( .A(sreg[1592]), .B(n25435), .Z(n25439) );
  NAND U26976 ( .A(n25437), .B(n25436), .Z(n25438) );
  NAND U26977 ( .A(n25439), .B(n25438), .Z(n25473) );
  XNOR U26978 ( .A(n25474), .B(n25473), .Z(c[1593]) );
  NANDN U26979 ( .A(n25441), .B(n25440), .Z(n25445) );
  NANDN U26980 ( .A(n25443), .B(n25442), .Z(n25444) );
  AND U26981 ( .A(n25445), .B(n25444), .Z(n25480) );
  NANDN U26982 ( .A(n25447), .B(n25446), .Z(n25451) );
  NANDN U26983 ( .A(n25449), .B(n25448), .Z(n25450) );
  AND U26984 ( .A(n25451), .B(n25450), .Z(n25478) );
  NAND U26985 ( .A(n42143), .B(n25452), .Z(n25454) );
  XNOR U26986 ( .A(a[572]), .B(n4153), .Z(n25489) );
  NAND U26987 ( .A(n42144), .B(n25489), .Z(n25453) );
  AND U26988 ( .A(n25454), .B(n25453), .Z(n25504) );
  XOR U26989 ( .A(a[576]), .B(n42012), .Z(n25492) );
  XNOR U26990 ( .A(n25504), .B(n25503), .Z(n25506) );
  AND U26991 ( .A(a[578]), .B(b[0]), .Z(n25456) );
  XNOR U26992 ( .A(n25456), .B(n4071), .Z(n25458) );
  NANDN U26993 ( .A(b[0]), .B(a[577]), .Z(n25457) );
  NAND U26994 ( .A(n25458), .B(n25457), .Z(n25500) );
  XOR U26995 ( .A(a[574]), .B(n42085), .Z(n25493) );
  AND U26996 ( .A(a[570]), .B(b[7]), .Z(n25497) );
  XNOR U26997 ( .A(n25498), .B(n25497), .Z(n25499) );
  XNOR U26998 ( .A(n25500), .B(n25499), .Z(n25505) );
  XOR U26999 ( .A(n25506), .B(n25505), .Z(n25484) );
  NANDN U27000 ( .A(n25461), .B(n25460), .Z(n25465) );
  NANDN U27001 ( .A(n25463), .B(n25462), .Z(n25464) );
  AND U27002 ( .A(n25465), .B(n25464), .Z(n25483) );
  XNOR U27003 ( .A(n25484), .B(n25483), .Z(n25485) );
  NANDN U27004 ( .A(n25467), .B(n25466), .Z(n25471) );
  NAND U27005 ( .A(n25469), .B(n25468), .Z(n25470) );
  NAND U27006 ( .A(n25471), .B(n25470), .Z(n25486) );
  XNOR U27007 ( .A(n25485), .B(n25486), .Z(n25477) );
  XNOR U27008 ( .A(n25478), .B(n25477), .Z(n25479) );
  XNOR U27009 ( .A(n25480), .B(n25479), .Z(n25509) );
  XNOR U27010 ( .A(sreg[1594]), .B(n25509), .Z(n25511) );
  NANDN U27011 ( .A(sreg[1593]), .B(n25472), .Z(n25476) );
  NAND U27012 ( .A(n25474), .B(n25473), .Z(n25475) );
  NAND U27013 ( .A(n25476), .B(n25475), .Z(n25510) );
  XNOR U27014 ( .A(n25511), .B(n25510), .Z(c[1594]) );
  NANDN U27015 ( .A(n25478), .B(n25477), .Z(n25482) );
  NANDN U27016 ( .A(n25480), .B(n25479), .Z(n25481) );
  AND U27017 ( .A(n25482), .B(n25481), .Z(n25517) );
  NANDN U27018 ( .A(n25484), .B(n25483), .Z(n25488) );
  NANDN U27019 ( .A(n25486), .B(n25485), .Z(n25487) );
  AND U27020 ( .A(n25488), .B(n25487), .Z(n25515) );
  NAND U27021 ( .A(n42143), .B(n25489), .Z(n25491) );
  XNOR U27022 ( .A(a[573]), .B(n4153), .Z(n25526) );
  NAND U27023 ( .A(n42144), .B(n25526), .Z(n25490) );
  AND U27024 ( .A(n25491), .B(n25490), .Z(n25541) );
  XOR U27025 ( .A(a[577]), .B(n42012), .Z(n25529) );
  XNOR U27026 ( .A(n25541), .B(n25540), .Z(n25543) );
  XOR U27027 ( .A(a[575]), .B(n42085), .Z(n25530) );
  AND U27028 ( .A(a[571]), .B(b[7]), .Z(n25534) );
  XNOR U27029 ( .A(n25535), .B(n25534), .Z(n25536) );
  AND U27030 ( .A(a[579]), .B(b[0]), .Z(n25494) );
  XNOR U27031 ( .A(n25494), .B(n4071), .Z(n25496) );
  NANDN U27032 ( .A(b[0]), .B(a[578]), .Z(n25495) );
  NAND U27033 ( .A(n25496), .B(n25495), .Z(n25537) );
  XNOR U27034 ( .A(n25536), .B(n25537), .Z(n25542) );
  XOR U27035 ( .A(n25543), .B(n25542), .Z(n25521) );
  NANDN U27036 ( .A(n25498), .B(n25497), .Z(n25502) );
  NANDN U27037 ( .A(n25500), .B(n25499), .Z(n25501) );
  AND U27038 ( .A(n25502), .B(n25501), .Z(n25520) );
  XNOR U27039 ( .A(n25521), .B(n25520), .Z(n25522) );
  NANDN U27040 ( .A(n25504), .B(n25503), .Z(n25508) );
  NAND U27041 ( .A(n25506), .B(n25505), .Z(n25507) );
  NAND U27042 ( .A(n25508), .B(n25507), .Z(n25523) );
  XNOR U27043 ( .A(n25522), .B(n25523), .Z(n25514) );
  XNOR U27044 ( .A(n25515), .B(n25514), .Z(n25516) );
  XNOR U27045 ( .A(n25517), .B(n25516), .Z(n25546) );
  XNOR U27046 ( .A(sreg[1595]), .B(n25546), .Z(n25548) );
  NANDN U27047 ( .A(sreg[1594]), .B(n25509), .Z(n25513) );
  NAND U27048 ( .A(n25511), .B(n25510), .Z(n25512) );
  NAND U27049 ( .A(n25513), .B(n25512), .Z(n25547) );
  XNOR U27050 ( .A(n25548), .B(n25547), .Z(c[1595]) );
  NANDN U27051 ( .A(n25515), .B(n25514), .Z(n25519) );
  NANDN U27052 ( .A(n25517), .B(n25516), .Z(n25518) );
  AND U27053 ( .A(n25519), .B(n25518), .Z(n25554) );
  NANDN U27054 ( .A(n25521), .B(n25520), .Z(n25525) );
  NANDN U27055 ( .A(n25523), .B(n25522), .Z(n25524) );
  AND U27056 ( .A(n25525), .B(n25524), .Z(n25552) );
  NAND U27057 ( .A(n42143), .B(n25526), .Z(n25528) );
  XNOR U27058 ( .A(a[574]), .B(n4153), .Z(n25563) );
  NAND U27059 ( .A(n42144), .B(n25563), .Z(n25527) );
  AND U27060 ( .A(n25528), .B(n25527), .Z(n25578) );
  XOR U27061 ( .A(a[578]), .B(n42012), .Z(n25566) );
  XNOR U27062 ( .A(n25578), .B(n25577), .Z(n25580) );
  XOR U27063 ( .A(a[576]), .B(n42085), .Z(n25567) );
  AND U27064 ( .A(a[572]), .B(b[7]), .Z(n25571) );
  XNOR U27065 ( .A(n25572), .B(n25571), .Z(n25573) );
  AND U27066 ( .A(a[580]), .B(b[0]), .Z(n25531) );
  XNOR U27067 ( .A(n25531), .B(n4071), .Z(n25533) );
  NANDN U27068 ( .A(b[0]), .B(a[579]), .Z(n25532) );
  NAND U27069 ( .A(n25533), .B(n25532), .Z(n25574) );
  XNOR U27070 ( .A(n25573), .B(n25574), .Z(n25579) );
  XOR U27071 ( .A(n25580), .B(n25579), .Z(n25558) );
  NANDN U27072 ( .A(n25535), .B(n25534), .Z(n25539) );
  NANDN U27073 ( .A(n25537), .B(n25536), .Z(n25538) );
  AND U27074 ( .A(n25539), .B(n25538), .Z(n25557) );
  XNOR U27075 ( .A(n25558), .B(n25557), .Z(n25559) );
  NANDN U27076 ( .A(n25541), .B(n25540), .Z(n25545) );
  NAND U27077 ( .A(n25543), .B(n25542), .Z(n25544) );
  NAND U27078 ( .A(n25545), .B(n25544), .Z(n25560) );
  XNOR U27079 ( .A(n25559), .B(n25560), .Z(n25551) );
  XNOR U27080 ( .A(n25552), .B(n25551), .Z(n25553) );
  XNOR U27081 ( .A(n25554), .B(n25553), .Z(n25583) );
  XNOR U27082 ( .A(sreg[1596]), .B(n25583), .Z(n25585) );
  NANDN U27083 ( .A(sreg[1595]), .B(n25546), .Z(n25550) );
  NAND U27084 ( .A(n25548), .B(n25547), .Z(n25549) );
  NAND U27085 ( .A(n25550), .B(n25549), .Z(n25584) );
  XNOR U27086 ( .A(n25585), .B(n25584), .Z(c[1596]) );
  NANDN U27087 ( .A(n25552), .B(n25551), .Z(n25556) );
  NANDN U27088 ( .A(n25554), .B(n25553), .Z(n25555) );
  AND U27089 ( .A(n25556), .B(n25555), .Z(n25591) );
  NANDN U27090 ( .A(n25558), .B(n25557), .Z(n25562) );
  NANDN U27091 ( .A(n25560), .B(n25559), .Z(n25561) );
  AND U27092 ( .A(n25562), .B(n25561), .Z(n25589) );
  NAND U27093 ( .A(n42143), .B(n25563), .Z(n25565) );
  XNOR U27094 ( .A(a[575]), .B(n4154), .Z(n25600) );
  NAND U27095 ( .A(n42144), .B(n25600), .Z(n25564) );
  AND U27096 ( .A(n25565), .B(n25564), .Z(n25615) );
  XOR U27097 ( .A(a[579]), .B(n42012), .Z(n25603) );
  XNOR U27098 ( .A(n25615), .B(n25614), .Z(n25617) );
  XOR U27099 ( .A(a[577]), .B(n42085), .Z(n25604) );
  AND U27100 ( .A(a[573]), .B(b[7]), .Z(n25608) );
  XNOR U27101 ( .A(n25609), .B(n25608), .Z(n25610) );
  AND U27102 ( .A(a[581]), .B(b[0]), .Z(n25568) );
  XNOR U27103 ( .A(n25568), .B(n4071), .Z(n25570) );
  NANDN U27104 ( .A(b[0]), .B(a[580]), .Z(n25569) );
  NAND U27105 ( .A(n25570), .B(n25569), .Z(n25611) );
  XNOR U27106 ( .A(n25610), .B(n25611), .Z(n25616) );
  XOR U27107 ( .A(n25617), .B(n25616), .Z(n25595) );
  NANDN U27108 ( .A(n25572), .B(n25571), .Z(n25576) );
  NANDN U27109 ( .A(n25574), .B(n25573), .Z(n25575) );
  AND U27110 ( .A(n25576), .B(n25575), .Z(n25594) );
  XNOR U27111 ( .A(n25595), .B(n25594), .Z(n25596) );
  NANDN U27112 ( .A(n25578), .B(n25577), .Z(n25582) );
  NAND U27113 ( .A(n25580), .B(n25579), .Z(n25581) );
  NAND U27114 ( .A(n25582), .B(n25581), .Z(n25597) );
  XNOR U27115 ( .A(n25596), .B(n25597), .Z(n25588) );
  XNOR U27116 ( .A(n25589), .B(n25588), .Z(n25590) );
  XNOR U27117 ( .A(n25591), .B(n25590), .Z(n25620) );
  XNOR U27118 ( .A(sreg[1597]), .B(n25620), .Z(n25622) );
  NANDN U27119 ( .A(sreg[1596]), .B(n25583), .Z(n25587) );
  NAND U27120 ( .A(n25585), .B(n25584), .Z(n25586) );
  NAND U27121 ( .A(n25587), .B(n25586), .Z(n25621) );
  XNOR U27122 ( .A(n25622), .B(n25621), .Z(c[1597]) );
  NANDN U27123 ( .A(n25589), .B(n25588), .Z(n25593) );
  NANDN U27124 ( .A(n25591), .B(n25590), .Z(n25592) );
  AND U27125 ( .A(n25593), .B(n25592), .Z(n25628) );
  NANDN U27126 ( .A(n25595), .B(n25594), .Z(n25599) );
  NANDN U27127 ( .A(n25597), .B(n25596), .Z(n25598) );
  AND U27128 ( .A(n25599), .B(n25598), .Z(n25626) );
  NAND U27129 ( .A(n42143), .B(n25600), .Z(n25602) );
  XNOR U27130 ( .A(a[576]), .B(n4154), .Z(n25637) );
  NAND U27131 ( .A(n42144), .B(n25637), .Z(n25601) );
  AND U27132 ( .A(n25602), .B(n25601), .Z(n25652) );
  XOR U27133 ( .A(a[580]), .B(n42012), .Z(n25640) );
  XNOR U27134 ( .A(n25652), .B(n25651), .Z(n25654) );
  XOR U27135 ( .A(a[578]), .B(n42085), .Z(n25644) );
  AND U27136 ( .A(a[574]), .B(b[7]), .Z(n25645) );
  XNOR U27137 ( .A(n25646), .B(n25645), .Z(n25647) );
  AND U27138 ( .A(a[582]), .B(b[0]), .Z(n25605) );
  XNOR U27139 ( .A(n25605), .B(n4071), .Z(n25607) );
  NANDN U27140 ( .A(b[0]), .B(a[581]), .Z(n25606) );
  NAND U27141 ( .A(n25607), .B(n25606), .Z(n25648) );
  XNOR U27142 ( .A(n25647), .B(n25648), .Z(n25653) );
  XOR U27143 ( .A(n25654), .B(n25653), .Z(n25632) );
  NANDN U27144 ( .A(n25609), .B(n25608), .Z(n25613) );
  NANDN U27145 ( .A(n25611), .B(n25610), .Z(n25612) );
  AND U27146 ( .A(n25613), .B(n25612), .Z(n25631) );
  XNOR U27147 ( .A(n25632), .B(n25631), .Z(n25633) );
  NANDN U27148 ( .A(n25615), .B(n25614), .Z(n25619) );
  NAND U27149 ( .A(n25617), .B(n25616), .Z(n25618) );
  NAND U27150 ( .A(n25619), .B(n25618), .Z(n25634) );
  XNOR U27151 ( .A(n25633), .B(n25634), .Z(n25625) );
  XNOR U27152 ( .A(n25626), .B(n25625), .Z(n25627) );
  XNOR U27153 ( .A(n25628), .B(n25627), .Z(n25657) );
  XNOR U27154 ( .A(sreg[1598]), .B(n25657), .Z(n25659) );
  NANDN U27155 ( .A(sreg[1597]), .B(n25620), .Z(n25624) );
  NAND U27156 ( .A(n25622), .B(n25621), .Z(n25623) );
  NAND U27157 ( .A(n25624), .B(n25623), .Z(n25658) );
  XNOR U27158 ( .A(n25659), .B(n25658), .Z(c[1598]) );
  NANDN U27159 ( .A(n25626), .B(n25625), .Z(n25630) );
  NANDN U27160 ( .A(n25628), .B(n25627), .Z(n25629) );
  AND U27161 ( .A(n25630), .B(n25629), .Z(n25665) );
  NANDN U27162 ( .A(n25632), .B(n25631), .Z(n25636) );
  NANDN U27163 ( .A(n25634), .B(n25633), .Z(n25635) );
  AND U27164 ( .A(n25636), .B(n25635), .Z(n25663) );
  NAND U27165 ( .A(n42143), .B(n25637), .Z(n25639) );
  XNOR U27166 ( .A(a[577]), .B(n4154), .Z(n25674) );
  NAND U27167 ( .A(n42144), .B(n25674), .Z(n25638) );
  AND U27168 ( .A(n25639), .B(n25638), .Z(n25689) );
  XOR U27169 ( .A(a[581]), .B(n42012), .Z(n25677) );
  XNOR U27170 ( .A(n25689), .B(n25688), .Z(n25691) );
  AND U27171 ( .A(a[583]), .B(b[0]), .Z(n25641) );
  XNOR U27172 ( .A(n25641), .B(n4071), .Z(n25643) );
  NANDN U27173 ( .A(b[0]), .B(a[582]), .Z(n25642) );
  NAND U27174 ( .A(n25643), .B(n25642), .Z(n25685) );
  XOR U27175 ( .A(a[579]), .B(n42085), .Z(n25681) );
  AND U27176 ( .A(a[575]), .B(b[7]), .Z(n25682) );
  XNOR U27177 ( .A(n25683), .B(n25682), .Z(n25684) );
  XNOR U27178 ( .A(n25685), .B(n25684), .Z(n25690) );
  XOR U27179 ( .A(n25691), .B(n25690), .Z(n25669) );
  NANDN U27180 ( .A(n25646), .B(n25645), .Z(n25650) );
  NANDN U27181 ( .A(n25648), .B(n25647), .Z(n25649) );
  AND U27182 ( .A(n25650), .B(n25649), .Z(n25668) );
  XNOR U27183 ( .A(n25669), .B(n25668), .Z(n25670) );
  NANDN U27184 ( .A(n25652), .B(n25651), .Z(n25656) );
  NAND U27185 ( .A(n25654), .B(n25653), .Z(n25655) );
  NAND U27186 ( .A(n25656), .B(n25655), .Z(n25671) );
  XNOR U27187 ( .A(n25670), .B(n25671), .Z(n25662) );
  XNOR U27188 ( .A(n25663), .B(n25662), .Z(n25664) );
  XNOR U27189 ( .A(n25665), .B(n25664), .Z(n25694) );
  XNOR U27190 ( .A(sreg[1599]), .B(n25694), .Z(n25696) );
  NANDN U27191 ( .A(sreg[1598]), .B(n25657), .Z(n25661) );
  NAND U27192 ( .A(n25659), .B(n25658), .Z(n25660) );
  NAND U27193 ( .A(n25661), .B(n25660), .Z(n25695) );
  XNOR U27194 ( .A(n25696), .B(n25695), .Z(c[1599]) );
  NANDN U27195 ( .A(n25663), .B(n25662), .Z(n25667) );
  NANDN U27196 ( .A(n25665), .B(n25664), .Z(n25666) );
  AND U27197 ( .A(n25667), .B(n25666), .Z(n25702) );
  NANDN U27198 ( .A(n25669), .B(n25668), .Z(n25673) );
  NANDN U27199 ( .A(n25671), .B(n25670), .Z(n25672) );
  AND U27200 ( .A(n25673), .B(n25672), .Z(n25700) );
  NAND U27201 ( .A(n42143), .B(n25674), .Z(n25676) );
  XNOR U27202 ( .A(a[578]), .B(n4154), .Z(n25711) );
  NAND U27203 ( .A(n42144), .B(n25711), .Z(n25675) );
  AND U27204 ( .A(n25676), .B(n25675), .Z(n25726) );
  XOR U27205 ( .A(a[582]), .B(n42012), .Z(n25714) );
  XNOR U27206 ( .A(n25726), .B(n25725), .Z(n25728) );
  AND U27207 ( .A(a[584]), .B(b[0]), .Z(n25678) );
  XNOR U27208 ( .A(n25678), .B(n4071), .Z(n25680) );
  NANDN U27209 ( .A(b[0]), .B(a[583]), .Z(n25679) );
  NAND U27210 ( .A(n25680), .B(n25679), .Z(n25722) );
  XOR U27211 ( .A(a[580]), .B(n42085), .Z(n25718) );
  AND U27212 ( .A(a[576]), .B(b[7]), .Z(n25719) );
  XNOR U27213 ( .A(n25720), .B(n25719), .Z(n25721) );
  XNOR U27214 ( .A(n25722), .B(n25721), .Z(n25727) );
  XOR U27215 ( .A(n25728), .B(n25727), .Z(n25706) );
  NANDN U27216 ( .A(n25683), .B(n25682), .Z(n25687) );
  NANDN U27217 ( .A(n25685), .B(n25684), .Z(n25686) );
  AND U27218 ( .A(n25687), .B(n25686), .Z(n25705) );
  XNOR U27219 ( .A(n25706), .B(n25705), .Z(n25707) );
  NANDN U27220 ( .A(n25689), .B(n25688), .Z(n25693) );
  NAND U27221 ( .A(n25691), .B(n25690), .Z(n25692) );
  NAND U27222 ( .A(n25693), .B(n25692), .Z(n25708) );
  XNOR U27223 ( .A(n25707), .B(n25708), .Z(n25699) );
  XNOR U27224 ( .A(n25700), .B(n25699), .Z(n25701) );
  XNOR U27225 ( .A(n25702), .B(n25701), .Z(n25731) );
  XNOR U27226 ( .A(sreg[1600]), .B(n25731), .Z(n25733) );
  NANDN U27227 ( .A(sreg[1599]), .B(n25694), .Z(n25698) );
  NAND U27228 ( .A(n25696), .B(n25695), .Z(n25697) );
  NAND U27229 ( .A(n25698), .B(n25697), .Z(n25732) );
  XNOR U27230 ( .A(n25733), .B(n25732), .Z(c[1600]) );
  NANDN U27231 ( .A(n25700), .B(n25699), .Z(n25704) );
  NANDN U27232 ( .A(n25702), .B(n25701), .Z(n25703) );
  AND U27233 ( .A(n25704), .B(n25703), .Z(n25739) );
  NANDN U27234 ( .A(n25706), .B(n25705), .Z(n25710) );
  NANDN U27235 ( .A(n25708), .B(n25707), .Z(n25709) );
  AND U27236 ( .A(n25710), .B(n25709), .Z(n25737) );
  NAND U27237 ( .A(n42143), .B(n25711), .Z(n25713) );
  XNOR U27238 ( .A(a[579]), .B(n4154), .Z(n25748) );
  NAND U27239 ( .A(n42144), .B(n25748), .Z(n25712) );
  AND U27240 ( .A(n25713), .B(n25712), .Z(n25763) );
  XOR U27241 ( .A(a[583]), .B(n42012), .Z(n25751) );
  XNOR U27242 ( .A(n25763), .B(n25762), .Z(n25765) );
  AND U27243 ( .A(a[585]), .B(b[0]), .Z(n25715) );
  XNOR U27244 ( .A(n25715), .B(n4071), .Z(n25717) );
  NANDN U27245 ( .A(b[0]), .B(a[584]), .Z(n25716) );
  NAND U27246 ( .A(n25717), .B(n25716), .Z(n25759) );
  XOR U27247 ( .A(a[581]), .B(n42085), .Z(n25755) );
  AND U27248 ( .A(a[577]), .B(b[7]), .Z(n25756) );
  XNOR U27249 ( .A(n25757), .B(n25756), .Z(n25758) );
  XNOR U27250 ( .A(n25759), .B(n25758), .Z(n25764) );
  XOR U27251 ( .A(n25765), .B(n25764), .Z(n25743) );
  NANDN U27252 ( .A(n25720), .B(n25719), .Z(n25724) );
  NANDN U27253 ( .A(n25722), .B(n25721), .Z(n25723) );
  AND U27254 ( .A(n25724), .B(n25723), .Z(n25742) );
  XNOR U27255 ( .A(n25743), .B(n25742), .Z(n25744) );
  NANDN U27256 ( .A(n25726), .B(n25725), .Z(n25730) );
  NAND U27257 ( .A(n25728), .B(n25727), .Z(n25729) );
  NAND U27258 ( .A(n25730), .B(n25729), .Z(n25745) );
  XNOR U27259 ( .A(n25744), .B(n25745), .Z(n25736) );
  XNOR U27260 ( .A(n25737), .B(n25736), .Z(n25738) );
  XNOR U27261 ( .A(n25739), .B(n25738), .Z(n25768) );
  XNOR U27262 ( .A(sreg[1601]), .B(n25768), .Z(n25770) );
  NANDN U27263 ( .A(sreg[1600]), .B(n25731), .Z(n25735) );
  NAND U27264 ( .A(n25733), .B(n25732), .Z(n25734) );
  NAND U27265 ( .A(n25735), .B(n25734), .Z(n25769) );
  XNOR U27266 ( .A(n25770), .B(n25769), .Z(c[1601]) );
  NANDN U27267 ( .A(n25737), .B(n25736), .Z(n25741) );
  NANDN U27268 ( .A(n25739), .B(n25738), .Z(n25740) );
  AND U27269 ( .A(n25741), .B(n25740), .Z(n25776) );
  NANDN U27270 ( .A(n25743), .B(n25742), .Z(n25747) );
  NANDN U27271 ( .A(n25745), .B(n25744), .Z(n25746) );
  AND U27272 ( .A(n25747), .B(n25746), .Z(n25774) );
  NAND U27273 ( .A(n42143), .B(n25748), .Z(n25750) );
  XNOR U27274 ( .A(a[580]), .B(n4154), .Z(n25785) );
  NAND U27275 ( .A(n42144), .B(n25785), .Z(n25749) );
  AND U27276 ( .A(n25750), .B(n25749), .Z(n25800) );
  XOR U27277 ( .A(a[584]), .B(n42012), .Z(n25788) );
  XNOR U27278 ( .A(n25800), .B(n25799), .Z(n25802) );
  AND U27279 ( .A(a[586]), .B(b[0]), .Z(n25752) );
  XNOR U27280 ( .A(n25752), .B(n4071), .Z(n25754) );
  NANDN U27281 ( .A(b[0]), .B(a[585]), .Z(n25753) );
  NAND U27282 ( .A(n25754), .B(n25753), .Z(n25796) );
  XOR U27283 ( .A(a[582]), .B(n42085), .Z(n25789) );
  AND U27284 ( .A(a[578]), .B(b[7]), .Z(n25793) );
  XNOR U27285 ( .A(n25794), .B(n25793), .Z(n25795) );
  XNOR U27286 ( .A(n25796), .B(n25795), .Z(n25801) );
  XOR U27287 ( .A(n25802), .B(n25801), .Z(n25780) );
  NANDN U27288 ( .A(n25757), .B(n25756), .Z(n25761) );
  NANDN U27289 ( .A(n25759), .B(n25758), .Z(n25760) );
  AND U27290 ( .A(n25761), .B(n25760), .Z(n25779) );
  XNOR U27291 ( .A(n25780), .B(n25779), .Z(n25781) );
  NANDN U27292 ( .A(n25763), .B(n25762), .Z(n25767) );
  NAND U27293 ( .A(n25765), .B(n25764), .Z(n25766) );
  NAND U27294 ( .A(n25767), .B(n25766), .Z(n25782) );
  XNOR U27295 ( .A(n25781), .B(n25782), .Z(n25773) );
  XNOR U27296 ( .A(n25774), .B(n25773), .Z(n25775) );
  XNOR U27297 ( .A(n25776), .B(n25775), .Z(n25805) );
  XNOR U27298 ( .A(sreg[1602]), .B(n25805), .Z(n25807) );
  NANDN U27299 ( .A(sreg[1601]), .B(n25768), .Z(n25772) );
  NAND U27300 ( .A(n25770), .B(n25769), .Z(n25771) );
  NAND U27301 ( .A(n25772), .B(n25771), .Z(n25806) );
  XNOR U27302 ( .A(n25807), .B(n25806), .Z(c[1602]) );
  NANDN U27303 ( .A(n25774), .B(n25773), .Z(n25778) );
  NANDN U27304 ( .A(n25776), .B(n25775), .Z(n25777) );
  AND U27305 ( .A(n25778), .B(n25777), .Z(n25813) );
  NANDN U27306 ( .A(n25780), .B(n25779), .Z(n25784) );
  NANDN U27307 ( .A(n25782), .B(n25781), .Z(n25783) );
  AND U27308 ( .A(n25784), .B(n25783), .Z(n25811) );
  NAND U27309 ( .A(n42143), .B(n25785), .Z(n25787) );
  XNOR U27310 ( .A(a[581]), .B(n4154), .Z(n25822) );
  NAND U27311 ( .A(n42144), .B(n25822), .Z(n25786) );
  AND U27312 ( .A(n25787), .B(n25786), .Z(n25837) );
  XOR U27313 ( .A(a[585]), .B(n42012), .Z(n25825) );
  XNOR U27314 ( .A(n25837), .B(n25836), .Z(n25839) );
  XOR U27315 ( .A(a[583]), .B(n42085), .Z(n25829) );
  AND U27316 ( .A(a[579]), .B(b[7]), .Z(n25830) );
  XNOR U27317 ( .A(n25831), .B(n25830), .Z(n25832) );
  AND U27318 ( .A(a[587]), .B(b[0]), .Z(n25790) );
  XNOR U27319 ( .A(n25790), .B(n4071), .Z(n25792) );
  NANDN U27320 ( .A(b[0]), .B(a[586]), .Z(n25791) );
  NAND U27321 ( .A(n25792), .B(n25791), .Z(n25833) );
  XNOR U27322 ( .A(n25832), .B(n25833), .Z(n25838) );
  XOR U27323 ( .A(n25839), .B(n25838), .Z(n25817) );
  NANDN U27324 ( .A(n25794), .B(n25793), .Z(n25798) );
  NANDN U27325 ( .A(n25796), .B(n25795), .Z(n25797) );
  AND U27326 ( .A(n25798), .B(n25797), .Z(n25816) );
  XNOR U27327 ( .A(n25817), .B(n25816), .Z(n25818) );
  NANDN U27328 ( .A(n25800), .B(n25799), .Z(n25804) );
  NAND U27329 ( .A(n25802), .B(n25801), .Z(n25803) );
  NAND U27330 ( .A(n25804), .B(n25803), .Z(n25819) );
  XNOR U27331 ( .A(n25818), .B(n25819), .Z(n25810) );
  XNOR U27332 ( .A(n25811), .B(n25810), .Z(n25812) );
  XNOR U27333 ( .A(n25813), .B(n25812), .Z(n25842) );
  XNOR U27334 ( .A(sreg[1603]), .B(n25842), .Z(n25844) );
  NANDN U27335 ( .A(sreg[1602]), .B(n25805), .Z(n25809) );
  NAND U27336 ( .A(n25807), .B(n25806), .Z(n25808) );
  NAND U27337 ( .A(n25809), .B(n25808), .Z(n25843) );
  XNOR U27338 ( .A(n25844), .B(n25843), .Z(c[1603]) );
  NANDN U27339 ( .A(n25811), .B(n25810), .Z(n25815) );
  NANDN U27340 ( .A(n25813), .B(n25812), .Z(n25814) );
  AND U27341 ( .A(n25815), .B(n25814), .Z(n25850) );
  NANDN U27342 ( .A(n25817), .B(n25816), .Z(n25821) );
  NANDN U27343 ( .A(n25819), .B(n25818), .Z(n25820) );
  AND U27344 ( .A(n25821), .B(n25820), .Z(n25848) );
  NAND U27345 ( .A(n42143), .B(n25822), .Z(n25824) );
  XNOR U27346 ( .A(a[582]), .B(n4155), .Z(n25859) );
  NAND U27347 ( .A(n42144), .B(n25859), .Z(n25823) );
  AND U27348 ( .A(n25824), .B(n25823), .Z(n25874) );
  XOR U27349 ( .A(a[586]), .B(n42012), .Z(n25862) );
  XNOR U27350 ( .A(n25874), .B(n25873), .Z(n25876) );
  NAND U27351 ( .A(a[588]), .B(b[0]), .Z(n25826) );
  XNOR U27352 ( .A(b[1]), .B(n25826), .Z(n25828) );
  NANDN U27353 ( .A(b[0]), .B(a[587]), .Z(n25827) );
  AND U27354 ( .A(n25828), .B(n25827), .Z(n25869) );
  XOR U27355 ( .A(a[584]), .B(n42085), .Z(n25866) );
  AND U27356 ( .A(a[580]), .B(b[7]), .Z(n25867) );
  XOR U27357 ( .A(n25868), .B(n25867), .Z(n25870) );
  XNOR U27358 ( .A(n25869), .B(n25870), .Z(n25875) );
  XOR U27359 ( .A(n25876), .B(n25875), .Z(n25854) );
  NANDN U27360 ( .A(n25831), .B(n25830), .Z(n25835) );
  NANDN U27361 ( .A(n25833), .B(n25832), .Z(n25834) );
  AND U27362 ( .A(n25835), .B(n25834), .Z(n25853) );
  XNOR U27363 ( .A(n25854), .B(n25853), .Z(n25855) );
  NANDN U27364 ( .A(n25837), .B(n25836), .Z(n25841) );
  NAND U27365 ( .A(n25839), .B(n25838), .Z(n25840) );
  NAND U27366 ( .A(n25841), .B(n25840), .Z(n25856) );
  XNOR U27367 ( .A(n25855), .B(n25856), .Z(n25847) );
  XNOR U27368 ( .A(n25848), .B(n25847), .Z(n25849) );
  XNOR U27369 ( .A(n25850), .B(n25849), .Z(n25879) );
  XNOR U27370 ( .A(sreg[1604]), .B(n25879), .Z(n25881) );
  NANDN U27371 ( .A(sreg[1603]), .B(n25842), .Z(n25846) );
  NAND U27372 ( .A(n25844), .B(n25843), .Z(n25845) );
  NAND U27373 ( .A(n25846), .B(n25845), .Z(n25880) );
  XNOR U27374 ( .A(n25881), .B(n25880), .Z(c[1604]) );
  NANDN U27375 ( .A(n25848), .B(n25847), .Z(n25852) );
  NANDN U27376 ( .A(n25850), .B(n25849), .Z(n25851) );
  AND U27377 ( .A(n25852), .B(n25851), .Z(n25887) );
  NANDN U27378 ( .A(n25854), .B(n25853), .Z(n25858) );
  NANDN U27379 ( .A(n25856), .B(n25855), .Z(n25857) );
  AND U27380 ( .A(n25858), .B(n25857), .Z(n25885) );
  NAND U27381 ( .A(n42143), .B(n25859), .Z(n25861) );
  XNOR U27382 ( .A(a[583]), .B(n4155), .Z(n25896) );
  NAND U27383 ( .A(n42144), .B(n25896), .Z(n25860) );
  AND U27384 ( .A(n25861), .B(n25860), .Z(n25911) );
  XOR U27385 ( .A(a[587]), .B(n42012), .Z(n25899) );
  XNOR U27386 ( .A(n25911), .B(n25910), .Z(n25913) );
  AND U27387 ( .A(a[589]), .B(b[0]), .Z(n25863) );
  XNOR U27388 ( .A(n25863), .B(n4071), .Z(n25865) );
  NANDN U27389 ( .A(b[0]), .B(a[588]), .Z(n25864) );
  NAND U27390 ( .A(n25865), .B(n25864), .Z(n25907) );
  XOR U27391 ( .A(a[585]), .B(n42085), .Z(n25900) );
  AND U27392 ( .A(a[581]), .B(b[7]), .Z(n25904) );
  XNOR U27393 ( .A(n25905), .B(n25904), .Z(n25906) );
  XNOR U27394 ( .A(n25907), .B(n25906), .Z(n25912) );
  XOR U27395 ( .A(n25913), .B(n25912), .Z(n25891) );
  NANDN U27396 ( .A(n25868), .B(n25867), .Z(n25872) );
  NANDN U27397 ( .A(n25870), .B(n25869), .Z(n25871) );
  AND U27398 ( .A(n25872), .B(n25871), .Z(n25890) );
  XNOR U27399 ( .A(n25891), .B(n25890), .Z(n25892) );
  NANDN U27400 ( .A(n25874), .B(n25873), .Z(n25878) );
  NAND U27401 ( .A(n25876), .B(n25875), .Z(n25877) );
  NAND U27402 ( .A(n25878), .B(n25877), .Z(n25893) );
  XNOR U27403 ( .A(n25892), .B(n25893), .Z(n25884) );
  XNOR U27404 ( .A(n25885), .B(n25884), .Z(n25886) );
  XNOR U27405 ( .A(n25887), .B(n25886), .Z(n25916) );
  XNOR U27406 ( .A(sreg[1605]), .B(n25916), .Z(n25918) );
  NANDN U27407 ( .A(sreg[1604]), .B(n25879), .Z(n25883) );
  NAND U27408 ( .A(n25881), .B(n25880), .Z(n25882) );
  NAND U27409 ( .A(n25883), .B(n25882), .Z(n25917) );
  XNOR U27410 ( .A(n25918), .B(n25917), .Z(c[1605]) );
  NANDN U27411 ( .A(n25885), .B(n25884), .Z(n25889) );
  NANDN U27412 ( .A(n25887), .B(n25886), .Z(n25888) );
  AND U27413 ( .A(n25889), .B(n25888), .Z(n25924) );
  NANDN U27414 ( .A(n25891), .B(n25890), .Z(n25895) );
  NANDN U27415 ( .A(n25893), .B(n25892), .Z(n25894) );
  AND U27416 ( .A(n25895), .B(n25894), .Z(n25922) );
  NAND U27417 ( .A(n42143), .B(n25896), .Z(n25898) );
  XNOR U27418 ( .A(a[584]), .B(n4155), .Z(n25933) );
  NAND U27419 ( .A(n42144), .B(n25933), .Z(n25897) );
  AND U27420 ( .A(n25898), .B(n25897), .Z(n25948) );
  XOR U27421 ( .A(a[588]), .B(n42012), .Z(n25936) );
  XNOR U27422 ( .A(n25948), .B(n25947), .Z(n25950) );
  XOR U27423 ( .A(a[586]), .B(n42085), .Z(n25940) );
  AND U27424 ( .A(a[582]), .B(b[7]), .Z(n25941) );
  XNOR U27425 ( .A(n25942), .B(n25941), .Z(n25943) );
  AND U27426 ( .A(a[590]), .B(b[0]), .Z(n25901) );
  XNOR U27427 ( .A(n25901), .B(n4071), .Z(n25903) );
  NANDN U27428 ( .A(b[0]), .B(a[589]), .Z(n25902) );
  NAND U27429 ( .A(n25903), .B(n25902), .Z(n25944) );
  XNOR U27430 ( .A(n25943), .B(n25944), .Z(n25949) );
  XOR U27431 ( .A(n25950), .B(n25949), .Z(n25928) );
  NANDN U27432 ( .A(n25905), .B(n25904), .Z(n25909) );
  NANDN U27433 ( .A(n25907), .B(n25906), .Z(n25908) );
  AND U27434 ( .A(n25909), .B(n25908), .Z(n25927) );
  XNOR U27435 ( .A(n25928), .B(n25927), .Z(n25929) );
  NANDN U27436 ( .A(n25911), .B(n25910), .Z(n25915) );
  NAND U27437 ( .A(n25913), .B(n25912), .Z(n25914) );
  NAND U27438 ( .A(n25915), .B(n25914), .Z(n25930) );
  XNOR U27439 ( .A(n25929), .B(n25930), .Z(n25921) );
  XNOR U27440 ( .A(n25922), .B(n25921), .Z(n25923) );
  XNOR U27441 ( .A(n25924), .B(n25923), .Z(n25953) );
  XNOR U27442 ( .A(sreg[1606]), .B(n25953), .Z(n25955) );
  NANDN U27443 ( .A(sreg[1605]), .B(n25916), .Z(n25920) );
  NAND U27444 ( .A(n25918), .B(n25917), .Z(n25919) );
  NAND U27445 ( .A(n25920), .B(n25919), .Z(n25954) );
  XNOR U27446 ( .A(n25955), .B(n25954), .Z(c[1606]) );
  NANDN U27447 ( .A(n25922), .B(n25921), .Z(n25926) );
  NANDN U27448 ( .A(n25924), .B(n25923), .Z(n25925) );
  AND U27449 ( .A(n25926), .B(n25925), .Z(n25961) );
  NANDN U27450 ( .A(n25928), .B(n25927), .Z(n25932) );
  NANDN U27451 ( .A(n25930), .B(n25929), .Z(n25931) );
  AND U27452 ( .A(n25932), .B(n25931), .Z(n25959) );
  NAND U27453 ( .A(n42143), .B(n25933), .Z(n25935) );
  XNOR U27454 ( .A(a[585]), .B(n4155), .Z(n25970) );
  NAND U27455 ( .A(n42144), .B(n25970), .Z(n25934) );
  AND U27456 ( .A(n25935), .B(n25934), .Z(n25985) );
  XOR U27457 ( .A(a[589]), .B(n42012), .Z(n25973) );
  XNOR U27458 ( .A(n25985), .B(n25984), .Z(n25987) );
  AND U27459 ( .A(a[591]), .B(b[0]), .Z(n25937) );
  XNOR U27460 ( .A(n25937), .B(n4071), .Z(n25939) );
  NANDN U27461 ( .A(b[0]), .B(a[590]), .Z(n25938) );
  NAND U27462 ( .A(n25939), .B(n25938), .Z(n25981) );
  XOR U27463 ( .A(a[587]), .B(n42085), .Z(n25974) );
  AND U27464 ( .A(a[583]), .B(b[7]), .Z(n25978) );
  XNOR U27465 ( .A(n25979), .B(n25978), .Z(n25980) );
  XNOR U27466 ( .A(n25981), .B(n25980), .Z(n25986) );
  XOR U27467 ( .A(n25987), .B(n25986), .Z(n25965) );
  NANDN U27468 ( .A(n25942), .B(n25941), .Z(n25946) );
  NANDN U27469 ( .A(n25944), .B(n25943), .Z(n25945) );
  AND U27470 ( .A(n25946), .B(n25945), .Z(n25964) );
  XNOR U27471 ( .A(n25965), .B(n25964), .Z(n25966) );
  NANDN U27472 ( .A(n25948), .B(n25947), .Z(n25952) );
  NAND U27473 ( .A(n25950), .B(n25949), .Z(n25951) );
  NAND U27474 ( .A(n25952), .B(n25951), .Z(n25967) );
  XNOR U27475 ( .A(n25966), .B(n25967), .Z(n25958) );
  XNOR U27476 ( .A(n25959), .B(n25958), .Z(n25960) );
  XNOR U27477 ( .A(n25961), .B(n25960), .Z(n25990) );
  XNOR U27478 ( .A(sreg[1607]), .B(n25990), .Z(n25992) );
  NANDN U27479 ( .A(sreg[1606]), .B(n25953), .Z(n25957) );
  NAND U27480 ( .A(n25955), .B(n25954), .Z(n25956) );
  NAND U27481 ( .A(n25957), .B(n25956), .Z(n25991) );
  XNOR U27482 ( .A(n25992), .B(n25991), .Z(c[1607]) );
  NANDN U27483 ( .A(n25959), .B(n25958), .Z(n25963) );
  NANDN U27484 ( .A(n25961), .B(n25960), .Z(n25962) );
  AND U27485 ( .A(n25963), .B(n25962), .Z(n25998) );
  NANDN U27486 ( .A(n25965), .B(n25964), .Z(n25969) );
  NANDN U27487 ( .A(n25967), .B(n25966), .Z(n25968) );
  AND U27488 ( .A(n25969), .B(n25968), .Z(n25996) );
  NAND U27489 ( .A(n42143), .B(n25970), .Z(n25972) );
  XNOR U27490 ( .A(a[586]), .B(n4155), .Z(n26007) );
  NAND U27491 ( .A(n42144), .B(n26007), .Z(n25971) );
  AND U27492 ( .A(n25972), .B(n25971), .Z(n26022) );
  XOR U27493 ( .A(a[590]), .B(n42012), .Z(n26010) );
  XNOR U27494 ( .A(n26022), .B(n26021), .Z(n26024) );
  XOR U27495 ( .A(a[588]), .B(n42085), .Z(n26014) );
  AND U27496 ( .A(a[584]), .B(b[7]), .Z(n26015) );
  XNOR U27497 ( .A(n26016), .B(n26015), .Z(n26017) );
  AND U27498 ( .A(a[592]), .B(b[0]), .Z(n25975) );
  XNOR U27499 ( .A(n25975), .B(n4071), .Z(n25977) );
  NANDN U27500 ( .A(b[0]), .B(a[591]), .Z(n25976) );
  NAND U27501 ( .A(n25977), .B(n25976), .Z(n26018) );
  XNOR U27502 ( .A(n26017), .B(n26018), .Z(n26023) );
  XOR U27503 ( .A(n26024), .B(n26023), .Z(n26002) );
  NANDN U27504 ( .A(n25979), .B(n25978), .Z(n25983) );
  NANDN U27505 ( .A(n25981), .B(n25980), .Z(n25982) );
  AND U27506 ( .A(n25983), .B(n25982), .Z(n26001) );
  XNOR U27507 ( .A(n26002), .B(n26001), .Z(n26003) );
  NANDN U27508 ( .A(n25985), .B(n25984), .Z(n25989) );
  NAND U27509 ( .A(n25987), .B(n25986), .Z(n25988) );
  NAND U27510 ( .A(n25989), .B(n25988), .Z(n26004) );
  XNOR U27511 ( .A(n26003), .B(n26004), .Z(n25995) );
  XNOR U27512 ( .A(n25996), .B(n25995), .Z(n25997) );
  XNOR U27513 ( .A(n25998), .B(n25997), .Z(n26027) );
  XNOR U27514 ( .A(sreg[1608]), .B(n26027), .Z(n26029) );
  NANDN U27515 ( .A(sreg[1607]), .B(n25990), .Z(n25994) );
  NAND U27516 ( .A(n25992), .B(n25991), .Z(n25993) );
  NAND U27517 ( .A(n25994), .B(n25993), .Z(n26028) );
  XNOR U27518 ( .A(n26029), .B(n26028), .Z(c[1608]) );
  NANDN U27519 ( .A(n25996), .B(n25995), .Z(n26000) );
  NANDN U27520 ( .A(n25998), .B(n25997), .Z(n25999) );
  AND U27521 ( .A(n26000), .B(n25999), .Z(n26035) );
  NANDN U27522 ( .A(n26002), .B(n26001), .Z(n26006) );
  NANDN U27523 ( .A(n26004), .B(n26003), .Z(n26005) );
  AND U27524 ( .A(n26006), .B(n26005), .Z(n26033) );
  NAND U27525 ( .A(n42143), .B(n26007), .Z(n26009) );
  XNOR U27526 ( .A(a[587]), .B(n4155), .Z(n26044) );
  NAND U27527 ( .A(n42144), .B(n26044), .Z(n26008) );
  AND U27528 ( .A(n26009), .B(n26008), .Z(n26059) );
  XOR U27529 ( .A(a[591]), .B(n42012), .Z(n26047) );
  XNOR U27530 ( .A(n26059), .B(n26058), .Z(n26061) );
  AND U27531 ( .A(a[593]), .B(b[0]), .Z(n26011) );
  XNOR U27532 ( .A(n26011), .B(n4071), .Z(n26013) );
  NANDN U27533 ( .A(b[0]), .B(a[592]), .Z(n26012) );
  NAND U27534 ( .A(n26013), .B(n26012), .Z(n26055) );
  XOR U27535 ( .A(a[589]), .B(n42085), .Z(n26051) );
  AND U27536 ( .A(a[585]), .B(b[7]), .Z(n26052) );
  XNOR U27537 ( .A(n26053), .B(n26052), .Z(n26054) );
  XNOR U27538 ( .A(n26055), .B(n26054), .Z(n26060) );
  XOR U27539 ( .A(n26061), .B(n26060), .Z(n26039) );
  NANDN U27540 ( .A(n26016), .B(n26015), .Z(n26020) );
  NANDN U27541 ( .A(n26018), .B(n26017), .Z(n26019) );
  AND U27542 ( .A(n26020), .B(n26019), .Z(n26038) );
  XNOR U27543 ( .A(n26039), .B(n26038), .Z(n26040) );
  NANDN U27544 ( .A(n26022), .B(n26021), .Z(n26026) );
  NAND U27545 ( .A(n26024), .B(n26023), .Z(n26025) );
  NAND U27546 ( .A(n26026), .B(n26025), .Z(n26041) );
  XNOR U27547 ( .A(n26040), .B(n26041), .Z(n26032) );
  XNOR U27548 ( .A(n26033), .B(n26032), .Z(n26034) );
  XNOR U27549 ( .A(n26035), .B(n26034), .Z(n26064) );
  XNOR U27550 ( .A(sreg[1609]), .B(n26064), .Z(n26066) );
  NANDN U27551 ( .A(sreg[1608]), .B(n26027), .Z(n26031) );
  NAND U27552 ( .A(n26029), .B(n26028), .Z(n26030) );
  NAND U27553 ( .A(n26031), .B(n26030), .Z(n26065) );
  XNOR U27554 ( .A(n26066), .B(n26065), .Z(c[1609]) );
  NANDN U27555 ( .A(n26033), .B(n26032), .Z(n26037) );
  NANDN U27556 ( .A(n26035), .B(n26034), .Z(n26036) );
  AND U27557 ( .A(n26037), .B(n26036), .Z(n26072) );
  NANDN U27558 ( .A(n26039), .B(n26038), .Z(n26043) );
  NANDN U27559 ( .A(n26041), .B(n26040), .Z(n26042) );
  AND U27560 ( .A(n26043), .B(n26042), .Z(n26070) );
  NAND U27561 ( .A(n42143), .B(n26044), .Z(n26046) );
  XNOR U27562 ( .A(a[588]), .B(n4155), .Z(n26081) );
  NAND U27563 ( .A(n42144), .B(n26081), .Z(n26045) );
  AND U27564 ( .A(n26046), .B(n26045), .Z(n26096) );
  XOR U27565 ( .A(a[592]), .B(n42012), .Z(n26084) );
  XNOR U27566 ( .A(n26096), .B(n26095), .Z(n26098) );
  AND U27567 ( .A(a[594]), .B(b[0]), .Z(n26048) );
  XNOR U27568 ( .A(n26048), .B(n4071), .Z(n26050) );
  NANDN U27569 ( .A(b[0]), .B(a[593]), .Z(n26049) );
  NAND U27570 ( .A(n26050), .B(n26049), .Z(n26092) );
  XOR U27571 ( .A(a[590]), .B(n42085), .Z(n26088) );
  AND U27572 ( .A(a[586]), .B(b[7]), .Z(n26089) );
  XNOR U27573 ( .A(n26090), .B(n26089), .Z(n26091) );
  XNOR U27574 ( .A(n26092), .B(n26091), .Z(n26097) );
  XOR U27575 ( .A(n26098), .B(n26097), .Z(n26076) );
  NANDN U27576 ( .A(n26053), .B(n26052), .Z(n26057) );
  NANDN U27577 ( .A(n26055), .B(n26054), .Z(n26056) );
  AND U27578 ( .A(n26057), .B(n26056), .Z(n26075) );
  XNOR U27579 ( .A(n26076), .B(n26075), .Z(n26077) );
  NANDN U27580 ( .A(n26059), .B(n26058), .Z(n26063) );
  NAND U27581 ( .A(n26061), .B(n26060), .Z(n26062) );
  NAND U27582 ( .A(n26063), .B(n26062), .Z(n26078) );
  XNOR U27583 ( .A(n26077), .B(n26078), .Z(n26069) );
  XNOR U27584 ( .A(n26070), .B(n26069), .Z(n26071) );
  XNOR U27585 ( .A(n26072), .B(n26071), .Z(n26101) );
  XNOR U27586 ( .A(sreg[1610]), .B(n26101), .Z(n26103) );
  NANDN U27587 ( .A(sreg[1609]), .B(n26064), .Z(n26068) );
  NAND U27588 ( .A(n26066), .B(n26065), .Z(n26067) );
  NAND U27589 ( .A(n26068), .B(n26067), .Z(n26102) );
  XNOR U27590 ( .A(n26103), .B(n26102), .Z(c[1610]) );
  NANDN U27591 ( .A(n26070), .B(n26069), .Z(n26074) );
  NANDN U27592 ( .A(n26072), .B(n26071), .Z(n26073) );
  AND U27593 ( .A(n26074), .B(n26073), .Z(n26109) );
  NANDN U27594 ( .A(n26076), .B(n26075), .Z(n26080) );
  NANDN U27595 ( .A(n26078), .B(n26077), .Z(n26079) );
  AND U27596 ( .A(n26080), .B(n26079), .Z(n26107) );
  NAND U27597 ( .A(n42143), .B(n26081), .Z(n26083) );
  XNOR U27598 ( .A(a[589]), .B(n4156), .Z(n26118) );
  NAND U27599 ( .A(n42144), .B(n26118), .Z(n26082) );
  AND U27600 ( .A(n26083), .B(n26082), .Z(n26133) );
  XOR U27601 ( .A(a[593]), .B(n42012), .Z(n26121) );
  XNOR U27602 ( .A(n26133), .B(n26132), .Z(n26135) );
  AND U27603 ( .A(a[595]), .B(b[0]), .Z(n26085) );
  XNOR U27604 ( .A(n26085), .B(n4071), .Z(n26087) );
  NANDN U27605 ( .A(b[0]), .B(a[594]), .Z(n26086) );
  NAND U27606 ( .A(n26087), .B(n26086), .Z(n26129) );
  XOR U27607 ( .A(a[591]), .B(n42085), .Z(n26125) );
  AND U27608 ( .A(a[587]), .B(b[7]), .Z(n26126) );
  XNOR U27609 ( .A(n26127), .B(n26126), .Z(n26128) );
  XNOR U27610 ( .A(n26129), .B(n26128), .Z(n26134) );
  XOR U27611 ( .A(n26135), .B(n26134), .Z(n26113) );
  NANDN U27612 ( .A(n26090), .B(n26089), .Z(n26094) );
  NANDN U27613 ( .A(n26092), .B(n26091), .Z(n26093) );
  AND U27614 ( .A(n26094), .B(n26093), .Z(n26112) );
  XNOR U27615 ( .A(n26113), .B(n26112), .Z(n26114) );
  NANDN U27616 ( .A(n26096), .B(n26095), .Z(n26100) );
  NAND U27617 ( .A(n26098), .B(n26097), .Z(n26099) );
  NAND U27618 ( .A(n26100), .B(n26099), .Z(n26115) );
  XNOR U27619 ( .A(n26114), .B(n26115), .Z(n26106) );
  XNOR U27620 ( .A(n26107), .B(n26106), .Z(n26108) );
  XNOR U27621 ( .A(n26109), .B(n26108), .Z(n26138) );
  XNOR U27622 ( .A(sreg[1611]), .B(n26138), .Z(n26140) );
  NANDN U27623 ( .A(sreg[1610]), .B(n26101), .Z(n26105) );
  NAND U27624 ( .A(n26103), .B(n26102), .Z(n26104) );
  NAND U27625 ( .A(n26105), .B(n26104), .Z(n26139) );
  XNOR U27626 ( .A(n26140), .B(n26139), .Z(c[1611]) );
  NANDN U27627 ( .A(n26107), .B(n26106), .Z(n26111) );
  NANDN U27628 ( .A(n26109), .B(n26108), .Z(n26110) );
  AND U27629 ( .A(n26111), .B(n26110), .Z(n26146) );
  NANDN U27630 ( .A(n26113), .B(n26112), .Z(n26117) );
  NANDN U27631 ( .A(n26115), .B(n26114), .Z(n26116) );
  AND U27632 ( .A(n26117), .B(n26116), .Z(n26144) );
  NAND U27633 ( .A(n42143), .B(n26118), .Z(n26120) );
  XNOR U27634 ( .A(a[590]), .B(n4156), .Z(n26155) );
  NAND U27635 ( .A(n42144), .B(n26155), .Z(n26119) );
  AND U27636 ( .A(n26120), .B(n26119), .Z(n26170) );
  XOR U27637 ( .A(a[594]), .B(n42012), .Z(n26158) );
  XNOR U27638 ( .A(n26170), .B(n26169), .Z(n26172) );
  AND U27639 ( .A(a[596]), .B(b[0]), .Z(n26122) );
  XNOR U27640 ( .A(n26122), .B(n4071), .Z(n26124) );
  NANDN U27641 ( .A(b[0]), .B(a[595]), .Z(n26123) );
  NAND U27642 ( .A(n26124), .B(n26123), .Z(n26166) );
  XOR U27643 ( .A(a[592]), .B(n42085), .Z(n26159) );
  AND U27644 ( .A(a[588]), .B(b[7]), .Z(n26163) );
  XNOR U27645 ( .A(n26164), .B(n26163), .Z(n26165) );
  XNOR U27646 ( .A(n26166), .B(n26165), .Z(n26171) );
  XOR U27647 ( .A(n26172), .B(n26171), .Z(n26150) );
  NANDN U27648 ( .A(n26127), .B(n26126), .Z(n26131) );
  NANDN U27649 ( .A(n26129), .B(n26128), .Z(n26130) );
  AND U27650 ( .A(n26131), .B(n26130), .Z(n26149) );
  XNOR U27651 ( .A(n26150), .B(n26149), .Z(n26151) );
  NANDN U27652 ( .A(n26133), .B(n26132), .Z(n26137) );
  NAND U27653 ( .A(n26135), .B(n26134), .Z(n26136) );
  NAND U27654 ( .A(n26137), .B(n26136), .Z(n26152) );
  XNOR U27655 ( .A(n26151), .B(n26152), .Z(n26143) );
  XNOR U27656 ( .A(n26144), .B(n26143), .Z(n26145) );
  XNOR U27657 ( .A(n26146), .B(n26145), .Z(n26175) );
  XNOR U27658 ( .A(sreg[1612]), .B(n26175), .Z(n26177) );
  NANDN U27659 ( .A(sreg[1611]), .B(n26138), .Z(n26142) );
  NAND U27660 ( .A(n26140), .B(n26139), .Z(n26141) );
  NAND U27661 ( .A(n26142), .B(n26141), .Z(n26176) );
  XNOR U27662 ( .A(n26177), .B(n26176), .Z(c[1612]) );
  NANDN U27663 ( .A(n26144), .B(n26143), .Z(n26148) );
  NANDN U27664 ( .A(n26146), .B(n26145), .Z(n26147) );
  AND U27665 ( .A(n26148), .B(n26147), .Z(n26183) );
  NANDN U27666 ( .A(n26150), .B(n26149), .Z(n26154) );
  NANDN U27667 ( .A(n26152), .B(n26151), .Z(n26153) );
  AND U27668 ( .A(n26154), .B(n26153), .Z(n26181) );
  NAND U27669 ( .A(n42143), .B(n26155), .Z(n26157) );
  XNOR U27670 ( .A(a[591]), .B(n4156), .Z(n26192) );
  NAND U27671 ( .A(n42144), .B(n26192), .Z(n26156) );
  AND U27672 ( .A(n26157), .B(n26156), .Z(n26207) );
  XOR U27673 ( .A(a[595]), .B(n42012), .Z(n26195) );
  XNOR U27674 ( .A(n26207), .B(n26206), .Z(n26209) );
  XOR U27675 ( .A(a[593]), .B(n42085), .Z(n26199) );
  AND U27676 ( .A(a[589]), .B(b[7]), .Z(n26200) );
  XNOR U27677 ( .A(n26201), .B(n26200), .Z(n26202) );
  AND U27678 ( .A(a[597]), .B(b[0]), .Z(n26160) );
  XNOR U27679 ( .A(n26160), .B(n4071), .Z(n26162) );
  NANDN U27680 ( .A(b[0]), .B(a[596]), .Z(n26161) );
  NAND U27681 ( .A(n26162), .B(n26161), .Z(n26203) );
  XNOR U27682 ( .A(n26202), .B(n26203), .Z(n26208) );
  XOR U27683 ( .A(n26209), .B(n26208), .Z(n26187) );
  NANDN U27684 ( .A(n26164), .B(n26163), .Z(n26168) );
  NANDN U27685 ( .A(n26166), .B(n26165), .Z(n26167) );
  AND U27686 ( .A(n26168), .B(n26167), .Z(n26186) );
  XNOR U27687 ( .A(n26187), .B(n26186), .Z(n26188) );
  NANDN U27688 ( .A(n26170), .B(n26169), .Z(n26174) );
  NAND U27689 ( .A(n26172), .B(n26171), .Z(n26173) );
  NAND U27690 ( .A(n26174), .B(n26173), .Z(n26189) );
  XNOR U27691 ( .A(n26188), .B(n26189), .Z(n26180) );
  XNOR U27692 ( .A(n26181), .B(n26180), .Z(n26182) );
  XNOR U27693 ( .A(n26183), .B(n26182), .Z(n26212) );
  XNOR U27694 ( .A(sreg[1613]), .B(n26212), .Z(n26214) );
  NANDN U27695 ( .A(sreg[1612]), .B(n26175), .Z(n26179) );
  NAND U27696 ( .A(n26177), .B(n26176), .Z(n26178) );
  NAND U27697 ( .A(n26179), .B(n26178), .Z(n26213) );
  XNOR U27698 ( .A(n26214), .B(n26213), .Z(c[1613]) );
  NANDN U27699 ( .A(n26181), .B(n26180), .Z(n26185) );
  NANDN U27700 ( .A(n26183), .B(n26182), .Z(n26184) );
  AND U27701 ( .A(n26185), .B(n26184), .Z(n26220) );
  NANDN U27702 ( .A(n26187), .B(n26186), .Z(n26191) );
  NANDN U27703 ( .A(n26189), .B(n26188), .Z(n26190) );
  AND U27704 ( .A(n26191), .B(n26190), .Z(n26218) );
  NAND U27705 ( .A(n42143), .B(n26192), .Z(n26194) );
  XNOR U27706 ( .A(a[592]), .B(n4156), .Z(n26229) );
  NAND U27707 ( .A(n42144), .B(n26229), .Z(n26193) );
  AND U27708 ( .A(n26194), .B(n26193), .Z(n26244) );
  XOR U27709 ( .A(a[596]), .B(n42012), .Z(n26232) );
  XNOR U27710 ( .A(n26244), .B(n26243), .Z(n26246) );
  AND U27711 ( .A(a[598]), .B(b[0]), .Z(n26196) );
  XNOR U27712 ( .A(n26196), .B(n4071), .Z(n26198) );
  NANDN U27713 ( .A(b[0]), .B(a[597]), .Z(n26197) );
  NAND U27714 ( .A(n26198), .B(n26197), .Z(n26240) );
  XOR U27715 ( .A(a[594]), .B(n42085), .Z(n26233) );
  AND U27716 ( .A(a[590]), .B(b[7]), .Z(n26237) );
  XNOR U27717 ( .A(n26238), .B(n26237), .Z(n26239) );
  XNOR U27718 ( .A(n26240), .B(n26239), .Z(n26245) );
  XOR U27719 ( .A(n26246), .B(n26245), .Z(n26224) );
  NANDN U27720 ( .A(n26201), .B(n26200), .Z(n26205) );
  NANDN U27721 ( .A(n26203), .B(n26202), .Z(n26204) );
  AND U27722 ( .A(n26205), .B(n26204), .Z(n26223) );
  XNOR U27723 ( .A(n26224), .B(n26223), .Z(n26225) );
  NANDN U27724 ( .A(n26207), .B(n26206), .Z(n26211) );
  NAND U27725 ( .A(n26209), .B(n26208), .Z(n26210) );
  NAND U27726 ( .A(n26211), .B(n26210), .Z(n26226) );
  XNOR U27727 ( .A(n26225), .B(n26226), .Z(n26217) );
  XNOR U27728 ( .A(n26218), .B(n26217), .Z(n26219) );
  XNOR U27729 ( .A(n26220), .B(n26219), .Z(n26249) );
  XNOR U27730 ( .A(sreg[1614]), .B(n26249), .Z(n26251) );
  NANDN U27731 ( .A(sreg[1613]), .B(n26212), .Z(n26216) );
  NAND U27732 ( .A(n26214), .B(n26213), .Z(n26215) );
  NAND U27733 ( .A(n26216), .B(n26215), .Z(n26250) );
  XNOR U27734 ( .A(n26251), .B(n26250), .Z(c[1614]) );
  NANDN U27735 ( .A(n26218), .B(n26217), .Z(n26222) );
  NANDN U27736 ( .A(n26220), .B(n26219), .Z(n26221) );
  AND U27737 ( .A(n26222), .B(n26221), .Z(n26257) );
  NANDN U27738 ( .A(n26224), .B(n26223), .Z(n26228) );
  NANDN U27739 ( .A(n26226), .B(n26225), .Z(n26227) );
  AND U27740 ( .A(n26228), .B(n26227), .Z(n26255) );
  NAND U27741 ( .A(n42143), .B(n26229), .Z(n26231) );
  XNOR U27742 ( .A(a[593]), .B(n4156), .Z(n26266) );
  NAND U27743 ( .A(n42144), .B(n26266), .Z(n26230) );
  AND U27744 ( .A(n26231), .B(n26230), .Z(n26281) );
  XOR U27745 ( .A(a[597]), .B(n42012), .Z(n26269) );
  XNOR U27746 ( .A(n26281), .B(n26280), .Z(n26283) );
  XOR U27747 ( .A(a[595]), .B(n42085), .Z(n26273) );
  AND U27748 ( .A(a[591]), .B(b[7]), .Z(n26274) );
  XNOR U27749 ( .A(n26275), .B(n26274), .Z(n26276) );
  AND U27750 ( .A(a[599]), .B(b[0]), .Z(n26234) );
  XNOR U27751 ( .A(n26234), .B(n4071), .Z(n26236) );
  NANDN U27752 ( .A(b[0]), .B(a[598]), .Z(n26235) );
  NAND U27753 ( .A(n26236), .B(n26235), .Z(n26277) );
  XNOR U27754 ( .A(n26276), .B(n26277), .Z(n26282) );
  XOR U27755 ( .A(n26283), .B(n26282), .Z(n26261) );
  NANDN U27756 ( .A(n26238), .B(n26237), .Z(n26242) );
  NANDN U27757 ( .A(n26240), .B(n26239), .Z(n26241) );
  AND U27758 ( .A(n26242), .B(n26241), .Z(n26260) );
  XNOR U27759 ( .A(n26261), .B(n26260), .Z(n26262) );
  NANDN U27760 ( .A(n26244), .B(n26243), .Z(n26248) );
  NAND U27761 ( .A(n26246), .B(n26245), .Z(n26247) );
  NAND U27762 ( .A(n26248), .B(n26247), .Z(n26263) );
  XNOR U27763 ( .A(n26262), .B(n26263), .Z(n26254) );
  XNOR U27764 ( .A(n26255), .B(n26254), .Z(n26256) );
  XNOR U27765 ( .A(n26257), .B(n26256), .Z(n26286) );
  XNOR U27766 ( .A(sreg[1615]), .B(n26286), .Z(n26288) );
  NANDN U27767 ( .A(sreg[1614]), .B(n26249), .Z(n26253) );
  NAND U27768 ( .A(n26251), .B(n26250), .Z(n26252) );
  NAND U27769 ( .A(n26253), .B(n26252), .Z(n26287) );
  XNOR U27770 ( .A(n26288), .B(n26287), .Z(c[1615]) );
  NANDN U27771 ( .A(n26255), .B(n26254), .Z(n26259) );
  NANDN U27772 ( .A(n26257), .B(n26256), .Z(n26258) );
  AND U27773 ( .A(n26259), .B(n26258), .Z(n26294) );
  NANDN U27774 ( .A(n26261), .B(n26260), .Z(n26265) );
  NANDN U27775 ( .A(n26263), .B(n26262), .Z(n26264) );
  AND U27776 ( .A(n26265), .B(n26264), .Z(n26292) );
  NAND U27777 ( .A(n42143), .B(n26266), .Z(n26268) );
  XNOR U27778 ( .A(a[594]), .B(n4156), .Z(n26303) );
  NAND U27779 ( .A(n42144), .B(n26303), .Z(n26267) );
  AND U27780 ( .A(n26268), .B(n26267), .Z(n26318) );
  XOR U27781 ( .A(a[598]), .B(n42012), .Z(n26306) );
  XNOR U27782 ( .A(n26318), .B(n26317), .Z(n26320) );
  AND U27783 ( .A(a[600]), .B(b[0]), .Z(n26270) );
  XNOR U27784 ( .A(n26270), .B(n4071), .Z(n26272) );
  NANDN U27785 ( .A(b[0]), .B(a[599]), .Z(n26271) );
  NAND U27786 ( .A(n26272), .B(n26271), .Z(n26314) );
  XOR U27787 ( .A(a[596]), .B(n42085), .Z(n26310) );
  AND U27788 ( .A(a[592]), .B(b[7]), .Z(n26311) );
  XNOR U27789 ( .A(n26312), .B(n26311), .Z(n26313) );
  XNOR U27790 ( .A(n26314), .B(n26313), .Z(n26319) );
  XOR U27791 ( .A(n26320), .B(n26319), .Z(n26298) );
  NANDN U27792 ( .A(n26275), .B(n26274), .Z(n26279) );
  NANDN U27793 ( .A(n26277), .B(n26276), .Z(n26278) );
  AND U27794 ( .A(n26279), .B(n26278), .Z(n26297) );
  XNOR U27795 ( .A(n26298), .B(n26297), .Z(n26299) );
  NANDN U27796 ( .A(n26281), .B(n26280), .Z(n26285) );
  NAND U27797 ( .A(n26283), .B(n26282), .Z(n26284) );
  NAND U27798 ( .A(n26285), .B(n26284), .Z(n26300) );
  XNOR U27799 ( .A(n26299), .B(n26300), .Z(n26291) );
  XNOR U27800 ( .A(n26292), .B(n26291), .Z(n26293) );
  XNOR U27801 ( .A(n26294), .B(n26293), .Z(n26323) );
  XNOR U27802 ( .A(sreg[1616]), .B(n26323), .Z(n26325) );
  NANDN U27803 ( .A(sreg[1615]), .B(n26286), .Z(n26290) );
  NAND U27804 ( .A(n26288), .B(n26287), .Z(n26289) );
  NAND U27805 ( .A(n26290), .B(n26289), .Z(n26324) );
  XNOR U27806 ( .A(n26325), .B(n26324), .Z(c[1616]) );
  NANDN U27807 ( .A(n26292), .B(n26291), .Z(n26296) );
  NANDN U27808 ( .A(n26294), .B(n26293), .Z(n26295) );
  AND U27809 ( .A(n26296), .B(n26295), .Z(n26331) );
  NANDN U27810 ( .A(n26298), .B(n26297), .Z(n26302) );
  NANDN U27811 ( .A(n26300), .B(n26299), .Z(n26301) );
  AND U27812 ( .A(n26302), .B(n26301), .Z(n26329) );
  NAND U27813 ( .A(n42143), .B(n26303), .Z(n26305) );
  XNOR U27814 ( .A(a[595]), .B(n4156), .Z(n26340) );
  NAND U27815 ( .A(n42144), .B(n26340), .Z(n26304) );
  AND U27816 ( .A(n26305), .B(n26304), .Z(n26355) );
  XOR U27817 ( .A(a[599]), .B(n42012), .Z(n26343) );
  XNOR U27818 ( .A(n26355), .B(n26354), .Z(n26357) );
  AND U27819 ( .A(b[0]), .B(a[601]), .Z(n26307) );
  XOR U27820 ( .A(b[1]), .B(n26307), .Z(n26309) );
  NANDN U27821 ( .A(b[0]), .B(a[600]), .Z(n26308) );
  AND U27822 ( .A(n26309), .B(n26308), .Z(n26350) );
  XOR U27823 ( .A(a[597]), .B(n42085), .Z(n26347) );
  AND U27824 ( .A(a[593]), .B(b[7]), .Z(n26348) );
  XOR U27825 ( .A(n26349), .B(n26348), .Z(n26351) );
  XNOR U27826 ( .A(n26350), .B(n26351), .Z(n26356) );
  XOR U27827 ( .A(n26357), .B(n26356), .Z(n26335) );
  NANDN U27828 ( .A(n26312), .B(n26311), .Z(n26316) );
  NANDN U27829 ( .A(n26314), .B(n26313), .Z(n26315) );
  AND U27830 ( .A(n26316), .B(n26315), .Z(n26334) );
  XNOR U27831 ( .A(n26335), .B(n26334), .Z(n26336) );
  NANDN U27832 ( .A(n26318), .B(n26317), .Z(n26322) );
  NAND U27833 ( .A(n26320), .B(n26319), .Z(n26321) );
  NAND U27834 ( .A(n26322), .B(n26321), .Z(n26337) );
  XNOR U27835 ( .A(n26336), .B(n26337), .Z(n26328) );
  XNOR U27836 ( .A(n26329), .B(n26328), .Z(n26330) );
  XNOR U27837 ( .A(n26331), .B(n26330), .Z(n26360) );
  XNOR U27838 ( .A(sreg[1617]), .B(n26360), .Z(n26362) );
  NANDN U27839 ( .A(sreg[1616]), .B(n26323), .Z(n26327) );
  NAND U27840 ( .A(n26325), .B(n26324), .Z(n26326) );
  NAND U27841 ( .A(n26327), .B(n26326), .Z(n26361) );
  XNOR U27842 ( .A(n26362), .B(n26361), .Z(c[1617]) );
  NANDN U27843 ( .A(n26329), .B(n26328), .Z(n26333) );
  NANDN U27844 ( .A(n26331), .B(n26330), .Z(n26332) );
  AND U27845 ( .A(n26333), .B(n26332), .Z(n26368) );
  NANDN U27846 ( .A(n26335), .B(n26334), .Z(n26339) );
  NANDN U27847 ( .A(n26337), .B(n26336), .Z(n26338) );
  AND U27848 ( .A(n26339), .B(n26338), .Z(n26366) );
  NAND U27849 ( .A(n42143), .B(n26340), .Z(n26342) );
  XNOR U27850 ( .A(a[596]), .B(n4157), .Z(n26377) );
  NAND U27851 ( .A(n42144), .B(n26377), .Z(n26341) );
  AND U27852 ( .A(n26342), .B(n26341), .Z(n26392) );
  XOR U27853 ( .A(a[600]), .B(n42012), .Z(n26380) );
  XNOR U27854 ( .A(n26392), .B(n26391), .Z(n26394) );
  AND U27855 ( .A(a[602]), .B(b[0]), .Z(n26344) );
  XNOR U27856 ( .A(n26344), .B(n4071), .Z(n26346) );
  NANDN U27857 ( .A(b[0]), .B(a[601]), .Z(n26345) );
  NAND U27858 ( .A(n26346), .B(n26345), .Z(n26388) );
  XOR U27859 ( .A(a[598]), .B(n42085), .Z(n26381) );
  AND U27860 ( .A(a[594]), .B(b[7]), .Z(n26385) );
  XNOR U27861 ( .A(n26386), .B(n26385), .Z(n26387) );
  XNOR U27862 ( .A(n26388), .B(n26387), .Z(n26393) );
  XOR U27863 ( .A(n26394), .B(n26393), .Z(n26372) );
  NANDN U27864 ( .A(n26349), .B(n26348), .Z(n26353) );
  NANDN U27865 ( .A(n26351), .B(n26350), .Z(n26352) );
  AND U27866 ( .A(n26353), .B(n26352), .Z(n26371) );
  XNOR U27867 ( .A(n26372), .B(n26371), .Z(n26373) );
  NANDN U27868 ( .A(n26355), .B(n26354), .Z(n26359) );
  NAND U27869 ( .A(n26357), .B(n26356), .Z(n26358) );
  NAND U27870 ( .A(n26359), .B(n26358), .Z(n26374) );
  XNOR U27871 ( .A(n26373), .B(n26374), .Z(n26365) );
  XNOR U27872 ( .A(n26366), .B(n26365), .Z(n26367) );
  XNOR U27873 ( .A(n26368), .B(n26367), .Z(n26397) );
  XNOR U27874 ( .A(sreg[1618]), .B(n26397), .Z(n26399) );
  NANDN U27875 ( .A(sreg[1617]), .B(n26360), .Z(n26364) );
  NAND U27876 ( .A(n26362), .B(n26361), .Z(n26363) );
  NAND U27877 ( .A(n26364), .B(n26363), .Z(n26398) );
  XNOR U27878 ( .A(n26399), .B(n26398), .Z(c[1618]) );
  NANDN U27879 ( .A(n26366), .B(n26365), .Z(n26370) );
  NANDN U27880 ( .A(n26368), .B(n26367), .Z(n26369) );
  AND U27881 ( .A(n26370), .B(n26369), .Z(n26405) );
  NANDN U27882 ( .A(n26372), .B(n26371), .Z(n26376) );
  NANDN U27883 ( .A(n26374), .B(n26373), .Z(n26375) );
  AND U27884 ( .A(n26376), .B(n26375), .Z(n26403) );
  NAND U27885 ( .A(n42143), .B(n26377), .Z(n26379) );
  XNOR U27886 ( .A(a[597]), .B(n4157), .Z(n26414) );
  NAND U27887 ( .A(n42144), .B(n26414), .Z(n26378) );
  AND U27888 ( .A(n26379), .B(n26378), .Z(n26429) );
  XOR U27889 ( .A(a[601]), .B(n42012), .Z(n26417) );
  XNOR U27890 ( .A(n26429), .B(n26428), .Z(n26431) );
  XOR U27891 ( .A(a[599]), .B(n42085), .Z(n26421) );
  AND U27892 ( .A(a[595]), .B(b[7]), .Z(n26422) );
  XNOR U27893 ( .A(n26423), .B(n26422), .Z(n26424) );
  AND U27894 ( .A(a[603]), .B(b[0]), .Z(n26382) );
  XNOR U27895 ( .A(n26382), .B(n4071), .Z(n26384) );
  NANDN U27896 ( .A(b[0]), .B(a[602]), .Z(n26383) );
  NAND U27897 ( .A(n26384), .B(n26383), .Z(n26425) );
  XNOR U27898 ( .A(n26424), .B(n26425), .Z(n26430) );
  XOR U27899 ( .A(n26431), .B(n26430), .Z(n26409) );
  NANDN U27900 ( .A(n26386), .B(n26385), .Z(n26390) );
  NANDN U27901 ( .A(n26388), .B(n26387), .Z(n26389) );
  AND U27902 ( .A(n26390), .B(n26389), .Z(n26408) );
  XNOR U27903 ( .A(n26409), .B(n26408), .Z(n26410) );
  NANDN U27904 ( .A(n26392), .B(n26391), .Z(n26396) );
  NAND U27905 ( .A(n26394), .B(n26393), .Z(n26395) );
  NAND U27906 ( .A(n26396), .B(n26395), .Z(n26411) );
  XNOR U27907 ( .A(n26410), .B(n26411), .Z(n26402) );
  XNOR U27908 ( .A(n26403), .B(n26402), .Z(n26404) );
  XNOR U27909 ( .A(n26405), .B(n26404), .Z(n26434) );
  XNOR U27910 ( .A(sreg[1619]), .B(n26434), .Z(n26436) );
  NANDN U27911 ( .A(sreg[1618]), .B(n26397), .Z(n26401) );
  NAND U27912 ( .A(n26399), .B(n26398), .Z(n26400) );
  NAND U27913 ( .A(n26401), .B(n26400), .Z(n26435) );
  XNOR U27914 ( .A(n26436), .B(n26435), .Z(c[1619]) );
  NANDN U27915 ( .A(n26403), .B(n26402), .Z(n26407) );
  NANDN U27916 ( .A(n26405), .B(n26404), .Z(n26406) );
  AND U27917 ( .A(n26407), .B(n26406), .Z(n26442) );
  NANDN U27918 ( .A(n26409), .B(n26408), .Z(n26413) );
  NANDN U27919 ( .A(n26411), .B(n26410), .Z(n26412) );
  AND U27920 ( .A(n26413), .B(n26412), .Z(n26440) );
  NAND U27921 ( .A(n42143), .B(n26414), .Z(n26416) );
  XNOR U27922 ( .A(a[598]), .B(n4157), .Z(n26451) );
  NAND U27923 ( .A(n42144), .B(n26451), .Z(n26415) );
  AND U27924 ( .A(n26416), .B(n26415), .Z(n26466) );
  XOR U27925 ( .A(a[602]), .B(n42012), .Z(n26454) );
  XNOR U27926 ( .A(n26466), .B(n26465), .Z(n26468) );
  AND U27927 ( .A(a[604]), .B(b[0]), .Z(n26418) );
  XNOR U27928 ( .A(n26418), .B(n4071), .Z(n26420) );
  NANDN U27929 ( .A(b[0]), .B(a[603]), .Z(n26419) );
  NAND U27930 ( .A(n26420), .B(n26419), .Z(n26462) );
  XOR U27931 ( .A(a[600]), .B(n42085), .Z(n26455) );
  AND U27932 ( .A(a[596]), .B(b[7]), .Z(n26459) );
  XNOR U27933 ( .A(n26460), .B(n26459), .Z(n26461) );
  XNOR U27934 ( .A(n26462), .B(n26461), .Z(n26467) );
  XOR U27935 ( .A(n26468), .B(n26467), .Z(n26446) );
  NANDN U27936 ( .A(n26423), .B(n26422), .Z(n26427) );
  NANDN U27937 ( .A(n26425), .B(n26424), .Z(n26426) );
  AND U27938 ( .A(n26427), .B(n26426), .Z(n26445) );
  XNOR U27939 ( .A(n26446), .B(n26445), .Z(n26447) );
  NANDN U27940 ( .A(n26429), .B(n26428), .Z(n26433) );
  NAND U27941 ( .A(n26431), .B(n26430), .Z(n26432) );
  NAND U27942 ( .A(n26433), .B(n26432), .Z(n26448) );
  XNOR U27943 ( .A(n26447), .B(n26448), .Z(n26439) );
  XNOR U27944 ( .A(n26440), .B(n26439), .Z(n26441) );
  XNOR U27945 ( .A(n26442), .B(n26441), .Z(n26471) );
  XNOR U27946 ( .A(sreg[1620]), .B(n26471), .Z(n26473) );
  NANDN U27947 ( .A(sreg[1619]), .B(n26434), .Z(n26438) );
  NAND U27948 ( .A(n26436), .B(n26435), .Z(n26437) );
  NAND U27949 ( .A(n26438), .B(n26437), .Z(n26472) );
  XNOR U27950 ( .A(n26473), .B(n26472), .Z(c[1620]) );
  NANDN U27951 ( .A(n26440), .B(n26439), .Z(n26444) );
  NANDN U27952 ( .A(n26442), .B(n26441), .Z(n26443) );
  AND U27953 ( .A(n26444), .B(n26443), .Z(n26479) );
  NANDN U27954 ( .A(n26446), .B(n26445), .Z(n26450) );
  NANDN U27955 ( .A(n26448), .B(n26447), .Z(n26449) );
  AND U27956 ( .A(n26450), .B(n26449), .Z(n26477) );
  NAND U27957 ( .A(n42143), .B(n26451), .Z(n26453) );
  XNOR U27958 ( .A(a[599]), .B(n4157), .Z(n26488) );
  NAND U27959 ( .A(n42144), .B(n26488), .Z(n26452) );
  AND U27960 ( .A(n26453), .B(n26452), .Z(n26503) );
  XOR U27961 ( .A(a[603]), .B(n42012), .Z(n26491) );
  XNOR U27962 ( .A(n26503), .B(n26502), .Z(n26505) );
  XOR U27963 ( .A(a[601]), .B(n42085), .Z(n26495) );
  AND U27964 ( .A(a[597]), .B(b[7]), .Z(n26496) );
  XNOR U27965 ( .A(n26497), .B(n26496), .Z(n26498) );
  AND U27966 ( .A(a[605]), .B(b[0]), .Z(n26456) );
  XNOR U27967 ( .A(n26456), .B(n4071), .Z(n26458) );
  NANDN U27968 ( .A(b[0]), .B(a[604]), .Z(n26457) );
  NAND U27969 ( .A(n26458), .B(n26457), .Z(n26499) );
  XNOR U27970 ( .A(n26498), .B(n26499), .Z(n26504) );
  XOR U27971 ( .A(n26505), .B(n26504), .Z(n26483) );
  NANDN U27972 ( .A(n26460), .B(n26459), .Z(n26464) );
  NANDN U27973 ( .A(n26462), .B(n26461), .Z(n26463) );
  AND U27974 ( .A(n26464), .B(n26463), .Z(n26482) );
  XNOR U27975 ( .A(n26483), .B(n26482), .Z(n26484) );
  NANDN U27976 ( .A(n26466), .B(n26465), .Z(n26470) );
  NAND U27977 ( .A(n26468), .B(n26467), .Z(n26469) );
  NAND U27978 ( .A(n26470), .B(n26469), .Z(n26485) );
  XNOR U27979 ( .A(n26484), .B(n26485), .Z(n26476) );
  XNOR U27980 ( .A(n26477), .B(n26476), .Z(n26478) );
  XNOR U27981 ( .A(n26479), .B(n26478), .Z(n26508) );
  XNOR U27982 ( .A(sreg[1621]), .B(n26508), .Z(n26510) );
  NANDN U27983 ( .A(sreg[1620]), .B(n26471), .Z(n26475) );
  NAND U27984 ( .A(n26473), .B(n26472), .Z(n26474) );
  NAND U27985 ( .A(n26475), .B(n26474), .Z(n26509) );
  XNOR U27986 ( .A(n26510), .B(n26509), .Z(c[1621]) );
  NANDN U27987 ( .A(n26477), .B(n26476), .Z(n26481) );
  NANDN U27988 ( .A(n26479), .B(n26478), .Z(n26480) );
  AND U27989 ( .A(n26481), .B(n26480), .Z(n26516) );
  NANDN U27990 ( .A(n26483), .B(n26482), .Z(n26487) );
  NANDN U27991 ( .A(n26485), .B(n26484), .Z(n26486) );
  AND U27992 ( .A(n26487), .B(n26486), .Z(n26514) );
  NAND U27993 ( .A(n42143), .B(n26488), .Z(n26490) );
  XNOR U27994 ( .A(a[600]), .B(n4157), .Z(n26525) );
  NAND U27995 ( .A(n42144), .B(n26525), .Z(n26489) );
  AND U27996 ( .A(n26490), .B(n26489), .Z(n26540) );
  XOR U27997 ( .A(a[604]), .B(n42012), .Z(n26528) );
  XNOR U27998 ( .A(n26540), .B(n26539), .Z(n26542) );
  AND U27999 ( .A(a[606]), .B(b[0]), .Z(n26492) );
  XNOR U28000 ( .A(n26492), .B(n4071), .Z(n26494) );
  NANDN U28001 ( .A(b[0]), .B(a[605]), .Z(n26493) );
  NAND U28002 ( .A(n26494), .B(n26493), .Z(n26536) );
  XOR U28003 ( .A(a[602]), .B(n42085), .Z(n26532) );
  AND U28004 ( .A(a[598]), .B(b[7]), .Z(n26533) );
  XNOR U28005 ( .A(n26534), .B(n26533), .Z(n26535) );
  XNOR U28006 ( .A(n26536), .B(n26535), .Z(n26541) );
  XOR U28007 ( .A(n26542), .B(n26541), .Z(n26520) );
  NANDN U28008 ( .A(n26497), .B(n26496), .Z(n26501) );
  NANDN U28009 ( .A(n26499), .B(n26498), .Z(n26500) );
  AND U28010 ( .A(n26501), .B(n26500), .Z(n26519) );
  XNOR U28011 ( .A(n26520), .B(n26519), .Z(n26521) );
  NANDN U28012 ( .A(n26503), .B(n26502), .Z(n26507) );
  NAND U28013 ( .A(n26505), .B(n26504), .Z(n26506) );
  NAND U28014 ( .A(n26507), .B(n26506), .Z(n26522) );
  XNOR U28015 ( .A(n26521), .B(n26522), .Z(n26513) );
  XNOR U28016 ( .A(n26514), .B(n26513), .Z(n26515) );
  XNOR U28017 ( .A(n26516), .B(n26515), .Z(n26545) );
  XNOR U28018 ( .A(sreg[1622]), .B(n26545), .Z(n26547) );
  NANDN U28019 ( .A(sreg[1621]), .B(n26508), .Z(n26512) );
  NAND U28020 ( .A(n26510), .B(n26509), .Z(n26511) );
  NAND U28021 ( .A(n26512), .B(n26511), .Z(n26546) );
  XNOR U28022 ( .A(n26547), .B(n26546), .Z(c[1622]) );
  NANDN U28023 ( .A(n26514), .B(n26513), .Z(n26518) );
  NANDN U28024 ( .A(n26516), .B(n26515), .Z(n26517) );
  AND U28025 ( .A(n26518), .B(n26517), .Z(n26553) );
  NANDN U28026 ( .A(n26520), .B(n26519), .Z(n26524) );
  NANDN U28027 ( .A(n26522), .B(n26521), .Z(n26523) );
  AND U28028 ( .A(n26524), .B(n26523), .Z(n26551) );
  NAND U28029 ( .A(n42143), .B(n26525), .Z(n26527) );
  XNOR U28030 ( .A(a[601]), .B(n4157), .Z(n26562) );
  NAND U28031 ( .A(n42144), .B(n26562), .Z(n26526) );
  AND U28032 ( .A(n26527), .B(n26526), .Z(n26577) );
  XOR U28033 ( .A(a[605]), .B(n42012), .Z(n26565) );
  XNOR U28034 ( .A(n26577), .B(n26576), .Z(n26579) );
  AND U28035 ( .A(a[607]), .B(b[0]), .Z(n26529) );
  XNOR U28036 ( .A(n26529), .B(n4071), .Z(n26531) );
  NANDN U28037 ( .A(b[0]), .B(a[606]), .Z(n26530) );
  NAND U28038 ( .A(n26531), .B(n26530), .Z(n26573) );
  XOR U28039 ( .A(a[603]), .B(n42085), .Z(n26569) );
  AND U28040 ( .A(a[599]), .B(b[7]), .Z(n26570) );
  XNOR U28041 ( .A(n26571), .B(n26570), .Z(n26572) );
  XNOR U28042 ( .A(n26573), .B(n26572), .Z(n26578) );
  XOR U28043 ( .A(n26579), .B(n26578), .Z(n26557) );
  NANDN U28044 ( .A(n26534), .B(n26533), .Z(n26538) );
  NANDN U28045 ( .A(n26536), .B(n26535), .Z(n26537) );
  AND U28046 ( .A(n26538), .B(n26537), .Z(n26556) );
  XNOR U28047 ( .A(n26557), .B(n26556), .Z(n26558) );
  NANDN U28048 ( .A(n26540), .B(n26539), .Z(n26544) );
  NAND U28049 ( .A(n26542), .B(n26541), .Z(n26543) );
  NAND U28050 ( .A(n26544), .B(n26543), .Z(n26559) );
  XNOR U28051 ( .A(n26558), .B(n26559), .Z(n26550) );
  XNOR U28052 ( .A(n26551), .B(n26550), .Z(n26552) );
  XNOR U28053 ( .A(n26553), .B(n26552), .Z(n26582) );
  XNOR U28054 ( .A(sreg[1623]), .B(n26582), .Z(n26584) );
  NANDN U28055 ( .A(sreg[1622]), .B(n26545), .Z(n26549) );
  NAND U28056 ( .A(n26547), .B(n26546), .Z(n26548) );
  NAND U28057 ( .A(n26549), .B(n26548), .Z(n26583) );
  XNOR U28058 ( .A(n26584), .B(n26583), .Z(c[1623]) );
  NANDN U28059 ( .A(n26551), .B(n26550), .Z(n26555) );
  NANDN U28060 ( .A(n26553), .B(n26552), .Z(n26554) );
  AND U28061 ( .A(n26555), .B(n26554), .Z(n26590) );
  NANDN U28062 ( .A(n26557), .B(n26556), .Z(n26561) );
  NANDN U28063 ( .A(n26559), .B(n26558), .Z(n26560) );
  AND U28064 ( .A(n26561), .B(n26560), .Z(n26588) );
  NAND U28065 ( .A(n42143), .B(n26562), .Z(n26564) );
  XNOR U28066 ( .A(a[602]), .B(n4157), .Z(n26599) );
  NAND U28067 ( .A(n42144), .B(n26599), .Z(n26563) );
  AND U28068 ( .A(n26564), .B(n26563), .Z(n26614) );
  XOR U28069 ( .A(a[606]), .B(n42012), .Z(n26602) );
  XNOR U28070 ( .A(n26614), .B(n26613), .Z(n26616) );
  AND U28071 ( .A(a[608]), .B(b[0]), .Z(n26566) );
  XNOR U28072 ( .A(n26566), .B(n4071), .Z(n26568) );
  NANDN U28073 ( .A(b[0]), .B(a[607]), .Z(n26567) );
  NAND U28074 ( .A(n26568), .B(n26567), .Z(n26610) );
  XOR U28075 ( .A(a[604]), .B(n42085), .Z(n26603) );
  AND U28076 ( .A(a[600]), .B(b[7]), .Z(n26607) );
  XNOR U28077 ( .A(n26608), .B(n26607), .Z(n26609) );
  XNOR U28078 ( .A(n26610), .B(n26609), .Z(n26615) );
  XOR U28079 ( .A(n26616), .B(n26615), .Z(n26594) );
  NANDN U28080 ( .A(n26571), .B(n26570), .Z(n26575) );
  NANDN U28081 ( .A(n26573), .B(n26572), .Z(n26574) );
  AND U28082 ( .A(n26575), .B(n26574), .Z(n26593) );
  XNOR U28083 ( .A(n26594), .B(n26593), .Z(n26595) );
  NANDN U28084 ( .A(n26577), .B(n26576), .Z(n26581) );
  NAND U28085 ( .A(n26579), .B(n26578), .Z(n26580) );
  NAND U28086 ( .A(n26581), .B(n26580), .Z(n26596) );
  XNOR U28087 ( .A(n26595), .B(n26596), .Z(n26587) );
  XNOR U28088 ( .A(n26588), .B(n26587), .Z(n26589) );
  XNOR U28089 ( .A(n26590), .B(n26589), .Z(n26619) );
  XNOR U28090 ( .A(sreg[1624]), .B(n26619), .Z(n26621) );
  NANDN U28091 ( .A(sreg[1623]), .B(n26582), .Z(n26586) );
  NAND U28092 ( .A(n26584), .B(n26583), .Z(n26585) );
  NAND U28093 ( .A(n26586), .B(n26585), .Z(n26620) );
  XNOR U28094 ( .A(n26621), .B(n26620), .Z(c[1624]) );
  NANDN U28095 ( .A(n26588), .B(n26587), .Z(n26592) );
  NANDN U28096 ( .A(n26590), .B(n26589), .Z(n26591) );
  AND U28097 ( .A(n26592), .B(n26591), .Z(n26627) );
  NANDN U28098 ( .A(n26594), .B(n26593), .Z(n26598) );
  NANDN U28099 ( .A(n26596), .B(n26595), .Z(n26597) );
  AND U28100 ( .A(n26598), .B(n26597), .Z(n26625) );
  NAND U28101 ( .A(n42143), .B(n26599), .Z(n26601) );
  XNOR U28102 ( .A(a[603]), .B(n4158), .Z(n26636) );
  NAND U28103 ( .A(n42144), .B(n26636), .Z(n26600) );
  AND U28104 ( .A(n26601), .B(n26600), .Z(n26651) );
  XOR U28105 ( .A(a[607]), .B(n42012), .Z(n26639) );
  XNOR U28106 ( .A(n26651), .B(n26650), .Z(n26653) );
  XOR U28107 ( .A(a[605]), .B(n42085), .Z(n26640) );
  AND U28108 ( .A(a[601]), .B(b[7]), .Z(n26644) );
  XNOR U28109 ( .A(n26645), .B(n26644), .Z(n26646) );
  AND U28110 ( .A(a[609]), .B(b[0]), .Z(n26604) );
  XNOR U28111 ( .A(n26604), .B(n4071), .Z(n26606) );
  NANDN U28112 ( .A(b[0]), .B(a[608]), .Z(n26605) );
  NAND U28113 ( .A(n26606), .B(n26605), .Z(n26647) );
  XNOR U28114 ( .A(n26646), .B(n26647), .Z(n26652) );
  XOR U28115 ( .A(n26653), .B(n26652), .Z(n26631) );
  NANDN U28116 ( .A(n26608), .B(n26607), .Z(n26612) );
  NANDN U28117 ( .A(n26610), .B(n26609), .Z(n26611) );
  AND U28118 ( .A(n26612), .B(n26611), .Z(n26630) );
  XNOR U28119 ( .A(n26631), .B(n26630), .Z(n26632) );
  NANDN U28120 ( .A(n26614), .B(n26613), .Z(n26618) );
  NAND U28121 ( .A(n26616), .B(n26615), .Z(n26617) );
  NAND U28122 ( .A(n26618), .B(n26617), .Z(n26633) );
  XNOR U28123 ( .A(n26632), .B(n26633), .Z(n26624) );
  XNOR U28124 ( .A(n26625), .B(n26624), .Z(n26626) );
  XNOR U28125 ( .A(n26627), .B(n26626), .Z(n26656) );
  XNOR U28126 ( .A(sreg[1625]), .B(n26656), .Z(n26658) );
  NANDN U28127 ( .A(sreg[1624]), .B(n26619), .Z(n26623) );
  NAND U28128 ( .A(n26621), .B(n26620), .Z(n26622) );
  NAND U28129 ( .A(n26623), .B(n26622), .Z(n26657) );
  XNOR U28130 ( .A(n26658), .B(n26657), .Z(c[1625]) );
  NANDN U28131 ( .A(n26625), .B(n26624), .Z(n26629) );
  NANDN U28132 ( .A(n26627), .B(n26626), .Z(n26628) );
  AND U28133 ( .A(n26629), .B(n26628), .Z(n26664) );
  NANDN U28134 ( .A(n26631), .B(n26630), .Z(n26635) );
  NANDN U28135 ( .A(n26633), .B(n26632), .Z(n26634) );
  AND U28136 ( .A(n26635), .B(n26634), .Z(n26662) );
  NAND U28137 ( .A(n42143), .B(n26636), .Z(n26638) );
  XNOR U28138 ( .A(a[604]), .B(n4158), .Z(n26673) );
  NAND U28139 ( .A(n42144), .B(n26673), .Z(n26637) );
  AND U28140 ( .A(n26638), .B(n26637), .Z(n26688) );
  XOR U28141 ( .A(a[608]), .B(n42012), .Z(n26676) );
  XNOR U28142 ( .A(n26688), .B(n26687), .Z(n26690) );
  XOR U28143 ( .A(a[606]), .B(n42085), .Z(n26680) );
  AND U28144 ( .A(a[602]), .B(b[7]), .Z(n26681) );
  XNOR U28145 ( .A(n26682), .B(n26681), .Z(n26683) );
  AND U28146 ( .A(a[610]), .B(b[0]), .Z(n26641) );
  XNOR U28147 ( .A(n26641), .B(n4071), .Z(n26643) );
  NANDN U28148 ( .A(b[0]), .B(a[609]), .Z(n26642) );
  NAND U28149 ( .A(n26643), .B(n26642), .Z(n26684) );
  XNOR U28150 ( .A(n26683), .B(n26684), .Z(n26689) );
  XOR U28151 ( .A(n26690), .B(n26689), .Z(n26668) );
  NANDN U28152 ( .A(n26645), .B(n26644), .Z(n26649) );
  NANDN U28153 ( .A(n26647), .B(n26646), .Z(n26648) );
  AND U28154 ( .A(n26649), .B(n26648), .Z(n26667) );
  XNOR U28155 ( .A(n26668), .B(n26667), .Z(n26669) );
  NANDN U28156 ( .A(n26651), .B(n26650), .Z(n26655) );
  NAND U28157 ( .A(n26653), .B(n26652), .Z(n26654) );
  NAND U28158 ( .A(n26655), .B(n26654), .Z(n26670) );
  XNOR U28159 ( .A(n26669), .B(n26670), .Z(n26661) );
  XNOR U28160 ( .A(n26662), .B(n26661), .Z(n26663) );
  XNOR U28161 ( .A(n26664), .B(n26663), .Z(n26693) );
  XNOR U28162 ( .A(sreg[1626]), .B(n26693), .Z(n26695) );
  NANDN U28163 ( .A(sreg[1625]), .B(n26656), .Z(n26660) );
  NAND U28164 ( .A(n26658), .B(n26657), .Z(n26659) );
  NAND U28165 ( .A(n26660), .B(n26659), .Z(n26694) );
  XNOR U28166 ( .A(n26695), .B(n26694), .Z(c[1626]) );
  NANDN U28167 ( .A(n26662), .B(n26661), .Z(n26666) );
  NANDN U28168 ( .A(n26664), .B(n26663), .Z(n26665) );
  AND U28169 ( .A(n26666), .B(n26665), .Z(n26701) );
  NANDN U28170 ( .A(n26668), .B(n26667), .Z(n26672) );
  NANDN U28171 ( .A(n26670), .B(n26669), .Z(n26671) );
  AND U28172 ( .A(n26672), .B(n26671), .Z(n26699) );
  NAND U28173 ( .A(n42143), .B(n26673), .Z(n26675) );
  XNOR U28174 ( .A(a[605]), .B(n4158), .Z(n26710) );
  NAND U28175 ( .A(n42144), .B(n26710), .Z(n26674) );
  AND U28176 ( .A(n26675), .B(n26674), .Z(n26725) );
  XOR U28177 ( .A(a[609]), .B(n42012), .Z(n26713) );
  XNOR U28178 ( .A(n26725), .B(n26724), .Z(n26727) );
  AND U28179 ( .A(a[611]), .B(b[0]), .Z(n26677) );
  XNOR U28180 ( .A(n26677), .B(n4071), .Z(n26679) );
  NANDN U28181 ( .A(b[0]), .B(a[610]), .Z(n26678) );
  NAND U28182 ( .A(n26679), .B(n26678), .Z(n26721) );
  XOR U28183 ( .A(a[607]), .B(n42085), .Z(n26717) );
  AND U28184 ( .A(a[603]), .B(b[7]), .Z(n26718) );
  XNOR U28185 ( .A(n26719), .B(n26718), .Z(n26720) );
  XNOR U28186 ( .A(n26721), .B(n26720), .Z(n26726) );
  XOR U28187 ( .A(n26727), .B(n26726), .Z(n26705) );
  NANDN U28188 ( .A(n26682), .B(n26681), .Z(n26686) );
  NANDN U28189 ( .A(n26684), .B(n26683), .Z(n26685) );
  AND U28190 ( .A(n26686), .B(n26685), .Z(n26704) );
  XNOR U28191 ( .A(n26705), .B(n26704), .Z(n26706) );
  NANDN U28192 ( .A(n26688), .B(n26687), .Z(n26692) );
  NAND U28193 ( .A(n26690), .B(n26689), .Z(n26691) );
  NAND U28194 ( .A(n26692), .B(n26691), .Z(n26707) );
  XNOR U28195 ( .A(n26706), .B(n26707), .Z(n26698) );
  XNOR U28196 ( .A(n26699), .B(n26698), .Z(n26700) );
  XNOR U28197 ( .A(n26701), .B(n26700), .Z(n26730) );
  XNOR U28198 ( .A(sreg[1627]), .B(n26730), .Z(n26732) );
  NANDN U28199 ( .A(sreg[1626]), .B(n26693), .Z(n26697) );
  NAND U28200 ( .A(n26695), .B(n26694), .Z(n26696) );
  NAND U28201 ( .A(n26697), .B(n26696), .Z(n26731) );
  XNOR U28202 ( .A(n26732), .B(n26731), .Z(c[1627]) );
  NANDN U28203 ( .A(n26699), .B(n26698), .Z(n26703) );
  NANDN U28204 ( .A(n26701), .B(n26700), .Z(n26702) );
  AND U28205 ( .A(n26703), .B(n26702), .Z(n26738) );
  NANDN U28206 ( .A(n26705), .B(n26704), .Z(n26709) );
  NANDN U28207 ( .A(n26707), .B(n26706), .Z(n26708) );
  AND U28208 ( .A(n26709), .B(n26708), .Z(n26736) );
  NAND U28209 ( .A(n42143), .B(n26710), .Z(n26712) );
  XNOR U28210 ( .A(a[606]), .B(n4158), .Z(n26747) );
  NAND U28211 ( .A(n42144), .B(n26747), .Z(n26711) );
  AND U28212 ( .A(n26712), .B(n26711), .Z(n26762) );
  XOR U28213 ( .A(a[610]), .B(n42012), .Z(n26750) );
  XNOR U28214 ( .A(n26762), .B(n26761), .Z(n26764) );
  AND U28215 ( .A(a[612]), .B(b[0]), .Z(n26714) );
  XNOR U28216 ( .A(n26714), .B(n4071), .Z(n26716) );
  NANDN U28217 ( .A(b[0]), .B(a[611]), .Z(n26715) );
  NAND U28218 ( .A(n26716), .B(n26715), .Z(n26758) );
  XOR U28219 ( .A(a[608]), .B(n42085), .Z(n26751) );
  AND U28220 ( .A(a[604]), .B(b[7]), .Z(n26755) );
  XNOR U28221 ( .A(n26756), .B(n26755), .Z(n26757) );
  XNOR U28222 ( .A(n26758), .B(n26757), .Z(n26763) );
  XOR U28223 ( .A(n26764), .B(n26763), .Z(n26742) );
  NANDN U28224 ( .A(n26719), .B(n26718), .Z(n26723) );
  NANDN U28225 ( .A(n26721), .B(n26720), .Z(n26722) );
  AND U28226 ( .A(n26723), .B(n26722), .Z(n26741) );
  XNOR U28227 ( .A(n26742), .B(n26741), .Z(n26743) );
  NANDN U28228 ( .A(n26725), .B(n26724), .Z(n26729) );
  NAND U28229 ( .A(n26727), .B(n26726), .Z(n26728) );
  NAND U28230 ( .A(n26729), .B(n26728), .Z(n26744) );
  XNOR U28231 ( .A(n26743), .B(n26744), .Z(n26735) );
  XNOR U28232 ( .A(n26736), .B(n26735), .Z(n26737) );
  XNOR U28233 ( .A(n26738), .B(n26737), .Z(n26767) );
  XNOR U28234 ( .A(sreg[1628]), .B(n26767), .Z(n26769) );
  NANDN U28235 ( .A(sreg[1627]), .B(n26730), .Z(n26734) );
  NAND U28236 ( .A(n26732), .B(n26731), .Z(n26733) );
  NAND U28237 ( .A(n26734), .B(n26733), .Z(n26768) );
  XNOR U28238 ( .A(n26769), .B(n26768), .Z(c[1628]) );
  NANDN U28239 ( .A(n26736), .B(n26735), .Z(n26740) );
  NANDN U28240 ( .A(n26738), .B(n26737), .Z(n26739) );
  AND U28241 ( .A(n26740), .B(n26739), .Z(n26775) );
  NANDN U28242 ( .A(n26742), .B(n26741), .Z(n26746) );
  NANDN U28243 ( .A(n26744), .B(n26743), .Z(n26745) );
  AND U28244 ( .A(n26746), .B(n26745), .Z(n26773) );
  NAND U28245 ( .A(n42143), .B(n26747), .Z(n26749) );
  XNOR U28246 ( .A(a[607]), .B(n4158), .Z(n26784) );
  NAND U28247 ( .A(n42144), .B(n26784), .Z(n26748) );
  AND U28248 ( .A(n26749), .B(n26748), .Z(n26799) );
  XOR U28249 ( .A(a[611]), .B(n42012), .Z(n26787) );
  XNOR U28250 ( .A(n26799), .B(n26798), .Z(n26801) );
  XOR U28251 ( .A(a[609]), .B(n42085), .Z(n26788) );
  AND U28252 ( .A(a[605]), .B(b[7]), .Z(n26792) );
  XNOR U28253 ( .A(n26793), .B(n26792), .Z(n26794) );
  AND U28254 ( .A(a[613]), .B(b[0]), .Z(n26752) );
  XNOR U28255 ( .A(n26752), .B(n4071), .Z(n26754) );
  NANDN U28256 ( .A(b[0]), .B(a[612]), .Z(n26753) );
  NAND U28257 ( .A(n26754), .B(n26753), .Z(n26795) );
  XNOR U28258 ( .A(n26794), .B(n26795), .Z(n26800) );
  XOR U28259 ( .A(n26801), .B(n26800), .Z(n26779) );
  NANDN U28260 ( .A(n26756), .B(n26755), .Z(n26760) );
  NANDN U28261 ( .A(n26758), .B(n26757), .Z(n26759) );
  AND U28262 ( .A(n26760), .B(n26759), .Z(n26778) );
  XNOR U28263 ( .A(n26779), .B(n26778), .Z(n26780) );
  NANDN U28264 ( .A(n26762), .B(n26761), .Z(n26766) );
  NAND U28265 ( .A(n26764), .B(n26763), .Z(n26765) );
  NAND U28266 ( .A(n26766), .B(n26765), .Z(n26781) );
  XNOR U28267 ( .A(n26780), .B(n26781), .Z(n26772) );
  XNOR U28268 ( .A(n26773), .B(n26772), .Z(n26774) );
  XNOR U28269 ( .A(n26775), .B(n26774), .Z(n26804) );
  XNOR U28270 ( .A(sreg[1629]), .B(n26804), .Z(n26806) );
  NANDN U28271 ( .A(sreg[1628]), .B(n26767), .Z(n26771) );
  NAND U28272 ( .A(n26769), .B(n26768), .Z(n26770) );
  NAND U28273 ( .A(n26771), .B(n26770), .Z(n26805) );
  XNOR U28274 ( .A(n26806), .B(n26805), .Z(c[1629]) );
  NANDN U28275 ( .A(n26773), .B(n26772), .Z(n26777) );
  NANDN U28276 ( .A(n26775), .B(n26774), .Z(n26776) );
  AND U28277 ( .A(n26777), .B(n26776), .Z(n26812) );
  NANDN U28278 ( .A(n26779), .B(n26778), .Z(n26783) );
  NANDN U28279 ( .A(n26781), .B(n26780), .Z(n26782) );
  AND U28280 ( .A(n26783), .B(n26782), .Z(n26810) );
  NAND U28281 ( .A(n42143), .B(n26784), .Z(n26786) );
  XNOR U28282 ( .A(a[608]), .B(n4158), .Z(n26821) );
  NAND U28283 ( .A(n42144), .B(n26821), .Z(n26785) );
  AND U28284 ( .A(n26786), .B(n26785), .Z(n26836) );
  XOR U28285 ( .A(a[612]), .B(n42012), .Z(n26824) );
  XNOR U28286 ( .A(n26836), .B(n26835), .Z(n26838) );
  XOR U28287 ( .A(a[610]), .B(n42085), .Z(n26828) );
  AND U28288 ( .A(a[606]), .B(b[7]), .Z(n26829) );
  XNOR U28289 ( .A(n26830), .B(n26829), .Z(n26831) );
  AND U28290 ( .A(a[614]), .B(b[0]), .Z(n26789) );
  XNOR U28291 ( .A(n26789), .B(n4071), .Z(n26791) );
  NANDN U28292 ( .A(b[0]), .B(a[613]), .Z(n26790) );
  NAND U28293 ( .A(n26791), .B(n26790), .Z(n26832) );
  XNOR U28294 ( .A(n26831), .B(n26832), .Z(n26837) );
  XOR U28295 ( .A(n26838), .B(n26837), .Z(n26816) );
  NANDN U28296 ( .A(n26793), .B(n26792), .Z(n26797) );
  NANDN U28297 ( .A(n26795), .B(n26794), .Z(n26796) );
  AND U28298 ( .A(n26797), .B(n26796), .Z(n26815) );
  XNOR U28299 ( .A(n26816), .B(n26815), .Z(n26817) );
  NANDN U28300 ( .A(n26799), .B(n26798), .Z(n26803) );
  NAND U28301 ( .A(n26801), .B(n26800), .Z(n26802) );
  NAND U28302 ( .A(n26803), .B(n26802), .Z(n26818) );
  XNOR U28303 ( .A(n26817), .B(n26818), .Z(n26809) );
  XNOR U28304 ( .A(n26810), .B(n26809), .Z(n26811) );
  XNOR U28305 ( .A(n26812), .B(n26811), .Z(n26841) );
  XNOR U28306 ( .A(sreg[1630]), .B(n26841), .Z(n26843) );
  NANDN U28307 ( .A(sreg[1629]), .B(n26804), .Z(n26808) );
  NAND U28308 ( .A(n26806), .B(n26805), .Z(n26807) );
  NAND U28309 ( .A(n26808), .B(n26807), .Z(n26842) );
  XNOR U28310 ( .A(n26843), .B(n26842), .Z(c[1630]) );
  NANDN U28311 ( .A(n26810), .B(n26809), .Z(n26814) );
  NANDN U28312 ( .A(n26812), .B(n26811), .Z(n26813) );
  AND U28313 ( .A(n26814), .B(n26813), .Z(n26849) );
  NANDN U28314 ( .A(n26816), .B(n26815), .Z(n26820) );
  NANDN U28315 ( .A(n26818), .B(n26817), .Z(n26819) );
  AND U28316 ( .A(n26820), .B(n26819), .Z(n26847) );
  NAND U28317 ( .A(n42143), .B(n26821), .Z(n26823) );
  XNOR U28318 ( .A(a[609]), .B(n4158), .Z(n26858) );
  NAND U28319 ( .A(n42144), .B(n26858), .Z(n26822) );
  AND U28320 ( .A(n26823), .B(n26822), .Z(n26873) );
  XOR U28321 ( .A(a[613]), .B(n42012), .Z(n26861) );
  XNOR U28322 ( .A(n26873), .B(n26872), .Z(n26875) );
  AND U28323 ( .A(a[615]), .B(b[0]), .Z(n26825) );
  XNOR U28324 ( .A(n26825), .B(n4071), .Z(n26827) );
  NANDN U28325 ( .A(b[0]), .B(a[614]), .Z(n26826) );
  NAND U28326 ( .A(n26827), .B(n26826), .Z(n26869) );
  XOR U28327 ( .A(a[611]), .B(n42085), .Z(n26865) );
  AND U28328 ( .A(a[607]), .B(b[7]), .Z(n26866) );
  XNOR U28329 ( .A(n26867), .B(n26866), .Z(n26868) );
  XNOR U28330 ( .A(n26869), .B(n26868), .Z(n26874) );
  XOR U28331 ( .A(n26875), .B(n26874), .Z(n26853) );
  NANDN U28332 ( .A(n26830), .B(n26829), .Z(n26834) );
  NANDN U28333 ( .A(n26832), .B(n26831), .Z(n26833) );
  AND U28334 ( .A(n26834), .B(n26833), .Z(n26852) );
  XNOR U28335 ( .A(n26853), .B(n26852), .Z(n26854) );
  NANDN U28336 ( .A(n26836), .B(n26835), .Z(n26840) );
  NAND U28337 ( .A(n26838), .B(n26837), .Z(n26839) );
  NAND U28338 ( .A(n26840), .B(n26839), .Z(n26855) );
  XNOR U28339 ( .A(n26854), .B(n26855), .Z(n26846) );
  XNOR U28340 ( .A(n26847), .B(n26846), .Z(n26848) );
  XNOR U28341 ( .A(n26849), .B(n26848), .Z(n26878) );
  XNOR U28342 ( .A(sreg[1631]), .B(n26878), .Z(n26880) );
  NANDN U28343 ( .A(sreg[1630]), .B(n26841), .Z(n26845) );
  NAND U28344 ( .A(n26843), .B(n26842), .Z(n26844) );
  NAND U28345 ( .A(n26845), .B(n26844), .Z(n26879) );
  XNOR U28346 ( .A(n26880), .B(n26879), .Z(c[1631]) );
  NANDN U28347 ( .A(n26847), .B(n26846), .Z(n26851) );
  NANDN U28348 ( .A(n26849), .B(n26848), .Z(n26850) );
  AND U28349 ( .A(n26851), .B(n26850), .Z(n26886) );
  NANDN U28350 ( .A(n26853), .B(n26852), .Z(n26857) );
  NANDN U28351 ( .A(n26855), .B(n26854), .Z(n26856) );
  AND U28352 ( .A(n26857), .B(n26856), .Z(n26884) );
  NAND U28353 ( .A(n42143), .B(n26858), .Z(n26860) );
  XNOR U28354 ( .A(a[610]), .B(n4159), .Z(n26895) );
  NAND U28355 ( .A(n42144), .B(n26895), .Z(n26859) );
  AND U28356 ( .A(n26860), .B(n26859), .Z(n26910) );
  XOR U28357 ( .A(a[614]), .B(n42012), .Z(n26898) );
  XNOR U28358 ( .A(n26910), .B(n26909), .Z(n26912) );
  NAND U28359 ( .A(a[616]), .B(b[0]), .Z(n26862) );
  XNOR U28360 ( .A(b[1]), .B(n26862), .Z(n26864) );
  NANDN U28361 ( .A(b[0]), .B(a[615]), .Z(n26863) );
  AND U28362 ( .A(n26864), .B(n26863), .Z(n26905) );
  XOR U28363 ( .A(a[612]), .B(n42085), .Z(n26902) );
  AND U28364 ( .A(a[608]), .B(b[7]), .Z(n26903) );
  XOR U28365 ( .A(n26904), .B(n26903), .Z(n26906) );
  XNOR U28366 ( .A(n26905), .B(n26906), .Z(n26911) );
  XOR U28367 ( .A(n26912), .B(n26911), .Z(n26890) );
  NANDN U28368 ( .A(n26867), .B(n26866), .Z(n26871) );
  NANDN U28369 ( .A(n26869), .B(n26868), .Z(n26870) );
  AND U28370 ( .A(n26871), .B(n26870), .Z(n26889) );
  XNOR U28371 ( .A(n26890), .B(n26889), .Z(n26891) );
  NANDN U28372 ( .A(n26873), .B(n26872), .Z(n26877) );
  NAND U28373 ( .A(n26875), .B(n26874), .Z(n26876) );
  NAND U28374 ( .A(n26877), .B(n26876), .Z(n26892) );
  XNOR U28375 ( .A(n26891), .B(n26892), .Z(n26883) );
  XNOR U28376 ( .A(n26884), .B(n26883), .Z(n26885) );
  XNOR U28377 ( .A(n26886), .B(n26885), .Z(n26915) );
  XNOR U28378 ( .A(sreg[1632]), .B(n26915), .Z(n26917) );
  NANDN U28379 ( .A(sreg[1631]), .B(n26878), .Z(n26882) );
  NAND U28380 ( .A(n26880), .B(n26879), .Z(n26881) );
  NAND U28381 ( .A(n26882), .B(n26881), .Z(n26916) );
  XNOR U28382 ( .A(n26917), .B(n26916), .Z(c[1632]) );
  NANDN U28383 ( .A(n26884), .B(n26883), .Z(n26888) );
  NANDN U28384 ( .A(n26886), .B(n26885), .Z(n26887) );
  AND U28385 ( .A(n26888), .B(n26887), .Z(n26923) );
  NANDN U28386 ( .A(n26890), .B(n26889), .Z(n26894) );
  NANDN U28387 ( .A(n26892), .B(n26891), .Z(n26893) );
  AND U28388 ( .A(n26894), .B(n26893), .Z(n26921) );
  NAND U28389 ( .A(n42143), .B(n26895), .Z(n26897) );
  XNOR U28390 ( .A(a[611]), .B(n4159), .Z(n26932) );
  NAND U28391 ( .A(n42144), .B(n26932), .Z(n26896) );
  AND U28392 ( .A(n26897), .B(n26896), .Z(n26947) );
  XOR U28393 ( .A(a[615]), .B(n42012), .Z(n26935) );
  XNOR U28394 ( .A(n26947), .B(n26946), .Z(n26949) );
  AND U28395 ( .A(a[617]), .B(b[0]), .Z(n26899) );
  XNOR U28396 ( .A(n26899), .B(n4071), .Z(n26901) );
  NANDN U28397 ( .A(b[0]), .B(a[616]), .Z(n26900) );
  NAND U28398 ( .A(n26901), .B(n26900), .Z(n26943) );
  XOR U28399 ( .A(a[613]), .B(n42085), .Z(n26939) );
  AND U28400 ( .A(a[609]), .B(b[7]), .Z(n26940) );
  XNOR U28401 ( .A(n26941), .B(n26940), .Z(n26942) );
  XNOR U28402 ( .A(n26943), .B(n26942), .Z(n26948) );
  XOR U28403 ( .A(n26949), .B(n26948), .Z(n26927) );
  NANDN U28404 ( .A(n26904), .B(n26903), .Z(n26908) );
  NANDN U28405 ( .A(n26906), .B(n26905), .Z(n26907) );
  AND U28406 ( .A(n26908), .B(n26907), .Z(n26926) );
  XNOR U28407 ( .A(n26927), .B(n26926), .Z(n26928) );
  NANDN U28408 ( .A(n26910), .B(n26909), .Z(n26914) );
  NAND U28409 ( .A(n26912), .B(n26911), .Z(n26913) );
  NAND U28410 ( .A(n26914), .B(n26913), .Z(n26929) );
  XNOR U28411 ( .A(n26928), .B(n26929), .Z(n26920) );
  XNOR U28412 ( .A(n26921), .B(n26920), .Z(n26922) );
  XNOR U28413 ( .A(n26923), .B(n26922), .Z(n26952) );
  XNOR U28414 ( .A(sreg[1633]), .B(n26952), .Z(n26954) );
  NANDN U28415 ( .A(sreg[1632]), .B(n26915), .Z(n26919) );
  NAND U28416 ( .A(n26917), .B(n26916), .Z(n26918) );
  NAND U28417 ( .A(n26919), .B(n26918), .Z(n26953) );
  XNOR U28418 ( .A(n26954), .B(n26953), .Z(c[1633]) );
  NANDN U28419 ( .A(n26921), .B(n26920), .Z(n26925) );
  NANDN U28420 ( .A(n26923), .B(n26922), .Z(n26924) );
  AND U28421 ( .A(n26925), .B(n26924), .Z(n26960) );
  NANDN U28422 ( .A(n26927), .B(n26926), .Z(n26931) );
  NANDN U28423 ( .A(n26929), .B(n26928), .Z(n26930) );
  AND U28424 ( .A(n26931), .B(n26930), .Z(n26958) );
  NAND U28425 ( .A(n42143), .B(n26932), .Z(n26934) );
  XNOR U28426 ( .A(a[612]), .B(n4159), .Z(n26969) );
  NAND U28427 ( .A(n42144), .B(n26969), .Z(n26933) );
  AND U28428 ( .A(n26934), .B(n26933), .Z(n26984) );
  XOR U28429 ( .A(a[616]), .B(n42012), .Z(n26972) );
  XNOR U28430 ( .A(n26984), .B(n26983), .Z(n26986) );
  AND U28431 ( .A(a[618]), .B(b[0]), .Z(n26936) );
  XNOR U28432 ( .A(n26936), .B(n4071), .Z(n26938) );
  NANDN U28433 ( .A(b[0]), .B(a[617]), .Z(n26937) );
  NAND U28434 ( .A(n26938), .B(n26937), .Z(n26980) );
  XOR U28435 ( .A(a[614]), .B(n42085), .Z(n26976) );
  AND U28436 ( .A(a[610]), .B(b[7]), .Z(n26977) );
  XNOR U28437 ( .A(n26978), .B(n26977), .Z(n26979) );
  XNOR U28438 ( .A(n26980), .B(n26979), .Z(n26985) );
  XOR U28439 ( .A(n26986), .B(n26985), .Z(n26964) );
  NANDN U28440 ( .A(n26941), .B(n26940), .Z(n26945) );
  NANDN U28441 ( .A(n26943), .B(n26942), .Z(n26944) );
  AND U28442 ( .A(n26945), .B(n26944), .Z(n26963) );
  XNOR U28443 ( .A(n26964), .B(n26963), .Z(n26965) );
  NANDN U28444 ( .A(n26947), .B(n26946), .Z(n26951) );
  NAND U28445 ( .A(n26949), .B(n26948), .Z(n26950) );
  NAND U28446 ( .A(n26951), .B(n26950), .Z(n26966) );
  XNOR U28447 ( .A(n26965), .B(n26966), .Z(n26957) );
  XNOR U28448 ( .A(n26958), .B(n26957), .Z(n26959) );
  XNOR U28449 ( .A(n26960), .B(n26959), .Z(n26989) );
  XNOR U28450 ( .A(sreg[1634]), .B(n26989), .Z(n26991) );
  NANDN U28451 ( .A(sreg[1633]), .B(n26952), .Z(n26956) );
  NAND U28452 ( .A(n26954), .B(n26953), .Z(n26955) );
  NAND U28453 ( .A(n26956), .B(n26955), .Z(n26990) );
  XNOR U28454 ( .A(n26991), .B(n26990), .Z(c[1634]) );
  NANDN U28455 ( .A(n26958), .B(n26957), .Z(n26962) );
  NANDN U28456 ( .A(n26960), .B(n26959), .Z(n26961) );
  AND U28457 ( .A(n26962), .B(n26961), .Z(n26997) );
  NANDN U28458 ( .A(n26964), .B(n26963), .Z(n26968) );
  NANDN U28459 ( .A(n26966), .B(n26965), .Z(n26967) );
  AND U28460 ( .A(n26968), .B(n26967), .Z(n26995) );
  NAND U28461 ( .A(n42143), .B(n26969), .Z(n26971) );
  XNOR U28462 ( .A(a[613]), .B(n4159), .Z(n27006) );
  NAND U28463 ( .A(n42144), .B(n27006), .Z(n26970) );
  AND U28464 ( .A(n26971), .B(n26970), .Z(n27021) );
  XOR U28465 ( .A(a[617]), .B(n42012), .Z(n27009) );
  XNOR U28466 ( .A(n27021), .B(n27020), .Z(n27023) );
  AND U28467 ( .A(a[619]), .B(b[0]), .Z(n26973) );
  XNOR U28468 ( .A(n26973), .B(n4071), .Z(n26975) );
  NANDN U28469 ( .A(b[0]), .B(a[618]), .Z(n26974) );
  NAND U28470 ( .A(n26975), .B(n26974), .Z(n27017) );
  XOR U28471 ( .A(a[615]), .B(n42085), .Z(n27010) );
  AND U28472 ( .A(a[611]), .B(b[7]), .Z(n27014) );
  XNOR U28473 ( .A(n27015), .B(n27014), .Z(n27016) );
  XNOR U28474 ( .A(n27017), .B(n27016), .Z(n27022) );
  XOR U28475 ( .A(n27023), .B(n27022), .Z(n27001) );
  NANDN U28476 ( .A(n26978), .B(n26977), .Z(n26982) );
  NANDN U28477 ( .A(n26980), .B(n26979), .Z(n26981) );
  AND U28478 ( .A(n26982), .B(n26981), .Z(n27000) );
  XNOR U28479 ( .A(n27001), .B(n27000), .Z(n27002) );
  NANDN U28480 ( .A(n26984), .B(n26983), .Z(n26988) );
  NAND U28481 ( .A(n26986), .B(n26985), .Z(n26987) );
  NAND U28482 ( .A(n26988), .B(n26987), .Z(n27003) );
  XNOR U28483 ( .A(n27002), .B(n27003), .Z(n26994) );
  XNOR U28484 ( .A(n26995), .B(n26994), .Z(n26996) );
  XNOR U28485 ( .A(n26997), .B(n26996), .Z(n27026) );
  XNOR U28486 ( .A(sreg[1635]), .B(n27026), .Z(n27028) );
  NANDN U28487 ( .A(sreg[1634]), .B(n26989), .Z(n26993) );
  NAND U28488 ( .A(n26991), .B(n26990), .Z(n26992) );
  NAND U28489 ( .A(n26993), .B(n26992), .Z(n27027) );
  XNOR U28490 ( .A(n27028), .B(n27027), .Z(c[1635]) );
  NANDN U28491 ( .A(n26995), .B(n26994), .Z(n26999) );
  NANDN U28492 ( .A(n26997), .B(n26996), .Z(n26998) );
  AND U28493 ( .A(n26999), .B(n26998), .Z(n27034) );
  NANDN U28494 ( .A(n27001), .B(n27000), .Z(n27005) );
  NANDN U28495 ( .A(n27003), .B(n27002), .Z(n27004) );
  AND U28496 ( .A(n27005), .B(n27004), .Z(n27032) );
  NAND U28497 ( .A(n42143), .B(n27006), .Z(n27008) );
  XNOR U28498 ( .A(a[614]), .B(n4159), .Z(n27043) );
  NAND U28499 ( .A(n42144), .B(n27043), .Z(n27007) );
  AND U28500 ( .A(n27008), .B(n27007), .Z(n27058) );
  XOR U28501 ( .A(a[618]), .B(n42012), .Z(n27046) );
  XNOR U28502 ( .A(n27058), .B(n27057), .Z(n27060) );
  XOR U28503 ( .A(a[616]), .B(n42085), .Z(n27050) );
  AND U28504 ( .A(a[612]), .B(b[7]), .Z(n27051) );
  XNOR U28505 ( .A(n27052), .B(n27051), .Z(n27053) );
  AND U28506 ( .A(a[620]), .B(b[0]), .Z(n27011) );
  XNOR U28507 ( .A(n27011), .B(n4071), .Z(n27013) );
  NANDN U28508 ( .A(b[0]), .B(a[619]), .Z(n27012) );
  NAND U28509 ( .A(n27013), .B(n27012), .Z(n27054) );
  XNOR U28510 ( .A(n27053), .B(n27054), .Z(n27059) );
  XOR U28511 ( .A(n27060), .B(n27059), .Z(n27038) );
  NANDN U28512 ( .A(n27015), .B(n27014), .Z(n27019) );
  NANDN U28513 ( .A(n27017), .B(n27016), .Z(n27018) );
  AND U28514 ( .A(n27019), .B(n27018), .Z(n27037) );
  XNOR U28515 ( .A(n27038), .B(n27037), .Z(n27039) );
  NANDN U28516 ( .A(n27021), .B(n27020), .Z(n27025) );
  NAND U28517 ( .A(n27023), .B(n27022), .Z(n27024) );
  NAND U28518 ( .A(n27025), .B(n27024), .Z(n27040) );
  XNOR U28519 ( .A(n27039), .B(n27040), .Z(n27031) );
  XNOR U28520 ( .A(n27032), .B(n27031), .Z(n27033) );
  XNOR U28521 ( .A(n27034), .B(n27033), .Z(n27063) );
  XNOR U28522 ( .A(sreg[1636]), .B(n27063), .Z(n27065) );
  NANDN U28523 ( .A(sreg[1635]), .B(n27026), .Z(n27030) );
  NAND U28524 ( .A(n27028), .B(n27027), .Z(n27029) );
  NAND U28525 ( .A(n27030), .B(n27029), .Z(n27064) );
  XNOR U28526 ( .A(n27065), .B(n27064), .Z(c[1636]) );
  NANDN U28527 ( .A(n27032), .B(n27031), .Z(n27036) );
  NANDN U28528 ( .A(n27034), .B(n27033), .Z(n27035) );
  AND U28529 ( .A(n27036), .B(n27035), .Z(n27071) );
  NANDN U28530 ( .A(n27038), .B(n27037), .Z(n27042) );
  NANDN U28531 ( .A(n27040), .B(n27039), .Z(n27041) );
  AND U28532 ( .A(n27042), .B(n27041), .Z(n27069) );
  NAND U28533 ( .A(n42143), .B(n27043), .Z(n27045) );
  XNOR U28534 ( .A(a[615]), .B(n4159), .Z(n27080) );
  NAND U28535 ( .A(n42144), .B(n27080), .Z(n27044) );
  AND U28536 ( .A(n27045), .B(n27044), .Z(n27095) );
  XOR U28537 ( .A(a[619]), .B(n42012), .Z(n27083) );
  XNOR U28538 ( .A(n27095), .B(n27094), .Z(n27097) );
  AND U28539 ( .A(a[621]), .B(b[0]), .Z(n27047) );
  XNOR U28540 ( .A(n27047), .B(n4071), .Z(n27049) );
  NANDN U28541 ( .A(b[0]), .B(a[620]), .Z(n27048) );
  NAND U28542 ( .A(n27049), .B(n27048), .Z(n27091) );
  XOR U28543 ( .A(a[617]), .B(n42085), .Z(n27084) );
  AND U28544 ( .A(a[613]), .B(b[7]), .Z(n27088) );
  XNOR U28545 ( .A(n27089), .B(n27088), .Z(n27090) );
  XNOR U28546 ( .A(n27091), .B(n27090), .Z(n27096) );
  XOR U28547 ( .A(n27097), .B(n27096), .Z(n27075) );
  NANDN U28548 ( .A(n27052), .B(n27051), .Z(n27056) );
  NANDN U28549 ( .A(n27054), .B(n27053), .Z(n27055) );
  AND U28550 ( .A(n27056), .B(n27055), .Z(n27074) );
  XNOR U28551 ( .A(n27075), .B(n27074), .Z(n27076) );
  NANDN U28552 ( .A(n27058), .B(n27057), .Z(n27062) );
  NAND U28553 ( .A(n27060), .B(n27059), .Z(n27061) );
  NAND U28554 ( .A(n27062), .B(n27061), .Z(n27077) );
  XNOR U28555 ( .A(n27076), .B(n27077), .Z(n27068) );
  XNOR U28556 ( .A(n27069), .B(n27068), .Z(n27070) );
  XNOR U28557 ( .A(n27071), .B(n27070), .Z(n27100) );
  XNOR U28558 ( .A(sreg[1637]), .B(n27100), .Z(n27102) );
  NANDN U28559 ( .A(sreg[1636]), .B(n27063), .Z(n27067) );
  NAND U28560 ( .A(n27065), .B(n27064), .Z(n27066) );
  NAND U28561 ( .A(n27067), .B(n27066), .Z(n27101) );
  XNOR U28562 ( .A(n27102), .B(n27101), .Z(c[1637]) );
  NANDN U28563 ( .A(n27069), .B(n27068), .Z(n27073) );
  NANDN U28564 ( .A(n27071), .B(n27070), .Z(n27072) );
  AND U28565 ( .A(n27073), .B(n27072), .Z(n27108) );
  NANDN U28566 ( .A(n27075), .B(n27074), .Z(n27079) );
  NANDN U28567 ( .A(n27077), .B(n27076), .Z(n27078) );
  AND U28568 ( .A(n27079), .B(n27078), .Z(n27106) );
  NAND U28569 ( .A(n42143), .B(n27080), .Z(n27082) );
  XNOR U28570 ( .A(a[616]), .B(n4159), .Z(n27117) );
  NAND U28571 ( .A(n42144), .B(n27117), .Z(n27081) );
  AND U28572 ( .A(n27082), .B(n27081), .Z(n27132) );
  XOR U28573 ( .A(a[620]), .B(n42012), .Z(n27120) );
  XNOR U28574 ( .A(n27132), .B(n27131), .Z(n27134) );
  XOR U28575 ( .A(a[618]), .B(n42085), .Z(n27124) );
  AND U28576 ( .A(a[614]), .B(b[7]), .Z(n27125) );
  XNOR U28577 ( .A(n27126), .B(n27125), .Z(n27127) );
  AND U28578 ( .A(a[622]), .B(b[0]), .Z(n27085) );
  XNOR U28579 ( .A(n27085), .B(n4071), .Z(n27087) );
  NANDN U28580 ( .A(b[0]), .B(a[621]), .Z(n27086) );
  NAND U28581 ( .A(n27087), .B(n27086), .Z(n27128) );
  XNOR U28582 ( .A(n27127), .B(n27128), .Z(n27133) );
  XOR U28583 ( .A(n27134), .B(n27133), .Z(n27112) );
  NANDN U28584 ( .A(n27089), .B(n27088), .Z(n27093) );
  NANDN U28585 ( .A(n27091), .B(n27090), .Z(n27092) );
  AND U28586 ( .A(n27093), .B(n27092), .Z(n27111) );
  XNOR U28587 ( .A(n27112), .B(n27111), .Z(n27113) );
  NANDN U28588 ( .A(n27095), .B(n27094), .Z(n27099) );
  NAND U28589 ( .A(n27097), .B(n27096), .Z(n27098) );
  NAND U28590 ( .A(n27099), .B(n27098), .Z(n27114) );
  XNOR U28591 ( .A(n27113), .B(n27114), .Z(n27105) );
  XNOR U28592 ( .A(n27106), .B(n27105), .Z(n27107) );
  XNOR U28593 ( .A(n27108), .B(n27107), .Z(n27137) );
  XNOR U28594 ( .A(sreg[1638]), .B(n27137), .Z(n27139) );
  NANDN U28595 ( .A(sreg[1637]), .B(n27100), .Z(n27104) );
  NAND U28596 ( .A(n27102), .B(n27101), .Z(n27103) );
  NAND U28597 ( .A(n27104), .B(n27103), .Z(n27138) );
  XNOR U28598 ( .A(n27139), .B(n27138), .Z(c[1638]) );
  NANDN U28599 ( .A(n27106), .B(n27105), .Z(n27110) );
  NANDN U28600 ( .A(n27108), .B(n27107), .Z(n27109) );
  AND U28601 ( .A(n27110), .B(n27109), .Z(n27145) );
  NANDN U28602 ( .A(n27112), .B(n27111), .Z(n27116) );
  NANDN U28603 ( .A(n27114), .B(n27113), .Z(n27115) );
  AND U28604 ( .A(n27116), .B(n27115), .Z(n27143) );
  NAND U28605 ( .A(n42143), .B(n27117), .Z(n27119) );
  XNOR U28606 ( .A(a[617]), .B(n4160), .Z(n27154) );
  NAND U28607 ( .A(n42144), .B(n27154), .Z(n27118) );
  AND U28608 ( .A(n27119), .B(n27118), .Z(n27169) );
  XOR U28609 ( .A(a[621]), .B(n42012), .Z(n27157) );
  XNOR U28610 ( .A(n27169), .B(n27168), .Z(n27171) );
  AND U28611 ( .A(a[623]), .B(b[0]), .Z(n27121) );
  XNOR U28612 ( .A(n27121), .B(n4071), .Z(n27123) );
  NANDN U28613 ( .A(b[0]), .B(a[622]), .Z(n27122) );
  NAND U28614 ( .A(n27123), .B(n27122), .Z(n27165) );
  XOR U28615 ( .A(a[619]), .B(n42085), .Z(n27158) );
  AND U28616 ( .A(a[615]), .B(b[7]), .Z(n27162) );
  XNOR U28617 ( .A(n27163), .B(n27162), .Z(n27164) );
  XNOR U28618 ( .A(n27165), .B(n27164), .Z(n27170) );
  XOR U28619 ( .A(n27171), .B(n27170), .Z(n27149) );
  NANDN U28620 ( .A(n27126), .B(n27125), .Z(n27130) );
  NANDN U28621 ( .A(n27128), .B(n27127), .Z(n27129) );
  AND U28622 ( .A(n27130), .B(n27129), .Z(n27148) );
  XNOR U28623 ( .A(n27149), .B(n27148), .Z(n27150) );
  NANDN U28624 ( .A(n27132), .B(n27131), .Z(n27136) );
  NAND U28625 ( .A(n27134), .B(n27133), .Z(n27135) );
  NAND U28626 ( .A(n27136), .B(n27135), .Z(n27151) );
  XNOR U28627 ( .A(n27150), .B(n27151), .Z(n27142) );
  XNOR U28628 ( .A(n27143), .B(n27142), .Z(n27144) );
  XNOR U28629 ( .A(n27145), .B(n27144), .Z(n27174) );
  XNOR U28630 ( .A(sreg[1639]), .B(n27174), .Z(n27176) );
  NANDN U28631 ( .A(sreg[1638]), .B(n27137), .Z(n27141) );
  NAND U28632 ( .A(n27139), .B(n27138), .Z(n27140) );
  NAND U28633 ( .A(n27141), .B(n27140), .Z(n27175) );
  XNOR U28634 ( .A(n27176), .B(n27175), .Z(c[1639]) );
  NANDN U28635 ( .A(n27143), .B(n27142), .Z(n27147) );
  NANDN U28636 ( .A(n27145), .B(n27144), .Z(n27146) );
  AND U28637 ( .A(n27147), .B(n27146), .Z(n27182) );
  NANDN U28638 ( .A(n27149), .B(n27148), .Z(n27153) );
  NANDN U28639 ( .A(n27151), .B(n27150), .Z(n27152) );
  AND U28640 ( .A(n27153), .B(n27152), .Z(n27180) );
  NAND U28641 ( .A(n42143), .B(n27154), .Z(n27156) );
  XNOR U28642 ( .A(a[618]), .B(n4160), .Z(n27191) );
  NAND U28643 ( .A(n42144), .B(n27191), .Z(n27155) );
  AND U28644 ( .A(n27156), .B(n27155), .Z(n27206) );
  XOR U28645 ( .A(a[622]), .B(n42012), .Z(n27194) );
  XNOR U28646 ( .A(n27206), .B(n27205), .Z(n27208) );
  XOR U28647 ( .A(a[620]), .B(n42085), .Z(n27198) );
  AND U28648 ( .A(a[616]), .B(b[7]), .Z(n27199) );
  XNOR U28649 ( .A(n27200), .B(n27199), .Z(n27201) );
  AND U28650 ( .A(a[624]), .B(b[0]), .Z(n27159) );
  XNOR U28651 ( .A(n27159), .B(n4071), .Z(n27161) );
  NANDN U28652 ( .A(b[0]), .B(a[623]), .Z(n27160) );
  NAND U28653 ( .A(n27161), .B(n27160), .Z(n27202) );
  XNOR U28654 ( .A(n27201), .B(n27202), .Z(n27207) );
  XOR U28655 ( .A(n27208), .B(n27207), .Z(n27186) );
  NANDN U28656 ( .A(n27163), .B(n27162), .Z(n27167) );
  NANDN U28657 ( .A(n27165), .B(n27164), .Z(n27166) );
  AND U28658 ( .A(n27167), .B(n27166), .Z(n27185) );
  XNOR U28659 ( .A(n27186), .B(n27185), .Z(n27187) );
  NANDN U28660 ( .A(n27169), .B(n27168), .Z(n27173) );
  NAND U28661 ( .A(n27171), .B(n27170), .Z(n27172) );
  NAND U28662 ( .A(n27173), .B(n27172), .Z(n27188) );
  XNOR U28663 ( .A(n27187), .B(n27188), .Z(n27179) );
  XNOR U28664 ( .A(n27180), .B(n27179), .Z(n27181) );
  XNOR U28665 ( .A(n27182), .B(n27181), .Z(n27211) );
  XNOR U28666 ( .A(sreg[1640]), .B(n27211), .Z(n27213) );
  NANDN U28667 ( .A(sreg[1639]), .B(n27174), .Z(n27178) );
  NAND U28668 ( .A(n27176), .B(n27175), .Z(n27177) );
  NAND U28669 ( .A(n27178), .B(n27177), .Z(n27212) );
  XNOR U28670 ( .A(n27213), .B(n27212), .Z(c[1640]) );
  NANDN U28671 ( .A(n27180), .B(n27179), .Z(n27184) );
  NANDN U28672 ( .A(n27182), .B(n27181), .Z(n27183) );
  AND U28673 ( .A(n27184), .B(n27183), .Z(n27219) );
  NANDN U28674 ( .A(n27186), .B(n27185), .Z(n27190) );
  NANDN U28675 ( .A(n27188), .B(n27187), .Z(n27189) );
  AND U28676 ( .A(n27190), .B(n27189), .Z(n27217) );
  NAND U28677 ( .A(n42143), .B(n27191), .Z(n27193) );
  XNOR U28678 ( .A(a[619]), .B(n4160), .Z(n27228) );
  NAND U28679 ( .A(n42144), .B(n27228), .Z(n27192) );
  AND U28680 ( .A(n27193), .B(n27192), .Z(n27243) );
  XOR U28681 ( .A(a[623]), .B(n42012), .Z(n27231) );
  XNOR U28682 ( .A(n27243), .B(n27242), .Z(n27245) );
  AND U28683 ( .A(a[625]), .B(b[0]), .Z(n27195) );
  XNOR U28684 ( .A(n27195), .B(n4071), .Z(n27197) );
  NANDN U28685 ( .A(b[0]), .B(a[624]), .Z(n27196) );
  NAND U28686 ( .A(n27197), .B(n27196), .Z(n27239) );
  XOR U28687 ( .A(a[621]), .B(n42085), .Z(n27235) );
  AND U28688 ( .A(a[617]), .B(b[7]), .Z(n27236) );
  XNOR U28689 ( .A(n27237), .B(n27236), .Z(n27238) );
  XNOR U28690 ( .A(n27239), .B(n27238), .Z(n27244) );
  XOR U28691 ( .A(n27245), .B(n27244), .Z(n27223) );
  NANDN U28692 ( .A(n27200), .B(n27199), .Z(n27204) );
  NANDN U28693 ( .A(n27202), .B(n27201), .Z(n27203) );
  AND U28694 ( .A(n27204), .B(n27203), .Z(n27222) );
  XNOR U28695 ( .A(n27223), .B(n27222), .Z(n27224) );
  NANDN U28696 ( .A(n27206), .B(n27205), .Z(n27210) );
  NAND U28697 ( .A(n27208), .B(n27207), .Z(n27209) );
  NAND U28698 ( .A(n27210), .B(n27209), .Z(n27225) );
  XNOR U28699 ( .A(n27224), .B(n27225), .Z(n27216) );
  XNOR U28700 ( .A(n27217), .B(n27216), .Z(n27218) );
  XNOR U28701 ( .A(n27219), .B(n27218), .Z(n27248) );
  XNOR U28702 ( .A(sreg[1641]), .B(n27248), .Z(n27250) );
  NANDN U28703 ( .A(sreg[1640]), .B(n27211), .Z(n27215) );
  NAND U28704 ( .A(n27213), .B(n27212), .Z(n27214) );
  NAND U28705 ( .A(n27215), .B(n27214), .Z(n27249) );
  XNOR U28706 ( .A(n27250), .B(n27249), .Z(c[1641]) );
  NANDN U28707 ( .A(n27217), .B(n27216), .Z(n27221) );
  NANDN U28708 ( .A(n27219), .B(n27218), .Z(n27220) );
  AND U28709 ( .A(n27221), .B(n27220), .Z(n27256) );
  NANDN U28710 ( .A(n27223), .B(n27222), .Z(n27227) );
  NANDN U28711 ( .A(n27225), .B(n27224), .Z(n27226) );
  AND U28712 ( .A(n27227), .B(n27226), .Z(n27254) );
  NAND U28713 ( .A(n42143), .B(n27228), .Z(n27230) );
  XNOR U28714 ( .A(a[620]), .B(n4160), .Z(n27265) );
  NAND U28715 ( .A(n42144), .B(n27265), .Z(n27229) );
  AND U28716 ( .A(n27230), .B(n27229), .Z(n27280) );
  XOR U28717 ( .A(a[624]), .B(n42012), .Z(n27268) );
  XNOR U28718 ( .A(n27280), .B(n27279), .Z(n27282) );
  AND U28719 ( .A(a[626]), .B(b[0]), .Z(n27232) );
  XNOR U28720 ( .A(n27232), .B(n4071), .Z(n27234) );
  NANDN U28721 ( .A(b[0]), .B(a[625]), .Z(n27233) );
  NAND U28722 ( .A(n27234), .B(n27233), .Z(n27276) );
  XOR U28723 ( .A(a[622]), .B(n42085), .Z(n27272) );
  AND U28724 ( .A(a[618]), .B(b[7]), .Z(n27273) );
  XNOR U28725 ( .A(n27274), .B(n27273), .Z(n27275) );
  XNOR U28726 ( .A(n27276), .B(n27275), .Z(n27281) );
  XOR U28727 ( .A(n27282), .B(n27281), .Z(n27260) );
  NANDN U28728 ( .A(n27237), .B(n27236), .Z(n27241) );
  NANDN U28729 ( .A(n27239), .B(n27238), .Z(n27240) );
  AND U28730 ( .A(n27241), .B(n27240), .Z(n27259) );
  XNOR U28731 ( .A(n27260), .B(n27259), .Z(n27261) );
  NANDN U28732 ( .A(n27243), .B(n27242), .Z(n27247) );
  NAND U28733 ( .A(n27245), .B(n27244), .Z(n27246) );
  NAND U28734 ( .A(n27247), .B(n27246), .Z(n27262) );
  XNOR U28735 ( .A(n27261), .B(n27262), .Z(n27253) );
  XNOR U28736 ( .A(n27254), .B(n27253), .Z(n27255) );
  XNOR U28737 ( .A(n27256), .B(n27255), .Z(n27285) );
  XNOR U28738 ( .A(sreg[1642]), .B(n27285), .Z(n27287) );
  NANDN U28739 ( .A(sreg[1641]), .B(n27248), .Z(n27252) );
  NAND U28740 ( .A(n27250), .B(n27249), .Z(n27251) );
  NAND U28741 ( .A(n27252), .B(n27251), .Z(n27286) );
  XNOR U28742 ( .A(n27287), .B(n27286), .Z(c[1642]) );
  NANDN U28743 ( .A(n27254), .B(n27253), .Z(n27258) );
  NANDN U28744 ( .A(n27256), .B(n27255), .Z(n27257) );
  AND U28745 ( .A(n27258), .B(n27257), .Z(n27293) );
  NANDN U28746 ( .A(n27260), .B(n27259), .Z(n27264) );
  NANDN U28747 ( .A(n27262), .B(n27261), .Z(n27263) );
  AND U28748 ( .A(n27264), .B(n27263), .Z(n27291) );
  NAND U28749 ( .A(n42143), .B(n27265), .Z(n27267) );
  XNOR U28750 ( .A(a[621]), .B(n4160), .Z(n27302) );
  NAND U28751 ( .A(n42144), .B(n27302), .Z(n27266) );
  AND U28752 ( .A(n27267), .B(n27266), .Z(n27317) );
  XOR U28753 ( .A(a[625]), .B(n42012), .Z(n27305) );
  XNOR U28754 ( .A(n27317), .B(n27316), .Z(n27319) );
  AND U28755 ( .A(a[627]), .B(b[0]), .Z(n27269) );
  XNOR U28756 ( .A(n27269), .B(n4071), .Z(n27271) );
  NANDN U28757 ( .A(b[0]), .B(a[626]), .Z(n27270) );
  NAND U28758 ( .A(n27271), .B(n27270), .Z(n27313) );
  XOR U28759 ( .A(a[623]), .B(n42085), .Z(n27306) );
  AND U28760 ( .A(a[619]), .B(b[7]), .Z(n27310) );
  XNOR U28761 ( .A(n27311), .B(n27310), .Z(n27312) );
  XNOR U28762 ( .A(n27313), .B(n27312), .Z(n27318) );
  XOR U28763 ( .A(n27319), .B(n27318), .Z(n27297) );
  NANDN U28764 ( .A(n27274), .B(n27273), .Z(n27278) );
  NANDN U28765 ( .A(n27276), .B(n27275), .Z(n27277) );
  AND U28766 ( .A(n27278), .B(n27277), .Z(n27296) );
  XNOR U28767 ( .A(n27297), .B(n27296), .Z(n27298) );
  NANDN U28768 ( .A(n27280), .B(n27279), .Z(n27284) );
  NAND U28769 ( .A(n27282), .B(n27281), .Z(n27283) );
  NAND U28770 ( .A(n27284), .B(n27283), .Z(n27299) );
  XNOR U28771 ( .A(n27298), .B(n27299), .Z(n27290) );
  XNOR U28772 ( .A(n27291), .B(n27290), .Z(n27292) );
  XNOR U28773 ( .A(n27293), .B(n27292), .Z(n27322) );
  XNOR U28774 ( .A(sreg[1643]), .B(n27322), .Z(n27324) );
  NANDN U28775 ( .A(sreg[1642]), .B(n27285), .Z(n27289) );
  NAND U28776 ( .A(n27287), .B(n27286), .Z(n27288) );
  NAND U28777 ( .A(n27289), .B(n27288), .Z(n27323) );
  XNOR U28778 ( .A(n27324), .B(n27323), .Z(c[1643]) );
  NANDN U28779 ( .A(n27291), .B(n27290), .Z(n27295) );
  NANDN U28780 ( .A(n27293), .B(n27292), .Z(n27294) );
  AND U28781 ( .A(n27295), .B(n27294), .Z(n27330) );
  NANDN U28782 ( .A(n27297), .B(n27296), .Z(n27301) );
  NANDN U28783 ( .A(n27299), .B(n27298), .Z(n27300) );
  AND U28784 ( .A(n27301), .B(n27300), .Z(n27328) );
  NAND U28785 ( .A(n42143), .B(n27302), .Z(n27304) );
  XNOR U28786 ( .A(a[622]), .B(n4160), .Z(n27339) );
  NAND U28787 ( .A(n42144), .B(n27339), .Z(n27303) );
  AND U28788 ( .A(n27304), .B(n27303), .Z(n27354) );
  XOR U28789 ( .A(a[626]), .B(n42012), .Z(n27342) );
  XNOR U28790 ( .A(n27354), .B(n27353), .Z(n27356) );
  XOR U28791 ( .A(a[624]), .B(n42085), .Z(n27346) );
  AND U28792 ( .A(a[620]), .B(b[7]), .Z(n27347) );
  XNOR U28793 ( .A(n27348), .B(n27347), .Z(n27349) );
  AND U28794 ( .A(a[628]), .B(b[0]), .Z(n27307) );
  XNOR U28795 ( .A(n27307), .B(n4071), .Z(n27309) );
  NANDN U28796 ( .A(b[0]), .B(a[627]), .Z(n27308) );
  NAND U28797 ( .A(n27309), .B(n27308), .Z(n27350) );
  XNOR U28798 ( .A(n27349), .B(n27350), .Z(n27355) );
  XOR U28799 ( .A(n27356), .B(n27355), .Z(n27334) );
  NANDN U28800 ( .A(n27311), .B(n27310), .Z(n27315) );
  NANDN U28801 ( .A(n27313), .B(n27312), .Z(n27314) );
  AND U28802 ( .A(n27315), .B(n27314), .Z(n27333) );
  XNOR U28803 ( .A(n27334), .B(n27333), .Z(n27335) );
  NANDN U28804 ( .A(n27317), .B(n27316), .Z(n27321) );
  NAND U28805 ( .A(n27319), .B(n27318), .Z(n27320) );
  NAND U28806 ( .A(n27321), .B(n27320), .Z(n27336) );
  XNOR U28807 ( .A(n27335), .B(n27336), .Z(n27327) );
  XNOR U28808 ( .A(n27328), .B(n27327), .Z(n27329) );
  XNOR U28809 ( .A(n27330), .B(n27329), .Z(n27359) );
  XNOR U28810 ( .A(sreg[1644]), .B(n27359), .Z(n27361) );
  NANDN U28811 ( .A(sreg[1643]), .B(n27322), .Z(n27326) );
  NAND U28812 ( .A(n27324), .B(n27323), .Z(n27325) );
  NAND U28813 ( .A(n27326), .B(n27325), .Z(n27360) );
  XNOR U28814 ( .A(n27361), .B(n27360), .Z(c[1644]) );
  NANDN U28815 ( .A(n27328), .B(n27327), .Z(n27332) );
  NANDN U28816 ( .A(n27330), .B(n27329), .Z(n27331) );
  AND U28817 ( .A(n27332), .B(n27331), .Z(n27367) );
  NANDN U28818 ( .A(n27334), .B(n27333), .Z(n27338) );
  NANDN U28819 ( .A(n27336), .B(n27335), .Z(n27337) );
  AND U28820 ( .A(n27338), .B(n27337), .Z(n27365) );
  NAND U28821 ( .A(n42143), .B(n27339), .Z(n27341) );
  XNOR U28822 ( .A(a[623]), .B(n4160), .Z(n27376) );
  NAND U28823 ( .A(n42144), .B(n27376), .Z(n27340) );
  AND U28824 ( .A(n27341), .B(n27340), .Z(n27391) );
  XOR U28825 ( .A(a[627]), .B(n42012), .Z(n27379) );
  XNOR U28826 ( .A(n27391), .B(n27390), .Z(n27393) );
  AND U28827 ( .A(a[629]), .B(b[0]), .Z(n27343) );
  XNOR U28828 ( .A(n27343), .B(n4071), .Z(n27345) );
  NANDN U28829 ( .A(b[0]), .B(a[628]), .Z(n27344) );
  NAND U28830 ( .A(n27345), .B(n27344), .Z(n27387) );
  XOR U28831 ( .A(a[625]), .B(n42085), .Z(n27383) );
  AND U28832 ( .A(a[621]), .B(b[7]), .Z(n27384) );
  XNOR U28833 ( .A(n27385), .B(n27384), .Z(n27386) );
  XNOR U28834 ( .A(n27387), .B(n27386), .Z(n27392) );
  XOR U28835 ( .A(n27393), .B(n27392), .Z(n27371) );
  NANDN U28836 ( .A(n27348), .B(n27347), .Z(n27352) );
  NANDN U28837 ( .A(n27350), .B(n27349), .Z(n27351) );
  AND U28838 ( .A(n27352), .B(n27351), .Z(n27370) );
  XNOR U28839 ( .A(n27371), .B(n27370), .Z(n27372) );
  NANDN U28840 ( .A(n27354), .B(n27353), .Z(n27358) );
  NAND U28841 ( .A(n27356), .B(n27355), .Z(n27357) );
  NAND U28842 ( .A(n27358), .B(n27357), .Z(n27373) );
  XNOR U28843 ( .A(n27372), .B(n27373), .Z(n27364) );
  XNOR U28844 ( .A(n27365), .B(n27364), .Z(n27366) );
  XNOR U28845 ( .A(n27367), .B(n27366), .Z(n27396) );
  XNOR U28846 ( .A(sreg[1645]), .B(n27396), .Z(n27398) );
  NANDN U28847 ( .A(sreg[1644]), .B(n27359), .Z(n27363) );
  NAND U28848 ( .A(n27361), .B(n27360), .Z(n27362) );
  NAND U28849 ( .A(n27363), .B(n27362), .Z(n27397) );
  XNOR U28850 ( .A(n27398), .B(n27397), .Z(c[1645]) );
  NANDN U28851 ( .A(n27365), .B(n27364), .Z(n27369) );
  NANDN U28852 ( .A(n27367), .B(n27366), .Z(n27368) );
  AND U28853 ( .A(n27369), .B(n27368), .Z(n27404) );
  NANDN U28854 ( .A(n27371), .B(n27370), .Z(n27375) );
  NANDN U28855 ( .A(n27373), .B(n27372), .Z(n27374) );
  AND U28856 ( .A(n27375), .B(n27374), .Z(n27402) );
  NAND U28857 ( .A(n42143), .B(n27376), .Z(n27378) );
  XNOR U28858 ( .A(a[624]), .B(n4161), .Z(n27413) );
  NAND U28859 ( .A(n42144), .B(n27413), .Z(n27377) );
  AND U28860 ( .A(n27378), .B(n27377), .Z(n27428) );
  XOR U28861 ( .A(a[628]), .B(n42012), .Z(n27416) );
  XNOR U28862 ( .A(n27428), .B(n27427), .Z(n27430) );
  AND U28863 ( .A(b[0]), .B(a[630]), .Z(n27380) );
  XOR U28864 ( .A(b[1]), .B(n27380), .Z(n27382) );
  NANDN U28865 ( .A(b[0]), .B(a[629]), .Z(n27381) );
  AND U28866 ( .A(n27382), .B(n27381), .Z(n27423) );
  XOR U28867 ( .A(a[626]), .B(n42085), .Z(n27420) );
  AND U28868 ( .A(a[622]), .B(b[7]), .Z(n27421) );
  XOR U28869 ( .A(n27422), .B(n27421), .Z(n27424) );
  XNOR U28870 ( .A(n27423), .B(n27424), .Z(n27429) );
  XOR U28871 ( .A(n27430), .B(n27429), .Z(n27408) );
  NANDN U28872 ( .A(n27385), .B(n27384), .Z(n27389) );
  NANDN U28873 ( .A(n27387), .B(n27386), .Z(n27388) );
  AND U28874 ( .A(n27389), .B(n27388), .Z(n27407) );
  XNOR U28875 ( .A(n27408), .B(n27407), .Z(n27409) );
  NANDN U28876 ( .A(n27391), .B(n27390), .Z(n27395) );
  NAND U28877 ( .A(n27393), .B(n27392), .Z(n27394) );
  NAND U28878 ( .A(n27395), .B(n27394), .Z(n27410) );
  XNOR U28879 ( .A(n27409), .B(n27410), .Z(n27401) );
  XNOR U28880 ( .A(n27402), .B(n27401), .Z(n27403) );
  XNOR U28881 ( .A(n27404), .B(n27403), .Z(n27433) );
  XNOR U28882 ( .A(sreg[1646]), .B(n27433), .Z(n27435) );
  NANDN U28883 ( .A(sreg[1645]), .B(n27396), .Z(n27400) );
  NAND U28884 ( .A(n27398), .B(n27397), .Z(n27399) );
  NAND U28885 ( .A(n27400), .B(n27399), .Z(n27434) );
  XNOR U28886 ( .A(n27435), .B(n27434), .Z(c[1646]) );
  NANDN U28887 ( .A(n27402), .B(n27401), .Z(n27406) );
  NANDN U28888 ( .A(n27404), .B(n27403), .Z(n27405) );
  AND U28889 ( .A(n27406), .B(n27405), .Z(n27441) );
  NANDN U28890 ( .A(n27408), .B(n27407), .Z(n27412) );
  NANDN U28891 ( .A(n27410), .B(n27409), .Z(n27411) );
  AND U28892 ( .A(n27412), .B(n27411), .Z(n27439) );
  NAND U28893 ( .A(n42143), .B(n27413), .Z(n27415) );
  XNOR U28894 ( .A(a[625]), .B(n4161), .Z(n27450) );
  NAND U28895 ( .A(n42144), .B(n27450), .Z(n27414) );
  AND U28896 ( .A(n27415), .B(n27414), .Z(n27465) );
  XOR U28897 ( .A(a[629]), .B(n42012), .Z(n27453) );
  XNOR U28898 ( .A(n27465), .B(n27464), .Z(n27467) );
  AND U28899 ( .A(a[631]), .B(b[0]), .Z(n27417) );
  XNOR U28900 ( .A(n27417), .B(n4071), .Z(n27419) );
  NANDN U28901 ( .A(b[0]), .B(a[630]), .Z(n27418) );
  NAND U28902 ( .A(n27419), .B(n27418), .Z(n27461) );
  XOR U28903 ( .A(a[627]), .B(n42085), .Z(n27457) );
  AND U28904 ( .A(a[623]), .B(b[7]), .Z(n27458) );
  XNOR U28905 ( .A(n27459), .B(n27458), .Z(n27460) );
  XNOR U28906 ( .A(n27461), .B(n27460), .Z(n27466) );
  XOR U28907 ( .A(n27467), .B(n27466), .Z(n27445) );
  NANDN U28908 ( .A(n27422), .B(n27421), .Z(n27426) );
  NANDN U28909 ( .A(n27424), .B(n27423), .Z(n27425) );
  AND U28910 ( .A(n27426), .B(n27425), .Z(n27444) );
  XNOR U28911 ( .A(n27445), .B(n27444), .Z(n27446) );
  NANDN U28912 ( .A(n27428), .B(n27427), .Z(n27432) );
  NAND U28913 ( .A(n27430), .B(n27429), .Z(n27431) );
  NAND U28914 ( .A(n27432), .B(n27431), .Z(n27447) );
  XNOR U28915 ( .A(n27446), .B(n27447), .Z(n27438) );
  XNOR U28916 ( .A(n27439), .B(n27438), .Z(n27440) );
  XNOR U28917 ( .A(n27441), .B(n27440), .Z(n27470) );
  XNOR U28918 ( .A(sreg[1647]), .B(n27470), .Z(n27472) );
  NANDN U28919 ( .A(sreg[1646]), .B(n27433), .Z(n27437) );
  NAND U28920 ( .A(n27435), .B(n27434), .Z(n27436) );
  NAND U28921 ( .A(n27437), .B(n27436), .Z(n27471) );
  XNOR U28922 ( .A(n27472), .B(n27471), .Z(c[1647]) );
  NANDN U28923 ( .A(n27439), .B(n27438), .Z(n27443) );
  NANDN U28924 ( .A(n27441), .B(n27440), .Z(n27442) );
  AND U28925 ( .A(n27443), .B(n27442), .Z(n27478) );
  NANDN U28926 ( .A(n27445), .B(n27444), .Z(n27449) );
  NANDN U28927 ( .A(n27447), .B(n27446), .Z(n27448) );
  AND U28928 ( .A(n27449), .B(n27448), .Z(n27476) );
  NAND U28929 ( .A(n42143), .B(n27450), .Z(n27452) );
  XNOR U28930 ( .A(a[626]), .B(n4161), .Z(n27487) );
  NAND U28931 ( .A(n42144), .B(n27487), .Z(n27451) );
  AND U28932 ( .A(n27452), .B(n27451), .Z(n27502) );
  XOR U28933 ( .A(a[630]), .B(n42012), .Z(n27490) );
  XNOR U28934 ( .A(n27502), .B(n27501), .Z(n27504) );
  AND U28935 ( .A(a[632]), .B(b[0]), .Z(n27454) );
  XNOR U28936 ( .A(n27454), .B(n4071), .Z(n27456) );
  NANDN U28937 ( .A(b[0]), .B(a[631]), .Z(n27455) );
  NAND U28938 ( .A(n27456), .B(n27455), .Z(n27498) );
  XOR U28939 ( .A(a[628]), .B(n42085), .Z(n27494) );
  AND U28940 ( .A(a[624]), .B(b[7]), .Z(n27495) );
  XNOR U28941 ( .A(n27496), .B(n27495), .Z(n27497) );
  XNOR U28942 ( .A(n27498), .B(n27497), .Z(n27503) );
  XOR U28943 ( .A(n27504), .B(n27503), .Z(n27482) );
  NANDN U28944 ( .A(n27459), .B(n27458), .Z(n27463) );
  NANDN U28945 ( .A(n27461), .B(n27460), .Z(n27462) );
  AND U28946 ( .A(n27463), .B(n27462), .Z(n27481) );
  XNOR U28947 ( .A(n27482), .B(n27481), .Z(n27483) );
  NANDN U28948 ( .A(n27465), .B(n27464), .Z(n27469) );
  NAND U28949 ( .A(n27467), .B(n27466), .Z(n27468) );
  NAND U28950 ( .A(n27469), .B(n27468), .Z(n27484) );
  XNOR U28951 ( .A(n27483), .B(n27484), .Z(n27475) );
  XNOR U28952 ( .A(n27476), .B(n27475), .Z(n27477) );
  XNOR U28953 ( .A(n27478), .B(n27477), .Z(n27507) );
  XNOR U28954 ( .A(sreg[1648]), .B(n27507), .Z(n27509) );
  NANDN U28955 ( .A(sreg[1647]), .B(n27470), .Z(n27474) );
  NAND U28956 ( .A(n27472), .B(n27471), .Z(n27473) );
  NAND U28957 ( .A(n27474), .B(n27473), .Z(n27508) );
  XNOR U28958 ( .A(n27509), .B(n27508), .Z(c[1648]) );
  NANDN U28959 ( .A(n27476), .B(n27475), .Z(n27480) );
  NANDN U28960 ( .A(n27478), .B(n27477), .Z(n27479) );
  AND U28961 ( .A(n27480), .B(n27479), .Z(n27515) );
  NANDN U28962 ( .A(n27482), .B(n27481), .Z(n27486) );
  NANDN U28963 ( .A(n27484), .B(n27483), .Z(n27485) );
  AND U28964 ( .A(n27486), .B(n27485), .Z(n27513) );
  NAND U28965 ( .A(n42143), .B(n27487), .Z(n27489) );
  XNOR U28966 ( .A(a[627]), .B(n4161), .Z(n27524) );
  NAND U28967 ( .A(n42144), .B(n27524), .Z(n27488) );
  AND U28968 ( .A(n27489), .B(n27488), .Z(n27539) );
  XOR U28969 ( .A(a[631]), .B(n42012), .Z(n27527) );
  XNOR U28970 ( .A(n27539), .B(n27538), .Z(n27541) );
  AND U28971 ( .A(a[633]), .B(b[0]), .Z(n27491) );
  XNOR U28972 ( .A(n27491), .B(n4071), .Z(n27493) );
  NANDN U28973 ( .A(b[0]), .B(a[632]), .Z(n27492) );
  NAND U28974 ( .A(n27493), .B(n27492), .Z(n27535) );
  XOR U28975 ( .A(a[629]), .B(n42085), .Z(n27531) );
  AND U28976 ( .A(a[625]), .B(b[7]), .Z(n27532) );
  XNOR U28977 ( .A(n27533), .B(n27532), .Z(n27534) );
  XNOR U28978 ( .A(n27535), .B(n27534), .Z(n27540) );
  XOR U28979 ( .A(n27541), .B(n27540), .Z(n27519) );
  NANDN U28980 ( .A(n27496), .B(n27495), .Z(n27500) );
  NANDN U28981 ( .A(n27498), .B(n27497), .Z(n27499) );
  AND U28982 ( .A(n27500), .B(n27499), .Z(n27518) );
  XNOR U28983 ( .A(n27519), .B(n27518), .Z(n27520) );
  NANDN U28984 ( .A(n27502), .B(n27501), .Z(n27506) );
  NAND U28985 ( .A(n27504), .B(n27503), .Z(n27505) );
  NAND U28986 ( .A(n27506), .B(n27505), .Z(n27521) );
  XNOR U28987 ( .A(n27520), .B(n27521), .Z(n27512) );
  XNOR U28988 ( .A(n27513), .B(n27512), .Z(n27514) );
  XNOR U28989 ( .A(n27515), .B(n27514), .Z(n27544) );
  XNOR U28990 ( .A(sreg[1649]), .B(n27544), .Z(n27546) );
  NANDN U28991 ( .A(sreg[1648]), .B(n27507), .Z(n27511) );
  NAND U28992 ( .A(n27509), .B(n27508), .Z(n27510) );
  NAND U28993 ( .A(n27511), .B(n27510), .Z(n27545) );
  XNOR U28994 ( .A(n27546), .B(n27545), .Z(c[1649]) );
  NANDN U28995 ( .A(n27513), .B(n27512), .Z(n27517) );
  NANDN U28996 ( .A(n27515), .B(n27514), .Z(n27516) );
  AND U28997 ( .A(n27517), .B(n27516), .Z(n27552) );
  NANDN U28998 ( .A(n27519), .B(n27518), .Z(n27523) );
  NANDN U28999 ( .A(n27521), .B(n27520), .Z(n27522) );
  AND U29000 ( .A(n27523), .B(n27522), .Z(n27550) );
  NAND U29001 ( .A(n42143), .B(n27524), .Z(n27526) );
  XNOR U29002 ( .A(a[628]), .B(n4161), .Z(n27561) );
  NAND U29003 ( .A(n42144), .B(n27561), .Z(n27525) );
  AND U29004 ( .A(n27526), .B(n27525), .Z(n27576) );
  XOR U29005 ( .A(a[632]), .B(n42012), .Z(n27564) );
  XNOR U29006 ( .A(n27576), .B(n27575), .Z(n27578) );
  AND U29007 ( .A(a[634]), .B(b[0]), .Z(n27528) );
  XNOR U29008 ( .A(n27528), .B(n4071), .Z(n27530) );
  NANDN U29009 ( .A(b[0]), .B(a[633]), .Z(n27529) );
  NAND U29010 ( .A(n27530), .B(n27529), .Z(n27572) );
  XOR U29011 ( .A(a[630]), .B(n42085), .Z(n27568) );
  AND U29012 ( .A(a[626]), .B(b[7]), .Z(n27569) );
  XNOR U29013 ( .A(n27570), .B(n27569), .Z(n27571) );
  XNOR U29014 ( .A(n27572), .B(n27571), .Z(n27577) );
  XOR U29015 ( .A(n27578), .B(n27577), .Z(n27556) );
  NANDN U29016 ( .A(n27533), .B(n27532), .Z(n27537) );
  NANDN U29017 ( .A(n27535), .B(n27534), .Z(n27536) );
  AND U29018 ( .A(n27537), .B(n27536), .Z(n27555) );
  XNOR U29019 ( .A(n27556), .B(n27555), .Z(n27557) );
  NANDN U29020 ( .A(n27539), .B(n27538), .Z(n27543) );
  NAND U29021 ( .A(n27541), .B(n27540), .Z(n27542) );
  NAND U29022 ( .A(n27543), .B(n27542), .Z(n27558) );
  XNOR U29023 ( .A(n27557), .B(n27558), .Z(n27549) );
  XNOR U29024 ( .A(n27550), .B(n27549), .Z(n27551) );
  XNOR U29025 ( .A(n27552), .B(n27551), .Z(n27581) );
  XNOR U29026 ( .A(sreg[1650]), .B(n27581), .Z(n27583) );
  NANDN U29027 ( .A(sreg[1649]), .B(n27544), .Z(n27548) );
  NAND U29028 ( .A(n27546), .B(n27545), .Z(n27547) );
  NAND U29029 ( .A(n27548), .B(n27547), .Z(n27582) );
  XNOR U29030 ( .A(n27583), .B(n27582), .Z(c[1650]) );
  NANDN U29031 ( .A(n27550), .B(n27549), .Z(n27554) );
  NANDN U29032 ( .A(n27552), .B(n27551), .Z(n27553) );
  AND U29033 ( .A(n27554), .B(n27553), .Z(n27589) );
  NANDN U29034 ( .A(n27556), .B(n27555), .Z(n27560) );
  NANDN U29035 ( .A(n27558), .B(n27557), .Z(n27559) );
  AND U29036 ( .A(n27560), .B(n27559), .Z(n27587) );
  NAND U29037 ( .A(n42143), .B(n27561), .Z(n27563) );
  XNOR U29038 ( .A(a[629]), .B(n4161), .Z(n27598) );
  NAND U29039 ( .A(n42144), .B(n27598), .Z(n27562) );
  AND U29040 ( .A(n27563), .B(n27562), .Z(n27613) );
  XOR U29041 ( .A(a[633]), .B(n42012), .Z(n27601) );
  XNOR U29042 ( .A(n27613), .B(n27612), .Z(n27615) );
  AND U29043 ( .A(a[635]), .B(b[0]), .Z(n27565) );
  XNOR U29044 ( .A(n27565), .B(n4071), .Z(n27567) );
  NANDN U29045 ( .A(b[0]), .B(a[634]), .Z(n27566) );
  NAND U29046 ( .A(n27567), .B(n27566), .Z(n27609) );
  XOR U29047 ( .A(a[631]), .B(n42085), .Z(n27605) );
  AND U29048 ( .A(a[627]), .B(b[7]), .Z(n27606) );
  XNOR U29049 ( .A(n27607), .B(n27606), .Z(n27608) );
  XNOR U29050 ( .A(n27609), .B(n27608), .Z(n27614) );
  XOR U29051 ( .A(n27615), .B(n27614), .Z(n27593) );
  NANDN U29052 ( .A(n27570), .B(n27569), .Z(n27574) );
  NANDN U29053 ( .A(n27572), .B(n27571), .Z(n27573) );
  AND U29054 ( .A(n27574), .B(n27573), .Z(n27592) );
  XNOR U29055 ( .A(n27593), .B(n27592), .Z(n27594) );
  NANDN U29056 ( .A(n27576), .B(n27575), .Z(n27580) );
  NAND U29057 ( .A(n27578), .B(n27577), .Z(n27579) );
  NAND U29058 ( .A(n27580), .B(n27579), .Z(n27595) );
  XNOR U29059 ( .A(n27594), .B(n27595), .Z(n27586) );
  XNOR U29060 ( .A(n27587), .B(n27586), .Z(n27588) );
  XNOR U29061 ( .A(n27589), .B(n27588), .Z(n27618) );
  XNOR U29062 ( .A(sreg[1651]), .B(n27618), .Z(n27620) );
  NANDN U29063 ( .A(sreg[1650]), .B(n27581), .Z(n27585) );
  NAND U29064 ( .A(n27583), .B(n27582), .Z(n27584) );
  NAND U29065 ( .A(n27585), .B(n27584), .Z(n27619) );
  XNOR U29066 ( .A(n27620), .B(n27619), .Z(c[1651]) );
  NANDN U29067 ( .A(n27587), .B(n27586), .Z(n27591) );
  NANDN U29068 ( .A(n27589), .B(n27588), .Z(n27590) );
  AND U29069 ( .A(n27591), .B(n27590), .Z(n27626) );
  NANDN U29070 ( .A(n27593), .B(n27592), .Z(n27597) );
  NANDN U29071 ( .A(n27595), .B(n27594), .Z(n27596) );
  AND U29072 ( .A(n27597), .B(n27596), .Z(n27624) );
  NAND U29073 ( .A(n42143), .B(n27598), .Z(n27600) );
  XNOR U29074 ( .A(a[630]), .B(n4161), .Z(n27635) );
  NAND U29075 ( .A(n42144), .B(n27635), .Z(n27599) );
  AND U29076 ( .A(n27600), .B(n27599), .Z(n27650) );
  XOR U29077 ( .A(a[634]), .B(n42012), .Z(n27638) );
  XNOR U29078 ( .A(n27650), .B(n27649), .Z(n27652) );
  AND U29079 ( .A(a[636]), .B(b[0]), .Z(n27602) );
  XNOR U29080 ( .A(n27602), .B(n4071), .Z(n27604) );
  NANDN U29081 ( .A(b[0]), .B(a[635]), .Z(n27603) );
  NAND U29082 ( .A(n27604), .B(n27603), .Z(n27646) );
  XOR U29083 ( .A(a[632]), .B(n42085), .Z(n27642) );
  AND U29084 ( .A(a[628]), .B(b[7]), .Z(n27643) );
  XNOR U29085 ( .A(n27644), .B(n27643), .Z(n27645) );
  XNOR U29086 ( .A(n27646), .B(n27645), .Z(n27651) );
  XOR U29087 ( .A(n27652), .B(n27651), .Z(n27630) );
  NANDN U29088 ( .A(n27607), .B(n27606), .Z(n27611) );
  NANDN U29089 ( .A(n27609), .B(n27608), .Z(n27610) );
  AND U29090 ( .A(n27611), .B(n27610), .Z(n27629) );
  XNOR U29091 ( .A(n27630), .B(n27629), .Z(n27631) );
  NANDN U29092 ( .A(n27613), .B(n27612), .Z(n27617) );
  NAND U29093 ( .A(n27615), .B(n27614), .Z(n27616) );
  NAND U29094 ( .A(n27617), .B(n27616), .Z(n27632) );
  XNOR U29095 ( .A(n27631), .B(n27632), .Z(n27623) );
  XNOR U29096 ( .A(n27624), .B(n27623), .Z(n27625) );
  XNOR U29097 ( .A(n27626), .B(n27625), .Z(n27655) );
  XNOR U29098 ( .A(sreg[1652]), .B(n27655), .Z(n27657) );
  NANDN U29099 ( .A(sreg[1651]), .B(n27618), .Z(n27622) );
  NAND U29100 ( .A(n27620), .B(n27619), .Z(n27621) );
  NAND U29101 ( .A(n27622), .B(n27621), .Z(n27656) );
  XNOR U29102 ( .A(n27657), .B(n27656), .Z(c[1652]) );
  NANDN U29103 ( .A(n27624), .B(n27623), .Z(n27628) );
  NANDN U29104 ( .A(n27626), .B(n27625), .Z(n27627) );
  AND U29105 ( .A(n27628), .B(n27627), .Z(n27663) );
  NANDN U29106 ( .A(n27630), .B(n27629), .Z(n27634) );
  NANDN U29107 ( .A(n27632), .B(n27631), .Z(n27633) );
  AND U29108 ( .A(n27634), .B(n27633), .Z(n27661) );
  NAND U29109 ( .A(n42143), .B(n27635), .Z(n27637) );
  XNOR U29110 ( .A(a[631]), .B(n4162), .Z(n27672) );
  NAND U29111 ( .A(n42144), .B(n27672), .Z(n27636) );
  AND U29112 ( .A(n27637), .B(n27636), .Z(n27687) );
  XOR U29113 ( .A(a[635]), .B(n42012), .Z(n27675) );
  XNOR U29114 ( .A(n27687), .B(n27686), .Z(n27689) );
  AND U29115 ( .A(a[637]), .B(b[0]), .Z(n27639) );
  XNOR U29116 ( .A(n27639), .B(n4071), .Z(n27641) );
  NANDN U29117 ( .A(b[0]), .B(a[636]), .Z(n27640) );
  NAND U29118 ( .A(n27641), .B(n27640), .Z(n27683) );
  XOR U29119 ( .A(a[633]), .B(n42085), .Z(n27676) );
  AND U29120 ( .A(a[629]), .B(b[7]), .Z(n27680) );
  XNOR U29121 ( .A(n27681), .B(n27680), .Z(n27682) );
  XNOR U29122 ( .A(n27683), .B(n27682), .Z(n27688) );
  XOR U29123 ( .A(n27689), .B(n27688), .Z(n27667) );
  NANDN U29124 ( .A(n27644), .B(n27643), .Z(n27648) );
  NANDN U29125 ( .A(n27646), .B(n27645), .Z(n27647) );
  AND U29126 ( .A(n27648), .B(n27647), .Z(n27666) );
  XNOR U29127 ( .A(n27667), .B(n27666), .Z(n27668) );
  NANDN U29128 ( .A(n27650), .B(n27649), .Z(n27654) );
  NAND U29129 ( .A(n27652), .B(n27651), .Z(n27653) );
  NAND U29130 ( .A(n27654), .B(n27653), .Z(n27669) );
  XNOR U29131 ( .A(n27668), .B(n27669), .Z(n27660) );
  XNOR U29132 ( .A(n27661), .B(n27660), .Z(n27662) );
  XNOR U29133 ( .A(n27663), .B(n27662), .Z(n27692) );
  XNOR U29134 ( .A(sreg[1653]), .B(n27692), .Z(n27694) );
  NANDN U29135 ( .A(sreg[1652]), .B(n27655), .Z(n27659) );
  NAND U29136 ( .A(n27657), .B(n27656), .Z(n27658) );
  NAND U29137 ( .A(n27659), .B(n27658), .Z(n27693) );
  XNOR U29138 ( .A(n27694), .B(n27693), .Z(c[1653]) );
  NANDN U29139 ( .A(n27661), .B(n27660), .Z(n27665) );
  NANDN U29140 ( .A(n27663), .B(n27662), .Z(n27664) );
  AND U29141 ( .A(n27665), .B(n27664), .Z(n27700) );
  NANDN U29142 ( .A(n27667), .B(n27666), .Z(n27671) );
  NANDN U29143 ( .A(n27669), .B(n27668), .Z(n27670) );
  AND U29144 ( .A(n27671), .B(n27670), .Z(n27698) );
  NAND U29145 ( .A(n42143), .B(n27672), .Z(n27674) );
  XNOR U29146 ( .A(a[632]), .B(n4162), .Z(n27709) );
  NAND U29147 ( .A(n42144), .B(n27709), .Z(n27673) );
  AND U29148 ( .A(n27674), .B(n27673), .Z(n27724) );
  XOR U29149 ( .A(a[636]), .B(n42012), .Z(n27712) );
  XNOR U29150 ( .A(n27724), .B(n27723), .Z(n27726) );
  XOR U29151 ( .A(a[634]), .B(n42085), .Z(n27716) );
  AND U29152 ( .A(a[630]), .B(b[7]), .Z(n27717) );
  XNOR U29153 ( .A(n27718), .B(n27717), .Z(n27719) );
  AND U29154 ( .A(a[638]), .B(b[0]), .Z(n27677) );
  XNOR U29155 ( .A(n27677), .B(n4071), .Z(n27679) );
  NANDN U29156 ( .A(b[0]), .B(a[637]), .Z(n27678) );
  NAND U29157 ( .A(n27679), .B(n27678), .Z(n27720) );
  XNOR U29158 ( .A(n27719), .B(n27720), .Z(n27725) );
  XOR U29159 ( .A(n27726), .B(n27725), .Z(n27704) );
  NANDN U29160 ( .A(n27681), .B(n27680), .Z(n27685) );
  NANDN U29161 ( .A(n27683), .B(n27682), .Z(n27684) );
  AND U29162 ( .A(n27685), .B(n27684), .Z(n27703) );
  XNOR U29163 ( .A(n27704), .B(n27703), .Z(n27705) );
  NANDN U29164 ( .A(n27687), .B(n27686), .Z(n27691) );
  NAND U29165 ( .A(n27689), .B(n27688), .Z(n27690) );
  NAND U29166 ( .A(n27691), .B(n27690), .Z(n27706) );
  XNOR U29167 ( .A(n27705), .B(n27706), .Z(n27697) );
  XNOR U29168 ( .A(n27698), .B(n27697), .Z(n27699) );
  XNOR U29169 ( .A(n27700), .B(n27699), .Z(n27729) );
  XNOR U29170 ( .A(sreg[1654]), .B(n27729), .Z(n27731) );
  NANDN U29171 ( .A(sreg[1653]), .B(n27692), .Z(n27696) );
  NAND U29172 ( .A(n27694), .B(n27693), .Z(n27695) );
  NAND U29173 ( .A(n27696), .B(n27695), .Z(n27730) );
  XNOR U29174 ( .A(n27731), .B(n27730), .Z(c[1654]) );
  NANDN U29175 ( .A(n27698), .B(n27697), .Z(n27702) );
  NANDN U29176 ( .A(n27700), .B(n27699), .Z(n27701) );
  AND U29177 ( .A(n27702), .B(n27701), .Z(n27737) );
  NANDN U29178 ( .A(n27704), .B(n27703), .Z(n27708) );
  NANDN U29179 ( .A(n27706), .B(n27705), .Z(n27707) );
  AND U29180 ( .A(n27708), .B(n27707), .Z(n27735) );
  NAND U29181 ( .A(n42143), .B(n27709), .Z(n27711) );
  XNOR U29182 ( .A(a[633]), .B(n4162), .Z(n27746) );
  NAND U29183 ( .A(n42144), .B(n27746), .Z(n27710) );
  AND U29184 ( .A(n27711), .B(n27710), .Z(n27761) );
  XOR U29185 ( .A(a[637]), .B(n42012), .Z(n27749) );
  XNOR U29186 ( .A(n27761), .B(n27760), .Z(n27763) );
  AND U29187 ( .A(a[639]), .B(b[0]), .Z(n27713) );
  XNOR U29188 ( .A(n27713), .B(n4071), .Z(n27715) );
  NANDN U29189 ( .A(b[0]), .B(a[638]), .Z(n27714) );
  NAND U29190 ( .A(n27715), .B(n27714), .Z(n27757) );
  XOR U29191 ( .A(a[635]), .B(n42085), .Z(n27750) );
  AND U29192 ( .A(a[631]), .B(b[7]), .Z(n27754) );
  XNOR U29193 ( .A(n27755), .B(n27754), .Z(n27756) );
  XNOR U29194 ( .A(n27757), .B(n27756), .Z(n27762) );
  XOR U29195 ( .A(n27763), .B(n27762), .Z(n27741) );
  NANDN U29196 ( .A(n27718), .B(n27717), .Z(n27722) );
  NANDN U29197 ( .A(n27720), .B(n27719), .Z(n27721) );
  AND U29198 ( .A(n27722), .B(n27721), .Z(n27740) );
  XNOR U29199 ( .A(n27741), .B(n27740), .Z(n27742) );
  NANDN U29200 ( .A(n27724), .B(n27723), .Z(n27728) );
  NAND U29201 ( .A(n27726), .B(n27725), .Z(n27727) );
  NAND U29202 ( .A(n27728), .B(n27727), .Z(n27743) );
  XNOR U29203 ( .A(n27742), .B(n27743), .Z(n27734) );
  XNOR U29204 ( .A(n27735), .B(n27734), .Z(n27736) );
  XNOR U29205 ( .A(n27737), .B(n27736), .Z(n27766) );
  XNOR U29206 ( .A(sreg[1655]), .B(n27766), .Z(n27768) );
  NANDN U29207 ( .A(sreg[1654]), .B(n27729), .Z(n27733) );
  NAND U29208 ( .A(n27731), .B(n27730), .Z(n27732) );
  NAND U29209 ( .A(n27733), .B(n27732), .Z(n27767) );
  XNOR U29210 ( .A(n27768), .B(n27767), .Z(c[1655]) );
  NANDN U29211 ( .A(n27735), .B(n27734), .Z(n27739) );
  NANDN U29212 ( .A(n27737), .B(n27736), .Z(n27738) );
  AND U29213 ( .A(n27739), .B(n27738), .Z(n27774) );
  NANDN U29214 ( .A(n27741), .B(n27740), .Z(n27745) );
  NANDN U29215 ( .A(n27743), .B(n27742), .Z(n27744) );
  AND U29216 ( .A(n27745), .B(n27744), .Z(n27772) );
  NAND U29217 ( .A(n42143), .B(n27746), .Z(n27748) );
  XNOR U29218 ( .A(a[634]), .B(n4162), .Z(n27783) );
  NAND U29219 ( .A(n42144), .B(n27783), .Z(n27747) );
  AND U29220 ( .A(n27748), .B(n27747), .Z(n27798) );
  XOR U29221 ( .A(a[638]), .B(n42012), .Z(n27786) );
  XNOR U29222 ( .A(n27798), .B(n27797), .Z(n27800) );
  XOR U29223 ( .A(a[636]), .B(n42085), .Z(n27790) );
  AND U29224 ( .A(a[632]), .B(b[7]), .Z(n27791) );
  XNOR U29225 ( .A(n27792), .B(n27791), .Z(n27793) );
  AND U29226 ( .A(a[640]), .B(b[0]), .Z(n27751) );
  XNOR U29227 ( .A(n27751), .B(n4071), .Z(n27753) );
  NANDN U29228 ( .A(b[0]), .B(a[639]), .Z(n27752) );
  NAND U29229 ( .A(n27753), .B(n27752), .Z(n27794) );
  XNOR U29230 ( .A(n27793), .B(n27794), .Z(n27799) );
  XOR U29231 ( .A(n27800), .B(n27799), .Z(n27778) );
  NANDN U29232 ( .A(n27755), .B(n27754), .Z(n27759) );
  NANDN U29233 ( .A(n27757), .B(n27756), .Z(n27758) );
  AND U29234 ( .A(n27759), .B(n27758), .Z(n27777) );
  XNOR U29235 ( .A(n27778), .B(n27777), .Z(n27779) );
  NANDN U29236 ( .A(n27761), .B(n27760), .Z(n27765) );
  NAND U29237 ( .A(n27763), .B(n27762), .Z(n27764) );
  NAND U29238 ( .A(n27765), .B(n27764), .Z(n27780) );
  XNOR U29239 ( .A(n27779), .B(n27780), .Z(n27771) );
  XNOR U29240 ( .A(n27772), .B(n27771), .Z(n27773) );
  XNOR U29241 ( .A(n27774), .B(n27773), .Z(n27803) );
  XNOR U29242 ( .A(sreg[1656]), .B(n27803), .Z(n27805) );
  NANDN U29243 ( .A(sreg[1655]), .B(n27766), .Z(n27770) );
  NAND U29244 ( .A(n27768), .B(n27767), .Z(n27769) );
  NAND U29245 ( .A(n27770), .B(n27769), .Z(n27804) );
  XNOR U29246 ( .A(n27805), .B(n27804), .Z(c[1656]) );
  NANDN U29247 ( .A(n27772), .B(n27771), .Z(n27776) );
  NANDN U29248 ( .A(n27774), .B(n27773), .Z(n27775) );
  AND U29249 ( .A(n27776), .B(n27775), .Z(n27811) );
  NANDN U29250 ( .A(n27778), .B(n27777), .Z(n27782) );
  NANDN U29251 ( .A(n27780), .B(n27779), .Z(n27781) );
  AND U29252 ( .A(n27782), .B(n27781), .Z(n27809) );
  NAND U29253 ( .A(n42143), .B(n27783), .Z(n27785) );
  XNOR U29254 ( .A(a[635]), .B(n4162), .Z(n27820) );
  NAND U29255 ( .A(n42144), .B(n27820), .Z(n27784) );
  AND U29256 ( .A(n27785), .B(n27784), .Z(n27835) );
  XOR U29257 ( .A(a[639]), .B(n42012), .Z(n27823) );
  XNOR U29258 ( .A(n27835), .B(n27834), .Z(n27837) );
  AND U29259 ( .A(a[641]), .B(b[0]), .Z(n27787) );
  XNOR U29260 ( .A(n27787), .B(n4071), .Z(n27789) );
  NANDN U29261 ( .A(b[0]), .B(a[640]), .Z(n27788) );
  NAND U29262 ( .A(n27789), .B(n27788), .Z(n27831) );
  XOR U29263 ( .A(a[637]), .B(n42085), .Z(n27827) );
  AND U29264 ( .A(a[633]), .B(b[7]), .Z(n27828) );
  XNOR U29265 ( .A(n27829), .B(n27828), .Z(n27830) );
  XNOR U29266 ( .A(n27831), .B(n27830), .Z(n27836) );
  XOR U29267 ( .A(n27837), .B(n27836), .Z(n27815) );
  NANDN U29268 ( .A(n27792), .B(n27791), .Z(n27796) );
  NANDN U29269 ( .A(n27794), .B(n27793), .Z(n27795) );
  AND U29270 ( .A(n27796), .B(n27795), .Z(n27814) );
  XNOR U29271 ( .A(n27815), .B(n27814), .Z(n27816) );
  NANDN U29272 ( .A(n27798), .B(n27797), .Z(n27802) );
  NAND U29273 ( .A(n27800), .B(n27799), .Z(n27801) );
  NAND U29274 ( .A(n27802), .B(n27801), .Z(n27817) );
  XNOR U29275 ( .A(n27816), .B(n27817), .Z(n27808) );
  XNOR U29276 ( .A(n27809), .B(n27808), .Z(n27810) );
  XNOR U29277 ( .A(n27811), .B(n27810), .Z(n27840) );
  XNOR U29278 ( .A(sreg[1657]), .B(n27840), .Z(n27842) );
  NANDN U29279 ( .A(sreg[1656]), .B(n27803), .Z(n27807) );
  NAND U29280 ( .A(n27805), .B(n27804), .Z(n27806) );
  NAND U29281 ( .A(n27807), .B(n27806), .Z(n27841) );
  XNOR U29282 ( .A(n27842), .B(n27841), .Z(c[1657]) );
  NANDN U29283 ( .A(n27809), .B(n27808), .Z(n27813) );
  NANDN U29284 ( .A(n27811), .B(n27810), .Z(n27812) );
  AND U29285 ( .A(n27813), .B(n27812), .Z(n27848) );
  NANDN U29286 ( .A(n27815), .B(n27814), .Z(n27819) );
  NANDN U29287 ( .A(n27817), .B(n27816), .Z(n27818) );
  AND U29288 ( .A(n27819), .B(n27818), .Z(n27846) );
  NAND U29289 ( .A(n42143), .B(n27820), .Z(n27822) );
  XNOR U29290 ( .A(a[636]), .B(n4162), .Z(n27857) );
  NAND U29291 ( .A(n42144), .B(n27857), .Z(n27821) );
  AND U29292 ( .A(n27822), .B(n27821), .Z(n27872) );
  XOR U29293 ( .A(a[640]), .B(n42012), .Z(n27860) );
  XNOR U29294 ( .A(n27872), .B(n27871), .Z(n27874) );
  AND U29295 ( .A(a[642]), .B(b[0]), .Z(n27824) );
  XNOR U29296 ( .A(n27824), .B(n4071), .Z(n27826) );
  NANDN U29297 ( .A(b[0]), .B(a[641]), .Z(n27825) );
  NAND U29298 ( .A(n27826), .B(n27825), .Z(n27868) );
  XOR U29299 ( .A(a[638]), .B(n42085), .Z(n27864) );
  AND U29300 ( .A(a[634]), .B(b[7]), .Z(n27865) );
  XNOR U29301 ( .A(n27866), .B(n27865), .Z(n27867) );
  XNOR U29302 ( .A(n27868), .B(n27867), .Z(n27873) );
  XOR U29303 ( .A(n27874), .B(n27873), .Z(n27852) );
  NANDN U29304 ( .A(n27829), .B(n27828), .Z(n27833) );
  NANDN U29305 ( .A(n27831), .B(n27830), .Z(n27832) );
  AND U29306 ( .A(n27833), .B(n27832), .Z(n27851) );
  XNOR U29307 ( .A(n27852), .B(n27851), .Z(n27853) );
  NANDN U29308 ( .A(n27835), .B(n27834), .Z(n27839) );
  NAND U29309 ( .A(n27837), .B(n27836), .Z(n27838) );
  NAND U29310 ( .A(n27839), .B(n27838), .Z(n27854) );
  XNOR U29311 ( .A(n27853), .B(n27854), .Z(n27845) );
  XNOR U29312 ( .A(n27846), .B(n27845), .Z(n27847) );
  XNOR U29313 ( .A(n27848), .B(n27847), .Z(n27877) );
  XNOR U29314 ( .A(sreg[1658]), .B(n27877), .Z(n27879) );
  NANDN U29315 ( .A(sreg[1657]), .B(n27840), .Z(n27844) );
  NAND U29316 ( .A(n27842), .B(n27841), .Z(n27843) );
  NAND U29317 ( .A(n27844), .B(n27843), .Z(n27878) );
  XNOR U29318 ( .A(n27879), .B(n27878), .Z(c[1658]) );
  NANDN U29319 ( .A(n27846), .B(n27845), .Z(n27850) );
  NANDN U29320 ( .A(n27848), .B(n27847), .Z(n27849) );
  AND U29321 ( .A(n27850), .B(n27849), .Z(n27885) );
  NANDN U29322 ( .A(n27852), .B(n27851), .Z(n27856) );
  NANDN U29323 ( .A(n27854), .B(n27853), .Z(n27855) );
  AND U29324 ( .A(n27856), .B(n27855), .Z(n27883) );
  NAND U29325 ( .A(n42143), .B(n27857), .Z(n27859) );
  XNOR U29326 ( .A(a[637]), .B(n4162), .Z(n27894) );
  NAND U29327 ( .A(n42144), .B(n27894), .Z(n27858) );
  AND U29328 ( .A(n27859), .B(n27858), .Z(n27909) );
  XOR U29329 ( .A(a[641]), .B(n42012), .Z(n27897) );
  XNOR U29330 ( .A(n27909), .B(n27908), .Z(n27911) );
  AND U29331 ( .A(a[643]), .B(b[0]), .Z(n27861) );
  XNOR U29332 ( .A(n27861), .B(n4071), .Z(n27863) );
  NANDN U29333 ( .A(b[0]), .B(a[642]), .Z(n27862) );
  NAND U29334 ( .A(n27863), .B(n27862), .Z(n27905) );
  XOR U29335 ( .A(a[639]), .B(n42085), .Z(n27898) );
  AND U29336 ( .A(a[635]), .B(b[7]), .Z(n27902) );
  XNOR U29337 ( .A(n27903), .B(n27902), .Z(n27904) );
  XNOR U29338 ( .A(n27905), .B(n27904), .Z(n27910) );
  XOR U29339 ( .A(n27911), .B(n27910), .Z(n27889) );
  NANDN U29340 ( .A(n27866), .B(n27865), .Z(n27870) );
  NANDN U29341 ( .A(n27868), .B(n27867), .Z(n27869) );
  AND U29342 ( .A(n27870), .B(n27869), .Z(n27888) );
  XNOR U29343 ( .A(n27889), .B(n27888), .Z(n27890) );
  NANDN U29344 ( .A(n27872), .B(n27871), .Z(n27876) );
  NAND U29345 ( .A(n27874), .B(n27873), .Z(n27875) );
  NAND U29346 ( .A(n27876), .B(n27875), .Z(n27891) );
  XNOR U29347 ( .A(n27890), .B(n27891), .Z(n27882) );
  XNOR U29348 ( .A(n27883), .B(n27882), .Z(n27884) );
  XNOR U29349 ( .A(n27885), .B(n27884), .Z(n27914) );
  XNOR U29350 ( .A(sreg[1659]), .B(n27914), .Z(n27916) );
  NANDN U29351 ( .A(sreg[1658]), .B(n27877), .Z(n27881) );
  NAND U29352 ( .A(n27879), .B(n27878), .Z(n27880) );
  NAND U29353 ( .A(n27881), .B(n27880), .Z(n27915) );
  XNOR U29354 ( .A(n27916), .B(n27915), .Z(c[1659]) );
  NANDN U29355 ( .A(n27883), .B(n27882), .Z(n27887) );
  NANDN U29356 ( .A(n27885), .B(n27884), .Z(n27886) );
  AND U29357 ( .A(n27887), .B(n27886), .Z(n27922) );
  NANDN U29358 ( .A(n27889), .B(n27888), .Z(n27893) );
  NANDN U29359 ( .A(n27891), .B(n27890), .Z(n27892) );
  AND U29360 ( .A(n27893), .B(n27892), .Z(n27920) );
  NAND U29361 ( .A(n42143), .B(n27894), .Z(n27896) );
  XNOR U29362 ( .A(a[638]), .B(n4163), .Z(n27931) );
  NAND U29363 ( .A(n42144), .B(n27931), .Z(n27895) );
  AND U29364 ( .A(n27896), .B(n27895), .Z(n27946) );
  XOR U29365 ( .A(a[642]), .B(n42012), .Z(n27934) );
  XNOR U29366 ( .A(n27946), .B(n27945), .Z(n27948) );
  XOR U29367 ( .A(a[640]), .B(n42085), .Z(n27935) );
  AND U29368 ( .A(a[636]), .B(b[7]), .Z(n27939) );
  XNOR U29369 ( .A(n27940), .B(n27939), .Z(n27941) );
  AND U29370 ( .A(a[644]), .B(b[0]), .Z(n27899) );
  XNOR U29371 ( .A(n27899), .B(n4071), .Z(n27901) );
  NANDN U29372 ( .A(b[0]), .B(a[643]), .Z(n27900) );
  NAND U29373 ( .A(n27901), .B(n27900), .Z(n27942) );
  XNOR U29374 ( .A(n27941), .B(n27942), .Z(n27947) );
  XOR U29375 ( .A(n27948), .B(n27947), .Z(n27926) );
  NANDN U29376 ( .A(n27903), .B(n27902), .Z(n27907) );
  NANDN U29377 ( .A(n27905), .B(n27904), .Z(n27906) );
  AND U29378 ( .A(n27907), .B(n27906), .Z(n27925) );
  XNOR U29379 ( .A(n27926), .B(n27925), .Z(n27927) );
  NANDN U29380 ( .A(n27909), .B(n27908), .Z(n27913) );
  NAND U29381 ( .A(n27911), .B(n27910), .Z(n27912) );
  NAND U29382 ( .A(n27913), .B(n27912), .Z(n27928) );
  XNOR U29383 ( .A(n27927), .B(n27928), .Z(n27919) );
  XNOR U29384 ( .A(n27920), .B(n27919), .Z(n27921) );
  XNOR U29385 ( .A(n27922), .B(n27921), .Z(n27951) );
  XNOR U29386 ( .A(sreg[1660]), .B(n27951), .Z(n27953) );
  NANDN U29387 ( .A(sreg[1659]), .B(n27914), .Z(n27918) );
  NAND U29388 ( .A(n27916), .B(n27915), .Z(n27917) );
  NAND U29389 ( .A(n27918), .B(n27917), .Z(n27952) );
  XNOR U29390 ( .A(n27953), .B(n27952), .Z(c[1660]) );
  NANDN U29391 ( .A(n27920), .B(n27919), .Z(n27924) );
  NANDN U29392 ( .A(n27922), .B(n27921), .Z(n27923) );
  AND U29393 ( .A(n27924), .B(n27923), .Z(n27959) );
  NANDN U29394 ( .A(n27926), .B(n27925), .Z(n27930) );
  NANDN U29395 ( .A(n27928), .B(n27927), .Z(n27929) );
  AND U29396 ( .A(n27930), .B(n27929), .Z(n27957) );
  NAND U29397 ( .A(n42143), .B(n27931), .Z(n27933) );
  XNOR U29398 ( .A(a[639]), .B(n4163), .Z(n27968) );
  NAND U29399 ( .A(n42144), .B(n27968), .Z(n27932) );
  AND U29400 ( .A(n27933), .B(n27932), .Z(n27983) );
  XOR U29401 ( .A(a[643]), .B(n42012), .Z(n27971) );
  XNOR U29402 ( .A(n27983), .B(n27982), .Z(n27985) );
  XOR U29403 ( .A(a[641]), .B(n42085), .Z(n27972) );
  AND U29404 ( .A(a[637]), .B(b[7]), .Z(n27976) );
  XNOR U29405 ( .A(n27977), .B(n27976), .Z(n27978) );
  AND U29406 ( .A(a[645]), .B(b[0]), .Z(n27936) );
  XNOR U29407 ( .A(n27936), .B(n4071), .Z(n27938) );
  NANDN U29408 ( .A(b[0]), .B(a[644]), .Z(n27937) );
  NAND U29409 ( .A(n27938), .B(n27937), .Z(n27979) );
  XNOR U29410 ( .A(n27978), .B(n27979), .Z(n27984) );
  XOR U29411 ( .A(n27985), .B(n27984), .Z(n27963) );
  NANDN U29412 ( .A(n27940), .B(n27939), .Z(n27944) );
  NANDN U29413 ( .A(n27942), .B(n27941), .Z(n27943) );
  AND U29414 ( .A(n27944), .B(n27943), .Z(n27962) );
  XNOR U29415 ( .A(n27963), .B(n27962), .Z(n27964) );
  NANDN U29416 ( .A(n27946), .B(n27945), .Z(n27950) );
  NAND U29417 ( .A(n27948), .B(n27947), .Z(n27949) );
  NAND U29418 ( .A(n27950), .B(n27949), .Z(n27965) );
  XNOR U29419 ( .A(n27964), .B(n27965), .Z(n27956) );
  XNOR U29420 ( .A(n27957), .B(n27956), .Z(n27958) );
  XNOR U29421 ( .A(n27959), .B(n27958), .Z(n27988) );
  XNOR U29422 ( .A(sreg[1661]), .B(n27988), .Z(n27990) );
  NANDN U29423 ( .A(sreg[1660]), .B(n27951), .Z(n27955) );
  NAND U29424 ( .A(n27953), .B(n27952), .Z(n27954) );
  NAND U29425 ( .A(n27955), .B(n27954), .Z(n27989) );
  XNOR U29426 ( .A(n27990), .B(n27989), .Z(c[1661]) );
  NANDN U29427 ( .A(n27957), .B(n27956), .Z(n27961) );
  NANDN U29428 ( .A(n27959), .B(n27958), .Z(n27960) );
  AND U29429 ( .A(n27961), .B(n27960), .Z(n27996) );
  NANDN U29430 ( .A(n27963), .B(n27962), .Z(n27967) );
  NANDN U29431 ( .A(n27965), .B(n27964), .Z(n27966) );
  AND U29432 ( .A(n27967), .B(n27966), .Z(n27994) );
  NAND U29433 ( .A(n42143), .B(n27968), .Z(n27970) );
  XNOR U29434 ( .A(a[640]), .B(n4163), .Z(n28005) );
  NAND U29435 ( .A(n42144), .B(n28005), .Z(n27969) );
  AND U29436 ( .A(n27970), .B(n27969), .Z(n28020) );
  XOR U29437 ( .A(a[644]), .B(n42012), .Z(n28008) );
  XNOR U29438 ( .A(n28020), .B(n28019), .Z(n28022) );
  XOR U29439 ( .A(a[642]), .B(n42085), .Z(n28012) );
  AND U29440 ( .A(a[638]), .B(b[7]), .Z(n28013) );
  XNOR U29441 ( .A(n28014), .B(n28013), .Z(n28015) );
  AND U29442 ( .A(a[646]), .B(b[0]), .Z(n27973) );
  XNOR U29443 ( .A(n27973), .B(n4071), .Z(n27975) );
  NANDN U29444 ( .A(b[0]), .B(a[645]), .Z(n27974) );
  NAND U29445 ( .A(n27975), .B(n27974), .Z(n28016) );
  XNOR U29446 ( .A(n28015), .B(n28016), .Z(n28021) );
  XOR U29447 ( .A(n28022), .B(n28021), .Z(n28000) );
  NANDN U29448 ( .A(n27977), .B(n27976), .Z(n27981) );
  NANDN U29449 ( .A(n27979), .B(n27978), .Z(n27980) );
  AND U29450 ( .A(n27981), .B(n27980), .Z(n27999) );
  XNOR U29451 ( .A(n28000), .B(n27999), .Z(n28001) );
  NANDN U29452 ( .A(n27983), .B(n27982), .Z(n27987) );
  NAND U29453 ( .A(n27985), .B(n27984), .Z(n27986) );
  NAND U29454 ( .A(n27987), .B(n27986), .Z(n28002) );
  XNOR U29455 ( .A(n28001), .B(n28002), .Z(n27993) );
  XNOR U29456 ( .A(n27994), .B(n27993), .Z(n27995) );
  XNOR U29457 ( .A(n27996), .B(n27995), .Z(n28025) );
  XNOR U29458 ( .A(sreg[1662]), .B(n28025), .Z(n28027) );
  NANDN U29459 ( .A(sreg[1661]), .B(n27988), .Z(n27992) );
  NAND U29460 ( .A(n27990), .B(n27989), .Z(n27991) );
  NAND U29461 ( .A(n27992), .B(n27991), .Z(n28026) );
  XNOR U29462 ( .A(n28027), .B(n28026), .Z(c[1662]) );
  NANDN U29463 ( .A(n27994), .B(n27993), .Z(n27998) );
  NANDN U29464 ( .A(n27996), .B(n27995), .Z(n27997) );
  AND U29465 ( .A(n27998), .B(n27997), .Z(n28033) );
  NANDN U29466 ( .A(n28000), .B(n27999), .Z(n28004) );
  NANDN U29467 ( .A(n28002), .B(n28001), .Z(n28003) );
  AND U29468 ( .A(n28004), .B(n28003), .Z(n28031) );
  NAND U29469 ( .A(n42143), .B(n28005), .Z(n28007) );
  XNOR U29470 ( .A(a[641]), .B(n4163), .Z(n28042) );
  NAND U29471 ( .A(n42144), .B(n28042), .Z(n28006) );
  AND U29472 ( .A(n28007), .B(n28006), .Z(n28057) );
  XOR U29473 ( .A(a[645]), .B(n42012), .Z(n28045) );
  XNOR U29474 ( .A(n28057), .B(n28056), .Z(n28059) );
  AND U29475 ( .A(a[647]), .B(b[0]), .Z(n28009) );
  XNOR U29476 ( .A(n28009), .B(n4071), .Z(n28011) );
  NANDN U29477 ( .A(b[0]), .B(a[646]), .Z(n28010) );
  NAND U29478 ( .A(n28011), .B(n28010), .Z(n28053) );
  XOR U29479 ( .A(a[643]), .B(n42085), .Z(n28046) );
  AND U29480 ( .A(a[639]), .B(b[7]), .Z(n28050) );
  XNOR U29481 ( .A(n28051), .B(n28050), .Z(n28052) );
  XNOR U29482 ( .A(n28053), .B(n28052), .Z(n28058) );
  XOR U29483 ( .A(n28059), .B(n28058), .Z(n28037) );
  NANDN U29484 ( .A(n28014), .B(n28013), .Z(n28018) );
  NANDN U29485 ( .A(n28016), .B(n28015), .Z(n28017) );
  AND U29486 ( .A(n28018), .B(n28017), .Z(n28036) );
  XNOR U29487 ( .A(n28037), .B(n28036), .Z(n28038) );
  NANDN U29488 ( .A(n28020), .B(n28019), .Z(n28024) );
  NAND U29489 ( .A(n28022), .B(n28021), .Z(n28023) );
  NAND U29490 ( .A(n28024), .B(n28023), .Z(n28039) );
  XNOR U29491 ( .A(n28038), .B(n28039), .Z(n28030) );
  XNOR U29492 ( .A(n28031), .B(n28030), .Z(n28032) );
  XNOR U29493 ( .A(n28033), .B(n28032), .Z(n28062) );
  XNOR U29494 ( .A(sreg[1663]), .B(n28062), .Z(n28064) );
  NANDN U29495 ( .A(sreg[1662]), .B(n28025), .Z(n28029) );
  NAND U29496 ( .A(n28027), .B(n28026), .Z(n28028) );
  NAND U29497 ( .A(n28029), .B(n28028), .Z(n28063) );
  XNOR U29498 ( .A(n28064), .B(n28063), .Z(c[1663]) );
  NANDN U29499 ( .A(n28031), .B(n28030), .Z(n28035) );
  NANDN U29500 ( .A(n28033), .B(n28032), .Z(n28034) );
  AND U29501 ( .A(n28035), .B(n28034), .Z(n28070) );
  NANDN U29502 ( .A(n28037), .B(n28036), .Z(n28041) );
  NANDN U29503 ( .A(n28039), .B(n28038), .Z(n28040) );
  AND U29504 ( .A(n28041), .B(n28040), .Z(n28068) );
  NAND U29505 ( .A(n42143), .B(n28042), .Z(n28044) );
  XNOR U29506 ( .A(a[642]), .B(n4163), .Z(n28079) );
  NAND U29507 ( .A(n42144), .B(n28079), .Z(n28043) );
  AND U29508 ( .A(n28044), .B(n28043), .Z(n28094) );
  XOR U29509 ( .A(a[646]), .B(n42012), .Z(n28082) );
  XNOR U29510 ( .A(n28094), .B(n28093), .Z(n28096) );
  XOR U29511 ( .A(a[644]), .B(n42085), .Z(n28086) );
  AND U29512 ( .A(a[640]), .B(b[7]), .Z(n28087) );
  XNOR U29513 ( .A(n28088), .B(n28087), .Z(n28089) );
  AND U29514 ( .A(a[648]), .B(b[0]), .Z(n28047) );
  XNOR U29515 ( .A(n28047), .B(n4071), .Z(n28049) );
  NANDN U29516 ( .A(b[0]), .B(a[647]), .Z(n28048) );
  NAND U29517 ( .A(n28049), .B(n28048), .Z(n28090) );
  XNOR U29518 ( .A(n28089), .B(n28090), .Z(n28095) );
  XOR U29519 ( .A(n28096), .B(n28095), .Z(n28074) );
  NANDN U29520 ( .A(n28051), .B(n28050), .Z(n28055) );
  NANDN U29521 ( .A(n28053), .B(n28052), .Z(n28054) );
  AND U29522 ( .A(n28055), .B(n28054), .Z(n28073) );
  XNOR U29523 ( .A(n28074), .B(n28073), .Z(n28075) );
  NANDN U29524 ( .A(n28057), .B(n28056), .Z(n28061) );
  NAND U29525 ( .A(n28059), .B(n28058), .Z(n28060) );
  NAND U29526 ( .A(n28061), .B(n28060), .Z(n28076) );
  XNOR U29527 ( .A(n28075), .B(n28076), .Z(n28067) );
  XNOR U29528 ( .A(n28068), .B(n28067), .Z(n28069) );
  XNOR U29529 ( .A(n28070), .B(n28069), .Z(n28099) );
  XNOR U29530 ( .A(sreg[1664]), .B(n28099), .Z(n28101) );
  NANDN U29531 ( .A(sreg[1663]), .B(n28062), .Z(n28066) );
  NAND U29532 ( .A(n28064), .B(n28063), .Z(n28065) );
  NAND U29533 ( .A(n28066), .B(n28065), .Z(n28100) );
  XNOR U29534 ( .A(n28101), .B(n28100), .Z(c[1664]) );
  NANDN U29535 ( .A(n28068), .B(n28067), .Z(n28072) );
  NANDN U29536 ( .A(n28070), .B(n28069), .Z(n28071) );
  AND U29537 ( .A(n28072), .B(n28071), .Z(n28107) );
  NANDN U29538 ( .A(n28074), .B(n28073), .Z(n28078) );
  NANDN U29539 ( .A(n28076), .B(n28075), .Z(n28077) );
  AND U29540 ( .A(n28078), .B(n28077), .Z(n28105) );
  NAND U29541 ( .A(n42143), .B(n28079), .Z(n28081) );
  XNOR U29542 ( .A(a[643]), .B(n4163), .Z(n28116) );
  NAND U29543 ( .A(n42144), .B(n28116), .Z(n28080) );
  AND U29544 ( .A(n28081), .B(n28080), .Z(n28131) );
  XOR U29545 ( .A(a[647]), .B(n42012), .Z(n28119) );
  XNOR U29546 ( .A(n28131), .B(n28130), .Z(n28133) );
  AND U29547 ( .A(a[649]), .B(b[0]), .Z(n28083) );
  XNOR U29548 ( .A(n28083), .B(n4071), .Z(n28085) );
  NANDN U29549 ( .A(b[0]), .B(a[648]), .Z(n28084) );
  NAND U29550 ( .A(n28085), .B(n28084), .Z(n28127) );
  XOR U29551 ( .A(a[645]), .B(n42085), .Z(n28123) );
  AND U29552 ( .A(a[641]), .B(b[7]), .Z(n28124) );
  XNOR U29553 ( .A(n28125), .B(n28124), .Z(n28126) );
  XNOR U29554 ( .A(n28127), .B(n28126), .Z(n28132) );
  XOR U29555 ( .A(n28133), .B(n28132), .Z(n28111) );
  NANDN U29556 ( .A(n28088), .B(n28087), .Z(n28092) );
  NANDN U29557 ( .A(n28090), .B(n28089), .Z(n28091) );
  AND U29558 ( .A(n28092), .B(n28091), .Z(n28110) );
  XNOR U29559 ( .A(n28111), .B(n28110), .Z(n28112) );
  NANDN U29560 ( .A(n28094), .B(n28093), .Z(n28098) );
  NAND U29561 ( .A(n28096), .B(n28095), .Z(n28097) );
  NAND U29562 ( .A(n28098), .B(n28097), .Z(n28113) );
  XNOR U29563 ( .A(n28112), .B(n28113), .Z(n28104) );
  XNOR U29564 ( .A(n28105), .B(n28104), .Z(n28106) );
  XNOR U29565 ( .A(n28107), .B(n28106), .Z(n28136) );
  XNOR U29566 ( .A(sreg[1665]), .B(n28136), .Z(n28138) );
  NANDN U29567 ( .A(sreg[1664]), .B(n28099), .Z(n28103) );
  NAND U29568 ( .A(n28101), .B(n28100), .Z(n28102) );
  NAND U29569 ( .A(n28103), .B(n28102), .Z(n28137) );
  XNOR U29570 ( .A(n28138), .B(n28137), .Z(c[1665]) );
  NANDN U29571 ( .A(n28105), .B(n28104), .Z(n28109) );
  NANDN U29572 ( .A(n28107), .B(n28106), .Z(n28108) );
  AND U29573 ( .A(n28109), .B(n28108), .Z(n28144) );
  NANDN U29574 ( .A(n28111), .B(n28110), .Z(n28115) );
  NANDN U29575 ( .A(n28113), .B(n28112), .Z(n28114) );
  AND U29576 ( .A(n28115), .B(n28114), .Z(n28142) );
  NAND U29577 ( .A(n42143), .B(n28116), .Z(n28118) );
  XNOR U29578 ( .A(a[644]), .B(n4163), .Z(n28153) );
  NAND U29579 ( .A(n42144), .B(n28153), .Z(n28117) );
  AND U29580 ( .A(n28118), .B(n28117), .Z(n28168) );
  XOR U29581 ( .A(a[648]), .B(n42012), .Z(n28156) );
  XNOR U29582 ( .A(n28168), .B(n28167), .Z(n28170) );
  AND U29583 ( .A(a[650]), .B(b[0]), .Z(n28120) );
  XNOR U29584 ( .A(n28120), .B(n4071), .Z(n28122) );
  NANDN U29585 ( .A(b[0]), .B(a[649]), .Z(n28121) );
  NAND U29586 ( .A(n28122), .B(n28121), .Z(n28164) );
  XOR U29587 ( .A(a[646]), .B(n42085), .Z(n28160) );
  AND U29588 ( .A(a[642]), .B(b[7]), .Z(n28161) );
  XNOR U29589 ( .A(n28162), .B(n28161), .Z(n28163) );
  XNOR U29590 ( .A(n28164), .B(n28163), .Z(n28169) );
  XOR U29591 ( .A(n28170), .B(n28169), .Z(n28148) );
  NANDN U29592 ( .A(n28125), .B(n28124), .Z(n28129) );
  NANDN U29593 ( .A(n28127), .B(n28126), .Z(n28128) );
  AND U29594 ( .A(n28129), .B(n28128), .Z(n28147) );
  XNOR U29595 ( .A(n28148), .B(n28147), .Z(n28149) );
  NANDN U29596 ( .A(n28131), .B(n28130), .Z(n28135) );
  NAND U29597 ( .A(n28133), .B(n28132), .Z(n28134) );
  NAND U29598 ( .A(n28135), .B(n28134), .Z(n28150) );
  XNOR U29599 ( .A(n28149), .B(n28150), .Z(n28141) );
  XNOR U29600 ( .A(n28142), .B(n28141), .Z(n28143) );
  XNOR U29601 ( .A(n28144), .B(n28143), .Z(n28173) );
  XNOR U29602 ( .A(sreg[1666]), .B(n28173), .Z(n28175) );
  NANDN U29603 ( .A(sreg[1665]), .B(n28136), .Z(n28140) );
  NAND U29604 ( .A(n28138), .B(n28137), .Z(n28139) );
  NAND U29605 ( .A(n28140), .B(n28139), .Z(n28174) );
  XNOR U29606 ( .A(n28175), .B(n28174), .Z(c[1666]) );
  NANDN U29607 ( .A(n28142), .B(n28141), .Z(n28146) );
  NANDN U29608 ( .A(n28144), .B(n28143), .Z(n28145) );
  AND U29609 ( .A(n28146), .B(n28145), .Z(n28181) );
  NANDN U29610 ( .A(n28148), .B(n28147), .Z(n28152) );
  NANDN U29611 ( .A(n28150), .B(n28149), .Z(n28151) );
  AND U29612 ( .A(n28152), .B(n28151), .Z(n28179) );
  NAND U29613 ( .A(n42143), .B(n28153), .Z(n28155) );
  XNOR U29614 ( .A(a[645]), .B(n4164), .Z(n28190) );
  NAND U29615 ( .A(n42144), .B(n28190), .Z(n28154) );
  AND U29616 ( .A(n28155), .B(n28154), .Z(n28205) );
  XOR U29617 ( .A(a[649]), .B(n42012), .Z(n28193) );
  XNOR U29618 ( .A(n28205), .B(n28204), .Z(n28207) );
  AND U29619 ( .A(a[651]), .B(b[0]), .Z(n28157) );
  XNOR U29620 ( .A(n28157), .B(n4071), .Z(n28159) );
  NANDN U29621 ( .A(b[0]), .B(a[650]), .Z(n28158) );
  NAND U29622 ( .A(n28159), .B(n28158), .Z(n28201) );
  XOR U29623 ( .A(a[647]), .B(n42085), .Z(n28197) );
  AND U29624 ( .A(a[643]), .B(b[7]), .Z(n28198) );
  XNOR U29625 ( .A(n28199), .B(n28198), .Z(n28200) );
  XNOR U29626 ( .A(n28201), .B(n28200), .Z(n28206) );
  XOR U29627 ( .A(n28207), .B(n28206), .Z(n28185) );
  NANDN U29628 ( .A(n28162), .B(n28161), .Z(n28166) );
  NANDN U29629 ( .A(n28164), .B(n28163), .Z(n28165) );
  AND U29630 ( .A(n28166), .B(n28165), .Z(n28184) );
  XNOR U29631 ( .A(n28185), .B(n28184), .Z(n28186) );
  NANDN U29632 ( .A(n28168), .B(n28167), .Z(n28172) );
  NAND U29633 ( .A(n28170), .B(n28169), .Z(n28171) );
  NAND U29634 ( .A(n28172), .B(n28171), .Z(n28187) );
  XNOR U29635 ( .A(n28186), .B(n28187), .Z(n28178) );
  XNOR U29636 ( .A(n28179), .B(n28178), .Z(n28180) );
  XNOR U29637 ( .A(n28181), .B(n28180), .Z(n28210) );
  XNOR U29638 ( .A(sreg[1667]), .B(n28210), .Z(n28212) );
  NANDN U29639 ( .A(sreg[1666]), .B(n28173), .Z(n28177) );
  NAND U29640 ( .A(n28175), .B(n28174), .Z(n28176) );
  NAND U29641 ( .A(n28177), .B(n28176), .Z(n28211) );
  XNOR U29642 ( .A(n28212), .B(n28211), .Z(c[1667]) );
  NANDN U29643 ( .A(n28179), .B(n28178), .Z(n28183) );
  NANDN U29644 ( .A(n28181), .B(n28180), .Z(n28182) );
  AND U29645 ( .A(n28183), .B(n28182), .Z(n28218) );
  NANDN U29646 ( .A(n28185), .B(n28184), .Z(n28189) );
  NANDN U29647 ( .A(n28187), .B(n28186), .Z(n28188) );
  AND U29648 ( .A(n28189), .B(n28188), .Z(n28216) );
  NAND U29649 ( .A(n42143), .B(n28190), .Z(n28192) );
  XNOR U29650 ( .A(a[646]), .B(n4164), .Z(n28227) );
  NAND U29651 ( .A(n42144), .B(n28227), .Z(n28191) );
  AND U29652 ( .A(n28192), .B(n28191), .Z(n28242) );
  XOR U29653 ( .A(a[650]), .B(n42012), .Z(n28230) );
  XNOR U29654 ( .A(n28242), .B(n28241), .Z(n28244) );
  AND U29655 ( .A(a[652]), .B(b[0]), .Z(n28194) );
  XNOR U29656 ( .A(n28194), .B(n4071), .Z(n28196) );
  NANDN U29657 ( .A(b[0]), .B(a[651]), .Z(n28195) );
  NAND U29658 ( .A(n28196), .B(n28195), .Z(n28238) );
  XOR U29659 ( .A(a[648]), .B(n42085), .Z(n28234) );
  AND U29660 ( .A(a[644]), .B(b[7]), .Z(n28235) );
  XNOR U29661 ( .A(n28236), .B(n28235), .Z(n28237) );
  XNOR U29662 ( .A(n28238), .B(n28237), .Z(n28243) );
  XOR U29663 ( .A(n28244), .B(n28243), .Z(n28222) );
  NANDN U29664 ( .A(n28199), .B(n28198), .Z(n28203) );
  NANDN U29665 ( .A(n28201), .B(n28200), .Z(n28202) );
  AND U29666 ( .A(n28203), .B(n28202), .Z(n28221) );
  XNOR U29667 ( .A(n28222), .B(n28221), .Z(n28223) );
  NANDN U29668 ( .A(n28205), .B(n28204), .Z(n28209) );
  NAND U29669 ( .A(n28207), .B(n28206), .Z(n28208) );
  NAND U29670 ( .A(n28209), .B(n28208), .Z(n28224) );
  XNOR U29671 ( .A(n28223), .B(n28224), .Z(n28215) );
  XNOR U29672 ( .A(n28216), .B(n28215), .Z(n28217) );
  XNOR U29673 ( .A(n28218), .B(n28217), .Z(n28247) );
  XNOR U29674 ( .A(sreg[1668]), .B(n28247), .Z(n28249) );
  NANDN U29675 ( .A(sreg[1667]), .B(n28210), .Z(n28214) );
  NAND U29676 ( .A(n28212), .B(n28211), .Z(n28213) );
  NAND U29677 ( .A(n28214), .B(n28213), .Z(n28248) );
  XNOR U29678 ( .A(n28249), .B(n28248), .Z(c[1668]) );
  NANDN U29679 ( .A(n28216), .B(n28215), .Z(n28220) );
  NANDN U29680 ( .A(n28218), .B(n28217), .Z(n28219) );
  AND U29681 ( .A(n28220), .B(n28219), .Z(n28255) );
  NANDN U29682 ( .A(n28222), .B(n28221), .Z(n28226) );
  NANDN U29683 ( .A(n28224), .B(n28223), .Z(n28225) );
  AND U29684 ( .A(n28226), .B(n28225), .Z(n28253) );
  NAND U29685 ( .A(n42143), .B(n28227), .Z(n28229) );
  XNOR U29686 ( .A(a[647]), .B(n4164), .Z(n28264) );
  NAND U29687 ( .A(n42144), .B(n28264), .Z(n28228) );
  AND U29688 ( .A(n28229), .B(n28228), .Z(n28279) );
  XOR U29689 ( .A(a[651]), .B(n42012), .Z(n28267) );
  XNOR U29690 ( .A(n28279), .B(n28278), .Z(n28281) );
  AND U29691 ( .A(a[653]), .B(b[0]), .Z(n28231) );
  XNOR U29692 ( .A(n28231), .B(n4071), .Z(n28233) );
  NANDN U29693 ( .A(b[0]), .B(a[652]), .Z(n28232) );
  NAND U29694 ( .A(n28233), .B(n28232), .Z(n28275) );
  XOR U29695 ( .A(a[649]), .B(n42085), .Z(n28271) );
  AND U29696 ( .A(a[645]), .B(b[7]), .Z(n28272) );
  XNOR U29697 ( .A(n28273), .B(n28272), .Z(n28274) );
  XNOR U29698 ( .A(n28275), .B(n28274), .Z(n28280) );
  XOR U29699 ( .A(n28281), .B(n28280), .Z(n28259) );
  NANDN U29700 ( .A(n28236), .B(n28235), .Z(n28240) );
  NANDN U29701 ( .A(n28238), .B(n28237), .Z(n28239) );
  AND U29702 ( .A(n28240), .B(n28239), .Z(n28258) );
  XNOR U29703 ( .A(n28259), .B(n28258), .Z(n28260) );
  NANDN U29704 ( .A(n28242), .B(n28241), .Z(n28246) );
  NAND U29705 ( .A(n28244), .B(n28243), .Z(n28245) );
  NAND U29706 ( .A(n28246), .B(n28245), .Z(n28261) );
  XNOR U29707 ( .A(n28260), .B(n28261), .Z(n28252) );
  XNOR U29708 ( .A(n28253), .B(n28252), .Z(n28254) );
  XNOR U29709 ( .A(n28255), .B(n28254), .Z(n28284) );
  XNOR U29710 ( .A(sreg[1669]), .B(n28284), .Z(n28286) );
  NANDN U29711 ( .A(sreg[1668]), .B(n28247), .Z(n28251) );
  NAND U29712 ( .A(n28249), .B(n28248), .Z(n28250) );
  NAND U29713 ( .A(n28251), .B(n28250), .Z(n28285) );
  XNOR U29714 ( .A(n28286), .B(n28285), .Z(c[1669]) );
  NANDN U29715 ( .A(n28253), .B(n28252), .Z(n28257) );
  NANDN U29716 ( .A(n28255), .B(n28254), .Z(n28256) );
  AND U29717 ( .A(n28257), .B(n28256), .Z(n28292) );
  NANDN U29718 ( .A(n28259), .B(n28258), .Z(n28263) );
  NANDN U29719 ( .A(n28261), .B(n28260), .Z(n28262) );
  AND U29720 ( .A(n28263), .B(n28262), .Z(n28290) );
  NAND U29721 ( .A(n42143), .B(n28264), .Z(n28266) );
  XNOR U29722 ( .A(a[648]), .B(n4164), .Z(n28301) );
  NAND U29723 ( .A(n42144), .B(n28301), .Z(n28265) );
  AND U29724 ( .A(n28266), .B(n28265), .Z(n28316) );
  XOR U29725 ( .A(a[652]), .B(n42012), .Z(n28304) );
  XNOR U29726 ( .A(n28316), .B(n28315), .Z(n28318) );
  AND U29727 ( .A(a[654]), .B(b[0]), .Z(n28268) );
  XNOR U29728 ( .A(n28268), .B(n4071), .Z(n28270) );
  NANDN U29729 ( .A(b[0]), .B(a[653]), .Z(n28269) );
  NAND U29730 ( .A(n28270), .B(n28269), .Z(n28312) );
  XOR U29731 ( .A(a[650]), .B(n42085), .Z(n28308) );
  AND U29732 ( .A(a[646]), .B(b[7]), .Z(n28309) );
  XNOR U29733 ( .A(n28310), .B(n28309), .Z(n28311) );
  XNOR U29734 ( .A(n28312), .B(n28311), .Z(n28317) );
  XOR U29735 ( .A(n28318), .B(n28317), .Z(n28296) );
  NANDN U29736 ( .A(n28273), .B(n28272), .Z(n28277) );
  NANDN U29737 ( .A(n28275), .B(n28274), .Z(n28276) );
  AND U29738 ( .A(n28277), .B(n28276), .Z(n28295) );
  XNOR U29739 ( .A(n28296), .B(n28295), .Z(n28297) );
  NANDN U29740 ( .A(n28279), .B(n28278), .Z(n28283) );
  NAND U29741 ( .A(n28281), .B(n28280), .Z(n28282) );
  NAND U29742 ( .A(n28283), .B(n28282), .Z(n28298) );
  XNOR U29743 ( .A(n28297), .B(n28298), .Z(n28289) );
  XNOR U29744 ( .A(n28290), .B(n28289), .Z(n28291) );
  XNOR U29745 ( .A(n28292), .B(n28291), .Z(n28321) );
  XNOR U29746 ( .A(sreg[1670]), .B(n28321), .Z(n28323) );
  NANDN U29747 ( .A(sreg[1669]), .B(n28284), .Z(n28288) );
  NAND U29748 ( .A(n28286), .B(n28285), .Z(n28287) );
  NAND U29749 ( .A(n28288), .B(n28287), .Z(n28322) );
  XNOR U29750 ( .A(n28323), .B(n28322), .Z(c[1670]) );
  NANDN U29751 ( .A(n28290), .B(n28289), .Z(n28294) );
  NANDN U29752 ( .A(n28292), .B(n28291), .Z(n28293) );
  AND U29753 ( .A(n28294), .B(n28293), .Z(n28329) );
  NANDN U29754 ( .A(n28296), .B(n28295), .Z(n28300) );
  NANDN U29755 ( .A(n28298), .B(n28297), .Z(n28299) );
  AND U29756 ( .A(n28300), .B(n28299), .Z(n28327) );
  NAND U29757 ( .A(n42143), .B(n28301), .Z(n28303) );
  XNOR U29758 ( .A(a[649]), .B(n4164), .Z(n28338) );
  NAND U29759 ( .A(n42144), .B(n28338), .Z(n28302) );
  AND U29760 ( .A(n28303), .B(n28302), .Z(n28353) );
  XOR U29761 ( .A(a[653]), .B(n42012), .Z(n28341) );
  XNOR U29762 ( .A(n28353), .B(n28352), .Z(n28355) );
  AND U29763 ( .A(a[655]), .B(b[0]), .Z(n28305) );
  XNOR U29764 ( .A(n28305), .B(n4071), .Z(n28307) );
  NANDN U29765 ( .A(b[0]), .B(a[654]), .Z(n28306) );
  NAND U29766 ( .A(n28307), .B(n28306), .Z(n28349) );
  XOR U29767 ( .A(a[651]), .B(n42085), .Z(n28345) );
  AND U29768 ( .A(a[647]), .B(b[7]), .Z(n28346) );
  XNOR U29769 ( .A(n28347), .B(n28346), .Z(n28348) );
  XNOR U29770 ( .A(n28349), .B(n28348), .Z(n28354) );
  XOR U29771 ( .A(n28355), .B(n28354), .Z(n28333) );
  NANDN U29772 ( .A(n28310), .B(n28309), .Z(n28314) );
  NANDN U29773 ( .A(n28312), .B(n28311), .Z(n28313) );
  AND U29774 ( .A(n28314), .B(n28313), .Z(n28332) );
  XNOR U29775 ( .A(n28333), .B(n28332), .Z(n28334) );
  NANDN U29776 ( .A(n28316), .B(n28315), .Z(n28320) );
  NAND U29777 ( .A(n28318), .B(n28317), .Z(n28319) );
  NAND U29778 ( .A(n28320), .B(n28319), .Z(n28335) );
  XNOR U29779 ( .A(n28334), .B(n28335), .Z(n28326) );
  XNOR U29780 ( .A(n28327), .B(n28326), .Z(n28328) );
  XNOR U29781 ( .A(n28329), .B(n28328), .Z(n28358) );
  XNOR U29782 ( .A(sreg[1671]), .B(n28358), .Z(n28360) );
  NANDN U29783 ( .A(sreg[1670]), .B(n28321), .Z(n28325) );
  NAND U29784 ( .A(n28323), .B(n28322), .Z(n28324) );
  NAND U29785 ( .A(n28325), .B(n28324), .Z(n28359) );
  XNOR U29786 ( .A(n28360), .B(n28359), .Z(c[1671]) );
  NANDN U29787 ( .A(n28327), .B(n28326), .Z(n28331) );
  NANDN U29788 ( .A(n28329), .B(n28328), .Z(n28330) );
  AND U29789 ( .A(n28331), .B(n28330), .Z(n28366) );
  NANDN U29790 ( .A(n28333), .B(n28332), .Z(n28337) );
  NANDN U29791 ( .A(n28335), .B(n28334), .Z(n28336) );
  AND U29792 ( .A(n28337), .B(n28336), .Z(n28364) );
  NAND U29793 ( .A(n42143), .B(n28338), .Z(n28340) );
  XNOR U29794 ( .A(a[650]), .B(n4164), .Z(n28375) );
  NAND U29795 ( .A(n42144), .B(n28375), .Z(n28339) );
  AND U29796 ( .A(n28340), .B(n28339), .Z(n28390) );
  XOR U29797 ( .A(a[654]), .B(n42012), .Z(n28378) );
  XNOR U29798 ( .A(n28390), .B(n28389), .Z(n28392) );
  AND U29799 ( .A(a[656]), .B(b[0]), .Z(n28342) );
  XNOR U29800 ( .A(n28342), .B(n4071), .Z(n28344) );
  NANDN U29801 ( .A(b[0]), .B(a[655]), .Z(n28343) );
  NAND U29802 ( .A(n28344), .B(n28343), .Z(n28386) );
  XOR U29803 ( .A(a[652]), .B(n42085), .Z(n28382) );
  AND U29804 ( .A(a[648]), .B(b[7]), .Z(n28383) );
  XNOR U29805 ( .A(n28384), .B(n28383), .Z(n28385) );
  XNOR U29806 ( .A(n28386), .B(n28385), .Z(n28391) );
  XOR U29807 ( .A(n28392), .B(n28391), .Z(n28370) );
  NANDN U29808 ( .A(n28347), .B(n28346), .Z(n28351) );
  NANDN U29809 ( .A(n28349), .B(n28348), .Z(n28350) );
  AND U29810 ( .A(n28351), .B(n28350), .Z(n28369) );
  XNOR U29811 ( .A(n28370), .B(n28369), .Z(n28371) );
  NANDN U29812 ( .A(n28353), .B(n28352), .Z(n28357) );
  NAND U29813 ( .A(n28355), .B(n28354), .Z(n28356) );
  NAND U29814 ( .A(n28357), .B(n28356), .Z(n28372) );
  XNOR U29815 ( .A(n28371), .B(n28372), .Z(n28363) );
  XNOR U29816 ( .A(n28364), .B(n28363), .Z(n28365) );
  XNOR U29817 ( .A(n28366), .B(n28365), .Z(n28395) );
  XNOR U29818 ( .A(sreg[1672]), .B(n28395), .Z(n28397) );
  NANDN U29819 ( .A(sreg[1671]), .B(n28358), .Z(n28362) );
  NAND U29820 ( .A(n28360), .B(n28359), .Z(n28361) );
  NAND U29821 ( .A(n28362), .B(n28361), .Z(n28396) );
  XNOR U29822 ( .A(n28397), .B(n28396), .Z(c[1672]) );
  NANDN U29823 ( .A(n28364), .B(n28363), .Z(n28368) );
  NANDN U29824 ( .A(n28366), .B(n28365), .Z(n28367) );
  AND U29825 ( .A(n28368), .B(n28367), .Z(n28403) );
  NANDN U29826 ( .A(n28370), .B(n28369), .Z(n28374) );
  NANDN U29827 ( .A(n28372), .B(n28371), .Z(n28373) );
  AND U29828 ( .A(n28374), .B(n28373), .Z(n28401) );
  NAND U29829 ( .A(n42143), .B(n28375), .Z(n28377) );
  XNOR U29830 ( .A(a[651]), .B(n4164), .Z(n28412) );
  NAND U29831 ( .A(n42144), .B(n28412), .Z(n28376) );
  AND U29832 ( .A(n28377), .B(n28376), .Z(n28427) );
  XOR U29833 ( .A(a[655]), .B(n42012), .Z(n28415) );
  XNOR U29834 ( .A(n28427), .B(n28426), .Z(n28429) );
  AND U29835 ( .A(a[657]), .B(b[0]), .Z(n28379) );
  XNOR U29836 ( .A(n28379), .B(n4071), .Z(n28381) );
  NANDN U29837 ( .A(b[0]), .B(a[656]), .Z(n28380) );
  NAND U29838 ( .A(n28381), .B(n28380), .Z(n28423) );
  XOR U29839 ( .A(a[653]), .B(n42085), .Z(n28416) );
  AND U29840 ( .A(a[649]), .B(b[7]), .Z(n28420) );
  XNOR U29841 ( .A(n28421), .B(n28420), .Z(n28422) );
  XNOR U29842 ( .A(n28423), .B(n28422), .Z(n28428) );
  XOR U29843 ( .A(n28429), .B(n28428), .Z(n28407) );
  NANDN U29844 ( .A(n28384), .B(n28383), .Z(n28388) );
  NANDN U29845 ( .A(n28386), .B(n28385), .Z(n28387) );
  AND U29846 ( .A(n28388), .B(n28387), .Z(n28406) );
  XNOR U29847 ( .A(n28407), .B(n28406), .Z(n28408) );
  NANDN U29848 ( .A(n28390), .B(n28389), .Z(n28394) );
  NAND U29849 ( .A(n28392), .B(n28391), .Z(n28393) );
  NAND U29850 ( .A(n28394), .B(n28393), .Z(n28409) );
  XNOR U29851 ( .A(n28408), .B(n28409), .Z(n28400) );
  XNOR U29852 ( .A(n28401), .B(n28400), .Z(n28402) );
  XNOR U29853 ( .A(n28403), .B(n28402), .Z(n28432) );
  XNOR U29854 ( .A(sreg[1673]), .B(n28432), .Z(n28434) );
  NANDN U29855 ( .A(sreg[1672]), .B(n28395), .Z(n28399) );
  NAND U29856 ( .A(n28397), .B(n28396), .Z(n28398) );
  NAND U29857 ( .A(n28399), .B(n28398), .Z(n28433) );
  XNOR U29858 ( .A(n28434), .B(n28433), .Z(c[1673]) );
  NANDN U29859 ( .A(n28401), .B(n28400), .Z(n28405) );
  NANDN U29860 ( .A(n28403), .B(n28402), .Z(n28404) );
  AND U29861 ( .A(n28405), .B(n28404), .Z(n28440) );
  NANDN U29862 ( .A(n28407), .B(n28406), .Z(n28411) );
  NANDN U29863 ( .A(n28409), .B(n28408), .Z(n28410) );
  AND U29864 ( .A(n28411), .B(n28410), .Z(n28438) );
  NAND U29865 ( .A(n42143), .B(n28412), .Z(n28414) );
  XNOR U29866 ( .A(a[652]), .B(n4165), .Z(n28449) );
  NAND U29867 ( .A(n42144), .B(n28449), .Z(n28413) );
  AND U29868 ( .A(n28414), .B(n28413), .Z(n28464) );
  XOR U29869 ( .A(a[656]), .B(n42012), .Z(n28452) );
  XNOR U29870 ( .A(n28464), .B(n28463), .Z(n28466) );
  XOR U29871 ( .A(a[654]), .B(n42085), .Z(n28453) );
  AND U29872 ( .A(a[650]), .B(b[7]), .Z(n28457) );
  XNOR U29873 ( .A(n28458), .B(n28457), .Z(n28459) );
  AND U29874 ( .A(a[658]), .B(b[0]), .Z(n28417) );
  XNOR U29875 ( .A(n28417), .B(n4071), .Z(n28419) );
  NANDN U29876 ( .A(b[0]), .B(a[657]), .Z(n28418) );
  NAND U29877 ( .A(n28419), .B(n28418), .Z(n28460) );
  XNOR U29878 ( .A(n28459), .B(n28460), .Z(n28465) );
  XOR U29879 ( .A(n28466), .B(n28465), .Z(n28444) );
  NANDN U29880 ( .A(n28421), .B(n28420), .Z(n28425) );
  NANDN U29881 ( .A(n28423), .B(n28422), .Z(n28424) );
  AND U29882 ( .A(n28425), .B(n28424), .Z(n28443) );
  XNOR U29883 ( .A(n28444), .B(n28443), .Z(n28445) );
  NANDN U29884 ( .A(n28427), .B(n28426), .Z(n28431) );
  NAND U29885 ( .A(n28429), .B(n28428), .Z(n28430) );
  NAND U29886 ( .A(n28431), .B(n28430), .Z(n28446) );
  XNOR U29887 ( .A(n28445), .B(n28446), .Z(n28437) );
  XNOR U29888 ( .A(n28438), .B(n28437), .Z(n28439) );
  XNOR U29889 ( .A(n28440), .B(n28439), .Z(n28469) );
  XNOR U29890 ( .A(sreg[1674]), .B(n28469), .Z(n28471) );
  NANDN U29891 ( .A(sreg[1673]), .B(n28432), .Z(n28436) );
  NAND U29892 ( .A(n28434), .B(n28433), .Z(n28435) );
  NAND U29893 ( .A(n28436), .B(n28435), .Z(n28470) );
  XNOR U29894 ( .A(n28471), .B(n28470), .Z(c[1674]) );
  NANDN U29895 ( .A(n28438), .B(n28437), .Z(n28442) );
  NANDN U29896 ( .A(n28440), .B(n28439), .Z(n28441) );
  AND U29897 ( .A(n28442), .B(n28441), .Z(n28477) );
  NANDN U29898 ( .A(n28444), .B(n28443), .Z(n28448) );
  NANDN U29899 ( .A(n28446), .B(n28445), .Z(n28447) );
  AND U29900 ( .A(n28448), .B(n28447), .Z(n28475) );
  NAND U29901 ( .A(n42143), .B(n28449), .Z(n28451) );
  XNOR U29902 ( .A(a[653]), .B(n4165), .Z(n28486) );
  NAND U29903 ( .A(n42144), .B(n28486), .Z(n28450) );
  AND U29904 ( .A(n28451), .B(n28450), .Z(n28501) );
  XOR U29905 ( .A(a[657]), .B(n42012), .Z(n28489) );
  XNOR U29906 ( .A(n28501), .B(n28500), .Z(n28503) );
  XOR U29907 ( .A(a[655]), .B(n42085), .Z(n28493) );
  AND U29908 ( .A(a[651]), .B(b[7]), .Z(n28494) );
  XNOR U29909 ( .A(n28495), .B(n28494), .Z(n28496) );
  AND U29910 ( .A(a[659]), .B(b[0]), .Z(n28454) );
  XNOR U29911 ( .A(n28454), .B(n4071), .Z(n28456) );
  NANDN U29912 ( .A(b[0]), .B(a[658]), .Z(n28455) );
  NAND U29913 ( .A(n28456), .B(n28455), .Z(n28497) );
  XNOR U29914 ( .A(n28496), .B(n28497), .Z(n28502) );
  XOR U29915 ( .A(n28503), .B(n28502), .Z(n28481) );
  NANDN U29916 ( .A(n28458), .B(n28457), .Z(n28462) );
  NANDN U29917 ( .A(n28460), .B(n28459), .Z(n28461) );
  AND U29918 ( .A(n28462), .B(n28461), .Z(n28480) );
  XNOR U29919 ( .A(n28481), .B(n28480), .Z(n28482) );
  NANDN U29920 ( .A(n28464), .B(n28463), .Z(n28468) );
  NAND U29921 ( .A(n28466), .B(n28465), .Z(n28467) );
  NAND U29922 ( .A(n28468), .B(n28467), .Z(n28483) );
  XNOR U29923 ( .A(n28482), .B(n28483), .Z(n28474) );
  XNOR U29924 ( .A(n28475), .B(n28474), .Z(n28476) );
  XNOR U29925 ( .A(n28477), .B(n28476), .Z(n28506) );
  XNOR U29926 ( .A(sreg[1675]), .B(n28506), .Z(n28508) );
  NANDN U29927 ( .A(sreg[1674]), .B(n28469), .Z(n28473) );
  NAND U29928 ( .A(n28471), .B(n28470), .Z(n28472) );
  NAND U29929 ( .A(n28473), .B(n28472), .Z(n28507) );
  XNOR U29930 ( .A(n28508), .B(n28507), .Z(c[1675]) );
  NANDN U29931 ( .A(n28475), .B(n28474), .Z(n28479) );
  NANDN U29932 ( .A(n28477), .B(n28476), .Z(n28478) );
  AND U29933 ( .A(n28479), .B(n28478), .Z(n28514) );
  NANDN U29934 ( .A(n28481), .B(n28480), .Z(n28485) );
  NANDN U29935 ( .A(n28483), .B(n28482), .Z(n28484) );
  AND U29936 ( .A(n28485), .B(n28484), .Z(n28512) );
  NAND U29937 ( .A(n42143), .B(n28486), .Z(n28488) );
  XNOR U29938 ( .A(a[654]), .B(n4165), .Z(n28523) );
  NAND U29939 ( .A(n42144), .B(n28523), .Z(n28487) );
  AND U29940 ( .A(n28488), .B(n28487), .Z(n28538) );
  XOR U29941 ( .A(a[658]), .B(n42012), .Z(n28526) );
  XNOR U29942 ( .A(n28538), .B(n28537), .Z(n28540) );
  AND U29943 ( .A(a[660]), .B(b[0]), .Z(n28490) );
  XNOR U29944 ( .A(n28490), .B(n4071), .Z(n28492) );
  NANDN U29945 ( .A(b[0]), .B(a[659]), .Z(n28491) );
  NAND U29946 ( .A(n28492), .B(n28491), .Z(n28534) );
  XOR U29947 ( .A(a[656]), .B(n42085), .Z(n28530) );
  AND U29948 ( .A(a[652]), .B(b[7]), .Z(n28531) );
  XNOR U29949 ( .A(n28532), .B(n28531), .Z(n28533) );
  XNOR U29950 ( .A(n28534), .B(n28533), .Z(n28539) );
  XOR U29951 ( .A(n28540), .B(n28539), .Z(n28518) );
  NANDN U29952 ( .A(n28495), .B(n28494), .Z(n28499) );
  NANDN U29953 ( .A(n28497), .B(n28496), .Z(n28498) );
  AND U29954 ( .A(n28499), .B(n28498), .Z(n28517) );
  XNOR U29955 ( .A(n28518), .B(n28517), .Z(n28519) );
  NANDN U29956 ( .A(n28501), .B(n28500), .Z(n28505) );
  NAND U29957 ( .A(n28503), .B(n28502), .Z(n28504) );
  NAND U29958 ( .A(n28505), .B(n28504), .Z(n28520) );
  XNOR U29959 ( .A(n28519), .B(n28520), .Z(n28511) );
  XNOR U29960 ( .A(n28512), .B(n28511), .Z(n28513) );
  XNOR U29961 ( .A(n28514), .B(n28513), .Z(n28543) );
  XNOR U29962 ( .A(sreg[1676]), .B(n28543), .Z(n28545) );
  NANDN U29963 ( .A(sreg[1675]), .B(n28506), .Z(n28510) );
  NAND U29964 ( .A(n28508), .B(n28507), .Z(n28509) );
  NAND U29965 ( .A(n28510), .B(n28509), .Z(n28544) );
  XNOR U29966 ( .A(n28545), .B(n28544), .Z(c[1676]) );
  NANDN U29967 ( .A(n28512), .B(n28511), .Z(n28516) );
  NANDN U29968 ( .A(n28514), .B(n28513), .Z(n28515) );
  AND U29969 ( .A(n28516), .B(n28515), .Z(n28551) );
  NANDN U29970 ( .A(n28518), .B(n28517), .Z(n28522) );
  NANDN U29971 ( .A(n28520), .B(n28519), .Z(n28521) );
  AND U29972 ( .A(n28522), .B(n28521), .Z(n28549) );
  NAND U29973 ( .A(n42143), .B(n28523), .Z(n28525) );
  XNOR U29974 ( .A(a[655]), .B(n4165), .Z(n28560) );
  NAND U29975 ( .A(n42144), .B(n28560), .Z(n28524) );
  AND U29976 ( .A(n28525), .B(n28524), .Z(n28575) );
  XOR U29977 ( .A(a[659]), .B(n42012), .Z(n28563) );
  XNOR U29978 ( .A(n28575), .B(n28574), .Z(n28577) );
  AND U29979 ( .A(a[661]), .B(b[0]), .Z(n28527) );
  XNOR U29980 ( .A(n28527), .B(n4071), .Z(n28529) );
  NANDN U29981 ( .A(b[0]), .B(a[660]), .Z(n28528) );
  NAND U29982 ( .A(n28529), .B(n28528), .Z(n28571) );
  XOR U29983 ( .A(a[657]), .B(n42085), .Z(n28564) );
  AND U29984 ( .A(a[653]), .B(b[7]), .Z(n28568) );
  XNOR U29985 ( .A(n28569), .B(n28568), .Z(n28570) );
  XNOR U29986 ( .A(n28571), .B(n28570), .Z(n28576) );
  XOR U29987 ( .A(n28577), .B(n28576), .Z(n28555) );
  NANDN U29988 ( .A(n28532), .B(n28531), .Z(n28536) );
  NANDN U29989 ( .A(n28534), .B(n28533), .Z(n28535) );
  AND U29990 ( .A(n28536), .B(n28535), .Z(n28554) );
  XNOR U29991 ( .A(n28555), .B(n28554), .Z(n28556) );
  NANDN U29992 ( .A(n28538), .B(n28537), .Z(n28542) );
  NAND U29993 ( .A(n28540), .B(n28539), .Z(n28541) );
  NAND U29994 ( .A(n28542), .B(n28541), .Z(n28557) );
  XNOR U29995 ( .A(n28556), .B(n28557), .Z(n28548) );
  XNOR U29996 ( .A(n28549), .B(n28548), .Z(n28550) );
  XNOR U29997 ( .A(n28551), .B(n28550), .Z(n28580) );
  XNOR U29998 ( .A(sreg[1677]), .B(n28580), .Z(n28582) );
  NANDN U29999 ( .A(sreg[1676]), .B(n28543), .Z(n28547) );
  NAND U30000 ( .A(n28545), .B(n28544), .Z(n28546) );
  NAND U30001 ( .A(n28547), .B(n28546), .Z(n28581) );
  XNOR U30002 ( .A(n28582), .B(n28581), .Z(c[1677]) );
  NANDN U30003 ( .A(n28549), .B(n28548), .Z(n28553) );
  NANDN U30004 ( .A(n28551), .B(n28550), .Z(n28552) );
  AND U30005 ( .A(n28553), .B(n28552), .Z(n28588) );
  NANDN U30006 ( .A(n28555), .B(n28554), .Z(n28559) );
  NANDN U30007 ( .A(n28557), .B(n28556), .Z(n28558) );
  AND U30008 ( .A(n28559), .B(n28558), .Z(n28586) );
  NAND U30009 ( .A(n42143), .B(n28560), .Z(n28562) );
  XNOR U30010 ( .A(a[656]), .B(n4165), .Z(n28597) );
  NAND U30011 ( .A(n42144), .B(n28597), .Z(n28561) );
  AND U30012 ( .A(n28562), .B(n28561), .Z(n28612) );
  XOR U30013 ( .A(a[660]), .B(n42012), .Z(n28600) );
  XNOR U30014 ( .A(n28612), .B(n28611), .Z(n28614) );
  XOR U30015 ( .A(a[658]), .B(n42085), .Z(n28604) );
  AND U30016 ( .A(a[654]), .B(b[7]), .Z(n28605) );
  XNOR U30017 ( .A(n28606), .B(n28605), .Z(n28607) );
  AND U30018 ( .A(a[662]), .B(b[0]), .Z(n28565) );
  XNOR U30019 ( .A(n28565), .B(n4071), .Z(n28567) );
  NANDN U30020 ( .A(b[0]), .B(a[661]), .Z(n28566) );
  NAND U30021 ( .A(n28567), .B(n28566), .Z(n28608) );
  XNOR U30022 ( .A(n28607), .B(n28608), .Z(n28613) );
  XOR U30023 ( .A(n28614), .B(n28613), .Z(n28592) );
  NANDN U30024 ( .A(n28569), .B(n28568), .Z(n28573) );
  NANDN U30025 ( .A(n28571), .B(n28570), .Z(n28572) );
  AND U30026 ( .A(n28573), .B(n28572), .Z(n28591) );
  XNOR U30027 ( .A(n28592), .B(n28591), .Z(n28593) );
  NANDN U30028 ( .A(n28575), .B(n28574), .Z(n28579) );
  NAND U30029 ( .A(n28577), .B(n28576), .Z(n28578) );
  NAND U30030 ( .A(n28579), .B(n28578), .Z(n28594) );
  XNOR U30031 ( .A(n28593), .B(n28594), .Z(n28585) );
  XNOR U30032 ( .A(n28586), .B(n28585), .Z(n28587) );
  XNOR U30033 ( .A(n28588), .B(n28587), .Z(n28617) );
  XNOR U30034 ( .A(sreg[1678]), .B(n28617), .Z(n28619) );
  NANDN U30035 ( .A(sreg[1677]), .B(n28580), .Z(n28584) );
  NAND U30036 ( .A(n28582), .B(n28581), .Z(n28583) );
  NAND U30037 ( .A(n28584), .B(n28583), .Z(n28618) );
  XNOR U30038 ( .A(n28619), .B(n28618), .Z(c[1678]) );
  NANDN U30039 ( .A(n28586), .B(n28585), .Z(n28590) );
  NANDN U30040 ( .A(n28588), .B(n28587), .Z(n28589) );
  AND U30041 ( .A(n28590), .B(n28589), .Z(n28625) );
  NANDN U30042 ( .A(n28592), .B(n28591), .Z(n28596) );
  NANDN U30043 ( .A(n28594), .B(n28593), .Z(n28595) );
  AND U30044 ( .A(n28596), .B(n28595), .Z(n28623) );
  NAND U30045 ( .A(n42143), .B(n28597), .Z(n28599) );
  XNOR U30046 ( .A(a[657]), .B(n4165), .Z(n28634) );
  NAND U30047 ( .A(n42144), .B(n28634), .Z(n28598) );
  AND U30048 ( .A(n28599), .B(n28598), .Z(n28649) );
  XOR U30049 ( .A(a[661]), .B(n42012), .Z(n28637) );
  XNOR U30050 ( .A(n28649), .B(n28648), .Z(n28651) );
  AND U30051 ( .A(a[663]), .B(b[0]), .Z(n28601) );
  XNOR U30052 ( .A(n28601), .B(n4071), .Z(n28603) );
  NANDN U30053 ( .A(b[0]), .B(a[662]), .Z(n28602) );
  NAND U30054 ( .A(n28603), .B(n28602), .Z(n28645) );
  XOR U30055 ( .A(a[659]), .B(n42085), .Z(n28641) );
  AND U30056 ( .A(a[655]), .B(b[7]), .Z(n28642) );
  XNOR U30057 ( .A(n28643), .B(n28642), .Z(n28644) );
  XNOR U30058 ( .A(n28645), .B(n28644), .Z(n28650) );
  XOR U30059 ( .A(n28651), .B(n28650), .Z(n28629) );
  NANDN U30060 ( .A(n28606), .B(n28605), .Z(n28610) );
  NANDN U30061 ( .A(n28608), .B(n28607), .Z(n28609) );
  AND U30062 ( .A(n28610), .B(n28609), .Z(n28628) );
  XNOR U30063 ( .A(n28629), .B(n28628), .Z(n28630) );
  NANDN U30064 ( .A(n28612), .B(n28611), .Z(n28616) );
  NAND U30065 ( .A(n28614), .B(n28613), .Z(n28615) );
  NAND U30066 ( .A(n28616), .B(n28615), .Z(n28631) );
  XNOR U30067 ( .A(n28630), .B(n28631), .Z(n28622) );
  XNOR U30068 ( .A(n28623), .B(n28622), .Z(n28624) );
  XNOR U30069 ( .A(n28625), .B(n28624), .Z(n28654) );
  XNOR U30070 ( .A(sreg[1679]), .B(n28654), .Z(n28656) );
  NANDN U30071 ( .A(sreg[1678]), .B(n28617), .Z(n28621) );
  NAND U30072 ( .A(n28619), .B(n28618), .Z(n28620) );
  NAND U30073 ( .A(n28621), .B(n28620), .Z(n28655) );
  XNOR U30074 ( .A(n28656), .B(n28655), .Z(c[1679]) );
  NANDN U30075 ( .A(n28623), .B(n28622), .Z(n28627) );
  NANDN U30076 ( .A(n28625), .B(n28624), .Z(n28626) );
  AND U30077 ( .A(n28627), .B(n28626), .Z(n28662) );
  NANDN U30078 ( .A(n28629), .B(n28628), .Z(n28633) );
  NANDN U30079 ( .A(n28631), .B(n28630), .Z(n28632) );
  AND U30080 ( .A(n28633), .B(n28632), .Z(n28660) );
  NAND U30081 ( .A(n42143), .B(n28634), .Z(n28636) );
  XNOR U30082 ( .A(a[658]), .B(n4165), .Z(n28671) );
  NAND U30083 ( .A(n42144), .B(n28671), .Z(n28635) );
  AND U30084 ( .A(n28636), .B(n28635), .Z(n28686) );
  XOR U30085 ( .A(a[662]), .B(n42012), .Z(n28674) );
  XNOR U30086 ( .A(n28686), .B(n28685), .Z(n28688) );
  AND U30087 ( .A(a[664]), .B(b[0]), .Z(n28638) );
  XNOR U30088 ( .A(n28638), .B(n4071), .Z(n28640) );
  NANDN U30089 ( .A(b[0]), .B(a[663]), .Z(n28639) );
  NAND U30090 ( .A(n28640), .B(n28639), .Z(n28682) );
  XOR U30091 ( .A(a[660]), .B(n42085), .Z(n28678) );
  AND U30092 ( .A(a[656]), .B(b[7]), .Z(n28679) );
  XNOR U30093 ( .A(n28680), .B(n28679), .Z(n28681) );
  XNOR U30094 ( .A(n28682), .B(n28681), .Z(n28687) );
  XOR U30095 ( .A(n28688), .B(n28687), .Z(n28666) );
  NANDN U30096 ( .A(n28643), .B(n28642), .Z(n28647) );
  NANDN U30097 ( .A(n28645), .B(n28644), .Z(n28646) );
  AND U30098 ( .A(n28647), .B(n28646), .Z(n28665) );
  XNOR U30099 ( .A(n28666), .B(n28665), .Z(n28667) );
  NANDN U30100 ( .A(n28649), .B(n28648), .Z(n28653) );
  NAND U30101 ( .A(n28651), .B(n28650), .Z(n28652) );
  NAND U30102 ( .A(n28653), .B(n28652), .Z(n28668) );
  XNOR U30103 ( .A(n28667), .B(n28668), .Z(n28659) );
  XNOR U30104 ( .A(n28660), .B(n28659), .Z(n28661) );
  XNOR U30105 ( .A(n28662), .B(n28661), .Z(n28691) );
  XNOR U30106 ( .A(sreg[1680]), .B(n28691), .Z(n28693) );
  NANDN U30107 ( .A(sreg[1679]), .B(n28654), .Z(n28658) );
  NAND U30108 ( .A(n28656), .B(n28655), .Z(n28657) );
  NAND U30109 ( .A(n28658), .B(n28657), .Z(n28692) );
  XNOR U30110 ( .A(n28693), .B(n28692), .Z(c[1680]) );
  NANDN U30111 ( .A(n28660), .B(n28659), .Z(n28664) );
  NANDN U30112 ( .A(n28662), .B(n28661), .Z(n28663) );
  AND U30113 ( .A(n28664), .B(n28663), .Z(n28699) );
  NANDN U30114 ( .A(n28666), .B(n28665), .Z(n28670) );
  NANDN U30115 ( .A(n28668), .B(n28667), .Z(n28669) );
  AND U30116 ( .A(n28670), .B(n28669), .Z(n28697) );
  NAND U30117 ( .A(n42143), .B(n28671), .Z(n28673) );
  XNOR U30118 ( .A(a[659]), .B(n4166), .Z(n28708) );
  NAND U30119 ( .A(n42144), .B(n28708), .Z(n28672) );
  AND U30120 ( .A(n28673), .B(n28672), .Z(n28723) );
  XOR U30121 ( .A(a[663]), .B(n42012), .Z(n28711) );
  XNOR U30122 ( .A(n28723), .B(n28722), .Z(n28725) );
  AND U30123 ( .A(a[665]), .B(b[0]), .Z(n28675) );
  XNOR U30124 ( .A(n28675), .B(n4071), .Z(n28677) );
  NANDN U30125 ( .A(b[0]), .B(a[664]), .Z(n28676) );
  NAND U30126 ( .A(n28677), .B(n28676), .Z(n28719) );
  XOR U30127 ( .A(a[661]), .B(n42085), .Z(n28715) );
  AND U30128 ( .A(a[657]), .B(b[7]), .Z(n28716) );
  XNOR U30129 ( .A(n28717), .B(n28716), .Z(n28718) );
  XNOR U30130 ( .A(n28719), .B(n28718), .Z(n28724) );
  XOR U30131 ( .A(n28725), .B(n28724), .Z(n28703) );
  NANDN U30132 ( .A(n28680), .B(n28679), .Z(n28684) );
  NANDN U30133 ( .A(n28682), .B(n28681), .Z(n28683) );
  AND U30134 ( .A(n28684), .B(n28683), .Z(n28702) );
  XNOR U30135 ( .A(n28703), .B(n28702), .Z(n28704) );
  NANDN U30136 ( .A(n28686), .B(n28685), .Z(n28690) );
  NAND U30137 ( .A(n28688), .B(n28687), .Z(n28689) );
  NAND U30138 ( .A(n28690), .B(n28689), .Z(n28705) );
  XNOR U30139 ( .A(n28704), .B(n28705), .Z(n28696) );
  XNOR U30140 ( .A(n28697), .B(n28696), .Z(n28698) );
  XNOR U30141 ( .A(n28699), .B(n28698), .Z(n28728) );
  XNOR U30142 ( .A(sreg[1681]), .B(n28728), .Z(n28730) );
  NANDN U30143 ( .A(sreg[1680]), .B(n28691), .Z(n28695) );
  NAND U30144 ( .A(n28693), .B(n28692), .Z(n28694) );
  NAND U30145 ( .A(n28695), .B(n28694), .Z(n28729) );
  XNOR U30146 ( .A(n28730), .B(n28729), .Z(c[1681]) );
  NANDN U30147 ( .A(n28697), .B(n28696), .Z(n28701) );
  NANDN U30148 ( .A(n28699), .B(n28698), .Z(n28700) );
  AND U30149 ( .A(n28701), .B(n28700), .Z(n28736) );
  NANDN U30150 ( .A(n28703), .B(n28702), .Z(n28707) );
  NANDN U30151 ( .A(n28705), .B(n28704), .Z(n28706) );
  AND U30152 ( .A(n28707), .B(n28706), .Z(n28734) );
  NAND U30153 ( .A(n42143), .B(n28708), .Z(n28710) );
  XNOR U30154 ( .A(a[660]), .B(n4166), .Z(n28745) );
  NAND U30155 ( .A(n42144), .B(n28745), .Z(n28709) );
  AND U30156 ( .A(n28710), .B(n28709), .Z(n28760) );
  XOR U30157 ( .A(a[664]), .B(n42012), .Z(n28748) );
  XNOR U30158 ( .A(n28760), .B(n28759), .Z(n28762) );
  AND U30159 ( .A(a[666]), .B(b[0]), .Z(n28712) );
  XNOR U30160 ( .A(n28712), .B(n4071), .Z(n28714) );
  NANDN U30161 ( .A(b[0]), .B(a[665]), .Z(n28713) );
  NAND U30162 ( .A(n28714), .B(n28713), .Z(n28756) );
  XOR U30163 ( .A(a[662]), .B(n42085), .Z(n28752) );
  AND U30164 ( .A(a[658]), .B(b[7]), .Z(n28753) );
  XNOR U30165 ( .A(n28754), .B(n28753), .Z(n28755) );
  XNOR U30166 ( .A(n28756), .B(n28755), .Z(n28761) );
  XOR U30167 ( .A(n28762), .B(n28761), .Z(n28740) );
  NANDN U30168 ( .A(n28717), .B(n28716), .Z(n28721) );
  NANDN U30169 ( .A(n28719), .B(n28718), .Z(n28720) );
  AND U30170 ( .A(n28721), .B(n28720), .Z(n28739) );
  XNOR U30171 ( .A(n28740), .B(n28739), .Z(n28741) );
  NANDN U30172 ( .A(n28723), .B(n28722), .Z(n28727) );
  NAND U30173 ( .A(n28725), .B(n28724), .Z(n28726) );
  NAND U30174 ( .A(n28727), .B(n28726), .Z(n28742) );
  XNOR U30175 ( .A(n28741), .B(n28742), .Z(n28733) );
  XNOR U30176 ( .A(n28734), .B(n28733), .Z(n28735) );
  XNOR U30177 ( .A(n28736), .B(n28735), .Z(n28765) );
  XNOR U30178 ( .A(sreg[1682]), .B(n28765), .Z(n28767) );
  NANDN U30179 ( .A(sreg[1681]), .B(n28728), .Z(n28732) );
  NAND U30180 ( .A(n28730), .B(n28729), .Z(n28731) );
  NAND U30181 ( .A(n28732), .B(n28731), .Z(n28766) );
  XNOR U30182 ( .A(n28767), .B(n28766), .Z(c[1682]) );
  NANDN U30183 ( .A(n28734), .B(n28733), .Z(n28738) );
  NANDN U30184 ( .A(n28736), .B(n28735), .Z(n28737) );
  AND U30185 ( .A(n28738), .B(n28737), .Z(n28773) );
  NANDN U30186 ( .A(n28740), .B(n28739), .Z(n28744) );
  NANDN U30187 ( .A(n28742), .B(n28741), .Z(n28743) );
  AND U30188 ( .A(n28744), .B(n28743), .Z(n28771) );
  NAND U30189 ( .A(n42143), .B(n28745), .Z(n28747) );
  XNOR U30190 ( .A(a[661]), .B(n4166), .Z(n28782) );
  NAND U30191 ( .A(n42144), .B(n28782), .Z(n28746) );
  AND U30192 ( .A(n28747), .B(n28746), .Z(n28797) );
  XOR U30193 ( .A(a[665]), .B(n42012), .Z(n28785) );
  XNOR U30194 ( .A(n28797), .B(n28796), .Z(n28799) );
  AND U30195 ( .A(a[667]), .B(b[0]), .Z(n28749) );
  XNOR U30196 ( .A(n28749), .B(n4071), .Z(n28751) );
  NANDN U30197 ( .A(b[0]), .B(a[666]), .Z(n28750) );
  NAND U30198 ( .A(n28751), .B(n28750), .Z(n28793) );
  XOR U30199 ( .A(a[663]), .B(n42085), .Z(n28789) );
  AND U30200 ( .A(a[659]), .B(b[7]), .Z(n28790) );
  XNOR U30201 ( .A(n28791), .B(n28790), .Z(n28792) );
  XNOR U30202 ( .A(n28793), .B(n28792), .Z(n28798) );
  XOR U30203 ( .A(n28799), .B(n28798), .Z(n28777) );
  NANDN U30204 ( .A(n28754), .B(n28753), .Z(n28758) );
  NANDN U30205 ( .A(n28756), .B(n28755), .Z(n28757) );
  AND U30206 ( .A(n28758), .B(n28757), .Z(n28776) );
  XNOR U30207 ( .A(n28777), .B(n28776), .Z(n28778) );
  NANDN U30208 ( .A(n28760), .B(n28759), .Z(n28764) );
  NAND U30209 ( .A(n28762), .B(n28761), .Z(n28763) );
  NAND U30210 ( .A(n28764), .B(n28763), .Z(n28779) );
  XNOR U30211 ( .A(n28778), .B(n28779), .Z(n28770) );
  XNOR U30212 ( .A(n28771), .B(n28770), .Z(n28772) );
  XNOR U30213 ( .A(n28773), .B(n28772), .Z(n28802) );
  XNOR U30214 ( .A(sreg[1683]), .B(n28802), .Z(n28804) );
  NANDN U30215 ( .A(sreg[1682]), .B(n28765), .Z(n28769) );
  NAND U30216 ( .A(n28767), .B(n28766), .Z(n28768) );
  NAND U30217 ( .A(n28769), .B(n28768), .Z(n28803) );
  XNOR U30218 ( .A(n28804), .B(n28803), .Z(c[1683]) );
  NANDN U30219 ( .A(n28771), .B(n28770), .Z(n28775) );
  NANDN U30220 ( .A(n28773), .B(n28772), .Z(n28774) );
  AND U30221 ( .A(n28775), .B(n28774), .Z(n28810) );
  NANDN U30222 ( .A(n28777), .B(n28776), .Z(n28781) );
  NANDN U30223 ( .A(n28779), .B(n28778), .Z(n28780) );
  AND U30224 ( .A(n28781), .B(n28780), .Z(n28808) );
  NAND U30225 ( .A(n42143), .B(n28782), .Z(n28784) );
  XNOR U30226 ( .A(a[662]), .B(n4166), .Z(n28819) );
  NAND U30227 ( .A(n42144), .B(n28819), .Z(n28783) );
  AND U30228 ( .A(n28784), .B(n28783), .Z(n28834) );
  XOR U30229 ( .A(a[666]), .B(n42012), .Z(n28822) );
  XNOR U30230 ( .A(n28834), .B(n28833), .Z(n28836) );
  AND U30231 ( .A(a[668]), .B(b[0]), .Z(n28786) );
  XNOR U30232 ( .A(n28786), .B(n4071), .Z(n28788) );
  NANDN U30233 ( .A(b[0]), .B(a[667]), .Z(n28787) );
  NAND U30234 ( .A(n28788), .B(n28787), .Z(n28830) );
  XOR U30235 ( .A(a[664]), .B(n42085), .Z(n28823) );
  AND U30236 ( .A(a[660]), .B(b[7]), .Z(n28827) );
  XNOR U30237 ( .A(n28828), .B(n28827), .Z(n28829) );
  XNOR U30238 ( .A(n28830), .B(n28829), .Z(n28835) );
  XOR U30239 ( .A(n28836), .B(n28835), .Z(n28814) );
  NANDN U30240 ( .A(n28791), .B(n28790), .Z(n28795) );
  NANDN U30241 ( .A(n28793), .B(n28792), .Z(n28794) );
  AND U30242 ( .A(n28795), .B(n28794), .Z(n28813) );
  XNOR U30243 ( .A(n28814), .B(n28813), .Z(n28815) );
  NANDN U30244 ( .A(n28797), .B(n28796), .Z(n28801) );
  NAND U30245 ( .A(n28799), .B(n28798), .Z(n28800) );
  NAND U30246 ( .A(n28801), .B(n28800), .Z(n28816) );
  XNOR U30247 ( .A(n28815), .B(n28816), .Z(n28807) );
  XNOR U30248 ( .A(n28808), .B(n28807), .Z(n28809) );
  XNOR U30249 ( .A(n28810), .B(n28809), .Z(n28839) );
  XNOR U30250 ( .A(sreg[1684]), .B(n28839), .Z(n28841) );
  NANDN U30251 ( .A(sreg[1683]), .B(n28802), .Z(n28806) );
  NAND U30252 ( .A(n28804), .B(n28803), .Z(n28805) );
  NAND U30253 ( .A(n28806), .B(n28805), .Z(n28840) );
  XNOR U30254 ( .A(n28841), .B(n28840), .Z(c[1684]) );
  NANDN U30255 ( .A(n28808), .B(n28807), .Z(n28812) );
  NANDN U30256 ( .A(n28810), .B(n28809), .Z(n28811) );
  AND U30257 ( .A(n28812), .B(n28811), .Z(n28847) );
  NANDN U30258 ( .A(n28814), .B(n28813), .Z(n28818) );
  NANDN U30259 ( .A(n28816), .B(n28815), .Z(n28817) );
  AND U30260 ( .A(n28818), .B(n28817), .Z(n28845) );
  NAND U30261 ( .A(n42143), .B(n28819), .Z(n28821) );
  XNOR U30262 ( .A(a[663]), .B(n4166), .Z(n28856) );
  NAND U30263 ( .A(n42144), .B(n28856), .Z(n28820) );
  AND U30264 ( .A(n28821), .B(n28820), .Z(n28871) );
  XOR U30265 ( .A(a[667]), .B(n42012), .Z(n28859) );
  XNOR U30266 ( .A(n28871), .B(n28870), .Z(n28873) );
  XOR U30267 ( .A(a[665]), .B(n42085), .Z(n28860) );
  AND U30268 ( .A(a[661]), .B(b[7]), .Z(n28864) );
  XNOR U30269 ( .A(n28865), .B(n28864), .Z(n28866) );
  AND U30270 ( .A(a[669]), .B(b[0]), .Z(n28824) );
  XNOR U30271 ( .A(n28824), .B(n4071), .Z(n28826) );
  NANDN U30272 ( .A(b[0]), .B(a[668]), .Z(n28825) );
  NAND U30273 ( .A(n28826), .B(n28825), .Z(n28867) );
  XNOR U30274 ( .A(n28866), .B(n28867), .Z(n28872) );
  XOR U30275 ( .A(n28873), .B(n28872), .Z(n28851) );
  NANDN U30276 ( .A(n28828), .B(n28827), .Z(n28832) );
  NANDN U30277 ( .A(n28830), .B(n28829), .Z(n28831) );
  AND U30278 ( .A(n28832), .B(n28831), .Z(n28850) );
  XNOR U30279 ( .A(n28851), .B(n28850), .Z(n28852) );
  NANDN U30280 ( .A(n28834), .B(n28833), .Z(n28838) );
  NAND U30281 ( .A(n28836), .B(n28835), .Z(n28837) );
  NAND U30282 ( .A(n28838), .B(n28837), .Z(n28853) );
  XNOR U30283 ( .A(n28852), .B(n28853), .Z(n28844) );
  XNOR U30284 ( .A(n28845), .B(n28844), .Z(n28846) );
  XNOR U30285 ( .A(n28847), .B(n28846), .Z(n28876) );
  XNOR U30286 ( .A(sreg[1685]), .B(n28876), .Z(n28878) );
  NANDN U30287 ( .A(sreg[1684]), .B(n28839), .Z(n28843) );
  NAND U30288 ( .A(n28841), .B(n28840), .Z(n28842) );
  NAND U30289 ( .A(n28843), .B(n28842), .Z(n28877) );
  XNOR U30290 ( .A(n28878), .B(n28877), .Z(c[1685]) );
  NANDN U30291 ( .A(n28845), .B(n28844), .Z(n28849) );
  NANDN U30292 ( .A(n28847), .B(n28846), .Z(n28848) );
  AND U30293 ( .A(n28849), .B(n28848), .Z(n28884) );
  NANDN U30294 ( .A(n28851), .B(n28850), .Z(n28855) );
  NANDN U30295 ( .A(n28853), .B(n28852), .Z(n28854) );
  AND U30296 ( .A(n28855), .B(n28854), .Z(n28882) );
  NAND U30297 ( .A(n42143), .B(n28856), .Z(n28858) );
  XNOR U30298 ( .A(a[664]), .B(n4166), .Z(n28893) );
  NAND U30299 ( .A(n42144), .B(n28893), .Z(n28857) );
  AND U30300 ( .A(n28858), .B(n28857), .Z(n28908) );
  XOR U30301 ( .A(a[668]), .B(n42012), .Z(n28896) );
  XNOR U30302 ( .A(n28908), .B(n28907), .Z(n28910) );
  XOR U30303 ( .A(a[666]), .B(n42085), .Z(n28900) );
  AND U30304 ( .A(a[662]), .B(b[7]), .Z(n28901) );
  XNOR U30305 ( .A(n28902), .B(n28901), .Z(n28903) );
  AND U30306 ( .A(a[670]), .B(b[0]), .Z(n28861) );
  XNOR U30307 ( .A(n28861), .B(n4071), .Z(n28863) );
  NANDN U30308 ( .A(b[0]), .B(a[669]), .Z(n28862) );
  NAND U30309 ( .A(n28863), .B(n28862), .Z(n28904) );
  XNOR U30310 ( .A(n28903), .B(n28904), .Z(n28909) );
  XOR U30311 ( .A(n28910), .B(n28909), .Z(n28888) );
  NANDN U30312 ( .A(n28865), .B(n28864), .Z(n28869) );
  NANDN U30313 ( .A(n28867), .B(n28866), .Z(n28868) );
  AND U30314 ( .A(n28869), .B(n28868), .Z(n28887) );
  XNOR U30315 ( .A(n28888), .B(n28887), .Z(n28889) );
  NANDN U30316 ( .A(n28871), .B(n28870), .Z(n28875) );
  NAND U30317 ( .A(n28873), .B(n28872), .Z(n28874) );
  NAND U30318 ( .A(n28875), .B(n28874), .Z(n28890) );
  XNOR U30319 ( .A(n28889), .B(n28890), .Z(n28881) );
  XNOR U30320 ( .A(n28882), .B(n28881), .Z(n28883) );
  XNOR U30321 ( .A(n28884), .B(n28883), .Z(n28913) );
  XNOR U30322 ( .A(sreg[1686]), .B(n28913), .Z(n28915) );
  NANDN U30323 ( .A(sreg[1685]), .B(n28876), .Z(n28880) );
  NAND U30324 ( .A(n28878), .B(n28877), .Z(n28879) );
  NAND U30325 ( .A(n28880), .B(n28879), .Z(n28914) );
  XNOR U30326 ( .A(n28915), .B(n28914), .Z(c[1686]) );
  NANDN U30327 ( .A(n28882), .B(n28881), .Z(n28886) );
  NANDN U30328 ( .A(n28884), .B(n28883), .Z(n28885) );
  AND U30329 ( .A(n28886), .B(n28885), .Z(n28921) );
  NANDN U30330 ( .A(n28888), .B(n28887), .Z(n28892) );
  NANDN U30331 ( .A(n28890), .B(n28889), .Z(n28891) );
  AND U30332 ( .A(n28892), .B(n28891), .Z(n28919) );
  NAND U30333 ( .A(n42143), .B(n28893), .Z(n28895) );
  XNOR U30334 ( .A(a[665]), .B(n4166), .Z(n28930) );
  NAND U30335 ( .A(n42144), .B(n28930), .Z(n28894) );
  AND U30336 ( .A(n28895), .B(n28894), .Z(n28945) );
  XOR U30337 ( .A(a[669]), .B(n42012), .Z(n28933) );
  XNOR U30338 ( .A(n28945), .B(n28944), .Z(n28947) );
  AND U30339 ( .A(a[671]), .B(b[0]), .Z(n28897) );
  XNOR U30340 ( .A(n28897), .B(n4071), .Z(n28899) );
  NANDN U30341 ( .A(b[0]), .B(a[670]), .Z(n28898) );
  NAND U30342 ( .A(n28899), .B(n28898), .Z(n28941) );
  XOR U30343 ( .A(a[667]), .B(n42085), .Z(n28934) );
  AND U30344 ( .A(a[663]), .B(b[7]), .Z(n28938) );
  XNOR U30345 ( .A(n28939), .B(n28938), .Z(n28940) );
  XNOR U30346 ( .A(n28941), .B(n28940), .Z(n28946) );
  XOR U30347 ( .A(n28947), .B(n28946), .Z(n28925) );
  NANDN U30348 ( .A(n28902), .B(n28901), .Z(n28906) );
  NANDN U30349 ( .A(n28904), .B(n28903), .Z(n28905) );
  AND U30350 ( .A(n28906), .B(n28905), .Z(n28924) );
  XNOR U30351 ( .A(n28925), .B(n28924), .Z(n28926) );
  NANDN U30352 ( .A(n28908), .B(n28907), .Z(n28912) );
  NAND U30353 ( .A(n28910), .B(n28909), .Z(n28911) );
  NAND U30354 ( .A(n28912), .B(n28911), .Z(n28927) );
  XNOR U30355 ( .A(n28926), .B(n28927), .Z(n28918) );
  XNOR U30356 ( .A(n28919), .B(n28918), .Z(n28920) );
  XNOR U30357 ( .A(n28921), .B(n28920), .Z(n28950) );
  XNOR U30358 ( .A(sreg[1687]), .B(n28950), .Z(n28952) );
  NANDN U30359 ( .A(sreg[1686]), .B(n28913), .Z(n28917) );
  NAND U30360 ( .A(n28915), .B(n28914), .Z(n28916) );
  NAND U30361 ( .A(n28917), .B(n28916), .Z(n28951) );
  XNOR U30362 ( .A(n28952), .B(n28951), .Z(c[1687]) );
  NANDN U30363 ( .A(n28919), .B(n28918), .Z(n28923) );
  NANDN U30364 ( .A(n28921), .B(n28920), .Z(n28922) );
  AND U30365 ( .A(n28923), .B(n28922), .Z(n28958) );
  NANDN U30366 ( .A(n28925), .B(n28924), .Z(n28929) );
  NANDN U30367 ( .A(n28927), .B(n28926), .Z(n28928) );
  AND U30368 ( .A(n28929), .B(n28928), .Z(n28956) );
  NAND U30369 ( .A(n42143), .B(n28930), .Z(n28932) );
  XNOR U30370 ( .A(a[666]), .B(n4167), .Z(n28967) );
  NAND U30371 ( .A(n42144), .B(n28967), .Z(n28931) );
  AND U30372 ( .A(n28932), .B(n28931), .Z(n28982) );
  XOR U30373 ( .A(a[670]), .B(n42012), .Z(n28970) );
  XNOR U30374 ( .A(n28982), .B(n28981), .Z(n28984) );
  XOR U30375 ( .A(a[668]), .B(n42085), .Z(n28974) );
  AND U30376 ( .A(a[664]), .B(b[7]), .Z(n28975) );
  XNOR U30377 ( .A(n28976), .B(n28975), .Z(n28977) );
  AND U30378 ( .A(a[672]), .B(b[0]), .Z(n28935) );
  XNOR U30379 ( .A(n28935), .B(n4071), .Z(n28937) );
  NANDN U30380 ( .A(b[0]), .B(a[671]), .Z(n28936) );
  NAND U30381 ( .A(n28937), .B(n28936), .Z(n28978) );
  XNOR U30382 ( .A(n28977), .B(n28978), .Z(n28983) );
  XOR U30383 ( .A(n28984), .B(n28983), .Z(n28962) );
  NANDN U30384 ( .A(n28939), .B(n28938), .Z(n28943) );
  NANDN U30385 ( .A(n28941), .B(n28940), .Z(n28942) );
  AND U30386 ( .A(n28943), .B(n28942), .Z(n28961) );
  XNOR U30387 ( .A(n28962), .B(n28961), .Z(n28963) );
  NANDN U30388 ( .A(n28945), .B(n28944), .Z(n28949) );
  NAND U30389 ( .A(n28947), .B(n28946), .Z(n28948) );
  NAND U30390 ( .A(n28949), .B(n28948), .Z(n28964) );
  XNOR U30391 ( .A(n28963), .B(n28964), .Z(n28955) );
  XNOR U30392 ( .A(n28956), .B(n28955), .Z(n28957) );
  XNOR U30393 ( .A(n28958), .B(n28957), .Z(n28987) );
  XNOR U30394 ( .A(sreg[1688]), .B(n28987), .Z(n28989) );
  NANDN U30395 ( .A(sreg[1687]), .B(n28950), .Z(n28954) );
  NAND U30396 ( .A(n28952), .B(n28951), .Z(n28953) );
  NAND U30397 ( .A(n28954), .B(n28953), .Z(n28988) );
  XNOR U30398 ( .A(n28989), .B(n28988), .Z(c[1688]) );
  NANDN U30399 ( .A(n28956), .B(n28955), .Z(n28960) );
  NANDN U30400 ( .A(n28958), .B(n28957), .Z(n28959) );
  AND U30401 ( .A(n28960), .B(n28959), .Z(n28995) );
  NANDN U30402 ( .A(n28962), .B(n28961), .Z(n28966) );
  NANDN U30403 ( .A(n28964), .B(n28963), .Z(n28965) );
  AND U30404 ( .A(n28966), .B(n28965), .Z(n28993) );
  NAND U30405 ( .A(n42143), .B(n28967), .Z(n28969) );
  XNOR U30406 ( .A(a[667]), .B(n4167), .Z(n29004) );
  NAND U30407 ( .A(n42144), .B(n29004), .Z(n28968) );
  AND U30408 ( .A(n28969), .B(n28968), .Z(n29019) );
  XOR U30409 ( .A(a[671]), .B(n42012), .Z(n29007) );
  XNOR U30410 ( .A(n29019), .B(n29018), .Z(n29021) );
  AND U30411 ( .A(a[673]), .B(b[0]), .Z(n28971) );
  XNOR U30412 ( .A(n28971), .B(n4071), .Z(n28973) );
  NANDN U30413 ( .A(b[0]), .B(a[672]), .Z(n28972) );
  NAND U30414 ( .A(n28973), .B(n28972), .Z(n29015) );
  XOR U30415 ( .A(a[669]), .B(n42085), .Z(n29011) );
  AND U30416 ( .A(a[665]), .B(b[7]), .Z(n29012) );
  XNOR U30417 ( .A(n29013), .B(n29012), .Z(n29014) );
  XNOR U30418 ( .A(n29015), .B(n29014), .Z(n29020) );
  XOR U30419 ( .A(n29021), .B(n29020), .Z(n28999) );
  NANDN U30420 ( .A(n28976), .B(n28975), .Z(n28980) );
  NANDN U30421 ( .A(n28978), .B(n28977), .Z(n28979) );
  AND U30422 ( .A(n28980), .B(n28979), .Z(n28998) );
  XNOR U30423 ( .A(n28999), .B(n28998), .Z(n29000) );
  NANDN U30424 ( .A(n28982), .B(n28981), .Z(n28986) );
  NAND U30425 ( .A(n28984), .B(n28983), .Z(n28985) );
  NAND U30426 ( .A(n28986), .B(n28985), .Z(n29001) );
  XNOR U30427 ( .A(n29000), .B(n29001), .Z(n28992) );
  XNOR U30428 ( .A(n28993), .B(n28992), .Z(n28994) );
  XNOR U30429 ( .A(n28995), .B(n28994), .Z(n29024) );
  XNOR U30430 ( .A(sreg[1689]), .B(n29024), .Z(n29026) );
  NANDN U30431 ( .A(sreg[1688]), .B(n28987), .Z(n28991) );
  NAND U30432 ( .A(n28989), .B(n28988), .Z(n28990) );
  NAND U30433 ( .A(n28991), .B(n28990), .Z(n29025) );
  XNOR U30434 ( .A(n29026), .B(n29025), .Z(c[1689]) );
  NANDN U30435 ( .A(n28993), .B(n28992), .Z(n28997) );
  NANDN U30436 ( .A(n28995), .B(n28994), .Z(n28996) );
  AND U30437 ( .A(n28997), .B(n28996), .Z(n29032) );
  NANDN U30438 ( .A(n28999), .B(n28998), .Z(n29003) );
  NANDN U30439 ( .A(n29001), .B(n29000), .Z(n29002) );
  AND U30440 ( .A(n29003), .B(n29002), .Z(n29030) );
  NAND U30441 ( .A(n42143), .B(n29004), .Z(n29006) );
  XNOR U30442 ( .A(a[668]), .B(n4167), .Z(n29041) );
  NAND U30443 ( .A(n42144), .B(n29041), .Z(n29005) );
  AND U30444 ( .A(n29006), .B(n29005), .Z(n29056) );
  XOR U30445 ( .A(a[672]), .B(n42012), .Z(n29044) );
  XNOR U30446 ( .A(n29056), .B(n29055), .Z(n29058) );
  AND U30447 ( .A(a[674]), .B(b[0]), .Z(n29008) );
  XNOR U30448 ( .A(n29008), .B(n4071), .Z(n29010) );
  NANDN U30449 ( .A(b[0]), .B(a[673]), .Z(n29009) );
  NAND U30450 ( .A(n29010), .B(n29009), .Z(n29052) );
  XOR U30451 ( .A(a[670]), .B(n42085), .Z(n29045) );
  AND U30452 ( .A(a[666]), .B(b[7]), .Z(n29049) );
  XNOR U30453 ( .A(n29050), .B(n29049), .Z(n29051) );
  XNOR U30454 ( .A(n29052), .B(n29051), .Z(n29057) );
  XOR U30455 ( .A(n29058), .B(n29057), .Z(n29036) );
  NANDN U30456 ( .A(n29013), .B(n29012), .Z(n29017) );
  NANDN U30457 ( .A(n29015), .B(n29014), .Z(n29016) );
  AND U30458 ( .A(n29017), .B(n29016), .Z(n29035) );
  XNOR U30459 ( .A(n29036), .B(n29035), .Z(n29037) );
  NANDN U30460 ( .A(n29019), .B(n29018), .Z(n29023) );
  NAND U30461 ( .A(n29021), .B(n29020), .Z(n29022) );
  NAND U30462 ( .A(n29023), .B(n29022), .Z(n29038) );
  XNOR U30463 ( .A(n29037), .B(n29038), .Z(n29029) );
  XNOR U30464 ( .A(n29030), .B(n29029), .Z(n29031) );
  XNOR U30465 ( .A(n29032), .B(n29031), .Z(n29061) );
  XNOR U30466 ( .A(sreg[1690]), .B(n29061), .Z(n29063) );
  NANDN U30467 ( .A(sreg[1689]), .B(n29024), .Z(n29028) );
  NAND U30468 ( .A(n29026), .B(n29025), .Z(n29027) );
  NAND U30469 ( .A(n29028), .B(n29027), .Z(n29062) );
  XNOR U30470 ( .A(n29063), .B(n29062), .Z(c[1690]) );
  NANDN U30471 ( .A(n29030), .B(n29029), .Z(n29034) );
  NANDN U30472 ( .A(n29032), .B(n29031), .Z(n29033) );
  AND U30473 ( .A(n29034), .B(n29033), .Z(n29069) );
  NANDN U30474 ( .A(n29036), .B(n29035), .Z(n29040) );
  NANDN U30475 ( .A(n29038), .B(n29037), .Z(n29039) );
  AND U30476 ( .A(n29040), .B(n29039), .Z(n29067) );
  NAND U30477 ( .A(n42143), .B(n29041), .Z(n29043) );
  XNOR U30478 ( .A(a[669]), .B(n4167), .Z(n29078) );
  NAND U30479 ( .A(n42144), .B(n29078), .Z(n29042) );
  AND U30480 ( .A(n29043), .B(n29042), .Z(n29093) );
  XOR U30481 ( .A(a[673]), .B(n42012), .Z(n29081) );
  XNOR U30482 ( .A(n29093), .B(n29092), .Z(n29095) );
  XOR U30483 ( .A(a[671]), .B(n42085), .Z(n29082) );
  AND U30484 ( .A(a[667]), .B(b[7]), .Z(n29086) );
  XNOR U30485 ( .A(n29087), .B(n29086), .Z(n29088) );
  AND U30486 ( .A(a[675]), .B(b[0]), .Z(n29046) );
  XNOR U30487 ( .A(n29046), .B(n4071), .Z(n29048) );
  NANDN U30488 ( .A(b[0]), .B(a[674]), .Z(n29047) );
  NAND U30489 ( .A(n29048), .B(n29047), .Z(n29089) );
  XNOR U30490 ( .A(n29088), .B(n29089), .Z(n29094) );
  XOR U30491 ( .A(n29095), .B(n29094), .Z(n29073) );
  NANDN U30492 ( .A(n29050), .B(n29049), .Z(n29054) );
  NANDN U30493 ( .A(n29052), .B(n29051), .Z(n29053) );
  AND U30494 ( .A(n29054), .B(n29053), .Z(n29072) );
  XNOR U30495 ( .A(n29073), .B(n29072), .Z(n29074) );
  NANDN U30496 ( .A(n29056), .B(n29055), .Z(n29060) );
  NAND U30497 ( .A(n29058), .B(n29057), .Z(n29059) );
  NAND U30498 ( .A(n29060), .B(n29059), .Z(n29075) );
  XNOR U30499 ( .A(n29074), .B(n29075), .Z(n29066) );
  XNOR U30500 ( .A(n29067), .B(n29066), .Z(n29068) );
  XNOR U30501 ( .A(n29069), .B(n29068), .Z(n29098) );
  XNOR U30502 ( .A(sreg[1691]), .B(n29098), .Z(n29100) );
  NANDN U30503 ( .A(sreg[1690]), .B(n29061), .Z(n29065) );
  NAND U30504 ( .A(n29063), .B(n29062), .Z(n29064) );
  NAND U30505 ( .A(n29065), .B(n29064), .Z(n29099) );
  XNOR U30506 ( .A(n29100), .B(n29099), .Z(c[1691]) );
  NANDN U30507 ( .A(n29067), .B(n29066), .Z(n29071) );
  NANDN U30508 ( .A(n29069), .B(n29068), .Z(n29070) );
  AND U30509 ( .A(n29071), .B(n29070), .Z(n29106) );
  NANDN U30510 ( .A(n29073), .B(n29072), .Z(n29077) );
  NANDN U30511 ( .A(n29075), .B(n29074), .Z(n29076) );
  AND U30512 ( .A(n29077), .B(n29076), .Z(n29104) );
  NAND U30513 ( .A(n42143), .B(n29078), .Z(n29080) );
  XNOR U30514 ( .A(a[670]), .B(n4167), .Z(n29115) );
  NAND U30515 ( .A(n42144), .B(n29115), .Z(n29079) );
  AND U30516 ( .A(n29080), .B(n29079), .Z(n29130) );
  XOR U30517 ( .A(a[674]), .B(n42012), .Z(n29118) );
  XNOR U30518 ( .A(n29130), .B(n29129), .Z(n29132) );
  XOR U30519 ( .A(a[672]), .B(n42085), .Z(n29122) );
  AND U30520 ( .A(a[668]), .B(b[7]), .Z(n29123) );
  XNOR U30521 ( .A(n29124), .B(n29123), .Z(n29125) );
  AND U30522 ( .A(a[676]), .B(b[0]), .Z(n29083) );
  XNOR U30523 ( .A(n29083), .B(n4071), .Z(n29085) );
  NANDN U30524 ( .A(b[0]), .B(a[675]), .Z(n29084) );
  NAND U30525 ( .A(n29085), .B(n29084), .Z(n29126) );
  XNOR U30526 ( .A(n29125), .B(n29126), .Z(n29131) );
  XOR U30527 ( .A(n29132), .B(n29131), .Z(n29110) );
  NANDN U30528 ( .A(n29087), .B(n29086), .Z(n29091) );
  NANDN U30529 ( .A(n29089), .B(n29088), .Z(n29090) );
  AND U30530 ( .A(n29091), .B(n29090), .Z(n29109) );
  XNOR U30531 ( .A(n29110), .B(n29109), .Z(n29111) );
  NANDN U30532 ( .A(n29093), .B(n29092), .Z(n29097) );
  NAND U30533 ( .A(n29095), .B(n29094), .Z(n29096) );
  NAND U30534 ( .A(n29097), .B(n29096), .Z(n29112) );
  XNOR U30535 ( .A(n29111), .B(n29112), .Z(n29103) );
  XNOR U30536 ( .A(n29104), .B(n29103), .Z(n29105) );
  XNOR U30537 ( .A(n29106), .B(n29105), .Z(n29135) );
  XNOR U30538 ( .A(sreg[1692]), .B(n29135), .Z(n29137) );
  NANDN U30539 ( .A(sreg[1691]), .B(n29098), .Z(n29102) );
  NAND U30540 ( .A(n29100), .B(n29099), .Z(n29101) );
  NAND U30541 ( .A(n29102), .B(n29101), .Z(n29136) );
  XNOR U30542 ( .A(n29137), .B(n29136), .Z(c[1692]) );
  NANDN U30543 ( .A(n29104), .B(n29103), .Z(n29108) );
  NANDN U30544 ( .A(n29106), .B(n29105), .Z(n29107) );
  AND U30545 ( .A(n29108), .B(n29107), .Z(n29143) );
  NANDN U30546 ( .A(n29110), .B(n29109), .Z(n29114) );
  NANDN U30547 ( .A(n29112), .B(n29111), .Z(n29113) );
  AND U30548 ( .A(n29114), .B(n29113), .Z(n29141) );
  NAND U30549 ( .A(n42143), .B(n29115), .Z(n29117) );
  XNOR U30550 ( .A(a[671]), .B(n4167), .Z(n29152) );
  NAND U30551 ( .A(n42144), .B(n29152), .Z(n29116) );
  AND U30552 ( .A(n29117), .B(n29116), .Z(n29167) );
  XOR U30553 ( .A(a[675]), .B(n42012), .Z(n29155) );
  XNOR U30554 ( .A(n29167), .B(n29166), .Z(n29169) );
  AND U30555 ( .A(a[677]), .B(b[0]), .Z(n29119) );
  XNOR U30556 ( .A(n29119), .B(n4071), .Z(n29121) );
  NANDN U30557 ( .A(b[0]), .B(a[676]), .Z(n29120) );
  NAND U30558 ( .A(n29121), .B(n29120), .Z(n29163) );
  XOR U30559 ( .A(a[673]), .B(n42085), .Z(n29159) );
  AND U30560 ( .A(a[669]), .B(b[7]), .Z(n29160) );
  XNOR U30561 ( .A(n29161), .B(n29160), .Z(n29162) );
  XNOR U30562 ( .A(n29163), .B(n29162), .Z(n29168) );
  XOR U30563 ( .A(n29169), .B(n29168), .Z(n29147) );
  NANDN U30564 ( .A(n29124), .B(n29123), .Z(n29128) );
  NANDN U30565 ( .A(n29126), .B(n29125), .Z(n29127) );
  AND U30566 ( .A(n29128), .B(n29127), .Z(n29146) );
  XNOR U30567 ( .A(n29147), .B(n29146), .Z(n29148) );
  NANDN U30568 ( .A(n29130), .B(n29129), .Z(n29134) );
  NAND U30569 ( .A(n29132), .B(n29131), .Z(n29133) );
  NAND U30570 ( .A(n29134), .B(n29133), .Z(n29149) );
  XNOR U30571 ( .A(n29148), .B(n29149), .Z(n29140) );
  XNOR U30572 ( .A(n29141), .B(n29140), .Z(n29142) );
  XNOR U30573 ( .A(n29143), .B(n29142), .Z(n29172) );
  XNOR U30574 ( .A(sreg[1693]), .B(n29172), .Z(n29174) );
  NANDN U30575 ( .A(sreg[1692]), .B(n29135), .Z(n29139) );
  NAND U30576 ( .A(n29137), .B(n29136), .Z(n29138) );
  NAND U30577 ( .A(n29139), .B(n29138), .Z(n29173) );
  XNOR U30578 ( .A(n29174), .B(n29173), .Z(c[1693]) );
  NANDN U30579 ( .A(n29141), .B(n29140), .Z(n29145) );
  NANDN U30580 ( .A(n29143), .B(n29142), .Z(n29144) );
  AND U30581 ( .A(n29145), .B(n29144), .Z(n29180) );
  NANDN U30582 ( .A(n29147), .B(n29146), .Z(n29151) );
  NANDN U30583 ( .A(n29149), .B(n29148), .Z(n29150) );
  AND U30584 ( .A(n29151), .B(n29150), .Z(n29178) );
  NAND U30585 ( .A(n42143), .B(n29152), .Z(n29154) );
  XNOR U30586 ( .A(a[672]), .B(n4167), .Z(n29189) );
  NAND U30587 ( .A(n42144), .B(n29189), .Z(n29153) );
  AND U30588 ( .A(n29154), .B(n29153), .Z(n29204) );
  XOR U30589 ( .A(a[676]), .B(n42012), .Z(n29192) );
  XNOR U30590 ( .A(n29204), .B(n29203), .Z(n29206) );
  AND U30591 ( .A(a[678]), .B(b[0]), .Z(n29156) );
  XNOR U30592 ( .A(n29156), .B(n4071), .Z(n29158) );
  NANDN U30593 ( .A(b[0]), .B(a[677]), .Z(n29157) );
  NAND U30594 ( .A(n29158), .B(n29157), .Z(n29200) );
  XOR U30595 ( .A(a[674]), .B(n42085), .Z(n29196) );
  AND U30596 ( .A(a[670]), .B(b[7]), .Z(n29197) );
  XNOR U30597 ( .A(n29198), .B(n29197), .Z(n29199) );
  XNOR U30598 ( .A(n29200), .B(n29199), .Z(n29205) );
  XOR U30599 ( .A(n29206), .B(n29205), .Z(n29184) );
  NANDN U30600 ( .A(n29161), .B(n29160), .Z(n29165) );
  NANDN U30601 ( .A(n29163), .B(n29162), .Z(n29164) );
  AND U30602 ( .A(n29165), .B(n29164), .Z(n29183) );
  XNOR U30603 ( .A(n29184), .B(n29183), .Z(n29185) );
  NANDN U30604 ( .A(n29167), .B(n29166), .Z(n29171) );
  NAND U30605 ( .A(n29169), .B(n29168), .Z(n29170) );
  NAND U30606 ( .A(n29171), .B(n29170), .Z(n29186) );
  XNOR U30607 ( .A(n29185), .B(n29186), .Z(n29177) );
  XNOR U30608 ( .A(n29178), .B(n29177), .Z(n29179) );
  XNOR U30609 ( .A(n29180), .B(n29179), .Z(n29209) );
  XNOR U30610 ( .A(sreg[1694]), .B(n29209), .Z(n29211) );
  NANDN U30611 ( .A(sreg[1693]), .B(n29172), .Z(n29176) );
  NAND U30612 ( .A(n29174), .B(n29173), .Z(n29175) );
  NAND U30613 ( .A(n29176), .B(n29175), .Z(n29210) );
  XNOR U30614 ( .A(n29211), .B(n29210), .Z(c[1694]) );
  NANDN U30615 ( .A(n29178), .B(n29177), .Z(n29182) );
  NANDN U30616 ( .A(n29180), .B(n29179), .Z(n29181) );
  AND U30617 ( .A(n29182), .B(n29181), .Z(n29217) );
  NANDN U30618 ( .A(n29184), .B(n29183), .Z(n29188) );
  NANDN U30619 ( .A(n29186), .B(n29185), .Z(n29187) );
  AND U30620 ( .A(n29188), .B(n29187), .Z(n29215) );
  NAND U30621 ( .A(n42143), .B(n29189), .Z(n29191) );
  XNOR U30622 ( .A(a[673]), .B(n4168), .Z(n29226) );
  NAND U30623 ( .A(n42144), .B(n29226), .Z(n29190) );
  AND U30624 ( .A(n29191), .B(n29190), .Z(n29241) );
  XOR U30625 ( .A(a[677]), .B(n42012), .Z(n29229) );
  XNOR U30626 ( .A(n29241), .B(n29240), .Z(n29243) );
  AND U30627 ( .A(a[679]), .B(b[0]), .Z(n29193) );
  XNOR U30628 ( .A(n29193), .B(n4071), .Z(n29195) );
  NANDN U30629 ( .A(b[0]), .B(a[678]), .Z(n29194) );
  NAND U30630 ( .A(n29195), .B(n29194), .Z(n29237) );
  XOR U30631 ( .A(a[675]), .B(n42085), .Z(n29230) );
  AND U30632 ( .A(a[671]), .B(b[7]), .Z(n29234) );
  XNOR U30633 ( .A(n29235), .B(n29234), .Z(n29236) );
  XNOR U30634 ( .A(n29237), .B(n29236), .Z(n29242) );
  XOR U30635 ( .A(n29243), .B(n29242), .Z(n29221) );
  NANDN U30636 ( .A(n29198), .B(n29197), .Z(n29202) );
  NANDN U30637 ( .A(n29200), .B(n29199), .Z(n29201) );
  AND U30638 ( .A(n29202), .B(n29201), .Z(n29220) );
  XNOR U30639 ( .A(n29221), .B(n29220), .Z(n29222) );
  NANDN U30640 ( .A(n29204), .B(n29203), .Z(n29208) );
  NAND U30641 ( .A(n29206), .B(n29205), .Z(n29207) );
  NAND U30642 ( .A(n29208), .B(n29207), .Z(n29223) );
  XNOR U30643 ( .A(n29222), .B(n29223), .Z(n29214) );
  XNOR U30644 ( .A(n29215), .B(n29214), .Z(n29216) );
  XNOR U30645 ( .A(n29217), .B(n29216), .Z(n29246) );
  XNOR U30646 ( .A(sreg[1695]), .B(n29246), .Z(n29248) );
  NANDN U30647 ( .A(sreg[1694]), .B(n29209), .Z(n29213) );
  NAND U30648 ( .A(n29211), .B(n29210), .Z(n29212) );
  NAND U30649 ( .A(n29213), .B(n29212), .Z(n29247) );
  XNOR U30650 ( .A(n29248), .B(n29247), .Z(c[1695]) );
  NANDN U30651 ( .A(n29215), .B(n29214), .Z(n29219) );
  NANDN U30652 ( .A(n29217), .B(n29216), .Z(n29218) );
  AND U30653 ( .A(n29219), .B(n29218), .Z(n29254) );
  NANDN U30654 ( .A(n29221), .B(n29220), .Z(n29225) );
  NANDN U30655 ( .A(n29223), .B(n29222), .Z(n29224) );
  AND U30656 ( .A(n29225), .B(n29224), .Z(n29252) );
  NAND U30657 ( .A(n42143), .B(n29226), .Z(n29228) );
  XNOR U30658 ( .A(a[674]), .B(n4168), .Z(n29263) );
  NAND U30659 ( .A(n42144), .B(n29263), .Z(n29227) );
  AND U30660 ( .A(n29228), .B(n29227), .Z(n29278) );
  XOR U30661 ( .A(a[678]), .B(n42012), .Z(n29266) );
  XNOR U30662 ( .A(n29278), .B(n29277), .Z(n29280) );
  XOR U30663 ( .A(a[676]), .B(n42085), .Z(n29270) );
  AND U30664 ( .A(a[672]), .B(b[7]), .Z(n29271) );
  XNOR U30665 ( .A(n29272), .B(n29271), .Z(n29273) );
  AND U30666 ( .A(a[680]), .B(b[0]), .Z(n29231) );
  XNOR U30667 ( .A(n29231), .B(n4071), .Z(n29233) );
  NANDN U30668 ( .A(b[0]), .B(a[679]), .Z(n29232) );
  NAND U30669 ( .A(n29233), .B(n29232), .Z(n29274) );
  XNOR U30670 ( .A(n29273), .B(n29274), .Z(n29279) );
  XOR U30671 ( .A(n29280), .B(n29279), .Z(n29258) );
  NANDN U30672 ( .A(n29235), .B(n29234), .Z(n29239) );
  NANDN U30673 ( .A(n29237), .B(n29236), .Z(n29238) );
  AND U30674 ( .A(n29239), .B(n29238), .Z(n29257) );
  XNOR U30675 ( .A(n29258), .B(n29257), .Z(n29259) );
  NANDN U30676 ( .A(n29241), .B(n29240), .Z(n29245) );
  NAND U30677 ( .A(n29243), .B(n29242), .Z(n29244) );
  NAND U30678 ( .A(n29245), .B(n29244), .Z(n29260) );
  XNOR U30679 ( .A(n29259), .B(n29260), .Z(n29251) );
  XNOR U30680 ( .A(n29252), .B(n29251), .Z(n29253) );
  XNOR U30681 ( .A(n29254), .B(n29253), .Z(n29283) );
  XNOR U30682 ( .A(sreg[1696]), .B(n29283), .Z(n29285) );
  NANDN U30683 ( .A(sreg[1695]), .B(n29246), .Z(n29250) );
  NAND U30684 ( .A(n29248), .B(n29247), .Z(n29249) );
  NAND U30685 ( .A(n29250), .B(n29249), .Z(n29284) );
  XNOR U30686 ( .A(n29285), .B(n29284), .Z(c[1696]) );
  NANDN U30687 ( .A(n29252), .B(n29251), .Z(n29256) );
  NANDN U30688 ( .A(n29254), .B(n29253), .Z(n29255) );
  AND U30689 ( .A(n29256), .B(n29255), .Z(n29291) );
  NANDN U30690 ( .A(n29258), .B(n29257), .Z(n29262) );
  NANDN U30691 ( .A(n29260), .B(n29259), .Z(n29261) );
  AND U30692 ( .A(n29262), .B(n29261), .Z(n29289) );
  NAND U30693 ( .A(n42143), .B(n29263), .Z(n29265) );
  XNOR U30694 ( .A(a[675]), .B(n4168), .Z(n29300) );
  NAND U30695 ( .A(n42144), .B(n29300), .Z(n29264) );
  AND U30696 ( .A(n29265), .B(n29264), .Z(n29315) );
  XOR U30697 ( .A(a[679]), .B(n42012), .Z(n29303) );
  XNOR U30698 ( .A(n29315), .B(n29314), .Z(n29317) );
  AND U30699 ( .A(a[681]), .B(b[0]), .Z(n29267) );
  XNOR U30700 ( .A(n29267), .B(n4071), .Z(n29269) );
  NANDN U30701 ( .A(b[0]), .B(a[680]), .Z(n29268) );
  NAND U30702 ( .A(n29269), .B(n29268), .Z(n29311) );
  XOR U30703 ( .A(a[677]), .B(n42085), .Z(n29307) );
  AND U30704 ( .A(a[673]), .B(b[7]), .Z(n29308) );
  XNOR U30705 ( .A(n29309), .B(n29308), .Z(n29310) );
  XNOR U30706 ( .A(n29311), .B(n29310), .Z(n29316) );
  XOR U30707 ( .A(n29317), .B(n29316), .Z(n29295) );
  NANDN U30708 ( .A(n29272), .B(n29271), .Z(n29276) );
  NANDN U30709 ( .A(n29274), .B(n29273), .Z(n29275) );
  AND U30710 ( .A(n29276), .B(n29275), .Z(n29294) );
  XNOR U30711 ( .A(n29295), .B(n29294), .Z(n29296) );
  NANDN U30712 ( .A(n29278), .B(n29277), .Z(n29282) );
  NAND U30713 ( .A(n29280), .B(n29279), .Z(n29281) );
  NAND U30714 ( .A(n29282), .B(n29281), .Z(n29297) );
  XNOR U30715 ( .A(n29296), .B(n29297), .Z(n29288) );
  XNOR U30716 ( .A(n29289), .B(n29288), .Z(n29290) );
  XNOR U30717 ( .A(n29291), .B(n29290), .Z(n29320) );
  XNOR U30718 ( .A(sreg[1697]), .B(n29320), .Z(n29322) );
  NANDN U30719 ( .A(sreg[1696]), .B(n29283), .Z(n29287) );
  NAND U30720 ( .A(n29285), .B(n29284), .Z(n29286) );
  NAND U30721 ( .A(n29287), .B(n29286), .Z(n29321) );
  XNOR U30722 ( .A(n29322), .B(n29321), .Z(c[1697]) );
  NANDN U30723 ( .A(n29289), .B(n29288), .Z(n29293) );
  NANDN U30724 ( .A(n29291), .B(n29290), .Z(n29292) );
  AND U30725 ( .A(n29293), .B(n29292), .Z(n29328) );
  NANDN U30726 ( .A(n29295), .B(n29294), .Z(n29299) );
  NANDN U30727 ( .A(n29297), .B(n29296), .Z(n29298) );
  AND U30728 ( .A(n29299), .B(n29298), .Z(n29326) );
  NAND U30729 ( .A(n42143), .B(n29300), .Z(n29302) );
  XNOR U30730 ( .A(a[676]), .B(n4168), .Z(n29337) );
  NAND U30731 ( .A(n42144), .B(n29337), .Z(n29301) );
  AND U30732 ( .A(n29302), .B(n29301), .Z(n29352) );
  XOR U30733 ( .A(a[680]), .B(n42012), .Z(n29340) );
  XNOR U30734 ( .A(n29352), .B(n29351), .Z(n29354) );
  AND U30735 ( .A(a[682]), .B(b[0]), .Z(n29304) );
  XNOR U30736 ( .A(n29304), .B(n4071), .Z(n29306) );
  NANDN U30737 ( .A(b[0]), .B(a[681]), .Z(n29305) );
  NAND U30738 ( .A(n29306), .B(n29305), .Z(n29348) );
  XOR U30739 ( .A(a[678]), .B(n42085), .Z(n29344) );
  AND U30740 ( .A(a[674]), .B(b[7]), .Z(n29345) );
  XNOR U30741 ( .A(n29346), .B(n29345), .Z(n29347) );
  XNOR U30742 ( .A(n29348), .B(n29347), .Z(n29353) );
  XOR U30743 ( .A(n29354), .B(n29353), .Z(n29332) );
  NANDN U30744 ( .A(n29309), .B(n29308), .Z(n29313) );
  NANDN U30745 ( .A(n29311), .B(n29310), .Z(n29312) );
  AND U30746 ( .A(n29313), .B(n29312), .Z(n29331) );
  XNOR U30747 ( .A(n29332), .B(n29331), .Z(n29333) );
  NANDN U30748 ( .A(n29315), .B(n29314), .Z(n29319) );
  NAND U30749 ( .A(n29317), .B(n29316), .Z(n29318) );
  NAND U30750 ( .A(n29319), .B(n29318), .Z(n29334) );
  XNOR U30751 ( .A(n29333), .B(n29334), .Z(n29325) );
  XNOR U30752 ( .A(n29326), .B(n29325), .Z(n29327) );
  XNOR U30753 ( .A(n29328), .B(n29327), .Z(n29357) );
  XNOR U30754 ( .A(sreg[1698]), .B(n29357), .Z(n29359) );
  NANDN U30755 ( .A(sreg[1697]), .B(n29320), .Z(n29324) );
  NAND U30756 ( .A(n29322), .B(n29321), .Z(n29323) );
  NAND U30757 ( .A(n29324), .B(n29323), .Z(n29358) );
  XNOR U30758 ( .A(n29359), .B(n29358), .Z(c[1698]) );
  NANDN U30759 ( .A(n29326), .B(n29325), .Z(n29330) );
  NANDN U30760 ( .A(n29328), .B(n29327), .Z(n29329) );
  AND U30761 ( .A(n29330), .B(n29329), .Z(n29365) );
  NANDN U30762 ( .A(n29332), .B(n29331), .Z(n29336) );
  NANDN U30763 ( .A(n29334), .B(n29333), .Z(n29335) );
  AND U30764 ( .A(n29336), .B(n29335), .Z(n29363) );
  NAND U30765 ( .A(n42143), .B(n29337), .Z(n29339) );
  XNOR U30766 ( .A(a[677]), .B(n4168), .Z(n29374) );
  NAND U30767 ( .A(n42144), .B(n29374), .Z(n29338) );
  AND U30768 ( .A(n29339), .B(n29338), .Z(n29389) );
  XOR U30769 ( .A(a[681]), .B(n42012), .Z(n29377) );
  XNOR U30770 ( .A(n29389), .B(n29388), .Z(n29391) );
  AND U30771 ( .A(a[683]), .B(b[0]), .Z(n29341) );
  XNOR U30772 ( .A(n29341), .B(n4071), .Z(n29343) );
  NANDN U30773 ( .A(b[0]), .B(a[682]), .Z(n29342) );
  NAND U30774 ( .A(n29343), .B(n29342), .Z(n29385) );
  XOR U30775 ( .A(a[679]), .B(n42085), .Z(n29381) );
  AND U30776 ( .A(a[675]), .B(b[7]), .Z(n29382) );
  XNOR U30777 ( .A(n29383), .B(n29382), .Z(n29384) );
  XNOR U30778 ( .A(n29385), .B(n29384), .Z(n29390) );
  XOR U30779 ( .A(n29391), .B(n29390), .Z(n29369) );
  NANDN U30780 ( .A(n29346), .B(n29345), .Z(n29350) );
  NANDN U30781 ( .A(n29348), .B(n29347), .Z(n29349) );
  AND U30782 ( .A(n29350), .B(n29349), .Z(n29368) );
  XNOR U30783 ( .A(n29369), .B(n29368), .Z(n29370) );
  NANDN U30784 ( .A(n29352), .B(n29351), .Z(n29356) );
  NAND U30785 ( .A(n29354), .B(n29353), .Z(n29355) );
  NAND U30786 ( .A(n29356), .B(n29355), .Z(n29371) );
  XNOR U30787 ( .A(n29370), .B(n29371), .Z(n29362) );
  XNOR U30788 ( .A(n29363), .B(n29362), .Z(n29364) );
  XNOR U30789 ( .A(n29365), .B(n29364), .Z(n29394) );
  XNOR U30790 ( .A(sreg[1699]), .B(n29394), .Z(n29396) );
  NANDN U30791 ( .A(sreg[1698]), .B(n29357), .Z(n29361) );
  NAND U30792 ( .A(n29359), .B(n29358), .Z(n29360) );
  NAND U30793 ( .A(n29361), .B(n29360), .Z(n29395) );
  XNOR U30794 ( .A(n29396), .B(n29395), .Z(c[1699]) );
  NANDN U30795 ( .A(n29363), .B(n29362), .Z(n29367) );
  NANDN U30796 ( .A(n29365), .B(n29364), .Z(n29366) );
  AND U30797 ( .A(n29367), .B(n29366), .Z(n29402) );
  NANDN U30798 ( .A(n29369), .B(n29368), .Z(n29373) );
  NANDN U30799 ( .A(n29371), .B(n29370), .Z(n29372) );
  AND U30800 ( .A(n29373), .B(n29372), .Z(n29400) );
  NAND U30801 ( .A(n42143), .B(n29374), .Z(n29376) );
  XNOR U30802 ( .A(a[678]), .B(n4168), .Z(n29411) );
  NAND U30803 ( .A(n42144), .B(n29411), .Z(n29375) );
  AND U30804 ( .A(n29376), .B(n29375), .Z(n29426) );
  XOR U30805 ( .A(a[682]), .B(n42012), .Z(n29414) );
  XNOR U30806 ( .A(n29426), .B(n29425), .Z(n29428) );
  AND U30807 ( .A(b[0]), .B(a[684]), .Z(n29378) );
  XOR U30808 ( .A(b[1]), .B(n29378), .Z(n29380) );
  NANDN U30809 ( .A(b[0]), .B(a[683]), .Z(n29379) );
  AND U30810 ( .A(n29380), .B(n29379), .Z(n29421) );
  XOR U30811 ( .A(a[680]), .B(n42085), .Z(n29418) );
  AND U30812 ( .A(a[676]), .B(b[7]), .Z(n29419) );
  XOR U30813 ( .A(n29420), .B(n29419), .Z(n29422) );
  XNOR U30814 ( .A(n29421), .B(n29422), .Z(n29427) );
  XOR U30815 ( .A(n29428), .B(n29427), .Z(n29406) );
  NANDN U30816 ( .A(n29383), .B(n29382), .Z(n29387) );
  NANDN U30817 ( .A(n29385), .B(n29384), .Z(n29386) );
  AND U30818 ( .A(n29387), .B(n29386), .Z(n29405) );
  XNOR U30819 ( .A(n29406), .B(n29405), .Z(n29407) );
  NANDN U30820 ( .A(n29389), .B(n29388), .Z(n29393) );
  NAND U30821 ( .A(n29391), .B(n29390), .Z(n29392) );
  NAND U30822 ( .A(n29393), .B(n29392), .Z(n29408) );
  XNOR U30823 ( .A(n29407), .B(n29408), .Z(n29399) );
  XNOR U30824 ( .A(n29400), .B(n29399), .Z(n29401) );
  XNOR U30825 ( .A(n29402), .B(n29401), .Z(n29431) );
  XNOR U30826 ( .A(sreg[1700]), .B(n29431), .Z(n29433) );
  NANDN U30827 ( .A(sreg[1699]), .B(n29394), .Z(n29398) );
  NAND U30828 ( .A(n29396), .B(n29395), .Z(n29397) );
  NAND U30829 ( .A(n29398), .B(n29397), .Z(n29432) );
  XNOR U30830 ( .A(n29433), .B(n29432), .Z(c[1700]) );
  NANDN U30831 ( .A(n29400), .B(n29399), .Z(n29404) );
  NANDN U30832 ( .A(n29402), .B(n29401), .Z(n29403) );
  AND U30833 ( .A(n29404), .B(n29403), .Z(n29439) );
  NANDN U30834 ( .A(n29406), .B(n29405), .Z(n29410) );
  NANDN U30835 ( .A(n29408), .B(n29407), .Z(n29409) );
  AND U30836 ( .A(n29410), .B(n29409), .Z(n29437) );
  NAND U30837 ( .A(n42143), .B(n29411), .Z(n29413) );
  XNOR U30838 ( .A(a[679]), .B(n4168), .Z(n29448) );
  NAND U30839 ( .A(n42144), .B(n29448), .Z(n29412) );
  AND U30840 ( .A(n29413), .B(n29412), .Z(n29463) );
  XOR U30841 ( .A(a[683]), .B(n42012), .Z(n29451) );
  XNOR U30842 ( .A(n29463), .B(n29462), .Z(n29465) );
  AND U30843 ( .A(a[685]), .B(b[0]), .Z(n29415) );
  XNOR U30844 ( .A(n29415), .B(n4071), .Z(n29417) );
  NANDN U30845 ( .A(b[0]), .B(a[684]), .Z(n29416) );
  NAND U30846 ( .A(n29417), .B(n29416), .Z(n29459) );
  XOR U30847 ( .A(a[681]), .B(n42085), .Z(n29455) );
  AND U30848 ( .A(a[677]), .B(b[7]), .Z(n29456) );
  XNOR U30849 ( .A(n29457), .B(n29456), .Z(n29458) );
  XNOR U30850 ( .A(n29459), .B(n29458), .Z(n29464) );
  XOR U30851 ( .A(n29465), .B(n29464), .Z(n29443) );
  NANDN U30852 ( .A(n29420), .B(n29419), .Z(n29424) );
  NANDN U30853 ( .A(n29422), .B(n29421), .Z(n29423) );
  AND U30854 ( .A(n29424), .B(n29423), .Z(n29442) );
  XNOR U30855 ( .A(n29443), .B(n29442), .Z(n29444) );
  NANDN U30856 ( .A(n29426), .B(n29425), .Z(n29430) );
  NAND U30857 ( .A(n29428), .B(n29427), .Z(n29429) );
  NAND U30858 ( .A(n29430), .B(n29429), .Z(n29445) );
  XNOR U30859 ( .A(n29444), .B(n29445), .Z(n29436) );
  XNOR U30860 ( .A(n29437), .B(n29436), .Z(n29438) );
  XNOR U30861 ( .A(n29439), .B(n29438), .Z(n29468) );
  XNOR U30862 ( .A(sreg[1701]), .B(n29468), .Z(n29470) );
  NANDN U30863 ( .A(sreg[1700]), .B(n29431), .Z(n29435) );
  NAND U30864 ( .A(n29433), .B(n29432), .Z(n29434) );
  NAND U30865 ( .A(n29435), .B(n29434), .Z(n29469) );
  XNOR U30866 ( .A(n29470), .B(n29469), .Z(c[1701]) );
  NANDN U30867 ( .A(n29437), .B(n29436), .Z(n29441) );
  NANDN U30868 ( .A(n29439), .B(n29438), .Z(n29440) );
  AND U30869 ( .A(n29441), .B(n29440), .Z(n29476) );
  NANDN U30870 ( .A(n29443), .B(n29442), .Z(n29447) );
  NANDN U30871 ( .A(n29445), .B(n29444), .Z(n29446) );
  AND U30872 ( .A(n29447), .B(n29446), .Z(n29474) );
  NAND U30873 ( .A(n42143), .B(n29448), .Z(n29450) );
  XNOR U30874 ( .A(a[680]), .B(n4169), .Z(n29485) );
  NAND U30875 ( .A(n42144), .B(n29485), .Z(n29449) );
  AND U30876 ( .A(n29450), .B(n29449), .Z(n29500) );
  XOR U30877 ( .A(a[684]), .B(n42012), .Z(n29488) );
  XNOR U30878 ( .A(n29500), .B(n29499), .Z(n29502) );
  AND U30879 ( .A(a[686]), .B(b[0]), .Z(n29452) );
  XNOR U30880 ( .A(n29452), .B(n4071), .Z(n29454) );
  NANDN U30881 ( .A(b[0]), .B(a[685]), .Z(n29453) );
  NAND U30882 ( .A(n29454), .B(n29453), .Z(n29496) );
  XOR U30883 ( .A(a[682]), .B(n42085), .Z(n29489) );
  AND U30884 ( .A(a[678]), .B(b[7]), .Z(n29493) );
  XNOR U30885 ( .A(n29494), .B(n29493), .Z(n29495) );
  XNOR U30886 ( .A(n29496), .B(n29495), .Z(n29501) );
  XOR U30887 ( .A(n29502), .B(n29501), .Z(n29480) );
  NANDN U30888 ( .A(n29457), .B(n29456), .Z(n29461) );
  NANDN U30889 ( .A(n29459), .B(n29458), .Z(n29460) );
  AND U30890 ( .A(n29461), .B(n29460), .Z(n29479) );
  XNOR U30891 ( .A(n29480), .B(n29479), .Z(n29481) );
  NANDN U30892 ( .A(n29463), .B(n29462), .Z(n29467) );
  NAND U30893 ( .A(n29465), .B(n29464), .Z(n29466) );
  NAND U30894 ( .A(n29467), .B(n29466), .Z(n29482) );
  XNOR U30895 ( .A(n29481), .B(n29482), .Z(n29473) );
  XNOR U30896 ( .A(n29474), .B(n29473), .Z(n29475) );
  XNOR U30897 ( .A(n29476), .B(n29475), .Z(n29505) );
  XNOR U30898 ( .A(sreg[1702]), .B(n29505), .Z(n29507) );
  NANDN U30899 ( .A(sreg[1701]), .B(n29468), .Z(n29472) );
  NAND U30900 ( .A(n29470), .B(n29469), .Z(n29471) );
  NAND U30901 ( .A(n29472), .B(n29471), .Z(n29506) );
  XNOR U30902 ( .A(n29507), .B(n29506), .Z(c[1702]) );
  NANDN U30903 ( .A(n29474), .B(n29473), .Z(n29478) );
  NANDN U30904 ( .A(n29476), .B(n29475), .Z(n29477) );
  AND U30905 ( .A(n29478), .B(n29477), .Z(n29513) );
  NANDN U30906 ( .A(n29480), .B(n29479), .Z(n29484) );
  NANDN U30907 ( .A(n29482), .B(n29481), .Z(n29483) );
  AND U30908 ( .A(n29484), .B(n29483), .Z(n29511) );
  NAND U30909 ( .A(n42143), .B(n29485), .Z(n29487) );
  XNOR U30910 ( .A(a[681]), .B(n4169), .Z(n29522) );
  NAND U30911 ( .A(n42144), .B(n29522), .Z(n29486) );
  AND U30912 ( .A(n29487), .B(n29486), .Z(n29537) );
  XOR U30913 ( .A(a[685]), .B(n42012), .Z(n29525) );
  XNOR U30914 ( .A(n29537), .B(n29536), .Z(n29539) );
  XOR U30915 ( .A(a[683]), .B(n42085), .Z(n29526) );
  AND U30916 ( .A(a[679]), .B(b[7]), .Z(n29530) );
  XNOR U30917 ( .A(n29531), .B(n29530), .Z(n29532) );
  AND U30918 ( .A(a[687]), .B(b[0]), .Z(n29490) );
  XNOR U30919 ( .A(n29490), .B(n4071), .Z(n29492) );
  NANDN U30920 ( .A(b[0]), .B(a[686]), .Z(n29491) );
  NAND U30921 ( .A(n29492), .B(n29491), .Z(n29533) );
  XNOR U30922 ( .A(n29532), .B(n29533), .Z(n29538) );
  XOR U30923 ( .A(n29539), .B(n29538), .Z(n29517) );
  NANDN U30924 ( .A(n29494), .B(n29493), .Z(n29498) );
  NANDN U30925 ( .A(n29496), .B(n29495), .Z(n29497) );
  AND U30926 ( .A(n29498), .B(n29497), .Z(n29516) );
  XNOR U30927 ( .A(n29517), .B(n29516), .Z(n29518) );
  NANDN U30928 ( .A(n29500), .B(n29499), .Z(n29504) );
  NAND U30929 ( .A(n29502), .B(n29501), .Z(n29503) );
  NAND U30930 ( .A(n29504), .B(n29503), .Z(n29519) );
  XNOR U30931 ( .A(n29518), .B(n29519), .Z(n29510) );
  XNOR U30932 ( .A(n29511), .B(n29510), .Z(n29512) );
  XNOR U30933 ( .A(n29513), .B(n29512), .Z(n29542) );
  XNOR U30934 ( .A(sreg[1703]), .B(n29542), .Z(n29544) );
  NANDN U30935 ( .A(sreg[1702]), .B(n29505), .Z(n29509) );
  NAND U30936 ( .A(n29507), .B(n29506), .Z(n29508) );
  NAND U30937 ( .A(n29509), .B(n29508), .Z(n29543) );
  XNOR U30938 ( .A(n29544), .B(n29543), .Z(c[1703]) );
  NANDN U30939 ( .A(n29511), .B(n29510), .Z(n29515) );
  NANDN U30940 ( .A(n29513), .B(n29512), .Z(n29514) );
  AND U30941 ( .A(n29515), .B(n29514), .Z(n29550) );
  NANDN U30942 ( .A(n29517), .B(n29516), .Z(n29521) );
  NANDN U30943 ( .A(n29519), .B(n29518), .Z(n29520) );
  AND U30944 ( .A(n29521), .B(n29520), .Z(n29548) );
  NAND U30945 ( .A(n42143), .B(n29522), .Z(n29524) );
  XNOR U30946 ( .A(a[682]), .B(n4169), .Z(n29559) );
  NAND U30947 ( .A(n42144), .B(n29559), .Z(n29523) );
  AND U30948 ( .A(n29524), .B(n29523), .Z(n29575) );
  XOR U30949 ( .A(a[686]), .B(n42012), .Z(n29562) );
  XNOR U30950 ( .A(n29575), .B(n29574), .Z(n29577) );
  XOR U30951 ( .A(a[684]), .B(n42085), .Z(n29567) );
  AND U30952 ( .A(a[680]), .B(b[7]), .Z(n29568) );
  XNOR U30953 ( .A(n29569), .B(n29568), .Z(n29570) );
  AND U30954 ( .A(a[688]), .B(b[0]), .Z(n29527) );
  XNOR U30955 ( .A(n29527), .B(n4071), .Z(n29529) );
  NANDN U30956 ( .A(b[0]), .B(a[687]), .Z(n29528) );
  NAND U30957 ( .A(n29529), .B(n29528), .Z(n29571) );
  XNOR U30958 ( .A(n29570), .B(n29571), .Z(n29576) );
  XOR U30959 ( .A(n29577), .B(n29576), .Z(n29554) );
  NANDN U30960 ( .A(n29531), .B(n29530), .Z(n29535) );
  NANDN U30961 ( .A(n29533), .B(n29532), .Z(n29534) );
  AND U30962 ( .A(n29535), .B(n29534), .Z(n29553) );
  XNOR U30963 ( .A(n29554), .B(n29553), .Z(n29555) );
  NANDN U30964 ( .A(n29537), .B(n29536), .Z(n29541) );
  NAND U30965 ( .A(n29539), .B(n29538), .Z(n29540) );
  NAND U30966 ( .A(n29541), .B(n29540), .Z(n29556) );
  XNOR U30967 ( .A(n29555), .B(n29556), .Z(n29547) );
  XNOR U30968 ( .A(n29548), .B(n29547), .Z(n29549) );
  XNOR U30969 ( .A(n29550), .B(n29549), .Z(n29580) );
  XNOR U30970 ( .A(sreg[1704]), .B(n29580), .Z(n29582) );
  NANDN U30971 ( .A(sreg[1703]), .B(n29542), .Z(n29546) );
  NAND U30972 ( .A(n29544), .B(n29543), .Z(n29545) );
  NAND U30973 ( .A(n29546), .B(n29545), .Z(n29581) );
  XNOR U30974 ( .A(n29582), .B(n29581), .Z(c[1704]) );
  NANDN U30975 ( .A(n29548), .B(n29547), .Z(n29552) );
  NANDN U30976 ( .A(n29550), .B(n29549), .Z(n29551) );
  AND U30977 ( .A(n29552), .B(n29551), .Z(n29588) );
  NANDN U30978 ( .A(n29554), .B(n29553), .Z(n29558) );
  NANDN U30979 ( .A(n29556), .B(n29555), .Z(n29557) );
  AND U30980 ( .A(n29558), .B(n29557), .Z(n29586) );
  NAND U30981 ( .A(n42143), .B(n29559), .Z(n29561) );
  XNOR U30982 ( .A(a[683]), .B(n4169), .Z(n29597) );
  NAND U30983 ( .A(n42144), .B(n29597), .Z(n29560) );
  AND U30984 ( .A(n29561), .B(n29560), .Z(n29612) );
  XOR U30985 ( .A(a[687]), .B(n42012), .Z(n29600) );
  XNOR U30986 ( .A(n29612), .B(n29611), .Z(n29614) );
  AND U30987 ( .A(b[0]), .B(a[689]), .Z(n29563) );
  XOR U30988 ( .A(b[1]), .B(n29563), .Z(n29566) );
  NANDN U30989 ( .A(n29564), .B(a[688]), .Z(n29565) );
  AND U30990 ( .A(n29566), .B(n29565), .Z(n29607) );
  XOR U30991 ( .A(a[685]), .B(n42085), .Z(n29604) );
  AND U30992 ( .A(a[681]), .B(b[7]), .Z(n29605) );
  XOR U30993 ( .A(n29606), .B(n29605), .Z(n29608) );
  XNOR U30994 ( .A(n29607), .B(n29608), .Z(n29613) );
  XOR U30995 ( .A(n29614), .B(n29613), .Z(n29592) );
  NANDN U30996 ( .A(n29569), .B(n29568), .Z(n29573) );
  NANDN U30997 ( .A(n29571), .B(n29570), .Z(n29572) );
  AND U30998 ( .A(n29573), .B(n29572), .Z(n29591) );
  XNOR U30999 ( .A(n29592), .B(n29591), .Z(n29593) );
  NANDN U31000 ( .A(n29575), .B(n29574), .Z(n29579) );
  NAND U31001 ( .A(n29577), .B(n29576), .Z(n29578) );
  NAND U31002 ( .A(n29579), .B(n29578), .Z(n29594) );
  XNOR U31003 ( .A(n29593), .B(n29594), .Z(n29585) );
  XNOR U31004 ( .A(n29586), .B(n29585), .Z(n29587) );
  XNOR U31005 ( .A(n29588), .B(n29587), .Z(n29617) );
  XNOR U31006 ( .A(sreg[1705]), .B(n29617), .Z(n29619) );
  NANDN U31007 ( .A(sreg[1704]), .B(n29580), .Z(n29584) );
  NAND U31008 ( .A(n29582), .B(n29581), .Z(n29583) );
  NAND U31009 ( .A(n29584), .B(n29583), .Z(n29618) );
  XNOR U31010 ( .A(n29619), .B(n29618), .Z(c[1705]) );
  NANDN U31011 ( .A(n29586), .B(n29585), .Z(n29590) );
  NANDN U31012 ( .A(n29588), .B(n29587), .Z(n29589) );
  AND U31013 ( .A(n29590), .B(n29589), .Z(n29625) );
  NANDN U31014 ( .A(n29592), .B(n29591), .Z(n29596) );
  NANDN U31015 ( .A(n29594), .B(n29593), .Z(n29595) );
  AND U31016 ( .A(n29596), .B(n29595), .Z(n29623) );
  NAND U31017 ( .A(n42143), .B(n29597), .Z(n29599) );
  XNOR U31018 ( .A(a[684]), .B(n4169), .Z(n29634) );
  NAND U31019 ( .A(n42144), .B(n29634), .Z(n29598) );
  AND U31020 ( .A(n29599), .B(n29598), .Z(n29649) );
  XOR U31021 ( .A(a[688]), .B(n42012), .Z(n29637) );
  XNOR U31022 ( .A(n29649), .B(n29648), .Z(n29651) );
  AND U31023 ( .A(a[690]), .B(b[0]), .Z(n29601) );
  XNOR U31024 ( .A(n29601), .B(n4071), .Z(n29603) );
  NANDN U31025 ( .A(b[0]), .B(a[689]), .Z(n29602) );
  NAND U31026 ( .A(n29603), .B(n29602), .Z(n29645) );
  XOR U31027 ( .A(a[686]), .B(n42085), .Z(n29641) );
  AND U31028 ( .A(a[682]), .B(b[7]), .Z(n29642) );
  XNOR U31029 ( .A(n29643), .B(n29642), .Z(n29644) );
  XNOR U31030 ( .A(n29645), .B(n29644), .Z(n29650) );
  XOR U31031 ( .A(n29651), .B(n29650), .Z(n29629) );
  NANDN U31032 ( .A(n29606), .B(n29605), .Z(n29610) );
  NANDN U31033 ( .A(n29608), .B(n29607), .Z(n29609) );
  AND U31034 ( .A(n29610), .B(n29609), .Z(n29628) );
  XNOR U31035 ( .A(n29629), .B(n29628), .Z(n29630) );
  NANDN U31036 ( .A(n29612), .B(n29611), .Z(n29616) );
  NAND U31037 ( .A(n29614), .B(n29613), .Z(n29615) );
  NAND U31038 ( .A(n29616), .B(n29615), .Z(n29631) );
  XNOR U31039 ( .A(n29630), .B(n29631), .Z(n29622) );
  XNOR U31040 ( .A(n29623), .B(n29622), .Z(n29624) );
  XNOR U31041 ( .A(n29625), .B(n29624), .Z(n29654) );
  XNOR U31042 ( .A(sreg[1706]), .B(n29654), .Z(n29656) );
  NANDN U31043 ( .A(sreg[1705]), .B(n29617), .Z(n29621) );
  NAND U31044 ( .A(n29619), .B(n29618), .Z(n29620) );
  NAND U31045 ( .A(n29621), .B(n29620), .Z(n29655) );
  XNOR U31046 ( .A(n29656), .B(n29655), .Z(c[1706]) );
  NANDN U31047 ( .A(n29623), .B(n29622), .Z(n29627) );
  NANDN U31048 ( .A(n29625), .B(n29624), .Z(n29626) );
  AND U31049 ( .A(n29627), .B(n29626), .Z(n29662) );
  NANDN U31050 ( .A(n29629), .B(n29628), .Z(n29633) );
  NANDN U31051 ( .A(n29631), .B(n29630), .Z(n29632) );
  AND U31052 ( .A(n29633), .B(n29632), .Z(n29660) );
  NAND U31053 ( .A(n42143), .B(n29634), .Z(n29636) );
  XNOR U31054 ( .A(a[685]), .B(n4169), .Z(n29671) );
  NAND U31055 ( .A(n42144), .B(n29671), .Z(n29635) );
  AND U31056 ( .A(n29636), .B(n29635), .Z(n29686) );
  XOR U31057 ( .A(a[689]), .B(n42012), .Z(n29674) );
  XNOR U31058 ( .A(n29686), .B(n29685), .Z(n29688) );
  AND U31059 ( .A(a[691]), .B(b[0]), .Z(n29638) );
  XNOR U31060 ( .A(n29638), .B(n4071), .Z(n29640) );
  NANDN U31061 ( .A(b[0]), .B(a[690]), .Z(n29639) );
  NAND U31062 ( .A(n29640), .B(n29639), .Z(n29682) );
  XOR U31063 ( .A(a[687]), .B(n42085), .Z(n29678) );
  AND U31064 ( .A(a[683]), .B(b[7]), .Z(n29679) );
  XNOR U31065 ( .A(n29680), .B(n29679), .Z(n29681) );
  XNOR U31066 ( .A(n29682), .B(n29681), .Z(n29687) );
  XOR U31067 ( .A(n29688), .B(n29687), .Z(n29666) );
  NANDN U31068 ( .A(n29643), .B(n29642), .Z(n29647) );
  NANDN U31069 ( .A(n29645), .B(n29644), .Z(n29646) );
  AND U31070 ( .A(n29647), .B(n29646), .Z(n29665) );
  XNOR U31071 ( .A(n29666), .B(n29665), .Z(n29667) );
  NANDN U31072 ( .A(n29649), .B(n29648), .Z(n29653) );
  NAND U31073 ( .A(n29651), .B(n29650), .Z(n29652) );
  NAND U31074 ( .A(n29653), .B(n29652), .Z(n29668) );
  XNOR U31075 ( .A(n29667), .B(n29668), .Z(n29659) );
  XNOR U31076 ( .A(n29660), .B(n29659), .Z(n29661) );
  XNOR U31077 ( .A(n29662), .B(n29661), .Z(n29691) );
  XNOR U31078 ( .A(sreg[1707]), .B(n29691), .Z(n29693) );
  NANDN U31079 ( .A(sreg[1706]), .B(n29654), .Z(n29658) );
  NAND U31080 ( .A(n29656), .B(n29655), .Z(n29657) );
  NAND U31081 ( .A(n29658), .B(n29657), .Z(n29692) );
  XNOR U31082 ( .A(n29693), .B(n29692), .Z(c[1707]) );
  NANDN U31083 ( .A(n29660), .B(n29659), .Z(n29664) );
  NANDN U31084 ( .A(n29662), .B(n29661), .Z(n29663) );
  AND U31085 ( .A(n29664), .B(n29663), .Z(n29699) );
  NANDN U31086 ( .A(n29666), .B(n29665), .Z(n29670) );
  NANDN U31087 ( .A(n29668), .B(n29667), .Z(n29669) );
  AND U31088 ( .A(n29670), .B(n29669), .Z(n29697) );
  NAND U31089 ( .A(n42143), .B(n29671), .Z(n29673) );
  XNOR U31090 ( .A(a[686]), .B(n4169), .Z(n29708) );
  NAND U31091 ( .A(n42144), .B(n29708), .Z(n29672) );
  AND U31092 ( .A(n29673), .B(n29672), .Z(n29723) );
  XOR U31093 ( .A(a[690]), .B(n42012), .Z(n29711) );
  XNOR U31094 ( .A(n29723), .B(n29722), .Z(n29725) );
  AND U31095 ( .A(a[692]), .B(b[0]), .Z(n29675) );
  XNOR U31096 ( .A(n29675), .B(n4071), .Z(n29677) );
  NANDN U31097 ( .A(b[0]), .B(a[691]), .Z(n29676) );
  NAND U31098 ( .A(n29677), .B(n29676), .Z(n29719) );
  XOR U31099 ( .A(a[688]), .B(n42085), .Z(n29712) );
  AND U31100 ( .A(a[684]), .B(b[7]), .Z(n29716) );
  XNOR U31101 ( .A(n29717), .B(n29716), .Z(n29718) );
  XNOR U31102 ( .A(n29719), .B(n29718), .Z(n29724) );
  XOR U31103 ( .A(n29725), .B(n29724), .Z(n29703) );
  NANDN U31104 ( .A(n29680), .B(n29679), .Z(n29684) );
  NANDN U31105 ( .A(n29682), .B(n29681), .Z(n29683) );
  AND U31106 ( .A(n29684), .B(n29683), .Z(n29702) );
  XNOR U31107 ( .A(n29703), .B(n29702), .Z(n29704) );
  NANDN U31108 ( .A(n29686), .B(n29685), .Z(n29690) );
  NAND U31109 ( .A(n29688), .B(n29687), .Z(n29689) );
  NAND U31110 ( .A(n29690), .B(n29689), .Z(n29705) );
  XNOR U31111 ( .A(n29704), .B(n29705), .Z(n29696) );
  XNOR U31112 ( .A(n29697), .B(n29696), .Z(n29698) );
  XNOR U31113 ( .A(n29699), .B(n29698), .Z(n29728) );
  XNOR U31114 ( .A(sreg[1708]), .B(n29728), .Z(n29730) );
  NANDN U31115 ( .A(sreg[1707]), .B(n29691), .Z(n29695) );
  NAND U31116 ( .A(n29693), .B(n29692), .Z(n29694) );
  NAND U31117 ( .A(n29695), .B(n29694), .Z(n29729) );
  XNOR U31118 ( .A(n29730), .B(n29729), .Z(c[1708]) );
  NANDN U31119 ( .A(n29697), .B(n29696), .Z(n29701) );
  NANDN U31120 ( .A(n29699), .B(n29698), .Z(n29700) );
  AND U31121 ( .A(n29701), .B(n29700), .Z(n29736) );
  NANDN U31122 ( .A(n29703), .B(n29702), .Z(n29707) );
  NANDN U31123 ( .A(n29705), .B(n29704), .Z(n29706) );
  AND U31124 ( .A(n29707), .B(n29706), .Z(n29734) );
  NAND U31125 ( .A(n42143), .B(n29708), .Z(n29710) );
  XNOR U31126 ( .A(a[687]), .B(n4170), .Z(n29745) );
  NAND U31127 ( .A(n42144), .B(n29745), .Z(n29709) );
  AND U31128 ( .A(n29710), .B(n29709), .Z(n29760) );
  XOR U31129 ( .A(a[691]), .B(n42012), .Z(n29748) );
  XNOR U31130 ( .A(n29760), .B(n29759), .Z(n29762) );
  XOR U31131 ( .A(a[689]), .B(n42085), .Z(n29752) );
  AND U31132 ( .A(a[685]), .B(b[7]), .Z(n29753) );
  XNOR U31133 ( .A(n29754), .B(n29753), .Z(n29755) );
  AND U31134 ( .A(a[693]), .B(b[0]), .Z(n29713) );
  XNOR U31135 ( .A(n29713), .B(n4071), .Z(n29715) );
  NANDN U31136 ( .A(b[0]), .B(a[692]), .Z(n29714) );
  NAND U31137 ( .A(n29715), .B(n29714), .Z(n29756) );
  XNOR U31138 ( .A(n29755), .B(n29756), .Z(n29761) );
  XOR U31139 ( .A(n29762), .B(n29761), .Z(n29740) );
  NANDN U31140 ( .A(n29717), .B(n29716), .Z(n29721) );
  NANDN U31141 ( .A(n29719), .B(n29718), .Z(n29720) );
  AND U31142 ( .A(n29721), .B(n29720), .Z(n29739) );
  XNOR U31143 ( .A(n29740), .B(n29739), .Z(n29741) );
  NANDN U31144 ( .A(n29723), .B(n29722), .Z(n29727) );
  NAND U31145 ( .A(n29725), .B(n29724), .Z(n29726) );
  NAND U31146 ( .A(n29727), .B(n29726), .Z(n29742) );
  XNOR U31147 ( .A(n29741), .B(n29742), .Z(n29733) );
  XNOR U31148 ( .A(n29734), .B(n29733), .Z(n29735) );
  XNOR U31149 ( .A(n29736), .B(n29735), .Z(n29765) );
  XNOR U31150 ( .A(sreg[1709]), .B(n29765), .Z(n29767) );
  NANDN U31151 ( .A(sreg[1708]), .B(n29728), .Z(n29732) );
  NAND U31152 ( .A(n29730), .B(n29729), .Z(n29731) );
  NAND U31153 ( .A(n29732), .B(n29731), .Z(n29766) );
  XNOR U31154 ( .A(n29767), .B(n29766), .Z(c[1709]) );
  NANDN U31155 ( .A(n29734), .B(n29733), .Z(n29738) );
  NANDN U31156 ( .A(n29736), .B(n29735), .Z(n29737) );
  AND U31157 ( .A(n29738), .B(n29737), .Z(n29773) );
  NANDN U31158 ( .A(n29740), .B(n29739), .Z(n29744) );
  NANDN U31159 ( .A(n29742), .B(n29741), .Z(n29743) );
  AND U31160 ( .A(n29744), .B(n29743), .Z(n29771) );
  NAND U31161 ( .A(n42143), .B(n29745), .Z(n29747) );
  XNOR U31162 ( .A(a[688]), .B(n4170), .Z(n29782) );
  NAND U31163 ( .A(n42144), .B(n29782), .Z(n29746) );
  AND U31164 ( .A(n29747), .B(n29746), .Z(n29797) );
  XOR U31165 ( .A(a[692]), .B(n42012), .Z(n29785) );
  XNOR U31166 ( .A(n29797), .B(n29796), .Z(n29799) );
  AND U31167 ( .A(a[694]), .B(b[0]), .Z(n29749) );
  XNOR U31168 ( .A(n29749), .B(n4071), .Z(n29751) );
  NANDN U31169 ( .A(b[0]), .B(a[693]), .Z(n29750) );
  NAND U31170 ( .A(n29751), .B(n29750), .Z(n29793) );
  XOR U31171 ( .A(a[690]), .B(n42085), .Z(n29786) );
  AND U31172 ( .A(a[686]), .B(b[7]), .Z(n29790) );
  XNOR U31173 ( .A(n29791), .B(n29790), .Z(n29792) );
  XNOR U31174 ( .A(n29793), .B(n29792), .Z(n29798) );
  XOR U31175 ( .A(n29799), .B(n29798), .Z(n29777) );
  NANDN U31176 ( .A(n29754), .B(n29753), .Z(n29758) );
  NANDN U31177 ( .A(n29756), .B(n29755), .Z(n29757) );
  AND U31178 ( .A(n29758), .B(n29757), .Z(n29776) );
  XNOR U31179 ( .A(n29777), .B(n29776), .Z(n29778) );
  NANDN U31180 ( .A(n29760), .B(n29759), .Z(n29764) );
  NAND U31181 ( .A(n29762), .B(n29761), .Z(n29763) );
  NAND U31182 ( .A(n29764), .B(n29763), .Z(n29779) );
  XNOR U31183 ( .A(n29778), .B(n29779), .Z(n29770) );
  XNOR U31184 ( .A(n29771), .B(n29770), .Z(n29772) );
  XNOR U31185 ( .A(n29773), .B(n29772), .Z(n29802) );
  XNOR U31186 ( .A(sreg[1710]), .B(n29802), .Z(n29804) );
  NANDN U31187 ( .A(sreg[1709]), .B(n29765), .Z(n29769) );
  NAND U31188 ( .A(n29767), .B(n29766), .Z(n29768) );
  NAND U31189 ( .A(n29769), .B(n29768), .Z(n29803) );
  XNOR U31190 ( .A(n29804), .B(n29803), .Z(c[1710]) );
  NANDN U31191 ( .A(n29771), .B(n29770), .Z(n29775) );
  NANDN U31192 ( .A(n29773), .B(n29772), .Z(n29774) );
  AND U31193 ( .A(n29775), .B(n29774), .Z(n29810) );
  NANDN U31194 ( .A(n29777), .B(n29776), .Z(n29781) );
  NANDN U31195 ( .A(n29779), .B(n29778), .Z(n29780) );
  AND U31196 ( .A(n29781), .B(n29780), .Z(n29808) );
  NAND U31197 ( .A(n42143), .B(n29782), .Z(n29784) );
  XNOR U31198 ( .A(a[689]), .B(n4170), .Z(n29819) );
  NAND U31199 ( .A(n42144), .B(n29819), .Z(n29783) );
  AND U31200 ( .A(n29784), .B(n29783), .Z(n29834) );
  XOR U31201 ( .A(a[693]), .B(n42012), .Z(n29822) );
  XNOR U31202 ( .A(n29834), .B(n29833), .Z(n29836) );
  XOR U31203 ( .A(a[691]), .B(n42085), .Z(n29826) );
  AND U31204 ( .A(a[687]), .B(b[7]), .Z(n29827) );
  XNOR U31205 ( .A(n29828), .B(n29827), .Z(n29829) );
  AND U31206 ( .A(a[695]), .B(b[0]), .Z(n29787) );
  XNOR U31207 ( .A(n29787), .B(n4071), .Z(n29789) );
  NANDN U31208 ( .A(b[0]), .B(a[694]), .Z(n29788) );
  NAND U31209 ( .A(n29789), .B(n29788), .Z(n29830) );
  XNOR U31210 ( .A(n29829), .B(n29830), .Z(n29835) );
  XOR U31211 ( .A(n29836), .B(n29835), .Z(n29814) );
  NANDN U31212 ( .A(n29791), .B(n29790), .Z(n29795) );
  NANDN U31213 ( .A(n29793), .B(n29792), .Z(n29794) );
  AND U31214 ( .A(n29795), .B(n29794), .Z(n29813) );
  XNOR U31215 ( .A(n29814), .B(n29813), .Z(n29815) );
  NANDN U31216 ( .A(n29797), .B(n29796), .Z(n29801) );
  NAND U31217 ( .A(n29799), .B(n29798), .Z(n29800) );
  NAND U31218 ( .A(n29801), .B(n29800), .Z(n29816) );
  XNOR U31219 ( .A(n29815), .B(n29816), .Z(n29807) );
  XNOR U31220 ( .A(n29808), .B(n29807), .Z(n29809) );
  XNOR U31221 ( .A(n29810), .B(n29809), .Z(n29839) );
  XNOR U31222 ( .A(sreg[1711]), .B(n29839), .Z(n29841) );
  NANDN U31223 ( .A(sreg[1710]), .B(n29802), .Z(n29806) );
  NAND U31224 ( .A(n29804), .B(n29803), .Z(n29805) );
  NAND U31225 ( .A(n29806), .B(n29805), .Z(n29840) );
  XNOR U31226 ( .A(n29841), .B(n29840), .Z(c[1711]) );
  NANDN U31227 ( .A(n29808), .B(n29807), .Z(n29812) );
  NANDN U31228 ( .A(n29810), .B(n29809), .Z(n29811) );
  AND U31229 ( .A(n29812), .B(n29811), .Z(n29847) );
  NANDN U31230 ( .A(n29814), .B(n29813), .Z(n29818) );
  NANDN U31231 ( .A(n29816), .B(n29815), .Z(n29817) );
  AND U31232 ( .A(n29818), .B(n29817), .Z(n29845) );
  NAND U31233 ( .A(n42143), .B(n29819), .Z(n29821) );
  XNOR U31234 ( .A(a[690]), .B(n4170), .Z(n29856) );
  NAND U31235 ( .A(n42144), .B(n29856), .Z(n29820) );
  AND U31236 ( .A(n29821), .B(n29820), .Z(n29871) );
  XOR U31237 ( .A(a[694]), .B(n42012), .Z(n29859) );
  XNOR U31238 ( .A(n29871), .B(n29870), .Z(n29873) );
  AND U31239 ( .A(a[696]), .B(b[0]), .Z(n29823) );
  XNOR U31240 ( .A(n29823), .B(n4071), .Z(n29825) );
  NANDN U31241 ( .A(b[0]), .B(a[695]), .Z(n29824) );
  NAND U31242 ( .A(n29825), .B(n29824), .Z(n29867) );
  XOR U31243 ( .A(a[692]), .B(n42085), .Z(n29863) );
  AND U31244 ( .A(a[688]), .B(b[7]), .Z(n29864) );
  XNOR U31245 ( .A(n29865), .B(n29864), .Z(n29866) );
  XNOR U31246 ( .A(n29867), .B(n29866), .Z(n29872) );
  XOR U31247 ( .A(n29873), .B(n29872), .Z(n29851) );
  NANDN U31248 ( .A(n29828), .B(n29827), .Z(n29832) );
  NANDN U31249 ( .A(n29830), .B(n29829), .Z(n29831) );
  AND U31250 ( .A(n29832), .B(n29831), .Z(n29850) );
  XNOR U31251 ( .A(n29851), .B(n29850), .Z(n29852) );
  NANDN U31252 ( .A(n29834), .B(n29833), .Z(n29838) );
  NAND U31253 ( .A(n29836), .B(n29835), .Z(n29837) );
  NAND U31254 ( .A(n29838), .B(n29837), .Z(n29853) );
  XNOR U31255 ( .A(n29852), .B(n29853), .Z(n29844) );
  XNOR U31256 ( .A(n29845), .B(n29844), .Z(n29846) );
  XNOR U31257 ( .A(n29847), .B(n29846), .Z(n29876) );
  XNOR U31258 ( .A(sreg[1712]), .B(n29876), .Z(n29878) );
  NANDN U31259 ( .A(sreg[1711]), .B(n29839), .Z(n29843) );
  NAND U31260 ( .A(n29841), .B(n29840), .Z(n29842) );
  NAND U31261 ( .A(n29843), .B(n29842), .Z(n29877) );
  XNOR U31262 ( .A(n29878), .B(n29877), .Z(c[1712]) );
  NANDN U31263 ( .A(n29845), .B(n29844), .Z(n29849) );
  NANDN U31264 ( .A(n29847), .B(n29846), .Z(n29848) );
  AND U31265 ( .A(n29849), .B(n29848), .Z(n29884) );
  NANDN U31266 ( .A(n29851), .B(n29850), .Z(n29855) );
  NANDN U31267 ( .A(n29853), .B(n29852), .Z(n29854) );
  AND U31268 ( .A(n29855), .B(n29854), .Z(n29882) );
  NAND U31269 ( .A(n42143), .B(n29856), .Z(n29858) );
  XNOR U31270 ( .A(a[691]), .B(n4170), .Z(n29893) );
  NAND U31271 ( .A(n42144), .B(n29893), .Z(n29857) );
  AND U31272 ( .A(n29858), .B(n29857), .Z(n29908) );
  XOR U31273 ( .A(a[695]), .B(n42012), .Z(n29896) );
  XNOR U31274 ( .A(n29908), .B(n29907), .Z(n29910) );
  AND U31275 ( .A(a[697]), .B(b[0]), .Z(n29860) );
  XNOR U31276 ( .A(n29860), .B(n4071), .Z(n29862) );
  NANDN U31277 ( .A(b[0]), .B(a[696]), .Z(n29861) );
  NAND U31278 ( .A(n29862), .B(n29861), .Z(n29904) );
  XOR U31279 ( .A(a[693]), .B(n42085), .Z(n29897) );
  AND U31280 ( .A(a[689]), .B(b[7]), .Z(n29901) );
  XNOR U31281 ( .A(n29902), .B(n29901), .Z(n29903) );
  XNOR U31282 ( .A(n29904), .B(n29903), .Z(n29909) );
  XOR U31283 ( .A(n29910), .B(n29909), .Z(n29888) );
  NANDN U31284 ( .A(n29865), .B(n29864), .Z(n29869) );
  NANDN U31285 ( .A(n29867), .B(n29866), .Z(n29868) );
  AND U31286 ( .A(n29869), .B(n29868), .Z(n29887) );
  XNOR U31287 ( .A(n29888), .B(n29887), .Z(n29889) );
  NANDN U31288 ( .A(n29871), .B(n29870), .Z(n29875) );
  NAND U31289 ( .A(n29873), .B(n29872), .Z(n29874) );
  NAND U31290 ( .A(n29875), .B(n29874), .Z(n29890) );
  XNOR U31291 ( .A(n29889), .B(n29890), .Z(n29881) );
  XNOR U31292 ( .A(n29882), .B(n29881), .Z(n29883) );
  XNOR U31293 ( .A(n29884), .B(n29883), .Z(n29913) );
  XNOR U31294 ( .A(sreg[1713]), .B(n29913), .Z(n29915) );
  NANDN U31295 ( .A(sreg[1712]), .B(n29876), .Z(n29880) );
  NAND U31296 ( .A(n29878), .B(n29877), .Z(n29879) );
  NAND U31297 ( .A(n29880), .B(n29879), .Z(n29914) );
  XNOR U31298 ( .A(n29915), .B(n29914), .Z(c[1713]) );
  NANDN U31299 ( .A(n29882), .B(n29881), .Z(n29886) );
  NANDN U31300 ( .A(n29884), .B(n29883), .Z(n29885) );
  AND U31301 ( .A(n29886), .B(n29885), .Z(n29921) );
  NANDN U31302 ( .A(n29888), .B(n29887), .Z(n29892) );
  NANDN U31303 ( .A(n29890), .B(n29889), .Z(n29891) );
  AND U31304 ( .A(n29892), .B(n29891), .Z(n29919) );
  NAND U31305 ( .A(n42143), .B(n29893), .Z(n29895) );
  XNOR U31306 ( .A(a[692]), .B(n4170), .Z(n29930) );
  NAND U31307 ( .A(n42144), .B(n29930), .Z(n29894) );
  AND U31308 ( .A(n29895), .B(n29894), .Z(n29945) );
  XOR U31309 ( .A(a[696]), .B(n42012), .Z(n29933) );
  XNOR U31310 ( .A(n29945), .B(n29944), .Z(n29947) );
  XOR U31311 ( .A(a[694]), .B(n42085), .Z(n29934) );
  AND U31312 ( .A(a[690]), .B(b[7]), .Z(n29938) );
  XNOR U31313 ( .A(n29939), .B(n29938), .Z(n29940) );
  AND U31314 ( .A(a[698]), .B(b[0]), .Z(n29898) );
  XNOR U31315 ( .A(n29898), .B(n4071), .Z(n29900) );
  NANDN U31316 ( .A(b[0]), .B(a[697]), .Z(n29899) );
  NAND U31317 ( .A(n29900), .B(n29899), .Z(n29941) );
  XNOR U31318 ( .A(n29940), .B(n29941), .Z(n29946) );
  XOR U31319 ( .A(n29947), .B(n29946), .Z(n29925) );
  NANDN U31320 ( .A(n29902), .B(n29901), .Z(n29906) );
  NANDN U31321 ( .A(n29904), .B(n29903), .Z(n29905) );
  AND U31322 ( .A(n29906), .B(n29905), .Z(n29924) );
  XNOR U31323 ( .A(n29925), .B(n29924), .Z(n29926) );
  NANDN U31324 ( .A(n29908), .B(n29907), .Z(n29912) );
  NAND U31325 ( .A(n29910), .B(n29909), .Z(n29911) );
  NAND U31326 ( .A(n29912), .B(n29911), .Z(n29927) );
  XNOR U31327 ( .A(n29926), .B(n29927), .Z(n29918) );
  XNOR U31328 ( .A(n29919), .B(n29918), .Z(n29920) );
  XNOR U31329 ( .A(n29921), .B(n29920), .Z(n29950) );
  XNOR U31330 ( .A(sreg[1714]), .B(n29950), .Z(n29952) );
  NANDN U31331 ( .A(sreg[1713]), .B(n29913), .Z(n29917) );
  NAND U31332 ( .A(n29915), .B(n29914), .Z(n29916) );
  NAND U31333 ( .A(n29917), .B(n29916), .Z(n29951) );
  XNOR U31334 ( .A(n29952), .B(n29951), .Z(c[1714]) );
  NANDN U31335 ( .A(n29919), .B(n29918), .Z(n29923) );
  NANDN U31336 ( .A(n29921), .B(n29920), .Z(n29922) );
  AND U31337 ( .A(n29923), .B(n29922), .Z(n29958) );
  NANDN U31338 ( .A(n29925), .B(n29924), .Z(n29929) );
  NANDN U31339 ( .A(n29927), .B(n29926), .Z(n29928) );
  AND U31340 ( .A(n29929), .B(n29928), .Z(n29956) );
  NAND U31341 ( .A(n42143), .B(n29930), .Z(n29932) );
  XNOR U31342 ( .A(a[693]), .B(n4170), .Z(n29967) );
  NAND U31343 ( .A(n42144), .B(n29967), .Z(n29931) );
  AND U31344 ( .A(n29932), .B(n29931), .Z(n29982) );
  XOR U31345 ( .A(a[697]), .B(n42012), .Z(n29970) );
  XNOR U31346 ( .A(n29982), .B(n29981), .Z(n29984) );
  XOR U31347 ( .A(a[695]), .B(n42085), .Z(n29974) );
  AND U31348 ( .A(a[691]), .B(b[7]), .Z(n29975) );
  XNOR U31349 ( .A(n29976), .B(n29975), .Z(n29977) );
  AND U31350 ( .A(a[699]), .B(b[0]), .Z(n29935) );
  XNOR U31351 ( .A(n29935), .B(n4071), .Z(n29937) );
  NANDN U31352 ( .A(b[0]), .B(a[698]), .Z(n29936) );
  NAND U31353 ( .A(n29937), .B(n29936), .Z(n29978) );
  XNOR U31354 ( .A(n29977), .B(n29978), .Z(n29983) );
  XOR U31355 ( .A(n29984), .B(n29983), .Z(n29962) );
  NANDN U31356 ( .A(n29939), .B(n29938), .Z(n29943) );
  NANDN U31357 ( .A(n29941), .B(n29940), .Z(n29942) );
  AND U31358 ( .A(n29943), .B(n29942), .Z(n29961) );
  XNOR U31359 ( .A(n29962), .B(n29961), .Z(n29963) );
  NANDN U31360 ( .A(n29945), .B(n29944), .Z(n29949) );
  NAND U31361 ( .A(n29947), .B(n29946), .Z(n29948) );
  NAND U31362 ( .A(n29949), .B(n29948), .Z(n29964) );
  XNOR U31363 ( .A(n29963), .B(n29964), .Z(n29955) );
  XNOR U31364 ( .A(n29956), .B(n29955), .Z(n29957) );
  XNOR U31365 ( .A(n29958), .B(n29957), .Z(n29987) );
  XNOR U31366 ( .A(sreg[1715]), .B(n29987), .Z(n29989) );
  NANDN U31367 ( .A(sreg[1714]), .B(n29950), .Z(n29954) );
  NAND U31368 ( .A(n29952), .B(n29951), .Z(n29953) );
  NAND U31369 ( .A(n29954), .B(n29953), .Z(n29988) );
  XNOR U31370 ( .A(n29989), .B(n29988), .Z(c[1715]) );
  NANDN U31371 ( .A(n29956), .B(n29955), .Z(n29960) );
  NANDN U31372 ( .A(n29958), .B(n29957), .Z(n29959) );
  AND U31373 ( .A(n29960), .B(n29959), .Z(n29995) );
  NANDN U31374 ( .A(n29962), .B(n29961), .Z(n29966) );
  NANDN U31375 ( .A(n29964), .B(n29963), .Z(n29965) );
  AND U31376 ( .A(n29966), .B(n29965), .Z(n29993) );
  NAND U31377 ( .A(n42143), .B(n29967), .Z(n29969) );
  XNOR U31378 ( .A(a[694]), .B(n4171), .Z(n30004) );
  NAND U31379 ( .A(n42144), .B(n30004), .Z(n29968) );
  AND U31380 ( .A(n29969), .B(n29968), .Z(n30019) );
  XOR U31381 ( .A(a[698]), .B(n42012), .Z(n30007) );
  XNOR U31382 ( .A(n30019), .B(n30018), .Z(n30021) );
  AND U31383 ( .A(a[700]), .B(b[0]), .Z(n29971) );
  XNOR U31384 ( .A(n29971), .B(n4071), .Z(n29973) );
  NANDN U31385 ( .A(b[0]), .B(a[699]), .Z(n29972) );
  NAND U31386 ( .A(n29973), .B(n29972), .Z(n30015) );
  XOR U31387 ( .A(a[696]), .B(n42085), .Z(n30011) );
  AND U31388 ( .A(a[692]), .B(b[7]), .Z(n30012) );
  XNOR U31389 ( .A(n30013), .B(n30012), .Z(n30014) );
  XNOR U31390 ( .A(n30015), .B(n30014), .Z(n30020) );
  XOR U31391 ( .A(n30021), .B(n30020), .Z(n29999) );
  NANDN U31392 ( .A(n29976), .B(n29975), .Z(n29980) );
  NANDN U31393 ( .A(n29978), .B(n29977), .Z(n29979) );
  AND U31394 ( .A(n29980), .B(n29979), .Z(n29998) );
  XNOR U31395 ( .A(n29999), .B(n29998), .Z(n30000) );
  NANDN U31396 ( .A(n29982), .B(n29981), .Z(n29986) );
  NAND U31397 ( .A(n29984), .B(n29983), .Z(n29985) );
  NAND U31398 ( .A(n29986), .B(n29985), .Z(n30001) );
  XNOR U31399 ( .A(n30000), .B(n30001), .Z(n29992) );
  XNOR U31400 ( .A(n29993), .B(n29992), .Z(n29994) );
  XNOR U31401 ( .A(n29995), .B(n29994), .Z(n30024) );
  XNOR U31402 ( .A(sreg[1716]), .B(n30024), .Z(n30026) );
  NANDN U31403 ( .A(sreg[1715]), .B(n29987), .Z(n29991) );
  NAND U31404 ( .A(n29989), .B(n29988), .Z(n29990) );
  NAND U31405 ( .A(n29991), .B(n29990), .Z(n30025) );
  XNOR U31406 ( .A(n30026), .B(n30025), .Z(c[1716]) );
  NANDN U31407 ( .A(n29993), .B(n29992), .Z(n29997) );
  NANDN U31408 ( .A(n29995), .B(n29994), .Z(n29996) );
  AND U31409 ( .A(n29997), .B(n29996), .Z(n30032) );
  NANDN U31410 ( .A(n29999), .B(n29998), .Z(n30003) );
  NANDN U31411 ( .A(n30001), .B(n30000), .Z(n30002) );
  AND U31412 ( .A(n30003), .B(n30002), .Z(n30030) );
  NAND U31413 ( .A(n42143), .B(n30004), .Z(n30006) );
  XNOR U31414 ( .A(a[695]), .B(n4171), .Z(n30041) );
  NAND U31415 ( .A(n42144), .B(n30041), .Z(n30005) );
  AND U31416 ( .A(n30006), .B(n30005), .Z(n30056) );
  XOR U31417 ( .A(a[699]), .B(n42012), .Z(n30044) );
  XNOR U31418 ( .A(n30056), .B(n30055), .Z(n30058) );
  AND U31419 ( .A(a[701]), .B(b[0]), .Z(n30008) );
  XNOR U31420 ( .A(n30008), .B(n4071), .Z(n30010) );
  NANDN U31421 ( .A(b[0]), .B(a[700]), .Z(n30009) );
  NAND U31422 ( .A(n30010), .B(n30009), .Z(n30052) );
  XOR U31423 ( .A(a[697]), .B(n42085), .Z(n30045) );
  AND U31424 ( .A(a[693]), .B(b[7]), .Z(n30049) );
  XNOR U31425 ( .A(n30050), .B(n30049), .Z(n30051) );
  XNOR U31426 ( .A(n30052), .B(n30051), .Z(n30057) );
  XOR U31427 ( .A(n30058), .B(n30057), .Z(n30036) );
  NANDN U31428 ( .A(n30013), .B(n30012), .Z(n30017) );
  NANDN U31429 ( .A(n30015), .B(n30014), .Z(n30016) );
  AND U31430 ( .A(n30017), .B(n30016), .Z(n30035) );
  XNOR U31431 ( .A(n30036), .B(n30035), .Z(n30037) );
  NANDN U31432 ( .A(n30019), .B(n30018), .Z(n30023) );
  NAND U31433 ( .A(n30021), .B(n30020), .Z(n30022) );
  NAND U31434 ( .A(n30023), .B(n30022), .Z(n30038) );
  XNOR U31435 ( .A(n30037), .B(n30038), .Z(n30029) );
  XNOR U31436 ( .A(n30030), .B(n30029), .Z(n30031) );
  XNOR U31437 ( .A(n30032), .B(n30031), .Z(n30061) );
  XNOR U31438 ( .A(sreg[1717]), .B(n30061), .Z(n30063) );
  NANDN U31439 ( .A(sreg[1716]), .B(n30024), .Z(n30028) );
  NAND U31440 ( .A(n30026), .B(n30025), .Z(n30027) );
  NAND U31441 ( .A(n30028), .B(n30027), .Z(n30062) );
  XNOR U31442 ( .A(n30063), .B(n30062), .Z(c[1717]) );
  NANDN U31443 ( .A(n30030), .B(n30029), .Z(n30034) );
  NANDN U31444 ( .A(n30032), .B(n30031), .Z(n30033) );
  AND U31445 ( .A(n30034), .B(n30033), .Z(n30069) );
  NANDN U31446 ( .A(n30036), .B(n30035), .Z(n30040) );
  NANDN U31447 ( .A(n30038), .B(n30037), .Z(n30039) );
  AND U31448 ( .A(n30040), .B(n30039), .Z(n30067) );
  NAND U31449 ( .A(n42143), .B(n30041), .Z(n30043) );
  XNOR U31450 ( .A(a[696]), .B(n4171), .Z(n30078) );
  NAND U31451 ( .A(n42144), .B(n30078), .Z(n30042) );
  AND U31452 ( .A(n30043), .B(n30042), .Z(n30093) );
  XOR U31453 ( .A(a[700]), .B(n42012), .Z(n30081) );
  XNOR U31454 ( .A(n30093), .B(n30092), .Z(n30095) );
  XOR U31455 ( .A(a[698]), .B(n42085), .Z(n30085) );
  AND U31456 ( .A(a[694]), .B(b[7]), .Z(n30086) );
  XNOR U31457 ( .A(n30087), .B(n30086), .Z(n30088) );
  AND U31458 ( .A(a[702]), .B(b[0]), .Z(n30046) );
  XNOR U31459 ( .A(n30046), .B(n4071), .Z(n30048) );
  NANDN U31460 ( .A(b[0]), .B(a[701]), .Z(n30047) );
  NAND U31461 ( .A(n30048), .B(n30047), .Z(n30089) );
  XNOR U31462 ( .A(n30088), .B(n30089), .Z(n30094) );
  XOR U31463 ( .A(n30095), .B(n30094), .Z(n30073) );
  NANDN U31464 ( .A(n30050), .B(n30049), .Z(n30054) );
  NANDN U31465 ( .A(n30052), .B(n30051), .Z(n30053) );
  AND U31466 ( .A(n30054), .B(n30053), .Z(n30072) );
  XNOR U31467 ( .A(n30073), .B(n30072), .Z(n30074) );
  NANDN U31468 ( .A(n30056), .B(n30055), .Z(n30060) );
  NAND U31469 ( .A(n30058), .B(n30057), .Z(n30059) );
  NAND U31470 ( .A(n30060), .B(n30059), .Z(n30075) );
  XNOR U31471 ( .A(n30074), .B(n30075), .Z(n30066) );
  XNOR U31472 ( .A(n30067), .B(n30066), .Z(n30068) );
  XNOR U31473 ( .A(n30069), .B(n30068), .Z(n30098) );
  XNOR U31474 ( .A(sreg[1718]), .B(n30098), .Z(n30100) );
  NANDN U31475 ( .A(sreg[1717]), .B(n30061), .Z(n30065) );
  NAND U31476 ( .A(n30063), .B(n30062), .Z(n30064) );
  NAND U31477 ( .A(n30065), .B(n30064), .Z(n30099) );
  XNOR U31478 ( .A(n30100), .B(n30099), .Z(c[1718]) );
  NANDN U31479 ( .A(n30067), .B(n30066), .Z(n30071) );
  NANDN U31480 ( .A(n30069), .B(n30068), .Z(n30070) );
  AND U31481 ( .A(n30071), .B(n30070), .Z(n30106) );
  NANDN U31482 ( .A(n30073), .B(n30072), .Z(n30077) );
  NANDN U31483 ( .A(n30075), .B(n30074), .Z(n30076) );
  AND U31484 ( .A(n30077), .B(n30076), .Z(n30104) );
  NAND U31485 ( .A(n42143), .B(n30078), .Z(n30080) );
  XNOR U31486 ( .A(a[697]), .B(n4171), .Z(n30115) );
  NAND U31487 ( .A(n42144), .B(n30115), .Z(n30079) );
  AND U31488 ( .A(n30080), .B(n30079), .Z(n30130) );
  XOR U31489 ( .A(a[701]), .B(n42012), .Z(n30118) );
  XNOR U31490 ( .A(n30130), .B(n30129), .Z(n30132) );
  AND U31491 ( .A(a[703]), .B(b[0]), .Z(n30082) );
  XNOR U31492 ( .A(n30082), .B(n4071), .Z(n30084) );
  NANDN U31493 ( .A(b[0]), .B(a[702]), .Z(n30083) );
  NAND U31494 ( .A(n30084), .B(n30083), .Z(n30126) );
  XOR U31495 ( .A(a[699]), .B(n42085), .Z(n30122) );
  AND U31496 ( .A(a[695]), .B(b[7]), .Z(n30123) );
  XNOR U31497 ( .A(n30124), .B(n30123), .Z(n30125) );
  XNOR U31498 ( .A(n30126), .B(n30125), .Z(n30131) );
  XOR U31499 ( .A(n30132), .B(n30131), .Z(n30110) );
  NANDN U31500 ( .A(n30087), .B(n30086), .Z(n30091) );
  NANDN U31501 ( .A(n30089), .B(n30088), .Z(n30090) );
  AND U31502 ( .A(n30091), .B(n30090), .Z(n30109) );
  XNOR U31503 ( .A(n30110), .B(n30109), .Z(n30111) );
  NANDN U31504 ( .A(n30093), .B(n30092), .Z(n30097) );
  NAND U31505 ( .A(n30095), .B(n30094), .Z(n30096) );
  NAND U31506 ( .A(n30097), .B(n30096), .Z(n30112) );
  XNOR U31507 ( .A(n30111), .B(n30112), .Z(n30103) );
  XNOR U31508 ( .A(n30104), .B(n30103), .Z(n30105) );
  XNOR U31509 ( .A(n30106), .B(n30105), .Z(n30135) );
  XNOR U31510 ( .A(sreg[1719]), .B(n30135), .Z(n30137) );
  NANDN U31511 ( .A(sreg[1718]), .B(n30098), .Z(n30102) );
  NAND U31512 ( .A(n30100), .B(n30099), .Z(n30101) );
  NAND U31513 ( .A(n30102), .B(n30101), .Z(n30136) );
  XNOR U31514 ( .A(n30137), .B(n30136), .Z(c[1719]) );
  NANDN U31515 ( .A(n30104), .B(n30103), .Z(n30108) );
  NANDN U31516 ( .A(n30106), .B(n30105), .Z(n30107) );
  AND U31517 ( .A(n30108), .B(n30107), .Z(n30143) );
  NANDN U31518 ( .A(n30110), .B(n30109), .Z(n30114) );
  NANDN U31519 ( .A(n30112), .B(n30111), .Z(n30113) );
  AND U31520 ( .A(n30114), .B(n30113), .Z(n30141) );
  NAND U31521 ( .A(n42143), .B(n30115), .Z(n30117) );
  XNOR U31522 ( .A(a[698]), .B(n4171), .Z(n30152) );
  NAND U31523 ( .A(n42144), .B(n30152), .Z(n30116) );
  AND U31524 ( .A(n30117), .B(n30116), .Z(n30167) );
  XOR U31525 ( .A(a[702]), .B(n42012), .Z(n30155) );
  XNOR U31526 ( .A(n30167), .B(n30166), .Z(n30169) );
  AND U31527 ( .A(a[704]), .B(b[0]), .Z(n30119) );
  XNOR U31528 ( .A(n30119), .B(n4071), .Z(n30121) );
  NANDN U31529 ( .A(b[0]), .B(a[703]), .Z(n30120) );
  NAND U31530 ( .A(n30121), .B(n30120), .Z(n30163) );
  XOR U31531 ( .A(a[700]), .B(n42085), .Z(n30159) );
  AND U31532 ( .A(a[696]), .B(b[7]), .Z(n30160) );
  XNOR U31533 ( .A(n30161), .B(n30160), .Z(n30162) );
  XNOR U31534 ( .A(n30163), .B(n30162), .Z(n30168) );
  XOR U31535 ( .A(n30169), .B(n30168), .Z(n30147) );
  NANDN U31536 ( .A(n30124), .B(n30123), .Z(n30128) );
  NANDN U31537 ( .A(n30126), .B(n30125), .Z(n30127) );
  AND U31538 ( .A(n30128), .B(n30127), .Z(n30146) );
  XNOR U31539 ( .A(n30147), .B(n30146), .Z(n30148) );
  NANDN U31540 ( .A(n30130), .B(n30129), .Z(n30134) );
  NAND U31541 ( .A(n30132), .B(n30131), .Z(n30133) );
  NAND U31542 ( .A(n30134), .B(n30133), .Z(n30149) );
  XNOR U31543 ( .A(n30148), .B(n30149), .Z(n30140) );
  XNOR U31544 ( .A(n30141), .B(n30140), .Z(n30142) );
  XNOR U31545 ( .A(n30143), .B(n30142), .Z(n30172) );
  XNOR U31546 ( .A(sreg[1720]), .B(n30172), .Z(n30174) );
  NANDN U31547 ( .A(sreg[1719]), .B(n30135), .Z(n30139) );
  NAND U31548 ( .A(n30137), .B(n30136), .Z(n30138) );
  NAND U31549 ( .A(n30139), .B(n30138), .Z(n30173) );
  XNOR U31550 ( .A(n30174), .B(n30173), .Z(c[1720]) );
  NANDN U31551 ( .A(n30141), .B(n30140), .Z(n30145) );
  NANDN U31552 ( .A(n30143), .B(n30142), .Z(n30144) );
  AND U31553 ( .A(n30145), .B(n30144), .Z(n30180) );
  NANDN U31554 ( .A(n30147), .B(n30146), .Z(n30151) );
  NANDN U31555 ( .A(n30149), .B(n30148), .Z(n30150) );
  AND U31556 ( .A(n30151), .B(n30150), .Z(n30178) );
  NAND U31557 ( .A(n42143), .B(n30152), .Z(n30154) );
  XNOR U31558 ( .A(a[699]), .B(n4171), .Z(n30189) );
  NAND U31559 ( .A(n42144), .B(n30189), .Z(n30153) );
  AND U31560 ( .A(n30154), .B(n30153), .Z(n30204) );
  XOR U31561 ( .A(a[703]), .B(n42012), .Z(n30192) );
  XNOR U31562 ( .A(n30204), .B(n30203), .Z(n30206) );
  AND U31563 ( .A(a[705]), .B(b[0]), .Z(n30156) );
  XNOR U31564 ( .A(n30156), .B(n4071), .Z(n30158) );
  NANDN U31565 ( .A(b[0]), .B(a[704]), .Z(n30157) );
  NAND U31566 ( .A(n30158), .B(n30157), .Z(n30200) );
  XOR U31567 ( .A(a[701]), .B(n42085), .Z(n30193) );
  AND U31568 ( .A(a[697]), .B(b[7]), .Z(n30197) );
  XNOR U31569 ( .A(n30198), .B(n30197), .Z(n30199) );
  XNOR U31570 ( .A(n30200), .B(n30199), .Z(n30205) );
  XOR U31571 ( .A(n30206), .B(n30205), .Z(n30184) );
  NANDN U31572 ( .A(n30161), .B(n30160), .Z(n30165) );
  NANDN U31573 ( .A(n30163), .B(n30162), .Z(n30164) );
  AND U31574 ( .A(n30165), .B(n30164), .Z(n30183) );
  XNOR U31575 ( .A(n30184), .B(n30183), .Z(n30185) );
  NANDN U31576 ( .A(n30167), .B(n30166), .Z(n30171) );
  NAND U31577 ( .A(n30169), .B(n30168), .Z(n30170) );
  NAND U31578 ( .A(n30171), .B(n30170), .Z(n30186) );
  XNOR U31579 ( .A(n30185), .B(n30186), .Z(n30177) );
  XNOR U31580 ( .A(n30178), .B(n30177), .Z(n30179) );
  XNOR U31581 ( .A(n30180), .B(n30179), .Z(n30209) );
  XNOR U31582 ( .A(sreg[1721]), .B(n30209), .Z(n30211) );
  NANDN U31583 ( .A(sreg[1720]), .B(n30172), .Z(n30176) );
  NAND U31584 ( .A(n30174), .B(n30173), .Z(n30175) );
  NAND U31585 ( .A(n30176), .B(n30175), .Z(n30210) );
  XNOR U31586 ( .A(n30211), .B(n30210), .Z(c[1721]) );
  NANDN U31587 ( .A(n30178), .B(n30177), .Z(n30182) );
  NANDN U31588 ( .A(n30180), .B(n30179), .Z(n30181) );
  AND U31589 ( .A(n30182), .B(n30181), .Z(n30217) );
  NANDN U31590 ( .A(n30184), .B(n30183), .Z(n30188) );
  NANDN U31591 ( .A(n30186), .B(n30185), .Z(n30187) );
  AND U31592 ( .A(n30188), .B(n30187), .Z(n30215) );
  NAND U31593 ( .A(n42143), .B(n30189), .Z(n30191) );
  XNOR U31594 ( .A(a[700]), .B(n4171), .Z(n30226) );
  NAND U31595 ( .A(n42144), .B(n30226), .Z(n30190) );
  AND U31596 ( .A(n30191), .B(n30190), .Z(n30241) );
  XOR U31597 ( .A(a[704]), .B(n42012), .Z(n30229) );
  XNOR U31598 ( .A(n30241), .B(n30240), .Z(n30243) );
  XOR U31599 ( .A(a[702]), .B(n42085), .Z(n30230) );
  AND U31600 ( .A(a[698]), .B(b[7]), .Z(n30234) );
  XNOR U31601 ( .A(n30235), .B(n30234), .Z(n30236) );
  AND U31602 ( .A(a[706]), .B(b[0]), .Z(n30194) );
  XNOR U31603 ( .A(n30194), .B(n4071), .Z(n30196) );
  NANDN U31604 ( .A(b[0]), .B(a[705]), .Z(n30195) );
  NAND U31605 ( .A(n30196), .B(n30195), .Z(n30237) );
  XNOR U31606 ( .A(n30236), .B(n30237), .Z(n30242) );
  XOR U31607 ( .A(n30243), .B(n30242), .Z(n30221) );
  NANDN U31608 ( .A(n30198), .B(n30197), .Z(n30202) );
  NANDN U31609 ( .A(n30200), .B(n30199), .Z(n30201) );
  AND U31610 ( .A(n30202), .B(n30201), .Z(n30220) );
  XNOR U31611 ( .A(n30221), .B(n30220), .Z(n30222) );
  NANDN U31612 ( .A(n30204), .B(n30203), .Z(n30208) );
  NAND U31613 ( .A(n30206), .B(n30205), .Z(n30207) );
  NAND U31614 ( .A(n30208), .B(n30207), .Z(n30223) );
  XNOR U31615 ( .A(n30222), .B(n30223), .Z(n30214) );
  XNOR U31616 ( .A(n30215), .B(n30214), .Z(n30216) );
  XNOR U31617 ( .A(n30217), .B(n30216), .Z(n30246) );
  XNOR U31618 ( .A(sreg[1722]), .B(n30246), .Z(n30248) );
  NANDN U31619 ( .A(sreg[1721]), .B(n30209), .Z(n30213) );
  NAND U31620 ( .A(n30211), .B(n30210), .Z(n30212) );
  NAND U31621 ( .A(n30213), .B(n30212), .Z(n30247) );
  XNOR U31622 ( .A(n30248), .B(n30247), .Z(c[1722]) );
  NANDN U31623 ( .A(n30215), .B(n30214), .Z(n30219) );
  NANDN U31624 ( .A(n30217), .B(n30216), .Z(n30218) );
  AND U31625 ( .A(n30219), .B(n30218), .Z(n30254) );
  NANDN U31626 ( .A(n30221), .B(n30220), .Z(n30225) );
  NANDN U31627 ( .A(n30223), .B(n30222), .Z(n30224) );
  AND U31628 ( .A(n30225), .B(n30224), .Z(n30252) );
  NAND U31629 ( .A(n42143), .B(n30226), .Z(n30228) );
  XNOR U31630 ( .A(a[701]), .B(n4172), .Z(n30263) );
  NAND U31631 ( .A(n42144), .B(n30263), .Z(n30227) );
  AND U31632 ( .A(n30228), .B(n30227), .Z(n30278) );
  XOR U31633 ( .A(a[705]), .B(n42012), .Z(n30266) );
  XNOR U31634 ( .A(n30278), .B(n30277), .Z(n30280) );
  XOR U31635 ( .A(a[703]), .B(n42085), .Z(n30270) );
  AND U31636 ( .A(a[699]), .B(b[7]), .Z(n30271) );
  XNOR U31637 ( .A(n30272), .B(n30271), .Z(n30273) );
  AND U31638 ( .A(a[707]), .B(b[0]), .Z(n30231) );
  XNOR U31639 ( .A(n30231), .B(n4071), .Z(n30233) );
  NANDN U31640 ( .A(b[0]), .B(a[706]), .Z(n30232) );
  NAND U31641 ( .A(n30233), .B(n30232), .Z(n30274) );
  XNOR U31642 ( .A(n30273), .B(n30274), .Z(n30279) );
  XOR U31643 ( .A(n30280), .B(n30279), .Z(n30258) );
  NANDN U31644 ( .A(n30235), .B(n30234), .Z(n30239) );
  NANDN U31645 ( .A(n30237), .B(n30236), .Z(n30238) );
  AND U31646 ( .A(n30239), .B(n30238), .Z(n30257) );
  XNOR U31647 ( .A(n30258), .B(n30257), .Z(n30259) );
  NANDN U31648 ( .A(n30241), .B(n30240), .Z(n30245) );
  NAND U31649 ( .A(n30243), .B(n30242), .Z(n30244) );
  NAND U31650 ( .A(n30245), .B(n30244), .Z(n30260) );
  XNOR U31651 ( .A(n30259), .B(n30260), .Z(n30251) );
  XNOR U31652 ( .A(n30252), .B(n30251), .Z(n30253) );
  XNOR U31653 ( .A(n30254), .B(n30253), .Z(n30283) );
  XNOR U31654 ( .A(sreg[1723]), .B(n30283), .Z(n30285) );
  NANDN U31655 ( .A(sreg[1722]), .B(n30246), .Z(n30250) );
  NAND U31656 ( .A(n30248), .B(n30247), .Z(n30249) );
  NAND U31657 ( .A(n30250), .B(n30249), .Z(n30284) );
  XNOR U31658 ( .A(n30285), .B(n30284), .Z(c[1723]) );
  NANDN U31659 ( .A(n30252), .B(n30251), .Z(n30256) );
  NANDN U31660 ( .A(n30254), .B(n30253), .Z(n30255) );
  AND U31661 ( .A(n30256), .B(n30255), .Z(n30291) );
  NANDN U31662 ( .A(n30258), .B(n30257), .Z(n30262) );
  NANDN U31663 ( .A(n30260), .B(n30259), .Z(n30261) );
  AND U31664 ( .A(n30262), .B(n30261), .Z(n30289) );
  NAND U31665 ( .A(n42143), .B(n30263), .Z(n30265) );
  XNOR U31666 ( .A(a[702]), .B(n4172), .Z(n30300) );
  NAND U31667 ( .A(n42144), .B(n30300), .Z(n30264) );
  AND U31668 ( .A(n30265), .B(n30264), .Z(n30315) );
  XOR U31669 ( .A(a[706]), .B(n42012), .Z(n30303) );
  XNOR U31670 ( .A(n30315), .B(n30314), .Z(n30317) );
  AND U31671 ( .A(a[708]), .B(b[0]), .Z(n30267) );
  XNOR U31672 ( .A(n30267), .B(n4071), .Z(n30269) );
  NANDN U31673 ( .A(b[0]), .B(a[707]), .Z(n30268) );
  NAND U31674 ( .A(n30269), .B(n30268), .Z(n30311) );
  XOR U31675 ( .A(a[704]), .B(n42085), .Z(n30304) );
  AND U31676 ( .A(a[700]), .B(b[7]), .Z(n30308) );
  XNOR U31677 ( .A(n30309), .B(n30308), .Z(n30310) );
  XNOR U31678 ( .A(n30311), .B(n30310), .Z(n30316) );
  XOR U31679 ( .A(n30317), .B(n30316), .Z(n30295) );
  NANDN U31680 ( .A(n30272), .B(n30271), .Z(n30276) );
  NANDN U31681 ( .A(n30274), .B(n30273), .Z(n30275) );
  AND U31682 ( .A(n30276), .B(n30275), .Z(n30294) );
  XNOR U31683 ( .A(n30295), .B(n30294), .Z(n30296) );
  NANDN U31684 ( .A(n30278), .B(n30277), .Z(n30282) );
  NAND U31685 ( .A(n30280), .B(n30279), .Z(n30281) );
  NAND U31686 ( .A(n30282), .B(n30281), .Z(n30297) );
  XNOR U31687 ( .A(n30296), .B(n30297), .Z(n30288) );
  XNOR U31688 ( .A(n30289), .B(n30288), .Z(n30290) );
  XNOR U31689 ( .A(n30291), .B(n30290), .Z(n30320) );
  XNOR U31690 ( .A(sreg[1724]), .B(n30320), .Z(n30322) );
  NANDN U31691 ( .A(sreg[1723]), .B(n30283), .Z(n30287) );
  NAND U31692 ( .A(n30285), .B(n30284), .Z(n30286) );
  NAND U31693 ( .A(n30287), .B(n30286), .Z(n30321) );
  XNOR U31694 ( .A(n30322), .B(n30321), .Z(c[1724]) );
  NANDN U31695 ( .A(n30289), .B(n30288), .Z(n30293) );
  NANDN U31696 ( .A(n30291), .B(n30290), .Z(n30292) );
  AND U31697 ( .A(n30293), .B(n30292), .Z(n30328) );
  NANDN U31698 ( .A(n30295), .B(n30294), .Z(n30299) );
  NANDN U31699 ( .A(n30297), .B(n30296), .Z(n30298) );
  AND U31700 ( .A(n30299), .B(n30298), .Z(n30326) );
  NAND U31701 ( .A(n42143), .B(n30300), .Z(n30302) );
  XNOR U31702 ( .A(a[703]), .B(n4172), .Z(n30337) );
  NAND U31703 ( .A(n42144), .B(n30337), .Z(n30301) );
  AND U31704 ( .A(n30302), .B(n30301), .Z(n30352) );
  XOR U31705 ( .A(a[707]), .B(n42012), .Z(n30340) );
  XNOR U31706 ( .A(n30352), .B(n30351), .Z(n30354) );
  XOR U31707 ( .A(a[705]), .B(n42085), .Z(n30344) );
  AND U31708 ( .A(a[701]), .B(b[7]), .Z(n30345) );
  XNOR U31709 ( .A(n30346), .B(n30345), .Z(n30347) );
  AND U31710 ( .A(a[709]), .B(b[0]), .Z(n30305) );
  XNOR U31711 ( .A(n30305), .B(n4071), .Z(n30307) );
  NANDN U31712 ( .A(b[0]), .B(a[708]), .Z(n30306) );
  NAND U31713 ( .A(n30307), .B(n30306), .Z(n30348) );
  XNOR U31714 ( .A(n30347), .B(n30348), .Z(n30353) );
  XOR U31715 ( .A(n30354), .B(n30353), .Z(n30332) );
  NANDN U31716 ( .A(n30309), .B(n30308), .Z(n30313) );
  NANDN U31717 ( .A(n30311), .B(n30310), .Z(n30312) );
  AND U31718 ( .A(n30313), .B(n30312), .Z(n30331) );
  XNOR U31719 ( .A(n30332), .B(n30331), .Z(n30333) );
  NANDN U31720 ( .A(n30315), .B(n30314), .Z(n30319) );
  NAND U31721 ( .A(n30317), .B(n30316), .Z(n30318) );
  NAND U31722 ( .A(n30319), .B(n30318), .Z(n30334) );
  XNOR U31723 ( .A(n30333), .B(n30334), .Z(n30325) );
  XNOR U31724 ( .A(n30326), .B(n30325), .Z(n30327) );
  XNOR U31725 ( .A(n30328), .B(n30327), .Z(n30357) );
  XNOR U31726 ( .A(sreg[1725]), .B(n30357), .Z(n30359) );
  NANDN U31727 ( .A(sreg[1724]), .B(n30320), .Z(n30324) );
  NAND U31728 ( .A(n30322), .B(n30321), .Z(n30323) );
  NAND U31729 ( .A(n30324), .B(n30323), .Z(n30358) );
  XNOR U31730 ( .A(n30359), .B(n30358), .Z(c[1725]) );
  NANDN U31731 ( .A(n30326), .B(n30325), .Z(n30330) );
  NANDN U31732 ( .A(n30328), .B(n30327), .Z(n30329) );
  AND U31733 ( .A(n30330), .B(n30329), .Z(n30365) );
  NANDN U31734 ( .A(n30332), .B(n30331), .Z(n30336) );
  NANDN U31735 ( .A(n30334), .B(n30333), .Z(n30335) );
  AND U31736 ( .A(n30336), .B(n30335), .Z(n30363) );
  NAND U31737 ( .A(n42143), .B(n30337), .Z(n30339) );
  XNOR U31738 ( .A(a[704]), .B(n4172), .Z(n30374) );
  NAND U31739 ( .A(n42144), .B(n30374), .Z(n30338) );
  AND U31740 ( .A(n30339), .B(n30338), .Z(n30389) );
  XOR U31741 ( .A(a[708]), .B(n42012), .Z(n30377) );
  XNOR U31742 ( .A(n30389), .B(n30388), .Z(n30391) );
  AND U31743 ( .A(a[710]), .B(b[0]), .Z(n30341) );
  XNOR U31744 ( .A(n30341), .B(n4071), .Z(n30343) );
  NANDN U31745 ( .A(b[0]), .B(a[709]), .Z(n30342) );
  NAND U31746 ( .A(n30343), .B(n30342), .Z(n30385) );
  XOR U31747 ( .A(a[706]), .B(n42085), .Z(n30381) );
  AND U31748 ( .A(a[702]), .B(b[7]), .Z(n30382) );
  XNOR U31749 ( .A(n30383), .B(n30382), .Z(n30384) );
  XNOR U31750 ( .A(n30385), .B(n30384), .Z(n30390) );
  XOR U31751 ( .A(n30391), .B(n30390), .Z(n30369) );
  NANDN U31752 ( .A(n30346), .B(n30345), .Z(n30350) );
  NANDN U31753 ( .A(n30348), .B(n30347), .Z(n30349) );
  AND U31754 ( .A(n30350), .B(n30349), .Z(n30368) );
  XNOR U31755 ( .A(n30369), .B(n30368), .Z(n30370) );
  NANDN U31756 ( .A(n30352), .B(n30351), .Z(n30356) );
  NAND U31757 ( .A(n30354), .B(n30353), .Z(n30355) );
  NAND U31758 ( .A(n30356), .B(n30355), .Z(n30371) );
  XNOR U31759 ( .A(n30370), .B(n30371), .Z(n30362) );
  XNOR U31760 ( .A(n30363), .B(n30362), .Z(n30364) );
  XNOR U31761 ( .A(n30365), .B(n30364), .Z(n30394) );
  XNOR U31762 ( .A(sreg[1726]), .B(n30394), .Z(n30396) );
  NANDN U31763 ( .A(sreg[1725]), .B(n30357), .Z(n30361) );
  NAND U31764 ( .A(n30359), .B(n30358), .Z(n30360) );
  NAND U31765 ( .A(n30361), .B(n30360), .Z(n30395) );
  XNOR U31766 ( .A(n30396), .B(n30395), .Z(c[1726]) );
  NANDN U31767 ( .A(n30363), .B(n30362), .Z(n30367) );
  NANDN U31768 ( .A(n30365), .B(n30364), .Z(n30366) );
  AND U31769 ( .A(n30367), .B(n30366), .Z(n30402) );
  NANDN U31770 ( .A(n30369), .B(n30368), .Z(n30373) );
  NANDN U31771 ( .A(n30371), .B(n30370), .Z(n30372) );
  AND U31772 ( .A(n30373), .B(n30372), .Z(n30400) );
  NAND U31773 ( .A(n42143), .B(n30374), .Z(n30376) );
  XNOR U31774 ( .A(a[705]), .B(n4172), .Z(n30411) );
  NAND U31775 ( .A(n42144), .B(n30411), .Z(n30375) );
  AND U31776 ( .A(n30376), .B(n30375), .Z(n30426) );
  XOR U31777 ( .A(a[709]), .B(n42012), .Z(n30414) );
  XNOR U31778 ( .A(n30426), .B(n30425), .Z(n30428) );
  AND U31779 ( .A(a[711]), .B(b[0]), .Z(n30378) );
  XNOR U31780 ( .A(n30378), .B(n4071), .Z(n30380) );
  NANDN U31781 ( .A(b[0]), .B(a[710]), .Z(n30379) );
  NAND U31782 ( .A(n30380), .B(n30379), .Z(n30422) );
  XOR U31783 ( .A(a[707]), .B(n42085), .Z(n30418) );
  AND U31784 ( .A(a[703]), .B(b[7]), .Z(n30419) );
  XNOR U31785 ( .A(n30420), .B(n30419), .Z(n30421) );
  XNOR U31786 ( .A(n30422), .B(n30421), .Z(n30427) );
  XOR U31787 ( .A(n30428), .B(n30427), .Z(n30406) );
  NANDN U31788 ( .A(n30383), .B(n30382), .Z(n30387) );
  NANDN U31789 ( .A(n30385), .B(n30384), .Z(n30386) );
  AND U31790 ( .A(n30387), .B(n30386), .Z(n30405) );
  XNOR U31791 ( .A(n30406), .B(n30405), .Z(n30407) );
  NANDN U31792 ( .A(n30389), .B(n30388), .Z(n30393) );
  NAND U31793 ( .A(n30391), .B(n30390), .Z(n30392) );
  NAND U31794 ( .A(n30393), .B(n30392), .Z(n30408) );
  XNOR U31795 ( .A(n30407), .B(n30408), .Z(n30399) );
  XNOR U31796 ( .A(n30400), .B(n30399), .Z(n30401) );
  XNOR U31797 ( .A(n30402), .B(n30401), .Z(n30431) );
  XNOR U31798 ( .A(sreg[1727]), .B(n30431), .Z(n30433) );
  NANDN U31799 ( .A(sreg[1726]), .B(n30394), .Z(n30398) );
  NAND U31800 ( .A(n30396), .B(n30395), .Z(n30397) );
  NAND U31801 ( .A(n30398), .B(n30397), .Z(n30432) );
  XNOR U31802 ( .A(n30433), .B(n30432), .Z(c[1727]) );
  NANDN U31803 ( .A(n30400), .B(n30399), .Z(n30404) );
  NANDN U31804 ( .A(n30402), .B(n30401), .Z(n30403) );
  AND U31805 ( .A(n30404), .B(n30403), .Z(n30439) );
  NANDN U31806 ( .A(n30406), .B(n30405), .Z(n30410) );
  NANDN U31807 ( .A(n30408), .B(n30407), .Z(n30409) );
  AND U31808 ( .A(n30410), .B(n30409), .Z(n30437) );
  NAND U31809 ( .A(n42143), .B(n30411), .Z(n30413) );
  XNOR U31810 ( .A(a[706]), .B(n4172), .Z(n30448) );
  NAND U31811 ( .A(n42144), .B(n30448), .Z(n30412) );
  AND U31812 ( .A(n30413), .B(n30412), .Z(n30463) );
  XOR U31813 ( .A(a[710]), .B(n42012), .Z(n30451) );
  XNOR U31814 ( .A(n30463), .B(n30462), .Z(n30465) );
  AND U31815 ( .A(a[712]), .B(b[0]), .Z(n30415) );
  XNOR U31816 ( .A(n30415), .B(n4071), .Z(n30417) );
  NANDN U31817 ( .A(b[0]), .B(a[711]), .Z(n30416) );
  NAND U31818 ( .A(n30417), .B(n30416), .Z(n30459) );
  XOR U31819 ( .A(a[708]), .B(n42085), .Z(n30452) );
  AND U31820 ( .A(a[704]), .B(b[7]), .Z(n30456) );
  XNOR U31821 ( .A(n30457), .B(n30456), .Z(n30458) );
  XNOR U31822 ( .A(n30459), .B(n30458), .Z(n30464) );
  XOR U31823 ( .A(n30465), .B(n30464), .Z(n30443) );
  NANDN U31824 ( .A(n30420), .B(n30419), .Z(n30424) );
  NANDN U31825 ( .A(n30422), .B(n30421), .Z(n30423) );
  AND U31826 ( .A(n30424), .B(n30423), .Z(n30442) );
  XNOR U31827 ( .A(n30443), .B(n30442), .Z(n30444) );
  NANDN U31828 ( .A(n30426), .B(n30425), .Z(n30430) );
  NAND U31829 ( .A(n30428), .B(n30427), .Z(n30429) );
  NAND U31830 ( .A(n30430), .B(n30429), .Z(n30445) );
  XNOR U31831 ( .A(n30444), .B(n30445), .Z(n30436) );
  XNOR U31832 ( .A(n30437), .B(n30436), .Z(n30438) );
  XNOR U31833 ( .A(n30439), .B(n30438), .Z(n30468) );
  XNOR U31834 ( .A(sreg[1728]), .B(n30468), .Z(n30470) );
  NANDN U31835 ( .A(sreg[1727]), .B(n30431), .Z(n30435) );
  NAND U31836 ( .A(n30433), .B(n30432), .Z(n30434) );
  NAND U31837 ( .A(n30435), .B(n30434), .Z(n30469) );
  XNOR U31838 ( .A(n30470), .B(n30469), .Z(c[1728]) );
  NANDN U31839 ( .A(n30437), .B(n30436), .Z(n30441) );
  NANDN U31840 ( .A(n30439), .B(n30438), .Z(n30440) );
  AND U31841 ( .A(n30441), .B(n30440), .Z(n30476) );
  NANDN U31842 ( .A(n30443), .B(n30442), .Z(n30447) );
  NANDN U31843 ( .A(n30445), .B(n30444), .Z(n30446) );
  AND U31844 ( .A(n30447), .B(n30446), .Z(n30474) );
  NAND U31845 ( .A(n42143), .B(n30448), .Z(n30450) );
  XNOR U31846 ( .A(a[707]), .B(n4172), .Z(n30485) );
  NAND U31847 ( .A(n42144), .B(n30485), .Z(n30449) );
  AND U31848 ( .A(n30450), .B(n30449), .Z(n30500) );
  XOR U31849 ( .A(a[711]), .B(n42012), .Z(n30488) );
  XNOR U31850 ( .A(n30500), .B(n30499), .Z(n30502) );
  XOR U31851 ( .A(a[709]), .B(n42085), .Z(n30492) );
  AND U31852 ( .A(a[705]), .B(b[7]), .Z(n30493) );
  XNOR U31853 ( .A(n30494), .B(n30493), .Z(n30495) );
  AND U31854 ( .A(a[713]), .B(b[0]), .Z(n30453) );
  XNOR U31855 ( .A(n30453), .B(n4071), .Z(n30455) );
  NANDN U31856 ( .A(b[0]), .B(a[712]), .Z(n30454) );
  NAND U31857 ( .A(n30455), .B(n30454), .Z(n30496) );
  XNOR U31858 ( .A(n30495), .B(n30496), .Z(n30501) );
  XOR U31859 ( .A(n30502), .B(n30501), .Z(n30480) );
  NANDN U31860 ( .A(n30457), .B(n30456), .Z(n30461) );
  NANDN U31861 ( .A(n30459), .B(n30458), .Z(n30460) );
  AND U31862 ( .A(n30461), .B(n30460), .Z(n30479) );
  XNOR U31863 ( .A(n30480), .B(n30479), .Z(n30481) );
  NANDN U31864 ( .A(n30463), .B(n30462), .Z(n30467) );
  NAND U31865 ( .A(n30465), .B(n30464), .Z(n30466) );
  NAND U31866 ( .A(n30467), .B(n30466), .Z(n30482) );
  XNOR U31867 ( .A(n30481), .B(n30482), .Z(n30473) );
  XNOR U31868 ( .A(n30474), .B(n30473), .Z(n30475) );
  XNOR U31869 ( .A(n30476), .B(n30475), .Z(n30505) );
  XNOR U31870 ( .A(sreg[1729]), .B(n30505), .Z(n30507) );
  NANDN U31871 ( .A(sreg[1728]), .B(n30468), .Z(n30472) );
  NAND U31872 ( .A(n30470), .B(n30469), .Z(n30471) );
  NAND U31873 ( .A(n30472), .B(n30471), .Z(n30506) );
  XNOR U31874 ( .A(n30507), .B(n30506), .Z(c[1729]) );
  NANDN U31875 ( .A(n30474), .B(n30473), .Z(n30478) );
  NANDN U31876 ( .A(n30476), .B(n30475), .Z(n30477) );
  AND U31877 ( .A(n30478), .B(n30477), .Z(n30513) );
  NANDN U31878 ( .A(n30480), .B(n30479), .Z(n30484) );
  NANDN U31879 ( .A(n30482), .B(n30481), .Z(n30483) );
  AND U31880 ( .A(n30484), .B(n30483), .Z(n30511) );
  NAND U31881 ( .A(n42143), .B(n30485), .Z(n30487) );
  XNOR U31882 ( .A(a[708]), .B(n4173), .Z(n30522) );
  NAND U31883 ( .A(n42144), .B(n30522), .Z(n30486) );
  AND U31884 ( .A(n30487), .B(n30486), .Z(n30537) );
  XOR U31885 ( .A(a[712]), .B(n42012), .Z(n30525) );
  XNOR U31886 ( .A(n30537), .B(n30536), .Z(n30539) );
  AND U31887 ( .A(a[714]), .B(b[0]), .Z(n30489) );
  XNOR U31888 ( .A(n30489), .B(n4071), .Z(n30491) );
  NANDN U31889 ( .A(b[0]), .B(a[713]), .Z(n30490) );
  NAND U31890 ( .A(n30491), .B(n30490), .Z(n30533) );
  XOR U31891 ( .A(a[710]), .B(n42085), .Z(n30529) );
  AND U31892 ( .A(a[706]), .B(b[7]), .Z(n30530) );
  XNOR U31893 ( .A(n30531), .B(n30530), .Z(n30532) );
  XNOR U31894 ( .A(n30533), .B(n30532), .Z(n30538) );
  XOR U31895 ( .A(n30539), .B(n30538), .Z(n30517) );
  NANDN U31896 ( .A(n30494), .B(n30493), .Z(n30498) );
  NANDN U31897 ( .A(n30496), .B(n30495), .Z(n30497) );
  AND U31898 ( .A(n30498), .B(n30497), .Z(n30516) );
  XNOR U31899 ( .A(n30517), .B(n30516), .Z(n30518) );
  NANDN U31900 ( .A(n30500), .B(n30499), .Z(n30504) );
  NAND U31901 ( .A(n30502), .B(n30501), .Z(n30503) );
  NAND U31902 ( .A(n30504), .B(n30503), .Z(n30519) );
  XNOR U31903 ( .A(n30518), .B(n30519), .Z(n30510) );
  XNOR U31904 ( .A(n30511), .B(n30510), .Z(n30512) );
  XNOR U31905 ( .A(n30513), .B(n30512), .Z(n30542) );
  XNOR U31906 ( .A(sreg[1730]), .B(n30542), .Z(n30544) );
  NANDN U31907 ( .A(sreg[1729]), .B(n30505), .Z(n30509) );
  NAND U31908 ( .A(n30507), .B(n30506), .Z(n30508) );
  NAND U31909 ( .A(n30509), .B(n30508), .Z(n30543) );
  XNOR U31910 ( .A(n30544), .B(n30543), .Z(c[1730]) );
  NANDN U31911 ( .A(n30511), .B(n30510), .Z(n30515) );
  NANDN U31912 ( .A(n30513), .B(n30512), .Z(n30514) );
  AND U31913 ( .A(n30515), .B(n30514), .Z(n30550) );
  NANDN U31914 ( .A(n30517), .B(n30516), .Z(n30521) );
  NANDN U31915 ( .A(n30519), .B(n30518), .Z(n30520) );
  AND U31916 ( .A(n30521), .B(n30520), .Z(n30548) );
  NAND U31917 ( .A(n42143), .B(n30522), .Z(n30524) );
  XNOR U31918 ( .A(a[709]), .B(n4173), .Z(n30559) );
  NAND U31919 ( .A(n42144), .B(n30559), .Z(n30523) );
  AND U31920 ( .A(n30524), .B(n30523), .Z(n30574) );
  XOR U31921 ( .A(a[713]), .B(n42012), .Z(n30562) );
  XNOR U31922 ( .A(n30574), .B(n30573), .Z(n30576) );
  AND U31923 ( .A(a[715]), .B(b[0]), .Z(n30526) );
  XNOR U31924 ( .A(n30526), .B(n4071), .Z(n30528) );
  NANDN U31925 ( .A(b[0]), .B(a[714]), .Z(n30527) );
  NAND U31926 ( .A(n30528), .B(n30527), .Z(n30570) );
  XOR U31927 ( .A(a[711]), .B(n42085), .Z(n30563) );
  AND U31928 ( .A(a[707]), .B(b[7]), .Z(n30567) );
  XNOR U31929 ( .A(n30568), .B(n30567), .Z(n30569) );
  XNOR U31930 ( .A(n30570), .B(n30569), .Z(n30575) );
  XOR U31931 ( .A(n30576), .B(n30575), .Z(n30554) );
  NANDN U31932 ( .A(n30531), .B(n30530), .Z(n30535) );
  NANDN U31933 ( .A(n30533), .B(n30532), .Z(n30534) );
  AND U31934 ( .A(n30535), .B(n30534), .Z(n30553) );
  XNOR U31935 ( .A(n30554), .B(n30553), .Z(n30555) );
  NANDN U31936 ( .A(n30537), .B(n30536), .Z(n30541) );
  NAND U31937 ( .A(n30539), .B(n30538), .Z(n30540) );
  NAND U31938 ( .A(n30541), .B(n30540), .Z(n30556) );
  XNOR U31939 ( .A(n30555), .B(n30556), .Z(n30547) );
  XNOR U31940 ( .A(n30548), .B(n30547), .Z(n30549) );
  XNOR U31941 ( .A(n30550), .B(n30549), .Z(n30579) );
  XNOR U31942 ( .A(sreg[1731]), .B(n30579), .Z(n30581) );
  NANDN U31943 ( .A(sreg[1730]), .B(n30542), .Z(n30546) );
  NAND U31944 ( .A(n30544), .B(n30543), .Z(n30545) );
  NAND U31945 ( .A(n30546), .B(n30545), .Z(n30580) );
  XNOR U31946 ( .A(n30581), .B(n30580), .Z(c[1731]) );
  NANDN U31947 ( .A(n30548), .B(n30547), .Z(n30552) );
  NANDN U31948 ( .A(n30550), .B(n30549), .Z(n30551) );
  AND U31949 ( .A(n30552), .B(n30551), .Z(n30587) );
  NANDN U31950 ( .A(n30554), .B(n30553), .Z(n30558) );
  NANDN U31951 ( .A(n30556), .B(n30555), .Z(n30557) );
  AND U31952 ( .A(n30558), .B(n30557), .Z(n30585) );
  NAND U31953 ( .A(n42143), .B(n30559), .Z(n30561) );
  XNOR U31954 ( .A(a[710]), .B(n4173), .Z(n30596) );
  NAND U31955 ( .A(n42144), .B(n30596), .Z(n30560) );
  AND U31956 ( .A(n30561), .B(n30560), .Z(n30611) );
  XOR U31957 ( .A(a[714]), .B(n42012), .Z(n30599) );
  XNOR U31958 ( .A(n30611), .B(n30610), .Z(n30613) );
  XOR U31959 ( .A(a[712]), .B(n42085), .Z(n30603) );
  AND U31960 ( .A(a[708]), .B(b[7]), .Z(n30604) );
  XNOR U31961 ( .A(n30605), .B(n30604), .Z(n30606) );
  AND U31962 ( .A(a[716]), .B(b[0]), .Z(n30564) );
  XNOR U31963 ( .A(n30564), .B(n4071), .Z(n30566) );
  NANDN U31964 ( .A(b[0]), .B(a[715]), .Z(n30565) );
  NAND U31965 ( .A(n30566), .B(n30565), .Z(n30607) );
  XNOR U31966 ( .A(n30606), .B(n30607), .Z(n30612) );
  XOR U31967 ( .A(n30613), .B(n30612), .Z(n30591) );
  NANDN U31968 ( .A(n30568), .B(n30567), .Z(n30572) );
  NANDN U31969 ( .A(n30570), .B(n30569), .Z(n30571) );
  AND U31970 ( .A(n30572), .B(n30571), .Z(n30590) );
  XNOR U31971 ( .A(n30591), .B(n30590), .Z(n30592) );
  NANDN U31972 ( .A(n30574), .B(n30573), .Z(n30578) );
  NAND U31973 ( .A(n30576), .B(n30575), .Z(n30577) );
  NAND U31974 ( .A(n30578), .B(n30577), .Z(n30593) );
  XNOR U31975 ( .A(n30592), .B(n30593), .Z(n30584) );
  XNOR U31976 ( .A(n30585), .B(n30584), .Z(n30586) );
  XNOR U31977 ( .A(n30587), .B(n30586), .Z(n30616) );
  XNOR U31978 ( .A(sreg[1732]), .B(n30616), .Z(n30618) );
  NANDN U31979 ( .A(sreg[1731]), .B(n30579), .Z(n30583) );
  NAND U31980 ( .A(n30581), .B(n30580), .Z(n30582) );
  NAND U31981 ( .A(n30583), .B(n30582), .Z(n30617) );
  XNOR U31982 ( .A(n30618), .B(n30617), .Z(c[1732]) );
  NANDN U31983 ( .A(n30585), .B(n30584), .Z(n30589) );
  NANDN U31984 ( .A(n30587), .B(n30586), .Z(n30588) );
  AND U31985 ( .A(n30589), .B(n30588), .Z(n30624) );
  NANDN U31986 ( .A(n30591), .B(n30590), .Z(n30595) );
  NANDN U31987 ( .A(n30593), .B(n30592), .Z(n30594) );
  AND U31988 ( .A(n30595), .B(n30594), .Z(n30622) );
  NAND U31989 ( .A(n42143), .B(n30596), .Z(n30598) );
  XNOR U31990 ( .A(a[711]), .B(n4173), .Z(n30633) );
  NAND U31991 ( .A(n42144), .B(n30633), .Z(n30597) );
  AND U31992 ( .A(n30598), .B(n30597), .Z(n30648) );
  XOR U31993 ( .A(a[715]), .B(n42012), .Z(n30636) );
  XNOR U31994 ( .A(n30648), .B(n30647), .Z(n30650) );
  AND U31995 ( .A(a[717]), .B(b[0]), .Z(n30600) );
  XNOR U31996 ( .A(n30600), .B(n4071), .Z(n30602) );
  NANDN U31997 ( .A(b[0]), .B(a[716]), .Z(n30601) );
  NAND U31998 ( .A(n30602), .B(n30601), .Z(n30644) );
  XOR U31999 ( .A(a[713]), .B(n42085), .Z(n30640) );
  AND U32000 ( .A(a[709]), .B(b[7]), .Z(n30641) );
  XNOR U32001 ( .A(n30642), .B(n30641), .Z(n30643) );
  XNOR U32002 ( .A(n30644), .B(n30643), .Z(n30649) );
  XOR U32003 ( .A(n30650), .B(n30649), .Z(n30628) );
  NANDN U32004 ( .A(n30605), .B(n30604), .Z(n30609) );
  NANDN U32005 ( .A(n30607), .B(n30606), .Z(n30608) );
  AND U32006 ( .A(n30609), .B(n30608), .Z(n30627) );
  XNOR U32007 ( .A(n30628), .B(n30627), .Z(n30629) );
  NANDN U32008 ( .A(n30611), .B(n30610), .Z(n30615) );
  NAND U32009 ( .A(n30613), .B(n30612), .Z(n30614) );
  NAND U32010 ( .A(n30615), .B(n30614), .Z(n30630) );
  XNOR U32011 ( .A(n30629), .B(n30630), .Z(n30621) );
  XNOR U32012 ( .A(n30622), .B(n30621), .Z(n30623) );
  XNOR U32013 ( .A(n30624), .B(n30623), .Z(n30653) );
  XNOR U32014 ( .A(sreg[1733]), .B(n30653), .Z(n30655) );
  NANDN U32015 ( .A(sreg[1732]), .B(n30616), .Z(n30620) );
  NAND U32016 ( .A(n30618), .B(n30617), .Z(n30619) );
  NAND U32017 ( .A(n30620), .B(n30619), .Z(n30654) );
  XNOR U32018 ( .A(n30655), .B(n30654), .Z(c[1733]) );
  NANDN U32019 ( .A(n30622), .B(n30621), .Z(n30626) );
  NANDN U32020 ( .A(n30624), .B(n30623), .Z(n30625) );
  AND U32021 ( .A(n30626), .B(n30625), .Z(n30661) );
  NANDN U32022 ( .A(n30628), .B(n30627), .Z(n30632) );
  NANDN U32023 ( .A(n30630), .B(n30629), .Z(n30631) );
  AND U32024 ( .A(n30632), .B(n30631), .Z(n30659) );
  NAND U32025 ( .A(n42143), .B(n30633), .Z(n30635) );
  XNOR U32026 ( .A(a[712]), .B(n4173), .Z(n30670) );
  NAND U32027 ( .A(n42144), .B(n30670), .Z(n30634) );
  AND U32028 ( .A(n30635), .B(n30634), .Z(n30685) );
  XOR U32029 ( .A(a[716]), .B(n42012), .Z(n30673) );
  XNOR U32030 ( .A(n30685), .B(n30684), .Z(n30687) );
  AND U32031 ( .A(a[718]), .B(b[0]), .Z(n30637) );
  XNOR U32032 ( .A(n30637), .B(n4071), .Z(n30639) );
  NANDN U32033 ( .A(b[0]), .B(a[717]), .Z(n30638) );
  NAND U32034 ( .A(n30639), .B(n30638), .Z(n30681) );
  XOR U32035 ( .A(a[714]), .B(n42085), .Z(n30677) );
  AND U32036 ( .A(a[710]), .B(b[7]), .Z(n30678) );
  XNOR U32037 ( .A(n30679), .B(n30678), .Z(n30680) );
  XNOR U32038 ( .A(n30681), .B(n30680), .Z(n30686) );
  XOR U32039 ( .A(n30687), .B(n30686), .Z(n30665) );
  NANDN U32040 ( .A(n30642), .B(n30641), .Z(n30646) );
  NANDN U32041 ( .A(n30644), .B(n30643), .Z(n30645) );
  AND U32042 ( .A(n30646), .B(n30645), .Z(n30664) );
  XNOR U32043 ( .A(n30665), .B(n30664), .Z(n30666) );
  NANDN U32044 ( .A(n30648), .B(n30647), .Z(n30652) );
  NAND U32045 ( .A(n30650), .B(n30649), .Z(n30651) );
  NAND U32046 ( .A(n30652), .B(n30651), .Z(n30667) );
  XNOR U32047 ( .A(n30666), .B(n30667), .Z(n30658) );
  XNOR U32048 ( .A(n30659), .B(n30658), .Z(n30660) );
  XNOR U32049 ( .A(n30661), .B(n30660), .Z(n30690) );
  XNOR U32050 ( .A(sreg[1734]), .B(n30690), .Z(n30692) );
  NANDN U32051 ( .A(sreg[1733]), .B(n30653), .Z(n30657) );
  NAND U32052 ( .A(n30655), .B(n30654), .Z(n30656) );
  NAND U32053 ( .A(n30657), .B(n30656), .Z(n30691) );
  XNOR U32054 ( .A(n30692), .B(n30691), .Z(c[1734]) );
  NANDN U32055 ( .A(n30659), .B(n30658), .Z(n30663) );
  NANDN U32056 ( .A(n30661), .B(n30660), .Z(n30662) );
  AND U32057 ( .A(n30663), .B(n30662), .Z(n30698) );
  NANDN U32058 ( .A(n30665), .B(n30664), .Z(n30669) );
  NANDN U32059 ( .A(n30667), .B(n30666), .Z(n30668) );
  AND U32060 ( .A(n30669), .B(n30668), .Z(n30696) );
  NAND U32061 ( .A(n42143), .B(n30670), .Z(n30672) );
  XNOR U32062 ( .A(a[713]), .B(n4173), .Z(n30707) );
  NAND U32063 ( .A(n42144), .B(n30707), .Z(n30671) );
  AND U32064 ( .A(n30672), .B(n30671), .Z(n30722) );
  XOR U32065 ( .A(a[717]), .B(n42012), .Z(n30710) );
  XNOR U32066 ( .A(n30722), .B(n30721), .Z(n30724) );
  AND U32067 ( .A(a[719]), .B(b[0]), .Z(n30674) );
  XNOR U32068 ( .A(n30674), .B(n4071), .Z(n30676) );
  NANDN U32069 ( .A(b[0]), .B(a[718]), .Z(n30675) );
  NAND U32070 ( .A(n30676), .B(n30675), .Z(n30718) );
  XOR U32071 ( .A(a[715]), .B(n42085), .Z(n30711) );
  AND U32072 ( .A(a[711]), .B(b[7]), .Z(n30715) );
  XNOR U32073 ( .A(n30716), .B(n30715), .Z(n30717) );
  XNOR U32074 ( .A(n30718), .B(n30717), .Z(n30723) );
  XOR U32075 ( .A(n30724), .B(n30723), .Z(n30702) );
  NANDN U32076 ( .A(n30679), .B(n30678), .Z(n30683) );
  NANDN U32077 ( .A(n30681), .B(n30680), .Z(n30682) );
  AND U32078 ( .A(n30683), .B(n30682), .Z(n30701) );
  XNOR U32079 ( .A(n30702), .B(n30701), .Z(n30703) );
  NANDN U32080 ( .A(n30685), .B(n30684), .Z(n30689) );
  NAND U32081 ( .A(n30687), .B(n30686), .Z(n30688) );
  NAND U32082 ( .A(n30689), .B(n30688), .Z(n30704) );
  XNOR U32083 ( .A(n30703), .B(n30704), .Z(n30695) );
  XNOR U32084 ( .A(n30696), .B(n30695), .Z(n30697) );
  XNOR U32085 ( .A(n30698), .B(n30697), .Z(n30727) );
  XNOR U32086 ( .A(sreg[1735]), .B(n30727), .Z(n30729) );
  NANDN U32087 ( .A(sreg[1734]), .B(n30690), .Z(n30694) );
  NAND U32088 ( .A(n30692), .B(n30691), .Z(n30693) );
  NAND U32089 ( .A(n30694), .B(n30693), .Z(n30728) );
  XNOR U32090 ( .A(n30729), .B(n30728), .Z(c[1735]) );
  NANDN U32091 ( .A(n30696), .B(n30695), .Z(n30700) );
  NANDN U32092 ( .A(n30698), .B(n30697), .Z(n30699) );
  AND U32093 ( .A(n30700), .B(n30699), .Z(n30735) );
  NANDN U32094 ( .A(n30702), .B(n30701), .Z(n30706) );
  NANDN U32095 ( .A(n30704), .B(n30703), .Z(n30705) );
  AND U32096 ( .A(n30706), .B(n30705), .Z(n30733) );
  NAND U32097 ( .A(n42143), .B(n30707), .Z(n30709) );
  XNOR U32098 ( .A(a[714]), .B(n4173), .Z(n30744) );
  NAND U32099 ( .A(n42144), .B(n30744), .Z(n30708) );
  AND U32100 ( .A(n30709), .B(n30708), .Z(n30759) );
  XOR U32101 ( .A(a[718]), .B(n42012), .Z(n30747) );
  XNOR U32102 ( .A(n30759), .B(n30758), .Z(n30761) );
  XOR U32103 ( .A(a[716]), .B(n42085), .Z(n30748) );
  AND U32104 ( .A(a[712]), .B(b[7]), .Z(n30752) );
  XNOR U32105 ( .A(n30753), .B(n30752), .Z(n30754) );
  AND U32106 ( .A(a[720]), .B(b[0]), .Z(n30712) );
  XNOR U32107 ( .A(n30712), .B(n4071), .Z(n30714) );
  NANDN U32108 ( .A(b[0]), .B(a[719]), .Z(n30713) );
  NAND U32109 ( .A(n30714), .B(n30713), .Z(n30755) );
  XNOR U32110 ( .A(n30754), .B(n30755), .Z(n30760) );
  XOR U32111 ( .A(n30761), .B(n30760), .Z(n30739) );
  NANDN U32112 ( .A(n30716), .B(n30715), .Z(n30720) );
  NANDN U32113 ( .A(n30718), .B(n30717), .Z(n30719) );
  AND U32114 ( .A(n30720), .B(n30719), .Z(n30738) );
  XNOR U32115 ( .A(n30739), .B(n30738), .Z(n30740) );
  NANDN U32116 ( .A(n30722), .B(n30721), .Z(n30726) );
  NAND U32117 ( .A(n30724), .B(n30723), .Z(n30725) );
  NAND U32118 ( .A(n30726), .B(n30725), .Z(n30741) );
  XNOR U32119 ( .A(n30740), .B(n30741), .Z(n30732) );
  XNOR U32120 ( .A(n30733), .B(n30732), .Z(n30734) );
  XNOR U32121 ( .A(n30735), .B(n30734), .Z(n30764) );
  XNOR U32122 ( .A(sreg[1736]), .B(n30764), .Z(n30766) );
  NANDN U32123 ( .A(sreg[1735]), .B(n30727), .Z(n30731) );
  NAND U32124 ( .A(n30729), .B(n30728), .Z(n30730) );
  NAND U32125 ( .A(n30731), .B(n30730), .Z(n30765) );
  XNOR U32126 ( .A(n30766), .B(n30765), .Z(c[1736]) );
  NANDN U32127 ( .A(n30733), .B(n30732), .Z(n30737) );
  NANDN U32128 ( .A(n30735), .B(n30734), .Z(n30736) );
  AND U32129 ( .A(n30737), .B(n30736), .Z(n30772) );
  NANDN U32130 ( .A(n30739), .B(n30738), .Z(n30743) );
  NANDN U32131 ( .A(n30741), .B(n30740), .Z(n30742) );
  AND U32132 ( .A(n30743), .B(n30742), .Z(n30770) );
  NAND U32133 ( .A(n42143), .B(n30744), .Z(n30746) );
  XNOR U32134 ( .A(a[715]), .B(n4174), .Z(n30781) );
  NAND U32135 ( .A(n42144), .B(n30781), .Z(n30745) );
  AND U32136 ( .A(n30746), .B(n30745), .Z(n30796) );
  XOR U32137 ( .A(a[719]), .B(n42012), .Z(n30784) );
  XNOR U32138 ( .A(n30796), .B(n30795), .Z(n30798) );
  XOR U32139 ( .A(a[717]), .B(n42085), .Z(n30788) );
  AND U32140 ( .A(a[713]), .B(b[7]), .Z(n30789) );
  XNOR U32141 ( .A(n30790), .B(n30789), .Z(n30791) );
  AND U32142 ( .A(a[721]), .B(b[0]), .Z(n30749) );
  XNOR U32143 ( .A(n30749), .B(n4071), .Z(n30751) );
  NANDN U32144 ( .A(b[0]), .B(a[720]), .Z(n30750) );
  NAND U32145 ( .A(n30751), .B(n30750), .Z(n30792) );
  XNOR U32146 ( .A(n30791), .B(n30792), .Z(n30797) );
  XOR U32147 ( .A(n30798), .B(n30797), .Z(n30776) );
  NANDN U32148 ( .A(n30753), .B(n30752), .Z(n30757) );
  NANDN U32149 ( .A(n30755), .B(n30754), .Z(n30756) );
  AND U32150 ( .A(n30757), .B(n30756), .Z(n30775) );
  XNOR U32151 ( .A(n30776), .B(n30775), .Z(n30777) );
  NANDN U32152 ( .A(n30759), .B(n30758), .Z(n30763) );
  NAND U32153 ( .A(n30761), .B(n30760), .Z(n30762) );
  NAND U32154 ( .A(n30763), .B(n30762), .Z(n30778) );
  XNOR U32155 ( .A(n30777), .B(n30778), .Z(n30769) );
  XNOR U32156 ( .A(n30770), .B(n30769), .Z(n30771) );
  XNOR U32157 ( .A(n30772), .B(n30771), .Z(n30801) );
  XNOR U32158 ( .A(sreg[1737]), .B(n30801), .Z(n30803) );
  NANDN U32159 ( .A(sreg[1736]), .B(n30764), .Z(n30768) );
  NAND U32160 ( .A(n30766), .B(n30765), .Z(n30767) );
  NAND U32161 ( .A(n30768), .B(n30767), .Z(n30802) );
  XNOR U32162 ( .A(n30803), .B(n30802), .Z(c[1737]) );
  NANDN U32163 ( .A(n30770), .B(n30769), .Z(n30774) );
  NANDN U32164 ( .A(n30772), .B(n30771), .Z(n30773) );
  AND U32165 ( .A(n30774), .B(n30773), .Z(n30809) );
  NANDN U32166 ( .A(n30776), .B(n30775), .Z(n30780) );
  NANDN U32167 ( .A(n30778), .B(n30777), .Z(n30779) );
  AND U32168 ( .A(n30780), .B(n30779), .Z(n30807) );
  NAND U32169 ( .A(n42143), .B(n30781), .Z(n30783) );
  XNOR U32170 ( .A(a[716]), .B(n4174), .Z(n30818) );
  NAND U32171 ( .A(n42144), .B(n30818), .Z(n30782) );
  AND U32172 ( .A(n30783), .B(n30782), .Z(n30833) );
  XOR U32173 ( .A(a[720]), .B(n42012), .Z(n30821) );
  XNOR U32174 ( .A(n30833), .B(n30832), .Z(n30835) );
  AND U32175 ( .A(a[722]), .B(b[0]), .Z(n30785) );
  XNOR U32176 ( .A(n30785), .B(n4071), .Z(n30787) );
  NANDN U32177 ( .A(b[0]), .B(a[721]), .Z(n30786) );
  NAND U32178 ( .A(n30787), .B(n30786), .Z(n30829) );
  XOR U32179 ( .A(a[718]), .B(n42085), .Z(n30822) );
  AND U32180 ( .A(a[714]), .B(b[7]), .Z(n30826) );
  XNOR U32181 ( .A(n30827), .B(n30826), .Z(n30828) );
  XNOR U32182 ( .A(n30829), .B(n30828), .Z(n30834) );
  XOR U32183 ( .A(n30835), .B(n30834), .Z(n30813) );
  NANDN U32184 ( .A(n30790), .B(n30789), .Z(n30794) );
  NANDN U32185 ( .A(n30792), .B(n30791), .Z(n30793) );
  AND U32186 ( .A(n30794), .B(n30793), .Z(n30812) );
  XNOR U32187 ( .A(n30813), .B(n30812), .Z(n30814) );
  NANDN U32188 ( .A(n30796), .B(n30795), .Z(n30800) );
  NAND U32189 ( .A(n30798), .B(n30797), .Z(n30799) );
  NAND U32190 ( .A(n30800), .B(n30799), .Z(n30815) );
  XNOR U32191 ( .A(n30814), .B(n30815), .Z(n30806) );
  XNOR U32192 ( .A(n30807), .B(n30806), .Z(n30808) );
  XNOR U32193 ( .A(n30809), .B(n30808), .Z(n30838) );
  XNOR U32194 ( .A(sreg[1738]), .B(n30838), .Z(n30840) );
  NANDN U32195 ( .A(sreg[1737]), .B(n30801), .Z(n30805) );
  NAND U32196 ( .A(n30803), .B(n30802), .Z(n30804) );
  NAND U32197 ( .A(n30805), .B(n30804), .Z(n30839) );
  XNOR U32198 ( .A(n30840), .B(n30839), .Z(c[1738]) );
  NANDN U32199 ( .A(n30807), .B(n30806), .Z(n30811) );
  NANDN U32200 ( .A(n30809), .B(n30808), .Z(n30810) );
  AND U32201 ( .A(n30811), .B(n30810), .Z(n30846) );
  NANDN U32202 ( .A(n30813), .B(n30812), .Z(n30817) );
  NANDN U32203 ( .A(n30815), .B(n30814), .Z(n30816) );
  AND U32204 ( .A(n30817), .B(n30816), .Z(n30844) );
  NAND U32205 ( .A(n42143), .B(n30818), .Z(n30820) );
  XNOR U32206 ( .A(a[717]), .B(n4174), .Z(n30855) );
  NAND U32207 ( .A(n42144), .B(n30855), .Z(n30819) );
  AND U32208 ( .A(n30820), .B(n30819), .Z(n30870) );
  XOR U32209 ( .A(a[721]), .B(n42012), .Z(n30858) );
  XNOR U32210 ( .A(n30870), .B(n30869), .Z(n30872) );
  XOR U32211 ( .A(a[719]), .B(n42085), .Z(n30862) );
  AND U32212 ( .A(a[715]), .B(b[7]), .Z(n30863) );
  XNOR U32213 ( .A(n30864), .B(n30863), .Z(n30865) );
  AND U32214 ( .A(a[723]), .B(b[0]), .Z(n30823) );
  XNOR U32215 ( .A(n30823), .B(n4071), .Z(n30825) );
  NANDN U32216 ( .A(b[0]), .B(a[722]), .Z(n30824) );
  NAND U32217 ( .A(n30825), .B(n30824), .Z(n30866) );
  XNOR U32218 ( .A(n30865), .B(n30866), .Z(n30871) );
  XOR U32219 ( .A(n30872), .B(n30871), .Z(n30850) );
  NANDN U32220 ( .A(n30827), .B(n30826), .Z(n30831) );
  NANDN U32221 ( .A(n30829), .B(n30828), .Z(n30830) );
  AND U32222 ( .A(n30831), .B(n30830), .Z(n30849) );
  XNOR U32223 ( .A(n30850), .B(n30849), .Z(n30851) );
  NANDN U32224 ( .A(n30833), .B(n30832), .Z(n30837) );
  NAND U32225 ( .A(n30835), .B(n30834), .Z(n30836) );
  NAND U32226 ( .A(n30837), .B(n30836), .Z(n30852) );
  XNOR U32227 ( .A(n30851), .B(n30852), .Z(n30843) );
  XNOR U32228 ( .A(n30844), .B(n30843), .Z(n30845) );
  XNOR U32229 ( .A(n30846), .B(n30845), .Z(n30875) );
  XNOR U32230 ( .A(sreg[1739]), .B(n30875), .Z(n30877) );
  NANDN U32231 ( .A(sreg[1738]), .B(n30838), .Z(n30842) );
  NAND U32232 ( .A(n30840), .B(n30839), .Z(n30841) );
  NAND U32233 ( .A(n30842), .B(n30841), .Z(n30876) );
  XNOR U32234 ( .A(n30877), .B(n30876), .Z(c[1739]) );
  NANDN U32235 ( .A(n30844), .B(n30843), .Z(n30848) );
  NANDN U32236 ( .A(n30846), .B(n30845), .Z(n30847) );
  AND U32237 ( .A(n30848), .B(n30847), .Z(n30883) );
  NANDN U32238 ( .A(n30850), .B(n30849), .Z(n30854) );
  NANDN U32239 ( .A(n30852), .B(n30851), .Z(n30853) );
  AND U32240 ( .A(n30854), .B(n30853), .Z(n30881) );
  NAND U32241 ( .A(n42143), .B(n30855), .Z(n30857) );
  XNOR U32242 ( .A(a[718]), .B(n4174), .Z(n30892) );
  NAND U32243 ( .A(n42144), .B(n30892), .Z(n30856) );
  AND U32244 ( .A(n30857), .B(n30856), .Z(n30907) );
  XOR U32245 ( .A(a[722]), .B(n42012), .Z(n30895) );
  XNOR U32246 ( .A(n30907), .B(n30906), .Z(n30909) );
  AND U32247 ( .A(a[724]), .B(b[0]), .Z(n30859) );
  XNOR U32248 ( .A(n30859), .B(n4071), .Z(n30861) );
  NANDN U32249 ( .A(b[0]), .B(a[723]), .Z(n30860) );
  NAND U32250 ( .A(n30861), .B(n30860), .Z(n30903) );
  XOR U32251 ( .A(a[720]), .B(n42085), .Z(n30899) );
  AND U32252 ( .A(a[716]), .B(b[7]), .Z(n30900) );
  XNOR U32253 ( .A(n30901), .B(n30900), .Z(n30902) );
  XNOR U32254 ( .A(n30903), .B(n30902), .Z(n30908) );
  XOR U32255 ( .A(n30909), .B(n30908), .Z(n30887) );
  NANDN U32256 ( .A(n30864), .B(n30863), .Z(n30868) );
  NANDN U32257 ( .A(n30866), .B(n30865), .Z(n30867) );
  AND U32258 ( .A(n30868), .B(n30867), .Z(n30886) );
  XNOR U32259 ( .A(n30887), .B(n30886), .Z(n30888) );
  NANDN U32260 ( .A(n30870), .B(n30869), .Z(n30874) );
  NAND U32261 ( .A(n30872), .B(n30871), .Z(n30873) );
  NAND U32262 ( .A(n30874), .B(n30873), .Z(n30889) );
  XNOR U32263 ( .A(n30888), .B(n30889), .Z(n30880) );
  XNOR U32264 ( .A(n30881), .B(n30880), .Z(n30882) );
  XNOR U32265 ( .A(n30883), .B(n30882), .Z(n30912) );
  XNOR U32266 ( .A(sreg[1740]), .B(n30912), .Z(n30914) );
  NANDN U32267 ( .A(sreg[1739]), .B(n30875), .Z(n30879) );
  NAND U32268 ( .A(n30877), .B(n30876), .Z(n30878) );
  NAND U32269 ( .A(n30879), .B(n30878), .Z(n30913) );
  XNOR U32270 ( .A(n30914), .B(n30913), .Z(c[1740]) );
  NANDN U32271 ( .A(n30881), .B(n30880), .Z(n30885) );
  NANDN U32272 ( .A(n30883), .B(n30882), .Z(n30884) );
  AND U32273 ( .A(n30885), .B(n30884), .Z(n30920) );
  NANDN U32274 ( .A(n30887), .B(n30886), .Z(n30891) );
  NANDN U32275 ( .A(n30889), .B(n30888), .Z(n30890) );
  AND U32276 ( .A(n30891), .B(n30890), .Z(n30918) );
  NAND U32277 ( .A(n42143), .B(n30892), .Z(n30894) );
  XNOR U32278 ( .A(a[719]), .B(n4174), .Z(n30929) );
  NAND U32279 ( .A(n42144), .B(n30929), .Z(n30893) );
  AND U32280 ( .A(n30894), .B(n30893), .Z(n30944) );
  XOR U32281 ( .A(a[723]), .B(n42012), .Z(n30932) );
  XNOR U32282 ( .A(n30944), .B(n30943), .Z(n30946) );
  AND U32283 ( .A(a[725]), .B(b[0]), .Z(n30896) );
  XNOR U32284 ( .A(n30896), .B(n4071), .Z(n30898) );
  NANDN U32285 ( .A(b[0]), .B(a[724]), .Z(n30897) );
  NAND U32286 ( .A(n30898), .B(n30897), .Z(n30940) );
  XOR U32287 ( .A(a[721]), .B(n42085), .Z(n30936) );
  AND U32288 ( .A(a[717]), .B(b[7]), .Z(n30937) );
  XNOR U32289 ( .A(n30938), .B(n30937), .Z(n30939) );
  XNOR U32290 ( .A(n30940), .B(n30939), .Z(n30945) );
  XOR U32291 ( .A(n30946), .B(n30945), .Z(n30924) );
  NANDN U32292 ( .A(n30901), .B(n30900), .Z(n30905) );
  NANDN U32293 ( .A(n30903), .B(n30902), .Z(n30904) );
  AND U32294 ( .A(n30905), .B(n30904), .Z(n30923) );
  XNOR U32295 ( .A(n30924), .B(n30923), .Z(n30925) );
  NANDN U32296 ( .A(n30907), .B(n30906), .Z(n30911) );
  NAND U32297 ( .A(n30909), .B(n30908), .Z(n30910) );
  NAND U32298 ( .A(n30911), .B(n30910), .Z(n30926) );
  XNOR U32299 ( .A(n30925), .B(n30926), .Z(n30917) );
  XNOR U32300 ( .A(n30918), .B(n30917), .Z(n30919) );
  XNOR U32301 ( .A(n30920), .B(n30919), .Z(n30949) );
  XNOR U32302 ( .A(sreg[1741]), .B(n30949), .Z(n30951) );
  NANDN U32303 ( .A(sreg[1740]), .B(n30912), .Z(n30916) );
  NAND U32304 ( .A(n30914), .B(n30913), .Z(n30915) );
  NAND U32305 ( .A(n30916), .B(n30915), .Z(n30950) );
  XNOR U32306 ( .A(n30951), .B(n30950), .Z(c[1741]) );
  NANDN U32307 ( .A(n30918), .B(n30917), .Z(n30922) );
  NANDN U32308 ( .A(n30920), .B(n30919), .Z(n30921) );
  AND U32309 ( .A(n30922), .B(n30921), .Z(n30957) );
  NANDN U32310 ( .A(n30924), .B(n30923), .Z(n30928) );
  NANDN U32311 ( .A(n30926), .B(n30925), .Z(n30927) );
  AND U32312 ( .A(n30928), .B(n30927), .Z(n30955) );
  NAND U32313 ( .A(n42143), .B(n30929), .Z(n30931) );
  XNOR U32314 ( .A(a[720]), .B(n4174), .Z(n30966) );
  NAND U32315 ( .A(n42144), .B(n30966), .Z(n30930) );
  AND U32316 ( .A(n30931), .B(n30930), .Z(n30981) );
  XOR U32317 ( .A(a[724]), .B(n42012), .Z(n30969) );
  XNOR U32318 ( .A(n30981), .B(n30980), .Z(n30983) );
  AND U32319 ( .A(a[726]), .B(b[0]), .Z(n30933) );
  XNOR U32320 ( .A(n30933), .B(n4071), .Z(n30935) );
  NANDN U32321 ( .A(b[0]), .B(a[725]), .Z(n30934) );
  NAND U32322 ( .A(n30935), .B(n30934), .Z(n30977) );
  XOR U32323 ( .A(a[722]), .B(n42085), .Z(n30970) );
  AND U32324 ( .A(a[718]), .B(b[7]), .Z(n30974) );
  XNOR U32325 ( .A(n30975), .B(n30974), .Z(n30976) );
  XNOR U32326 ( .A(n30977), .B(n30976), .Z(n30982) );
  XOR U32327 ( .A(n30983), .B(n30982), .Z(n30961) );
  NANDN U32328 ( .A(n30938), .B(n30937), .Z(n30942) );
  NANDN U32329 ( .A(n30940), .B(n30939), .Z(n30941) );
  AND U32330 ( .A(n30942), .B(n30941), .Z(n30960) );
  XNOR U32331 ( .A(n30961), .B(n30960), .Z(n30962) );
  NANDN U32332 ( .A(n30944), .B(n30943), .Z(n30948) );
  NAND U32333 ( .A(n30946), .B(n30945), .Z(n30947) );
  NAND U32334 ( .A(n30948), .B(n30947), .Z(n30963) );
  XNOR U32335 ( .A(n30962), .B(n30963), .Z(n30954) );
  XNOR U32336 ( .A(n30955), .B(n30954), .Z(n30956) );
  XNOR U32337 ( .A(n30957), .B(n30956), .Z(n30986) );
  XNOR U32338 ( .A(sreg[1742]), .B(n30986), .Z(n30988) );
  NANDN U32339 ( .A(sreg[1741]), .B(n30949), .Z(n30953) );
  NAND U32340 ( .A(n30951), .B(n30950), .Z(n30952) );
  NAND U32341 ( .A(n30953), .B(n30952), .Z(n30987) );
  XNOR U32342 ( .A(n30988), .B(n30987), .Z(c[1742]) );
  NANDN U32343 ( .A(n30955), .B(n30954), .Z(n30959) );
  NANDN U32344 ( .A(n30957), .B(n30956), .Z(n30958) );
  AND U32345 ( .A(n30959), .B(n30958), .Z(n30994) );
  NANDN U32346 ( .A(n30961), .B(n30960), .Z(n30965) );
  NANDN U32347 ( .A(n30963), .B(n30962), .Z(n30964) );
  AND U32348 ( .A(n30965), .B(n30964), .Z(n30992) );
  NAND U32349 ( .A(n42143), .B(n30966), .Z(n30968) );
  XNOR U32350 ( .A(a[721]), .B(n4174), .Z(n31003) );
  NAND U32351 ( .A(n42144), .B(n31003), .Z(n30967) );
  AND U32352 ( .A(n30968), .B(n30967), .Z(n31018) );
  XOR U32353 ( .A(a[725]), .B(n42012), .Z(n31006) );
  XNOR U32354 ( .A(n31018), .B(n31017), .Z(n31020) );
  XOR U32355 ( .A(a[723]), .B(n42085), .Z(n31010) );
  AND U32356 ( .A(a[719]), .B(b[7]), .Z(n31011) );
  XNOR U32357 ( .A(n31012), .B(n31011), .Z(n31013) );
  AND U32358 ( .A(a[727]), .B(b[0]), .Z(n30971) );
  XNOR U32359 ( .A(n30971), .B(n4071), .Z(n30973) );
  NANDN U32360 ( .A(b[0]), .B(a[726]), .Z(n30972) );
  NAND U32361 ( .A(n30973), .B(n30972), .Z(n31014) );
  XNOR U32362 ( .A(n31013), .B(n31014), .Z(n31019) );
  XOR U32363 ( .A(n31020), .B(n31019), .Z(n30998) );
  NANDN U32364 ( .A(n30975), .B(n30974), .Z(n30979) );
  NANDN U32365 ( .A(n30977), .B(n30976), .Z(n30978) );
  AND U32366 ( .A(n30979), .B(n30978), .Z(n30997) );
  XNOR U32367 ( .A(n30998), .B(n30997), .Z(n30999) );
  NANDN U32368 ( .A(n30981), .B(n30980), .Z(n30985) );
  NAND U32369 ( .A(n30983), .B(n30982), .Z(n30984) );
  NAND U32370 ( .A(n30985), .B(n30984), .Z(n31000) );
  XNOR U32371 ( .A(n30999), .B(n31000), .Z(n30991) );
  XNOR U32372 ( .A(n30992), .B(n30991), .Z(n30993) );
  XNOR U32373 ( .A(n30994), .B(n30993), .Z(n31023) );
  XNOR U32374 ( .A(sreg[1743]), .B(n31023), .Z(n31025) );
  NANDN U32375 ( .A(sreg[1742]), .B(n30986), .Z(n30990) );
  NAND U32376 ( .A(n30988), .B(n30987), .Z(n30989) );
  NAND U32377 ( .A(n30990), .B(n30989), .Z(n31024) );
  XNOR U32378 ( .A(n31025), .B(n31024), .Z(c[1743]) );
  NANDN U32379 ( .A(n30992), .B(n30991), .Z(n30996) );
  NANDN U32380 ( .A(n30994), .B(n30993), .Z(n30995) );
  AND U32381 ( .A(n30996), .B(n30995), .Z(n31031) );
  NANDN U32382 ( .A(n30998), .B(n30997), .Z(n31002) );
  NANDN U32383 ( .A(n31000), .B(n30999), .Z(n31001) );
  AND U32384 ( .A(n31002), .B(n31001), .Z(n31029) );
  NAND U32385 ( .A(n42143), .B(n31003), .Z(n31005) );
  XNOR U32386 ( .A(a[722]), .B(n4175), .Z(n31040) );
  NAND U32387 ( .A(n42144), .B(n31040), .Z(n31004) );
  AND U32388 ( .A(n31005), .B(n31004), .Z(n31055) );
  XOR U32389 ( .A(a[726]), .B(n42012), .Z(n31043) );
  XNOR U32390 ( .A(n31055), .B(n31054), .Z(n31057) );
  AND U32391 ( .A(a[728]), .B(b[0]), .Z(n31007) );
  XNOR U32392 ( .A(n31007), .B(n4071), .Z(n31009) );
  NANDN U32393 ( .A(b[0]), .B(a[727]), .Z(n31008) );
  NAND U32394 ( .A(n31009), .B(n31008), .Z(n31051) );
  XOR U32395 ( .A(a[724]), .B(n42085), .Z(n31047) );
  AND U32396 ( .A(a[720]), .B(b[7]), .Z(n31048) );
  XNOR U32397 ( .A(n31049), .B(n31048), .Z(n31050) );
  XNOR U32398 ( .A(n31051), .B(n31050), .Z(n31056) );
  XOR U32399 ( .A(n31057), .B(n31056), .Z(n31035) );
  NANDN U32400 ( .A(n31012), .B(n31011), .Z(n31016) );
  NANDN U32401 ( .A(n31014), .B(n31013), .Z(n31015) );
  AND U32402 ( .A(n31016), .B(n31015), .Z(n31034) );
  XNOR U32403 ( .A(n31035), .B(n31034), .Z(n31036) );
  NANDN U32404 ( .A(n31018), .B(n31017), .Z(n31022) );
  NAND U32405 ( .A(n31020), .B(n31019), .Z(n31021) );
  NAND U32406 ( .A(n31022), .B(n31021), .Z(n31037) );
  XNOR U32407 ( .A(n31036), .B(n31037), .Z(n31028) );
  XNOR U32408 ( .A(n31029), .B(n31028), .Z(n31030) );
  XNOR U32409 ( .A(n31031), .B(n31030), .Z(n31060) );
  XNOR U32410 ( .A(sreg[1744]), .B(n31060), .Z(n31062) );
  NANDN U32411 ( .A(sreg[1743]), .B(n31023), .Z(n31027) );
  NAND U32412 ( .A(n31025), .B(n31024), .Z(n31026) );
  NAND U32413 ( .A(n31027), .B(n31026), .Z(n31061) );
  XNOR U32414 ( .A(n31062), .B(n31061), .Z(c[1744]) );
  NANDN U32415 ( .A(n31029), .B(n31028), .Z(n31033) );
  NANDN U32416 ( .A(n31031), .B(n31030), .Z(n31032) );
  AND U32417 ( .A(n31033), .B(n31032), .Z(n31068) );
  NANDN U32418 ( .A(n31035), .B(n31034), .Z(n31039) );
  NANDN U32419 ( .A(n31037), .B(n31036), .Z(n31038) );
  AND U32420 ( .A(n31039), .B(n31038), .Z(n31066) );
  NAND U32421 ( .A(n42143), .B(n31040), .Z(n31042) );
  XNOR U32422 ( .A(a[723]), .B(n4175), .Z(n31077) );
  NAND U32423 ( .A(n42144), .B(n31077), .Z(n31041) );
  AND U32424 ( .A(n31042), .B(n31041), .Z(n31092) );
  XOR U32425 ( .A(a[727]), .B(n42012), .Z(n31080) );
  XNOR U32426 ( .A(n31092), .B(n31091), .Z(n31094) );
  AND U32427 ( .A(a[729]), .B(b[0]), .Z(n31044) );
  XNOR U32428 ( .A(n31044), .B(n4071), .Z(n31046) );
  NANDN U32429 ( .A(b[0]), .B(a[728]), .Z(n31045) );
  NAND U32430 ( .A(n31046), .B(n31045), .Z(n31088) );
  XOR U32431 ( .A(a[725]), .B(n42085), .Z(n31084) );
  AND U32432 ( .A(a[721]), .B(b[7]), .Z(n31085) );
  XNOR U32433 ( .A(n31086), .B(n31085), .Z(n31087) );
  XNOR U32434 ( .A(n31088), .B(n31087), .Z(n31093) );
  XOR U32435 ( .A(n31094), .B(n31093), .Z(n31072) );
  NANDN U32436 ( .A(n31049), .B(n31048), .Z(n31053) );
  NANDN U32437 ( .A(n31051), .B(n31050), .Z(n31052) );
  AND U32438 ( .A(n31053), .B(n31052), .Z(n31071) );
  XNOR U32439 ( .A(n31072), .B(n31071), .Z(n31073) );
  NANDN U32440 ( .A(n31055), .B(n31054), .Z(n31059) );
  NAND U32441 ( .A(n31057), .B(n31056), .Z(n31058) );
  NAND U32442 ( .A(n31059), .B(n31058), .Z(n31074) );
  XNOR U32443 ( .A(n31073), .B(n31074), .Z(n31065) );
  XNOR U32444 ( .A(n31066), .B(n31065), .Z(n31067) );
  XNOR U32445 ( .A(n31068), .B(n31067), .Z(n31097) );
  XNOR U32446 ( .A(sreg[1745]), .B(n31097), .Z(n31099) );
  NANDN U32447 ( .A(sreg[1744]), .B(n31060), .Z(n31064) );
  NAND U32448 ( .A(n31062), .B(n31061), .Z(n31063) );
  NAND U32449 ( .A(n31064), .B(n31063), .Z(n31098) );
  XNOR U32450 ( .A(n31099), .B(n31098), .Z(c[1745]) );
  NANDN U32451 ( .A(n31066), .B(n31065), .Z(n31070) );
  NANDN U32452 ( .A(n31068), .B(n31067), .Z(n31069) );
  AND U32453 ( .A(n31070), .B(n31069), .Z(n31105) );
  NANDN U32454 ( .A(n31072), .B(n31071), .Z(n31076) );
  NANDN U32455 ( .A(n31074), .B(n31073), .Z(n31075) );
  AND U32456 ( .A(n31076), .B(n31075), .Z(n31103) );
  NAND U32457 ( .A(n42143), .B(n31077), .Z(n31079) );
  XNOR U32458 ( .A(a[724]), .B(n4175), .Z(n31114) );
  NAND U32459 ( .A(n42144), .B(n31114), .Z(n31078) );
  AND U32460 ( .A(n31079), .B(n31078), .Z(n31129) );
  XOR U32461 ( .A(a[728]), .B(n42012), .Z(n31117) );
  XNOR U32462 ( .A(n31129), .B(n31128), .Z(n31131) );
  AND U32463 ( .A(a[730]), .B(b[0]), .Z(n31081) );
  XNOR U32464 ( .A(n31081), .B(n4071), .Z(n31083) );
  NANDN U32465 ( .A(b[0]), .B(a[729]), .Z(n31082) );
  NAND U32466 ( .A(n31083), .B(n31082), .Z(n31125) );
  XOR U32467 ( .A(a[726]), .B(n42085), .Z(n31121) );
  AND U32468 ( .A(a[722]), .B(b[7]), .Z(n31122) );
  XNOR U32469 ( .A(n31123), .B(n31122), .Z(n31124) );
  XNOR U32470 ( .A(n31125), .B(n31124), .Z(n31130) );
  XOR U32471 ( .A(n31131), .B(n31130), .Z(n31109) );
  NANDN U32472 ( .A(n31086), .B(n31085), .Z(n31090) );
  NANDN U32473 ( .A(n31088), .B(n31087), .Z(n31089) );
  AND U32474 ( .A(n31090), .B(n31089), .Z(n31108) );
  XNOR U32475 ( .A(n31109), .B(n31108), .Z(n31110) );
  NANDN U32476 ( .A(n31092), .B(n31091), .Z(n31096) );
  NAND U32477 ( .A(n31094), .B(n31093), .Z(n31095) );
  NAND U32478 ( .A(n31096), .B(n31095), .Z(n31111) );
  XNOR U32479 ( .A(n31110), .B(n31111), .Z(n31102) );
  XNOR U32480 ( .A(n31103), .B(n31102), .Z(n31104) );
  XNOR U32481 ( .A(n31105), .B(n31104), .Z(n31134) );
  XNOR U32482 ( .A(sreg[1746]), .B(n31134), .Z(n31136) );
  NANDN U32483 ( .A(sreg[1745]), .B(n31097), .Z(n31101) );
  NAND U32484 ( .A(n31099), .B(n31098), .Z(n31100) );
  NAND U32485 ( .A(n31101), .B(n31100), .Z(n31135) );
  XNOR U32486 ( .A(n31136), .B(n31135), .Z(c[1746]) );
  NANDN U32487 ( .A(n31103), .B(n31102), .Z(n31107) );
  NANDN U32488 ( .A(n31105), .B(n31104), .Z(n31106) );
  AND U32489 ( .A(n31107), .B(n31106), .Z(n31142) );
  NANDN U32490 ( .A(n31109), .B(n31108), .Z(n31113) );
  NANDN U32491 ( .A(n31111), .B(n31110), .Z(n31112) );
  AND U32492 ( .A(n31113), .B(n31112), .Z(n31140) );
  NAND U32493 ( .A(n42143), .B(n31114), .Z(n31116) );
  XNOR U32494 ( .A(a[725]), .B(n4175), .Z(n31151) );
  NAND U32495 ( .A(n42144), .B(n31151), .Z(n31115) );
  AND U32496 ( .A(n31116), .B(n31115), .Z(n31166) );
  XOR U32497 ( .A(a[729]), .B(n42012), .Z(n31154) );
  XNOR U32498 ( .A(n31166), .B(n31165), .Z(n31168) );
  AND U32499 ( .A(a[731]), .B(b[0]), .Z(n31118) );
  XNOR U32500 ( .A(n31118), .B(n4071), .Z(n31120) );
  NANDN U32501 ( .A(b[0]), .B(a[730]), .Z(n31119) );
  NAND U32502 ( .A(n31120), .B(n31119), .Z(n31162) );
  XOR U32503 ( .A(a[727]), .B(n42085), .Z(n31155) );
  AND U32504 ( .A(a[723]), .B(b[7]), .Z(n31159) );
  XNOR U32505 ( .A(n31160), .B(n31159), .Z(n31161) );
  XNOR U32506 ( .A(n31162), .B(n31161), .Z(n31167) );
  XOR U32507 ( .A(n31168), .B(n31167), .Z(n31146) );
  NANDN U32508 ( .A(n31123), .B(n31122), .Z(n31127) );
  NANDN U32509 ( .A(n31125), .B(n31124), .Z(n31126) );
  AND U32510 ( .A(n31127), .B(n31126), .Z(n31145) );
  XNOR U32511 ( .A(n31146), .B(n31145), .Z(n31147) );
  NANDN U32512 ( .A(n31129), .B(n31128), .Z(n31133) );
  NAND U32513 ( .A(n31131), .B(n31130), .Z(n31132) );
  NAND U32514 ( .A(n31133), .B(n31132), .Z(n31148) );
  XNOR U32515 ( .A(n31147), .B(n31148), .Z(n31139) );
  XNOR U32516 ( .A(n31140), .B(n31139), .Z(n31141) );
  XNOR U32517 ( .A(n31142), .B(n31141), .Z(n31171) );
  XNOR U32518 ( .A(sreg[1747]), .B(n31171), .Z(n31173) );
  NANDN U32519 ( .A(sreg[1746]), .B(n31134), .Z(n31138) );
  NAND U32520 ( .A(n31136), .B(n31135), .Z(n31137) );
  NAND U32521 ( .A(n31138), .B(n31137), .Z(n31172) );
  XNOR U32522 ( .A(n31173), .B(n31172), .Z(c[1747]) );
  NANDN U32523 ( .A(n31140), .B(n31139), .Z(n31144) );
  NANDN U32524 ( .A(n31142), .B(n31141), .Z(n31143) );
  AND U32525 ( .A(n31144), .B(n31143), .Z(n31179) );
  NANDN U32526 ( .A(n31146), .B(n31145), .Z(n31150) );
  NANDN U32527 ( .A(n31148), .B(n31147), .Z(n31149) );
  AND U32528 ( .A(n31150), .B(n31149), .Z(n31177) );
  NAND U32529 ( .A(n42143), .B(n31151), .Z(n31153) );
  XNOR U32530 ( .A(a[726]), .B(n4175), .Z(n31188) );
  NAND U32531 ( .A(n42144), .B(n31188), .Z(n31152) );
  AND U32532 ( .A(n31153), .B(n31152), .Z(n31203) );
  XOR U32533 ( .A(a[730]), .B(n42012), .Z(n31191) );
  XNOR U32534 ( .A(n31203), .B(n31202), .Z(n31205) );
  XOR U32535 ( .A(a[728]), .B(n42085), .Z(n31195) );
  AND U32536 ( .A(a[724]), .B(b[7]), .Z(n31196) );
  XNOR U32537 ( .A(n31197), .B(n31196), .Z(n31198) );
  AND U32538 ( .A(a[732]), .B(b[0]), .Z(n31156) );
  XNOR U32539 ( .A(n31156), .B(n4071), .Z(n31158) );
  NANDN U32540 ( .A(b[0]), .B(a[731]), .Z(n31157) );
  NAND U32541 ( .A(n31158), .B(n31157), .Z(n31199) );
  XNOR U32542 ( .A(n31198), .B(n31199), .Z(n31204) );
  XOR U32543 ( .A(n31205), .B(n31204), .Z(n31183) );
  NANDN U32544 ( .A(n31160), .B(n31159), .Z(n31164) );
  NANDN U32545 ( .A(n31162), .B(n31161), .Z(n31163) );
  AND U32546 ( .A(n31164), .B(n31163), .Z(n31182) );
  XNOR U32547 ( .A(n31183), .B(n31182), .Z(n31184) );
  NANDN U32548 ( .A(n31166), .B(n31165), .Z(n31170) );
  NAND U32549 ( .A(n31168), .B(n31167), .Z(n31169) );
  NAND U32550 ( .A(n31170), .B(n31169), .Z(n31185) );
  XNOR U32551 ( .A(n31184), .B(n31185), .Z(n31176) );
  XNOR U32552 ( .A(n31177), .B(n31176), .Z(n31178) );
  XNOR U32553 ( .A(n31179), .B(n31178), .Z(n31208) );
  XNOR U32554 ( .A(sreg[1748]), .B(n31208), .Z(n31210) );
  NANDN U32555 ( .A(sreg[1747]), .B(n31171), .Z(n31175) );
  NAND U32556 ( .A(n31173), .B(n31172), .Z(n31174) );
  NAND U32557 ( .A(n31175), .B(n31174), .Z(n31209) );
  XNOR U32558 ( .A(n31210), .B(n31209), .Z(c[1748]) );
  NANDN U32559 ( .A(n31177), .B(n31176), .Z(n31181) );
  NANDN U32560 ( .A(n31179), .B(n31178), .Z(n31180) );
  AND U32561 ( .A(n31181), .B(n31180), .Z(n31216) );
  NANDN U32562 ( .A(n31183), .B(n31182), .Z(n31187) );
  NANDN U32563 ( .A(n31185), .B(n31184), .Z(n31186) );
  AND U32564 ( .A(n31187), .B(n31186), .Z(n31214) );
  NAND U32565 ( .A(n42143), .B(n31188), .Z(n31190) );
  XNOR U32566 ( .A(a[727]), .B(n4175), .Z(n31225) );
  NAND U32567 ( .A(n42144), .B(n31225), .Z(n31189) );
  AND U32568 ( .A(n31190), .B(n31189), .Z(n31240) );
  XOR U32569 ( .A(a[731]), .B(n42012), .Z(n31228) );
  XNOR U32570 ( .A(n31240), .B(n31239), .Z(n31242) );
  AND U32571 ( .A(a[733]), .B(b[0]), .Z(n31192) );
  XNOR U32572 ( .A(n31192), .B(n4071), .Z(n31194) );
  NANDN U32573 ( .A(b[0]), .B(a[732]), .Z(n31193) );
  NAND U32574 ( .A(n31194), .B(n31193), .Z(n31236) );
  XOR U32575 ( .A(a[729]), .B(n42085), .Z(n31232) );
  AND U32576 ( .A(a[725]), .B(b[7]), .Z(n31233) );
  XNOR U32577 ( .A(n31234), .B(n31233), .Z(n31235) );
  XNOR U32578 ( .A(n31236), .B(n31235), .Z(n31241) );
  XOR U32579 ( .A(n31242), .B(n31241), .Z(n31220) );
  NANDN U32580 ( .A(n31197), .B(n31196), .Z(n31201) );
  NANDN U32581 ( .A(n31199), .B(n31198), .Z(n31200) );
  AND U32582 ( .A(n31201), .B(n31200), .Z(n31219) );
  XNOR U32583 ( .A(n31220), .B(n31219), .Z(n31221) );
  NANDN U32584 ( .A(n31203), .B(n31202), .Z(n31207) );
  NAND U32585 ( .A(n31205), .B(n31204), .Z(n31206) );
  NAND U32586 ( .A(n31207), .B(n31206), .Z(n31222) );
  XNOR U32587 ( .A(n31221), .B(n31222), .Z(n31213) );
  XNOR U32588 ( .A(n31214), .B(n31213), .Z(n31215) );
  XNOR U32589 ( .A(n31216), .B(n31215), .Z(n31245) );
  XNOR U32590 ( .A(sreg[1749]), .B(n31245), .Z(n31247) );
  NANDN U32591 ( .A(sreg[1748]), .B(n31208), .Z(n31212) );
  NAND U32592 ( .A(n31210), .B(n31209), .Z(n31211) );
  NAND U32593 ( .A(n31212), .B(n31211), .Z(n31246) );
  XNOR U32594 ( .A(n31247), .B(n31246), .Z(c[1749]) );
  NANDN U32595 ( .A(n31214), .B(n31213), .Z(n31218) );
  NANDN U32596 ( .A(n31216), .B(n31215), .Z(n31217) );
  AND U32597 ( .A(n31218), .B(n31217), .Z(n31253) );
  NANDN U32598 ( .A(n31220), .B(n31219), .Z(n31224) );
  NANDN U32599 ( .A(n31222), .B(n31221), .Z(n31223) );
  AND U32600 ( .A(n31224), .B(n31223), .Z(n31251) );
  NAND U32601 ( .A(n42143), .B(n31225), .Z(n31227) );
  XNOR U32602 ( .A(a[728]), .B(n4175), .Z(n31262) );
  NAND U32603 ( .A(n42144), .B(n31262), .Z(n31226) );
  AND U32604 ( .A(n31227), .B(n31226), .Z(n31277) );
  XOR U32605 ( .A(a[732]), .B(n42012), .Z(n31265) );
  XNOR U32606 ( .A(n31277), .B(n31276), .Z(n31279) );
  AND U32607 ( .A(a[734]), .B(b[0]), .Z(n31229) );
  XNOR U32608 ( .A(n31229), .B(n4071), .Z(n31231) );
  NANDN U32609 ( .A(b[0]), .B(a[733]), .Z(n31230) );
  NAND U32610 ( .A(n31231), .B(n31230), .Z(n31273) );
  XOR U32611 ( .A(a[730]), .B(n42085), .Z(n31269) );
  AND U32612 ( .A(a[726]), .B(b[7]), .Z(n31270) );
  XNOR U32613 ( .A(n31271), .B(n31270), .Z(n31272) );
  XNOR U32614 ( .A(n31273), .B(n31272), .Z(n31278) );
  XOR U32615 ( .A(n31279), .B(n31278), .Z(n31257) );
  NANDN U32616 ( .A(n31234), .B(n31233), .Z(n31238) );
  NANDN U32617 ( .A(n31236), .B(n31235), .Z(n31237) );
  AND U32618 ( .A(n31238), .B(n31237), .Z(n31256) );
  XNOR U32619 ( .A(n31257), .B(n31256), .Z(n31258) );
  NANDN U32620 ( .A(n31240), .B(n31239), .Z(n31244) );
  NAND U32621 ( .A(n31242), .B(n31241), .Z(n31243) );
  NAND U32622 ( .A(n31244), .B(n31243), .Z(n31259) );
  XNOR U32623 ( .A(n31258), .B(n31259), .Z(n31250) );
  XNOR U32624 ( .A(n31251), .B(n31250), .Z(n31252) );
  XNOR U32625 ( .A(n31253), .B(n31252), .Z(n31282) );
  XNOR U32626 ( .A(sreg[1750]), .B(n31282), .Z(n31284) );
  NANDN U32627 ( .A(sreg[1749]), .B(n31245), .Z(n31249) );
  NAND U32628 ( .A(n31247), .B(n31246), .Z(n31248) );
  NAND U32629 ( .A(n31249), .B(n31248), .Z(n31283) );
  XNOR U32630 ( .A(n31284), .B(n31283), .Z(c[1750]) );
  NANDN U32631 ( .A(n31251), .B(n31250), .Z(n31255) );
  NANDN U32632 ( .A(n31253), .B(n31252), .Z(n31254) );
  AND U32633 ( .A(n31255), .B(n31254), .Z(n31290) );
  NANDN U32634 ( .A(n31257), .B(n31256), .Z(n31261) );
  NANDN U32635 ( .A(n31259), .B(n31258), .Z(n31260) );
  AND U32636 ( .A(n31261), .B(n31260), .Z(n31288) );
  NAND U32637 ( .A(n42143), .B(n31262), .Z(n31264) );
  XNOR U32638 ( .A(a[729]), .B(n4176), .Z(n31299) );
  NAND U32639 ( .A(n42144), .B(n31299), .Z(n31263) );
  AND U32640 ( .A(n31264), .B(n31263), .Z(n31314) );
  XOR U32641 ( .A(a[733]), .B(n42012), .Z(n31302) );
  XNOR U32642 ( .A(n31314), .B(n31313), .Z(n31316) );
  AND U32643 ( .A(a[735]), .B(b[0]), .Z(n31266) );
  XNOR U32644 ( .A(n31266), .B(n4071), .Z(n31268) );
  NANDN U32645 ( .A(b[0]), .B(a[734]), .Z(n31267) );
  NAND U32646 ( .A(n31268), .B(n31267), .Z(n31310) );
  XOR U32647 ( .A(a[731]), .B(n42085), .Z(n31306) );
  AND U32648 ( .A(a[727]), .B(b[7]), .Z(n31307) );
  XNOR U32649 ( .A(n31308), .B(n31307), .Z(n31309) );
  XNOR U32650 ( .A(n31310), .B(n31309), .Z(n31315) );
  XOR U32651 ( .A(n31316), .B(n31315), .Z(n31294) );
  NANDN U32652 ( .A(n31271), .B(n31270), .Z(n31275) );
  NANDN U32653 ( .A(n31273), .B(n31272), .Z(n31274) );
  AND U32654 ( .A(n31275), .B(n31274), .Z(n31293) );
  XNOR U32655 ( .A(n31294), .B(n31293), .Z(n31295) );
  NANDN U32656 ( .A(n31277), .B(n31276), .Z(n31281) );
  NAND U32657 ( .A(n31279), .B(n31278), .Z(n31280) );
  NAND U32658 ( .A(n31281), .B(n31280), .Z(n31296) );
  XNOR U32659 ( .A(n31295), .B(n31296), .Z(n31287) );
  XNOR U32660 ( .A(n31288), .B(n31287), .Z(n31289) );
  XNOR U32661 ( .A(n31290), .B(n31289), .Z(n31319) );
  XNOR U32662 ( .A(sreg[1751]), .B(n31319), .Z(n31321) );
  NANDN U32663 ( .A(sreg[1750]), .B(n31282), .Z(n31286) );
  NAND U32664 ( .A(n31284), .B(n31283), .Z(n31285) );
  NAND U32665 ( .A(n31286), .B(n31285), .Z(n31320) );
  XNOR U32666 ( .A(n31321), .B(n31320), .Z(c[1751]) );
  NANDN U32667 ( .A(n31288), .B(n31287), .Z(n31292) );
  NANDN U32668 ( .A(n31290), .B(n31289), .Z(n31291) );
  AND U32669 ( .A(n31292), .B(n31291), .Z(n31327) );
  NANDN U32670 ( .A(n31294), .B(n31293), .Z(n31298) );
  NANDN U32671 ( .A(n31296), .B(n31295), .Z(n31297) );
  AND U32672 ( .A(n31298), .B(n31297), .Z(n31325) );
  NAND U32673 ( .A(n42143), .B(n31299), .Z(n31301) );
  XNOR U32674 ( .A(a[730]), .B(n4176), .Z(n31336) );
  NAND U32675 ( .A(n42144), .B(n31336), .Z(n31300) );
  AND U32676 ( .A(n31301), .B(n31300), .Z(n31351) );
  XOR U32677 ( .A(a[734]), .B(n42012), .Z(n31339) );
  XNOR U32678 ( .A(n31351), .B(n31350), .Z(n31353) );
  AND U32679 ( .A(a[736]), .B(b[0]), .Z(n31303) );
  XNOR U32680 ( .A(n31303), .B(n4071), .Z(n31305) );
  NANDN U32681 ( .A(b[0]), .B(a[735]), .Z(n31304) );
  NAND U32682 ( .A(n31305), .B(n31304), .Z(n31347) );
  XOR U32683 ( .A(a[732]), .B(n42085), .Z(n31340) );
  AND U32684 ( .A(a[728]), .B(b[7]), .Z(n31344) );
  XNOR U32685 ( .A(n31345), .B(n31344), .Z(n31346) );
  XNOR U32686 ( .A(n31347), .B(n31346), .Z(n31352) );
  XOR U32687 ( .A(n31353), .B(n31352), .Z(n31331) );
  NANDN U32688 ( .A(n31308), .B(n31307), .Z(n31312) );
  NANDN U32689 ( .A(n31310), .B(n31309), .Z(n31311) );
  AND U32690 ( .A(n31312), .B(n31311), .Z(n31330) );
  XNOR U32691 ( .A(n31331), .B(n31330), .Z(n31332) );
  NANDN U32692 ( .A(n31314), .B(n31313), .Z(n31318) );
  NAND U32693 ( .A(n31316), .B(n31315), .Z(n31317) );
  NAND U32694 ( .A(n31318), .B(n31317), .Z(n31333) );
  XNOR U32695 ( .A(n31332), .B(n31333), .Z(n31324) );
  XNOR U32696 ( .A(n31325), .B(n31324), .Z(n31326) );
  XNOR U32697 ( .A(n31327), .B(n31326), .Z(n31356) );
  XNOR U32698 ( .A(sreg[1752]), .B(n31356), .Z(n31358) );
  NANDN U32699 ( .A(sreg[1751]), .B(n31319), .Z(n31323) );
  NAND U32700 ( .A(n31321), .B(n31320), .Z(n31322) );
  NAND U32701 ( .A(n31323), .B(n31322), .Z(n31357) );
  XNOR U32702 ( .A(n31358), .B(n31357), .Z(c[1752]) );
  NANDN U32703 ( .A(n31325), .B(n31324), .Z(n31329) );
  NANDN U32704 ( .A(n31327), .B(n31326), .Z(n31328) );
  AND U32705 ( .A(n31329), .B(n31328), .Z(n31364) );
  NANDN U32706 ( .A(n31331), .B(n31330), .Z(n31335) );
  NANDN U32707 ( .A(n31333), .B(n31332), .Z(n31334) );
  AND U32708 ( .A(n31335), .B(n31334), .Z(n31362) );
  NAND U32709 ( .A(n42143), .B(n31336), .Z(n31338) );
  XNOR U32710 ( .A(a[731]), .B(n4176), .Z(n31373) );
  NAND U32711 ( .A(n42144), .B(n31373), .Z(n31337) );
  AND U32712 ( .A(n31338), .B(n31337), .Z(n31388) );
  XOR U32713 ( .A(a[735]), .B(n42012), .Z(n31376) );
  XNOR U32714 ( .A(n31388), .B(n31387), .Z(n31390) );
  XOR U32715 ( .A(a[733]), .B(n42085), .Z(n31380) );
  AND U32716 ( .A(a[729]), .B(b[7]), .Z(n31381) );
  XNOR U32717 ( .A(n31382), .B(n31381), .Z(n31383) );
  AND U32718 ( .A(a[737]), .B(b[0]), .Z(n31341) );
  XNOR U32719 ( .A(n31341), .B(n4071), .Z(n31343) );
  NANDN U32720 ( .A(b[0]), .B(a[736]), .Z(n31342) );
  NAND U32721 ( .A(n31343), .B(n31342), .Z(n31384) );
  XNOR U32722 ( .A(n31383), .B(n31384), .Z(n31389) );
  XOR U32723 ( .A(n31390), .B(n31389), .Z(n31368) );
  NANDN U32724 ( .A(n31345), .B(n31344), .Z(n31349) );
  NANDN U32725 ( .A(n31347), .B(n31346), .Z(n31348) );
  AND U32726 ( .A(n31349), .B(n31348), .Z(n31367) );
  XNOR U32727 ( .A(n31368), .B(n31367), .Z(n31369) );
  NANDN U32728 ( .A(n31351), .B(n31350), .Z(n31355) );
  NAND U32729 ( .A(n31353), .B(n31352), .Z(n31354) );
  NAND U32730 ( .A(n31355), .B(n31354), .Z(n31370) );
  XNOR U32731 ( .A(n31369), .B(n31370), .Z(n31361) );
  XNOR U32732 ( .A(n31362), .B(n31361), .Z(n31363) );
  XNOR U32733 ( .A(n31364), .B(n31363), .Z(n31393) );
  XNOR U32734 ( .A(sreg[1753]), .B(n31393), .Z(n31395) );
  NANDN U32735 ( .A(sreg[1752]), .B(n31356), .Z(n31360) );
  NAND U32736 ( .A(n31358), .B(n31357), .Z(n31359) );
  NAND U32737 ( .A(n31360), .B(n31359), .Z(n31394) );
  XNOR U32738 ( .A(n31395), .B(n31394), .Z(c[1753]) );
  NANDN U32739 ( .A(n31362), .B(n31361), .Z(n31366) );
  NANDN U32740 ( .A(n31364), .B(n31363), .Z(n31365) );
  AND U32741 ( .A(n31366), .B(n31365), .Z(n31401) );
  NANDN U32742 ( .A(n31368), .B(n31367), .Z(n31372) );
  NANDN U32743 ( .A(n31370), .B(n31369), .Z(n31371) );
  AND U32744 ( .A(n31372), .B(n31371), .Z(n31399) );
  NAND U32745 ( .A(n42143), .B(n31373), .Z(n31375) );
  XNOR U32746 ( .A(a[732]), .B(n4176), .Z(n31410) );
  NAND U32747 ( .A(n42144), .B(n31410), .Z(n31374) );
  AND U32748 ( .A(n31375), .B(n31374), .Z(n31425) );
  XOR U32749 ( .A(a[736]), .B(n42012), .Z(n31413) );
  XNOR U32750 ( .A(n31425), .B(n31424), .Z(n31427) );
  AND U32751 ( .A(a[738]), .B(b[0]), .Z(n31377) );
  XNOR U32752 ( .A(n31377), .B(n4071), .Z(n31379) );
  NANDN U32753 ( .A(b[0]), .B(a[737]), .Z(n31378) );
  NAND U32754 ( .A(n31379), .B(n31378), .Z(n31421) );
  XOR U32755 ( .A(a[734]), .B(n42085), .Z(n31417) );
  AND U32756 ( .A(a[730]), .B(b[7]), .Z(n31418) );
  XNOR U32757 ( .A(n31419), .B(n31418), .Z(n31420) );
  XNOR U32758 ( .A(n31421), .B(n31420), .Z(n31426) );
  XOR U32759 ( .A(n31427), .B(n31426), .Z(n31405) );
  NANDN U32760 ( .A(n31382), .B(n31381), .Z(n31386) );
  NANDN U32761 ( .A(n31384), .B(n31383), .Z(n31385) );
  AND U32762 ( .A(n31386), .B(n31385), .Z(n31404) );
  XNOR U32763 ( .A(n31405), .B(n31404), .Z(n31406) );
  NANDN U32764 ( .A(n31388), .B(n31387), .Z(n31392) );
  NAND U32765 ( .A(n31390), .B(n31389), .Z(n31391) );
  NAND U32766 ( .A(n31392), .B(n31391), .Z(n31407) );
  XNOR U32767 ( .A(n31406), .B(n31407), .Z(n31398) );
  XNOR U32768 ( .A(n31399), .B(n31398), .Z(n31400) );
  XNOR U32769 ( .A(n31401), .B(n31400), .Z(n31430) );
  XNOR U32770 ( .A(sreg[1754]), .B(n31430), .Z(n31432) );
  NANDN U32771 ( .A(sreg[1753]), .B(n31393), .Z(n31397) );
  NAND U32772 ( .A(n31395), .B(n31394), .Z(n31396) );
  NAND U32773 ( .A(n31397), .B(n31396), .Z(n31431) );
  XNOR U32774 ( .A(n31432), .B(n31431), .Z(c[1754]) );
  NANDN U32775 ( .A(n31399), .B(n31398), .Z(n31403) );
  NANDN U32776 ( .A(n31401), .B(n31400), .Z(n31402) );
  AND U32777 ( .A(n31403), .B(n31402), .Z(n31438) );
  NANDN U32778 ( .A(n31405), .B(n31404), .Z(n31409) );
  NANDN U32779 ( .A(n31407), .B(n31406), .Z(n31408) );
  AND U32780 ( .A(n31409), .B(n31408), .Z(n31436) );
  NAND U32781 ( .A(n42143), .B(n31410), .Z(n31412) );
  XNOR U32782 ( .A(a[733]), .B(n4176), .Z(n31447) );
  NAND U32783 ( .A(n42144), .B(n31447), .Z(n31411) );
  AND U32784 ( .A(n31412), .B(n31411), .Z(n31462) );
  XOR U32785 ( .A(a[737]), .B(n42012), .Z(n31450) );
  XNOR U32786 ( .A(n31462), .B(n31461), .Z(n31464) );
  AND U32787 ( .A(a[739]), .B(b[0]), .Z(n31414) );
  XNOR U32788 ( .A(n31414), .B(n4071), .Z(n31416) );
  NANDN U32789 ( .A(b[0]), .B(a[738]), .Z(n31415) );
  NAND U32790 ( .A(n31416), .B(n31415), .Z(n31458) );
  XOR U32791 ( .A(a[735]), .B(n42085), .Z(n31454) );
  AND U32792 ( .A(a[731]), .B(b[7]), .Z(n31455) );
  XNOR U32793 ( .A(n31456), .B(n31455), .Z(n31457) );
  XNOR U32794 ( .A(n31458), .B(n31457), .Z(n31463) );
  XOR U32795 ( .A(n31464), .B(n31463), .Z(n31442) );
  NANDN U32796 ( .A(n31419), .B(n31418), .Z(n31423) );
  NANDN U32797 ( .A(n31421), .B(n31420), .Z(n31422) );
  AND U32798 ( .A(n31423), .B(n31422), .Z(n31441) );
  XNOR U32799 ( .A(n31442), .B(n31441), .Z(n31443) );
  NANDN U32800 ( .A(n31425), .B(n31424), .Z(n31429) );
  NAND U32801 ( .A(n31427), .B(n31426), .Z(n31428) );
  NAND U32802 ( .A(n31429), .B(n31428), .Z(n31444) );
  XNOR U32803 ( .A(n31443), .B(n31444), .Z(n31435) );
  XNOR U32804 ( .A(n31436), .B(n31435), .Z(n31437) );
  XNOR U32805 ( .A(n31438), .B(n31437), .Z(n31467) );
  XNOR U32806 ( .A(sreg[1755]), .B(n31467), .Z(n31469) );
  NANDN U32807 ( .A(sreg[1754]), .B(n31430), .Z(n31434) );
  NAND U32808 ( .A(n31432), .B(n31431), .Z(n31433) );
  NAND U32809 ( .A(n31434), .B(n31433), .Z(n31468) );
  XNOR U32810 ( .A(n31469), .B(n31468), .Z(c[1755]) );
  NANDN U32811 ( .A(n31436), .B(n31435), .Z(n31440) );
  NANDN U32812 ( .A(n31438), .B(n31437), .Z(n31439) );
  AND U32813 ( .A(n31440), .B(n31439), .Z(n31475) );
  NANDN U32814 ( .A(n31442), .B(n31441), .Z(n31446) );
  NANDN U32815 ( .A(n31444), .B(n31443), .Z(n31445) );
  AND U32816 ( .A(n31446), .B(n31445), .Z(n31473) );
  NAND U32817 ( .A(n42143), .B(n31447), .Z(n31449) );
  XNOR U32818 ( .A(a[734]), .B(n4176), .Z(n31484) );
  NAND U32819 ( .A(n42144), .B(n31484), .Z(n31448) );
  AND U32820 ( .A(n31449), .B(n31448), .Z(n31499) );
  XOR U32821 ( .A(a[738]), .B(n42012), .Z(n31487) );
  XNOR U32822 ( .A(n31499), .B(n31498), .Z(n31501) );
  AND U32823 ( .A(a[740]), .B(b[0]), .Z(n31451) );
  XNOR U32824 ( .A(n31451), .B(n4071), .Z(n31453) );
  NANDN U32825 ( .A(b[0]), .B(a[739]), .Z(n31452) );
  NAND U32826 ( .A(n31453), .B(n31452), .Z(n31495) );
  XOR U32827 ( .A(a[736]), .B(n42085), .Z(n31491) );
  AND U32828 ( .A(a[732]), .B(b[7]), .Z(n31492) );
  XNOR U32829 ( .A(n31493), .B(n31492), .Z(n31494) );
  XNOR U32830 ( .A(n31495), .B(n31494), .Z(n31500) );
  XOR U32831 ( .A(n31501), .B(n31500), .Z(n31479) );
  NANDN U32832 ( .A(n31456), .B(n31455), .Z(n31460) );
  NANDN U32833 ( .A(n31458), .B(n31457), .Z(n31459) );
  AND U32834 ( .A(n31460), .B(n31459), .Z(n31478) );
  XNOR U32835 ( .A(n31479), .B(n31478), .Z(n31480) );
  NANDN U32836 ( .A(n31462), .B(n31461), .Z(n31466) );
  NAND U32837 ( .A(n31464), .B(n31463), .Z(n31465) );
  NAND U32838 ( .A(n31466), .B(n31465), .Z(n31481) );
  XNOR U32839 ( .A(n31480), .B(n31481), .Z(n31472) );
  XNOR U32840 ( .A(n31473), .B(n31472), .Z(n31474) );
  XNOR U32841 ( .A(n31475), .B(n31474), .Z(n31504) );
  XNOR U32842 ( .A(sreg[1756]), .B(n31504), .Z(n31506) );
  NANDN U32843 ( .A(sreg[1755]), .B(n31467), .Z(n31471) );
  NAND U32844 ( .A(n31469), .B(n31468), .Z(n31470) );
  NAND U32845 ( .A(n31471), .B(n31470), .Z(n31505) );
  XNOR U32846 ( .A(n31506), .B(n31505), .Z(c[1756]) );
  NANDN U32847 ( .A(n31473), .B(n31472), .Z(n31477) );
  NANDN U32848 ( .A(n31475), .B(n31474), .Z(n31476) );
  AND U32849 ( .A(n31477), .B(n31476), .Z(n31512) );
  NANDN U32850 ( .A(n31479), .B(n31478), .Z(n31483) );
  NANDN U32851 ( .A(n31481), .B(n31480), .Z(n31482) );
  AND U32852 ( .A(n31483), .B(n31482), .Z(n31510) );
  NAND U32853 ( .A(n42143), .B(n31484), .Z(n31486) );
  XNOR U32854 ( .A(a[735]), .B(n4176), .Z(n31521) );
  NAND U32855 ( .A(n42144), .B(n31521), .Z(n31485) );
  AND U32856 ( .A(n31486), .B(n31485), .Z(n31536) );
  XOR U32857 ( .A(a[739]), .B(n42012), .Z(n31524) );
  XNOR U32858 ( .A(n31536), .B(n31535), .Z(n31538) );
  AND U32859 ( .A(a[741]), .B(b[0]), .Z(n31488) );
  XNOR U32860 ( .A(n31488), .B(n4071), .Z(n31490) );
  NANDN U32861 ( .A(b[0]), .B(a[740]), .Z(n31489) );
  NAND U32862 ( .A(n31490), .B(n31489), .Z(n31532) );
  XOR U32863 ( .A(a[737]), .B(n42085), .Z(n31525) );
  AND U32864 ( .A(a[733]), .B(b[7]), .Z(n31529) );
  XNOR U32865 ( .A(n31530), .B(n31529), .Z(n31531) );
  XNOR U32866 ( .A(n31532), .B(n31531), .Z(n31537) );
  XOR U32867 ( .A(n31538), .B(n31537), .Z(n31516) );
  NANDN U32868 ( .A(n31493), .B(n31492), .Z(n31497) );
  NANDN U32869 ( .A(n31495), .B(n31494), .Z(n31496) );
  AND U32870 ( .A(n31497), .B(n31496), .Z(n31515) );
  XNOR U32871 ( .A(n31516), .B(n31515), .Z(n31517) );
  NANDN U32872 ( .A(n31499), .B(n31498), .Z(n31503) );
  NAND U32873 ( .A(n31501), .B(n31500), .Z(n31502) );
  NAND U32874 ( .A(n31503), .B(n31502), .Z(n31518) );
  XNOR U32875 ( .A(n31517), .B(n31518), .Z(n31509) );
  XNOR U32876 ( .A(n31510), .B(n31509), .Z(n31511) );
  XNOR U32877 ( .A(n31512), .B(n31511), .Z(n31541) );
  XNOR U32878 ( .A(sreg[1757]), .B(n31541), .Z(n31543) );
  NANDN U32879 ( .A(sreg[1756]), .B(n31504), .Z(n31508) );
  NAND U32880 ( .A(n31506), .B(n31505), .Z(n31507) );
  NAND U32881 ( .A(n31508), .B(n31507), .Z(n31542) );
  XNOR U32882 ( .A(n31543), .B(n31542), .Z(c[1757]) );
  NANDN U32883 ( .A(n31510), .B(n31509), .Z(n31514) );
  NANDN U32884 ( .A(n31512), .B(n31511), .Z(n31513) );
  AND U32885 ( .A(n31514), .B(n31513), .Z(n31549) );
  NANDN U32886 ( .A(n31516), .B(n31515), .Z(n31520) );
  NANDN U32887 ( .A(n31518), .B(n31517), .Z(n31519) );
  AND U32888 ( .A(n31520), .B(n31519), .Z(n31547) );
  NAND U32889 ( .A(n42143), .B(n31521), .Z(n31523) );
  XNOR U32890 ( .A(a[736]), .B(n4177), .Z(n31558) );
  NAND U32891 ( .A(n42144), .B(n31558), .Z(n31522) );
  AND U32892 ( .A(n31523), .B(n31522), .Z(n31573) );
  XOR U32893 ( .A(a[740]), .B(n42012), .Z(n31561) );
  XNOR U32894 ( .A(n31573), .B(n31572), .Z(n31575) );
  XOR U32895 ( .A(a[738]), .B(n42085), .Z(n31562) );
  AND U32896 ( .A(a[734]), .B(b[7]), .Z(n31566) );
  XNOR U32897 ( .A(n31567), .B(n31566), .Z(n31568) );
  AND U32898 ( .A(a[742]), .B(b[0]), .Z(n31526) );
  XNOR U32899 ( .A(n31526), .B(n4071), .Z(n31528) );
  NANDN U32900 ( .A(b[0]), .B(a[741]), .Z(n31527) );
  NAND U32901 ( .A(n31528), .B(n31527), .Z(n31569) );
  XNOR U32902 ( .A(n31568), .B(n31569), .Z(n31574) );
  XOR U32903 ( .A(n31575), .B(n31574), .Z(n31553) );
  NANDN U32904 ( .A(n31530), .B(n31529), .Z(n31534) );
  NANDN U32905 ( .A(n31532), .B(n31531), .Z(n31533) );
  AND U32906 ( .A(n31534), .B(n31533), .Z(n31552) );
  XNOR U32907 ( .A(n31553), .B(n31552), .Z(n31554) );
  NANDN U32908 ( .A(n31536), .B(n31535), .Z(n31540) );
  NAND U32909 ( .A(n31538), .B(n31537), .Z(n31539) );
  NAND U32910 ( .A(n31540), .B(n31539), .Z(n31555) );
  XNOR U32911 ( .A(n31554), .B(n31555), .Z(n31546) );
  XNOR U32912 ( .A(n31547), .B(n31546), .Z(n31548) );
  XNOR U32913 ( .A(n31549), .B(n31548), .Z(n31578) );
  XNOR U32914 ( .A(sreg[1758]), .B(n31578), .Z(n31580) );
  NANDN U32915 ( .A(sreg[1757]), .B(n31541), .Z(n31545) );
  NAND U32916 ( .A(n31543), .B(n31542), .Z(n31544) );
  NAND U32917 ( .A(n31545), .B(n31544), .Z(n31579) );
  XNOR U32918 ( .A(n31580), .B(n31579), .Z(c[1758]) );
  NANDN U32919 ( .A(n31547), .B(n31546), .Z(n31551) );
  NANDN U32920 ( .A(n31549), .B(n31548), .Z(n31550) );
  AND U32921 ( .A(n31551), .B(n31550), .Z(n31586) );
  NANDN U32922 ( .A(n31553), .B(n31552), .Z(n31557) );
  NANDN U32923 ( .A(n31555), .B(n31554), .Z(n31556) );
  AND U32924 ( .A(n31557), .B(n31556), .Z(n31584) );
  NAND U32925 ( .A(n42143), .B(n31558), .Z(n31560) );
  XNOR U32926 ( .A(a[737]), .B(n4177), .Z(n31595) );
  NAND U32927 ( .A(n42144), .B(n31595), .Z(n31559) );
  AND U32928 ( .A(n31560), .B(n31559), .Z(n31610) );
  XOR U32929 ( .A(a[741]), .B(n42012), .Z(n31598) );
  XNOR U32930 ( .A(n31610), .B(n31609), .Z(n31612) );
  XOR U32931 ( .A(a[739]), .B(n42085), .Z(n31602) );
  AND U32932 ( .A(a[735]), .B(b[7]), .Z(n31603) );
  XNOR U32933 ( .A(n31604), .B(n31603), .Z(n31605) );
  AND U32934 ( .A(a[743]), .B(b[0]), .Z(n31563) );
  XNOR U32935 ( .A(n31563), .B(n4071), .Z(n31565) );
  NANDN U32936 ( .A(b[0]), .B(a[742]), .Z(n31564) );
  NAND U32937 ( .A(n31565), .B(n31564), .Z(n31606) );
  XNOR U32938 ( .A(n31605), .B(n31606), .Z(n31611) );
  XOR U32939 ( .A(n31612), .B(n31611), .Z(n31590) );
  NANDN U32940 ( .A(n31567), .B(n31566), .Z(n31571) );
  NANDN U32941 ( .A(n31569), .B(n31568), .Z(n31570) );
  AND U32942 ( .A(n31571), .B(n31570), .Z(n31589) );
  XNOR U32943 ( .A(n31590), .B(n31589), .Z(n31591) );
  NANDN U32944 ( .A(n31573), .B(n31572), .Z(n31577) );
  NAND U32945 ( .A(n31575), .B(n31574), .Z(n31576) );
  NAND U32946 ( .A(n31577), .B(n31576), .Z(n31592) );
  XNOR U32947 ( .A(n31591), .B(n31592), .Z(n31583) );
  XNOR U32948 ( .A(n31584), .B(n31583), .Z(n31585) );
  XNOR U32949 ( .A(n31586), .B(n31585), .Z(n31615) );
  XNOR U32950 ( .A(sreg[1759]), .B(n31615), .Z(n31617) );
  NANDN U32951 ( .A(sreg[1758]), .B(n31578), .Z(n31582) );
  NAND U32952 ( .A(n31580), .B(n31579), .Z(n31581) );
  NAND U32953 ( .A(n31582), .B(n31581), .Z(n31616) );
  XNOR U32954 ( .A(n31617), .B(n31616), .Z(c[1759]) );
  NANDN U32955 ( .A(n31584), .B(n31583), .Z(n31588) );
  NANDN U32956 ( .A(n31586), .B(n31585), .Z(n31587) );
  AND U32957 ( .A(n31588), .B(n31587), .Z(n31623) );
  NANDN U32958 ( .A(n31590), .B(n31589), .Z(n31594) );
  NANDN U32959 ( .A(n31592), .B(n31591), .Z(n31593) );
  AND U32960 ( .A(n31594), .B(n31593), .Z(n31621) );
  NAND U32961 ( .A(n42143), .B(n31595), .Z(n31597) );
  XNOR U32962 ( .A(a[738]), .B(n4177), .Z(n31632) );
  NAND U32963 ( .A(n42144), .B(n31632), .Z(n31596) );
  AND U32964 ( .A(n31597), .B(n31596), .Z(n31647) );
  XOR U32965 ( .A(a[742]), .B(n42012), .Z(n31635) );
  XNOR U32966 ( .A(n31647), .B(n31646), .Z(n31649) );
  AND U32967 ( .A(a[744]), .B(b[0]), .Z(n31599) );
  XNOR U32968 ( .A(n31599), .B(n4071), .Z(n31601) );
  NANDN U32969 ( .A(b[0]), .B(a[743]), .Z(n31600) );
  NAND U32970 ( .A(n31601), .B(n31600), .Z(n31643) );
  XOR U32971 ( .A(a[740]), .B(n42085), .Z(n31639) );
  AND U32972 ( .A(a[736]), .B(b[7]), .Z(n31640) );
  XNOR U32973 ( .A(n31641), .B(n31640), .Z(n31642) );
  XNOR U32974 ( .A(n31643), .B(n31642), .Z(n31648) );
  XOR U32975 ( .A(n31649), .B(n31648), .Z(n31627) );
  NANDN U32976 ( .A(n31604), .B(n31603), .Z(n31608) );
  NANDN U32977 ( .A(n31606), .B(n31605), .Z(n31607) );
  AND U32978 ( .A(n31608), .B(n31607), .Z(n31626) );
  XNOR U32979 ( .A(n31627), .B(n31626), .Z(n31628) );
  NANDN U32980 ( .A(n31610), .B(n31609), .Z(n31614) );
  NAND U32981 ( .A(n31612), .B(n31611), .Z(n31613) );
  NAND U32982 ( .A(n31614), .B(n31613), .Z(n31629) );
  XNOR U32983 ( .A(n31628), .B(n31629), .Z(n31620) );
  XNOR U32984 ( .A(n31621), .B(n31620), .Z(n31622) );
  XNOR U32985 ( .A(n31623), .B(n31622), .Z(n31652) );
  XNOR U32986 ( .A(sreg[1760]), .B(n31652), .Z(n31654) );
  NANDN U32987 ( .A(sreg[1759]), .B(n31615), .Z(n31619) );
  NAND U32988 ( .A(n31617), .B(n31616), .Z(n31618) );
  NAND U32989 ( .A(n31619), .B(n31618), .Z(n31653) );
  XNOR U32990 ( .A(n31654), .B(n31653), .Z(c[1760]) );
  NANDN U32991 ( .A(n31621), .B(n31620), .Z(n31625) );
  NANDN U32992 ( .A(n31623), .B(n31622), .Z(n31624) );
  AND U32993 ( .A(n31625), .B(n31624), .Z(n31660) );
  NANDN U32994 ( .A(n31627), .B(n31626), .Z(n31631) );
  NANDN U32995 ( .A(n31629), .B(n31628), .Z(n31630) );
  AND U32996 ( .A(n31631), .B(n31630), .Z(n31658) );
  NAND U32997 ( .A(n42143), .B(n31632), .Z(n31634) );
  XNOR U32998 ( .A(a[739]), .B(n4177), .Z(n31669) );
  NAND U32999 ( .A(n42144), .B(n31669), .Z(n31633) );
  AND U33000 ( .A(n31634), .B(n31633), .Z(n31684) );
  XOR U33001 ( .A(a[743]), .B(n42012), .Z(n31672) );
  XNOR U33002 ( .A(n31684), .B(n31683), .Z(n31686) );
  AND U33003 ( .A(a[745]), .B(b[0]), .Z(n31636) );
  XNOR U33004 ( .A(n31636), .B(n4071), .Z(n31638) );
  NANDN U33005 ( .A(b[0]), .B(a[744]), .Z(n31637) );
  NAND U33006 ( .A(n31638), .B(n31637), .Z(n31680) );
  XOR U33007 ( .A(a[741]), .B(n42085), .Z(n31673) );
  AND U33008 ( .A(a[737]), .B(b[7]), .Z(n31677) );
  XNOR U33009 ( .A(n31678), .B(n31677), .Z(n31679) );
  XNOR U33010 ( .A(n31680), .B(n31679), .Z(n31685) );
  XOR U33011 ( .A(n31686), .B(n31685), .Z(n31664) );
  NANDN U33012 ( .A(n31641), .B(n31640), .Z(n31645) );
  NANDN U33013 ( .A(n31643), .B(n31642), .Z(n31644) );
  AND U33014 ( .A(n31645), .B(n31644), .Z(n31663) );
  XNOR U33015 ( .A(n31664), .B(n31663), .Z(n31665) );
  NANDN U33016 ( .A(n31647), .B(n31646), .Z(n31651) );
  NAND U33017 ( .A(n31649), .B(n31648), .Z(n31650) );
  NAND U33018 ( .A(n31651), .B(n31650), .Z(n31666) );
  XNOR U33019 ( .A(n31665), .B(n31666), .Z(n31657) );
  XNOR U33020 ( .A(n31658), .B(n31657), .Z(n31659) );
  XNOR U33021 ( .A(n31660), .B(n31659), .Z(n31689) );
  XNOR U33022 ( .A(sreg[1761]), .B(n31689), .Z(n31691) );
  NANDN U33023 ( .A(sreg[1760]), .B(n31652), .Z(n31656) );
  NAND U33024 ( .A(n31654), .B(n31653), .Z(n31655) );
  NAND U33025 ( .A(n31656), .B(n31655), .Z(n31690) );
  XNOR U33026 ( .A(n31691), .B(n31690), .Z(c[1761]) );
  NANDN U33027 ( .A(n31658), .B(n31657), .Z(n31662) );
  NANDN U33028 ( .A(n31660), .B(n31659), .Z(n31661) );
  AND U33029 ( .A(n31662), .B(n31661), .Z(n31697) );
  NANDN U33030 ( .A(n31664), .B(n31663), .Z(n31668) );
  NANDN U33031 ( .A(n31666), .B(n31665), .Z(n31667) );
  AND U33032 ( .A(n31668), .B(n31667), .Z(n31695) );
  NAND U33033 ( .A(n42143), .B(n31669), .Z(n31671) );
  XNOR U33034 ( .A(a[740]), .B(n4177), .Z(n31706) );
  NAND U33035 ( .A(n42144), .B(n31706), .Z(n31670) );
  AND U33036 ( .A(n31671), .B(n31670), .Z(n31721) );
  XOR U33037 ( .A(a[744]), .B(n42012), .Z(n31709) );
  XNOR U33038 ( .A(n31721), .B(n31720), .Z(n31723) );
  XOR U33039 ( .A(a[742]), .B(n42085), .Z(n31713) );
  AND U33040 ( .A(a[738]), .B(b[7]), .Z(n31714) );
  XNOR U33041 ( .A(n31715), .B(n31714), .Z(n31716) );
  AND U33042 ( .A(a[746]), .B(b[0]), .Z(n31674) );
  XNOR U33043 ( .A(n31674), .B(n4071), .Z(n31676) );
  NANDN U33044 ( .A(b[0]), .B(a[745]), .Z(n31675) );
  NAND U33045 ( .A(n31676), .B(n31675), .Z(n31717) );
  XNOR U33046 ( .A(n31716), .B(n31717), .Z(n31722) );
  XOR U33047 ( .A(n31723), .B(n31722), .Z(n31701) );
  NANDN U33048 ( .A(n31678), .B(n31677), .Z(n31682) );
  NANDN U33049 ( .A(n31680), .B(n31679), .Z(n31681) );
  AND U33050 ( .A(n31682), .B(n31681), .Z(n31700) );
  XNOR U33051 ( .A(n31701), .B(n31700), .Z(n31702) );
  NANDN U33052 ( .A(n31684), .B(n31683), .Z(n31688) );
  NAND U33053 ( .A(n31686), .B(n31685), .Z(n31687) );
  NAND U33054 ( .A(n31688), .B(n31687), .Z(n31703) );
  XNOR U33055 ( .A(n31702), .B(n31703), .Z(n31694) );
  XNOR U33056 ( .A(n31695), .B(n31694), .Z(n31696) );
  XNOR U33057 ( .A(n31697), .B(n31696), .Z(n31726) );
  XNOR U33058 ( .A(sreg[1762]), .B(n31726), .Z(n31728) );
  NANDN U33059 ( .A(sreg[1761]), .B(n31689), .Z(n31693) );
  NAND U33060 ( .A(n31691), .B(n31690), .Z(n31692) );
  NAND U33061 ( .A(n31693), .B(n31692), .Z(n31727) );
  XNOR U33062 ( .A(n31728), .B(n31727), .Z(c[1762]) );
  NANDN U33063 ( .A(n31695), .B(n31694), .Z(n31699) );
  NANDN U33064 ( .A(n31697), .B(n31696), .Z(n31698) );
  AND U33065 ( .A(n31699), .B(n31698), .Z(n31734) );
  NANDN U33066 ( .A(n31701), .B(n31700), .Z(n31705) );
  NANDN U33067 ( .A(n31703), .B(n31702), .Z(n31704) );
  AND U33068 ( .A(n31705), .B(n31704), .Z(n31732) );
  NAND U33069 ( .A(n42143), .B(n31706), .Z(n31708) );
  XNOR U33070 ( .A(a[741]), .B(n4177), .Z(n31743) );
  NAND U33071 ( .A(n42144), .B(n31743), .Z(n31707) );
  AND U33072 ( .A(n31708), .B(n31707), .Z(n31758) );
  XOR U33073 ( .A(a[745]), .B(n42012), .Z(n31746) );
  XNOR U33074 ( .A(n31758), .B(n31757), .Z(n31760) );
  AND U33075 ( .A(a[747]), .B(b[0]), .Z(n31710) );
  XNOR U33076 ( .A(n31710), .B(n4071), .Z(n31712) );
  NANDN U33077 ( .A(b[0]), .B(a[746]), .Z(n31711) );
  NAND U33078 ( .A(n31712), .B(n31711), .Z(n31754) );
  XOR U33079 ( .A(a[743]), .B(n42085), .Z(n31747) );
  AND U33080 ( .A(a[739]), .B(b[7]), .Z(n31751) );
  XNOR U33081 ( .A(n31752), .B(n31751), .Z(n31753) );
  XNOR U33082 ( .A(n31754), .B(n31753), .Z(n31759) );
  XOR U33083 ( .A(n31760), .B(n31759), .Z(n31738) );
  NANDN U33084 ( .A(n31715), .B(n31714), .Z(n31719) );
  NANDN U33085 ( .A(n31717), .B(n31716), .Z(n31718) );
  AND U33086 ( .A(n31719), .B(n31718), .Z(n31737) );
  XNOR U33087 ( .A(n31738), .B(n31737), .Z(n31739) );
  NANDN U33088 ( .A(n31721), .B(n31720), .Z(n31725) );
  NAND U33089 ( .A(n31723), .B(n31722), .Z(n31724) );
  NAND U33090 ( .A(n31725), .B(n31724), .Z(n31740) );
  XNOR U33091 ( .A(n31739), .B(n31740), .Z(n31731) );
  XNOR U33092 ( .A(n31732), .B(n31731), .Z(n31733) );
  XNOR U33093 ( .A(n31734), .B(n31733), .Z(n31763) );
  XNOR U33094 ( .A(sreg[1763]), .B(n31763), .Z(n31765) );
  NANDN U33095 ( .A(sreg[1762]), .B(n31726), .Z(n31730) );
  NAND U33096 ( .A(n31728), .B(n31727), .Z(n31729) );
  NAND U33097 ( .A(n31730), .B(n31729), .Z(n31764) );
  XNOR U33098 ( .A(n31765), .B(n31764), .Z(c[1763]) );
  NANDN U33099 ( .A(n31732), .B(n31731), .Z(n31736) );
  NANDN U33100 ( .A(n31734), .B(n31733), .Z(n31735) );
  AND U33101 ( .A(n31736), .B(n31735), .Z(n31771) );
  NANDN U33102 ( .A(n31738), .B(n31737), .Z(n31742) );
  NANDN U33103 ( .A(n31740), .B(n31739), .Z(n31741) );
  AND U33104 ( .A(n31742), .B(n31741), .Z(n31769) );
  NAND U33105 ( .A(n42143), .B(n31743), .Z(n31745) );
  XNOR U33106 ( .A(a[742]), .B(n4177), .Z(n31780) );
  NAND U33107 ( .A(n42144), .B(n31780), .Z(n31744) );
  AND U33108 ( .A(n31745), .B(n31744), .Z(n31795) );
  XOR U33109 ( .A(a[746]), .B(n42012), .Z(n31783) );
  XNOR U33110 ( .A(n31795), .B(n31794), .Z(n31797) );
  XOR U33111 ( .A(a[744]), .B(n42085), .Z(n31787) );
  AND U33112 ( .A(a[740]), .B(b[7]), .Z(n31788) );
  XNOR U33113 ( .A(n31789), .B(n31788), .Z(n31790) );
  AND U33114 ( .A(a[748]), .B(b[0]), .Z(n31748) );
  XNOR U33115 ( .A(n31748), .B(n4071), .Z(n31750) );
  NANDN U33116 ( .A(b[0]), .B(a[747]), .Z(n31749) );
  NAND U33117 ( .A(n31750), .B(n31749), .Z(n31791) );
  XNOR U33118 ( .A(n31790), .B(n31791), .Z(n31796) );
  XOR U33119 ( .A(n31797), .B(n31796), .Z(n31775) );
  NANDN U33120 ( .A(n31752), .B(n31751), .Z(n31756) );
  NANDN U33121 ( .A(n31754), .B(n31753), .Z(n31755) );
  AND U33122 ( .A(n31756), .B(n31755), .Z(n31774) );
  XNOR U33123 ( .A(n31775), .B(n31774), .Z(n31776) );
  NANDN U33124 ( .A(n31758), .B(n31757), .Z(n31762) );
  NAND U33125 ( .A(n31760), .B(n31759), .Z(n31761) );
  NAND U33126 ( .A(n31762), .B(n31761), .Z(n31777) );
  XNOR U33127 ( .A(n31776), .B(n31777), .Z(n31768) );
  XNOR U33128 ( .A(n31769), .B(n31768), .Z(n31770) );
  XNOR U33129 ( .A(n31771), .B(n31770), .Z(n31800) );
  XNOR U33130 ( .A(sreg[1764]), .B(n31800), .Z(n31802) );
  NANDN U33131 ( .A(sreg[1763]), .B(n31763), .Z(n31767) );
  NAND U33132 ( .A(n31765), .B(n31764), .Z(n31766) );
  NAND U33133 ( .A(n31767), .B(n31766), .Z(n31801) );
  XNOR U33134 ( .A(n31802), .B(n31801), .Z(c[1764]) );
  NANDN U33135 ( .A(n31769), .B(n31768), .Z(n31773) );
  NANDN U33136 ( .A(n31771), .B(n31770), .Z(n31772) );
  AND U33137 ( .A(n31773), .B(n31772), .Z(n31808) );
  NANDN U33138 ( .A(n31775), .B(n31774), .Z(n31779) );
  NANDN U33139 ( .A(n31777), .B(n31776), .Z(n31778) );
  AND U33140 ( .A(n31779), .B(n31778), .Z(n31806) );
  NAND U33141 ( .A(n42143), .B(n31780), .Z(n31782) );
  XNOR U33142 ( .A(a[743]), .B(n4178), .Z(n31817) );
  NAND U33143 ( .A(n42144), .B(n31817), .Z(n31781) );
  AND U33144 ( .A(n31782), .B(n31781), .Z(n31832) );
  XOR U33145 ( .A(a[747]), .B(n42012), .Z(n31820) );
  XNOR U33146 ( .A(n31832), .B(n31831), .Z(n31834) );
  AND U33147 ( .A(a[749]), .B(b[0]), .Z(n31784) );
  XNOR U33148 ( .A(n31784), .B(n4071), .Z(n31786) );
  NANDN U33149 ( .A(b[0]), .B(a[748]), .Z(n31785) );
  NAND U33150 ( .A(n31786), .B(n31785), .Z(n31828) );
  XOR U33151 ( .A(a[745]), .B(n42085), .Z(n31824) );
  AND U33152 ( .A(a[741]), .B(b[7]), .Z(n31825) );
  XNOR U33153 ( .A(n31826), .B(n31825), .Z(n31827) );
  XNOR U33154 ( .A(n31828), .B(n31827), .Z(n31833) );
  XOR U33155 ( .A(n31834), .B(n31833), .Z(n31812) );
  NANDN U33156 ( .A(n31789), .B(n31788), .Z(n31793) );
  NANDN U33157 ( .A(n31791), .B(n31790), .Z(n31792) );
  AND U33158 ( .A(n31793), .B(n31792), .Z(n31811) );
  XNOR U33159 ( .A(n31812), .B(n31811), .Z(n31813) );
  NANDN U33160 ( .A(n31795), .B(n31794), .Z(n31799) );
  NAND U33161 ( .A(n31797), .B(n31796), .Z(n31798) );
  NAND U33162 ( .A(n31799), .B(n31798), .Z(n31814) );
  XNOR U33163 ( .A(n31813), .B(n31814), .Z(n31805) );
  XNOR U33164 ( .A(n31806), .B(n31805), .Z(n31807) );
  XNOR U33165 ( .A(n31808), .B(n31807), .Z(n31837) );
  XNOR U33166 ( .A(sreg[1765]), .B(n31837), .Z(n31839) );
  NANDN U33167 ( .A(sreg[1764]), .B(n31800), .Z(n31804) );
  NAND U33168 ( .A(n31802), .B(n31801), .Z(n31803) );
  NAND U33169 ( .A(n31804), .B(n31803), .Z(n31838) );
  XNOR U33170 ( .A(n31839), .B(n31838), .Z(c[1765]) );
  NANDN U33171 ( .A(n31806), .B(n31805), .Z(n31810) );
  NANDN U33172 ( .A(n31808), .B(n31807), .Z(n31809) );
  AND U33173 ( .A(n31810), .B(n31809), .Z(n31845) );
  NANDN U33174 ( .A(n31812), .B(n31811), .Z(n31816) );
  NANDN U33175 ( .A(n31814), .B(n31813), .Z(n31815) );
  AND U33176 ( .A(n31816), .B(n31815), .Z(n31843) );
  NAND U33177 ( .A(n42143), .B(n31817), .Z(n31819) );
  XNOR U33178 ( .A(a[744]), .B(n4178), .Z(n31854) );
  NAND U33179 ( .A(n42144), .B(n31854), .Z(n31818) );
  AND U33180 ( .A(n31819), .B(n31818), .Z(n31869) );
  XOR U33181 ( .A(a[748]), .B(n42012), .Z(n31857) );
  XNOR U33182 ( .A(n31869), .B(n31868), .Z(n31871) );
  AND U33183 ( .A(a[750]), .B(b[0]), .Z(n31821) );
  XNOR U33184 ( .A(n31821), .B(n4071), .Z(n31823) );
  NANDN U33185 ( .A(b[0]), .B(a[749]), .Z(n31822) );
  NAND U33186 ( .A(n31823), .B(n31822), .Z(n31865) );
  XOR U33187 ( .A(a[746]), .B(n42085), .Z(n31858) );
  AND U33188 ( .A(a[742]), .B(b[7]), .Z(n31862) );
  XNOR U33189 ( .A(n31863), .B(n31862), .Z(n31864) );
  XNOR U33190 ( .A(n31865), .B(n31864), .Z(n31870) );
  XOR U33191 ( .A(n31871), .B(n31870), .Z(n31849) );
  NANDN U33192 ( .A(n31826), .B(n31825), .Z(n31830) );
  NANDN U33193 ( .A(n31828), .B(n31827), .Z(n31829) );
  AND U33194 ( .A(n31830), .B(n31829), .Z(n31848) );
  XNOR U33195 ( .A(n31849), .B(n31848), .Z(n31850) );
  NANDN U33196 ( .A(n31832), .B(n31831), .Z(n31836) );
  NAND U33197 ( .A(n31834), .B(n31833), .Z(n31835) );
  NAND U33198 ( .A(n31836), .B(n31835), .Z(n31851) );
  XNOR U33199 ( .A(n31850), .B(n31851), .Z(n31842) );
  XNOR U33200 ( .A(n31843), .B(n31842), .Z(n31844) );
  XNOR U33201 ( .A(n31845), .B(n31844), .Z(n31874) );
  XNOR U33202 ( .A(sreg[1766]), .B(n31874), .Z(n31876) );
  NANDN U33203 ( .A(sreg[1765]), .B(n31837), .Z(n31841) );
  NAND U33204 ( .A(n31839), .B(n31838), .Z(n31840) );
  NAND U33205 ( .A(n31841), .B(n31840), .Z(n31875) );
  XNOR U33206 ( .A(n31876), .B(n31875), .Z(c[1766]) );
  NANDN U33207 ( .A(n31843), .B(n31842), .Z(n31847) );
  NANDN U33208 ( .A(n31845), .B(n31844), .Z(n31846) );
  AND U33209 ( .A(n31847), .B(n31846), .Z(n31882) );
  NANDN U33210 ( .A(n31849), .B(n31848), .Z(n31853) );
  NANDN U33211 ( .A(n31851), .B(n31850), .Z(n31852) );
  AND U33212 ( .A(n31853), .B(n31852), .Z(n31880) );
  NAND U33213 ( .A(n42143), .B(n31854), .Z(n31856) );
  XNOR U33214 ( .A(a[745]), .B(n4178), .Z(n31891) );
  NAND U33215 ( .A(n42144), .B(n31891), .Z(n31855) );
  AND U33216 ( .A(n31856), .B(n31855), .Z(n31906) );
  XOR U33217 ( .A(a[749]), .B(n42012), .Z(n31894) );
  XNOR U33218 ( .A(n31906), .B(n31905), .Z(n31908) );
  XOR U33219 ( .A(a[747]), .B(n42085), .Z(n31898) );
  AND U33220 ( .A(a[743]), .B(b[7]), .Z(n31899) );
  XNOR U33221 ( .A(n31900), .B(n31899), .Z(n31901) );
  AND U33222 ( .A(a[751]), .B(b[0]), .Z(n31859) );
  XNOR U33223 ( .A(n31859), .B(n4071), .Z(n31861) );
  NANDN U33224 ( .A(b[0]), .B(a[750]), .Z(n31860) );
  NAND U33225 ( .A(n31861), .B(n31860), .Z(n31902) );
  XNOR U33226 ( .A(n31901), .B(n31902), .Z(n31907) );
  XOR U33227 ( .A(n31908), .B(n31907), .Z(n31886) );
  NANDN U33228 ( .A(n31863), .B(n31862), .Z(n31867) );
  NANDN U33229 ( .A(n31865), .B(n31864), .Z(n31866) );
  AND U33230 ( .A(n31867), .B(n31866), .Z(n31885) );
  XNOR U33231 ( .A(n31886), .B(n31885), .Z(n31887) );
  NANDN U33232 ( .A(n31869), .B(n31868), .Z(n31873) );
  NAND U33233 ( .A(n31871), .B(n31870), .Z(n31872) );
  NAND U33234 ( .A(n31873), .B(n31872), .Z(n31888) );
  XNOR U33235 ( .A(n31887), .B(n31888), .Z(n31879) );
  XNOR U33236 ( .A(n31880), .B(n31879), .Z(n31881) );
  XNOR U33237 ( .A(n31882), .B(n31881), .Z(n31911) );
  XNOR U33238 ( .A(sreg[1767]), .B(n31911), .Z(n31913) );
  NANDN U33239 ( .A(sreg[1766]), .B(n31874), .Z(n31878) );
  NAND U33240 ( .A(n31876), .B(n31875), .Z(n31877) );
  NAND U33241 ( .A(n31878), .B(n31877), .Z(n31912) );
  XNOR U33242 ( .A(n31913), .B(n31912), .Z(c[1767]) );
  NANDN U33243 ( .A(n31880), .B(n31879), .Z(n31884) );
  NANDN U33244 ( .A(n31882), .B(n31881), .Z(n31883) );
  AND U33245 ( .A(n31884), .B(n31883), .Z(n31919) );
  NANDN U33246 ( .A(n31886), .B(n31885), .Z(n31890) );
  NANDN U33247 ( .A(n31888), .B(n31887), .Z(n31889) );
  AND U33248 ( .A(n31890), .B(n31889), .Z(n31917) );
  NAND U33249 ( .A(n42143), .B(n31891), .Z(n31893) );
  XNOR U33250 ( .A(a[746]), .B(n4178), .Z(n31928) );
  NAND U33251 ( .A(n42144), .B(n31928), .Z(n31892) );
  AND U33252 ( .A(n31893), .B(n31892), .Z(n31943) );
  XOR U33253 ( .A(a[750]), .B(n42012), .Z(n31931) );
  XNOR U33254 ( .A(n31943), .B(n31942), .Z(n31945) );
  AND U33255 ( .A(a[752]), .B(b[0]), .Z(n31895) );
  XNOR U33256 ( .A(n31895), .B(n4071), .Z(n31897) );
  NANDN U33257 ( .A(b[0]), .B(a[751]), .Z(n31896) );
  NAND U33258 ( .A(n31897), .B(n31896), .Z(n31939) );
  XOR U33259 ( .A(a[748]), .B(n42085), .Z(n31935) );
  AND U33260 ( .A(a[744]), .B(b[7]), .Z(n31936) );
  XNOR U33261 ( .A(n31937), .B(n31936), .Z(n31938) );
  XNOR U33262 ( .A(n31939), .B(n31938), .Z(n31944) );
  XOR U33263 ( .A(n31945), .B(n31944), .Z(n31923) );
  NANDN U33264 ( .A(n31900), .B(n31899), .Z(n31904) );
  NANDN U33265 ( .A(n31902), .B(n31901), .Z(n31903) );
  AND U33266 ( .A(n31904), .B(n31903), .Z(n31922) );
  XNOR U33267 ( .A(n31923), .B(n31922), .Z(n31924) );
  NANDN U33268 ( .A(n31906), .B(n31905), .Z(n31910) );
  NAND U33269 ( .A(n31908), .B(n31907), .Z(n31909) );
  NAND U33270 ( .A(n31910), .B(n31909), .Z(n31925) );
  XNOR U33271 ( .A(n31924), .B(n31925), .Z(n31916) );
  XNOR U33272 ( .A(n31917), .B(n31916), .Z(n31918) );
  XNOR U33273 ( .A(n31919), .B(n31918), .Z(n31948) );
  XNOR U33274 ( .A(sreg[1768]), .B(n31948), .Z(n31950) );
  NANDN U33275 ( .A(sreg[1767]), .B(n31911), .Z(n31915) );
  NAND U33276 ( .A(n31913), .B(n31912), .Z(n31914) );
  NAND U33277 ( .A(n31915), .B(n31914), .Z(n31949) );
  XNOR U33278 ( .A(n31950), .B(n31949), .Z(c[1768]) );
  NANDN U33279 ( .A(n31917), .B(n31916), .Z(n31921) );
  NANDN U33280 ( .A(n31919), .B(n31918), .Z(n31920) );
  AND U33281 ( .A(n31921), .B(n31920), .Z(n31956) );
  NANDN U33282 ( .A(n31923), .B(n31922), .Z(n31927) );
  NANDN U33283 ( .A(n31925), .B(n31924), .Z(n31926) );
  AND U33284 ( .A(n31927), .B(n31926), .Z(n31954) );
  NAND U33285 ( .A(n42143), .B(n31928), .Z(n31930) );
  XNOR U33286 ( .A(a[747]), .B(n4178), .Z(n31965) );
  NAND U33287 ( .A(n42144), .B(n31965), .Z(n31929) );
  AND U33288 ( .A(n31930), .B(n31929), .Z(n31980) );
  XOR U33289 ( .A(a[751]), .B(n42012), .Z(n31968) );
  XNOR U33290 ( .A(n31980), .B(n31979), .Z(n31982) );
  AND U33291 ( .A(a[753]), .B(b[0]), .Z(n31932) );
  XNOR U33292 ( .A(n31932), .B(n4071), .Z(n31934) );
  NANDN U33293 ( .A(b[0]), .B(a[752]), .Z(n31933) );
  NAND U33294 ( .A(n31934), .B(n31933), .Z(n31976) );
  XOR U33295 ( .A(a[749]), .B(n42085), .Z(n31972) );
  AND U33296 ( .A(a[745]), .B(b[7]), .Z(n31973) );
  XNOR U33297 ( .A(n31974), .B(n31973), .Z(n31975) );
  XNOR U33298 ( .A(n31976), .B(n31975), .Z(n31981) );
  XOR U33299 ( .A(n31982), .B(n31981), .Z(n31960) );
  NANDN U33300 ( .A(n31937), .B(n31936), .Z(n31941) );
  NANDN U33301 ( .A(n31939), .B(n31938), .Z(n31940) );
  AND U33302 ( .A(n31941), .B(n31940), .Z(n31959) );
  XNOR U33303 ( .A(n31960), .B(n31959), .Z(n31961) );
  NANDN U33304 ( .A(n31943), .B(n31942), .Z(n31947) );
  NAND U33305 ( .A(n31945), .B(n31944), .Z(n31946) );
  NAND U33306 ( .A(n31947), .B(n31946), .Z(n31962) );
  XNOR U33307 ( .A(n31961), .B(n31962), .Z(n31953) );
  XNOR U33308 ( .A(n31954), .B(n31953), .Z(n31955) );
  XNOR U33309 ( .A(n31956), .B(n31955), .Z(n31985) );
  XNOR U33310 ( .A(sreg[1769]), .B(n31985), .Z(n31987) );
  NANDN U33311 ( .A(sreg[1768]), .B(n31948), .Z(n31952) );
  NAND U33312 ( .A(n31950), .B(n31949), .Z(n31951) );
  NAND U33313 ( .A(n31952), .B(n31951), .Z(n31986) );
  XNOR U33314 ( .A(n31987), .B(n31986), .Z(c[1769]) );
  NANDN U33315 ( .A(n31954), .B(n31953), .Z(n31958) );
  NANDN U33316 ( .A(n31956), .B(n31955), .Z(n31957) );
  AND U33317 ( .A(n31958), .B(n31957), .Z(n31993) );
  NANDN U33318 ( .A(n31960), .B(n31959), .Z(n31964) );
  NANDN U33319 ( .A(n31962), .B(n31961), .Z(n31963) );
  AND U33320 ( .A(n31964), .B(n31963), .Z(n31991) );
  NAND U33321 ( .A(n42143), .B(n31965), .Z(n31967) );
  XNOR U33322 ( .A(a[748]), .B(n4178), .Z(n32002) );
  NAND U33323 ( .A(n42144), .B(n32002), .Z(n31966) );
  AND U33324 ( .A(n31967), .B(n31966), .Z(n32017) );
  XOR U33325 ( .A(a[752]), .B(n42012), .Z(n32005) );
  XNOR U33326 ( .A(n32017), .B(n32016), .Z(n32019) );
  AND U33327 ( .A(a[754]), .B(b[0]), .Z(n31969) );
  XNOR U33328 ( .A(n31969), .B(n4071), .Z(n31971) );
  NANDN U33329 ( .A(b[0]), .B(a[753]), .Z(n31970) );
  NAND U33330 ( .A(n31971), .B(n31970), .Z(n32013) );
  XOR U33331 ( .A(a[750]), .B(n42085), .Z(n32006) );
  AND U33332 ( .A(a[746]), .B(b[7]), .Z(n32010) );
  XNOR U33333 ( .A(n32011), .B(n32010), .Z(n32012) );
  XNOR U33334 ( .A(n32013), .B(n32012), .Z(n32018) );
  XOR U33335 ( .A(n32019), .B(n32018), .Z(n31997) );
  NANDN U33336 ( .A(n31974), .B(n31973), .Z(n31978) );
  NANDN U33337 ( .A(n31976), .B(n31975), .Z(n31977) );
  AND U33338 ( .A(n31978), .B(n31977), .Z(n31996) );
  XNOR U33339 ( .A(n31997), .B(n31996), .Z(n31998) );
  NANDN U33340 ( .A(n31980), .B(n31979), .Z(n31984) );
  NAND U33341 ( .A(n31982), .B(n31981), .Z(n31983) );
  NAND U33342 ( .A(n31984), .B(n31983), .Z(n31999) );
  XNOR U33343 ( .A(n31998), .B(n31999), .Z(n31990) );
  XNOR U33344 ( .A(n31991), .B(n31990), .Z(n31992) );
  XNOR U33345 ( .A(n31993), .B(n31992), .Z(n32022) );
  XNOR U33346 ( .A(sreg[1770]), .B(n32022), .Z(n32024) );
  NANDN U33347 ( .A(sreg[1769]), .B(n31985), .Z(n31989) );
  NAND U33348 ( .A(n31987), .B(n31986), .Z(n31988) );
  NAND U33349 ( .A(n31989), .B(n31988), .Z(n32023) );
  XNOR U33350 ( .A(n32024), .B(n32023), .Z(c[1770]) );
  NANDN U33351 ( .A(n31991), .B(n31990), .Z(n31995) );
  NANDN U33352 ( .A(n31993), .B(n31992), .Z(n31994) );
  AND U33353 ( .A(n31995), .B(n31994), .Z(n32030) );
  NANDN U33354 ( .A(n31997), .B(n31996), .Z(n32001) );
  NANDN U33355 ( .A(n31999), .B(n31998), .Z(n32000) );
  AND U33356 ( .A(n32001), .B(n32000), .Z(n32028) );
  NAND U33357 ( .A(n42143), .B(n32002), .Z(n32004) );
  XNOR U33358 ( .A(a[749]), .B(n4178), .Z(n32039) );
  NAND U33359 ( .A(n42144), .B(n32039), .Z(n32003) );
  AND U33360 ( .A(n32004), .B(n32003), .Z(n32054) );
  XOR U33361 ( .A(a[753]), .B(n42012), .Z(n32042) );
  XNOR U33362 ( .A(n32054), .B(n32053), .Z(n32056) );
  XOR U33363 ( .A(a[751]), .B(n42085), .Z(n32046) );
  AND U33364 ( .A(a[747]), .B(b[7]), .Z(n32047) );
  XNOR U33365 ( .A(n32048), .B(n32047), .Z(n32049) );
  AND U33366 ( .A(a[755]), .B(b[0]), .Z(n32007) );
  XNOR U33367 ( .A(n32007), .B(n4071), .Z(n32009) );
  NANDN U33368 ( .A(b[0]), .B(a[754]), .Z(n32008) );
  NAND U33369 ( .A(n32009), .B(n32008), .Z(n32050) );
  XNOR U33370 ( .A(n32049), .B(n32050), .Z(n32055) );
  XOR U33371 ( .A(n32056), .B(n32055), .Z(n32034) );
  NANDN U33372 ( .A(n32011), .B(n32010), .Z(n32015) );
  NANDN U33373 ( .A(n32013), .B(n32012), .Z(n32014) );
  AND U33374 ( .A(n32015), .B(n32014), .Z(n32033) );
  XNOR U33375 ( .A(n32034), .B(n32033), .Z(n32035) );
  NANDN U33376 ( .A(n32017), .B(n32016), .Z(n32021) );
  NAND U33377 ( .A(n32019), .B(n32018), .Z(n32020) );
  NAND U33378 ( .A(n32021), .B(n32020), .Z(n32036) );
  XNOR U33379 ( .A(n32035), .B(n32036), .Z(n32027) );
  XNOR U33380 ( .A(n32028), .B(n32027), .Z(n32029) );
  XNOR U33381 ( .A(n32030), .B(n32029), .Z(n32059) );
  XNOR U33382 ( .A(sreg[1771]), .B(n32059), .Z(n32061) );
  NANDN U33383 ( .A(sreg[1770]), .B(n32022), .Z(n32026) );
  NAND U33384 ( .A(n32024), .B(n32023), .Z(n32025) );
  NAND U33385 ( .A(n32026), .B(n32025), .Z(n32060) );
  XNOR U33386 ( .A(n32061), .B(n32060), .Z(c[1771]) );
  NANDN U33387 ( .A(n32028), .B(n32027), .Z(n32032) );
  NANDN U33388 ( .A(n32030), .B(n32029), .Z(n32031) );
  AND U33389 ( .A(n32032), .B(n32031), .Z(n32067) );
  NANDN U33390 ( .A(n32034), .B(n32033), .Z(n32038) );
  NANDN U33391 ( .A(n32036), .B(n32035), .Z(n32037) );
  AND U33392 ( .A(n32038), .B(n32037), .Z(n32065) );
  NAND U33393 ( .A(n42143), .B(n32039), .Z(n32041) );
  XNOR U33394 ( .A(a[750]), .B(n4179), .Z(n32076) );
  NAND U33395 ( .A(n42144), .B(n32076), .Z(n32040) );
  AND U33396 ( .A(n32041), .B(n32040), .Z(n32091) );
  XOR U33397 ( .A(a[754]), .B(n42012), .Z(n32079) );
  XNOR U33398 ( .A(n32091), .B(n32090), .Z(n32093) );
  AND U33399 ( .A(a[756]), .B(b[0]), .Z(n32043) );
  XNOR U33400 ( .A(n32043), .B(n4071), .Z(n32045) );
  NANDN U33401 ( .A(b[0]), .B(a[755]), .Z(n32044) );
  NAND U33402 ( .A(n32045), .B(n32044), .Z(n32087) );
  XOR U33403 ( .A(a[752]), .B(n42085), .Z(n32083) );
  AND U33404 ( .A(a[748]), .B(b[7]), .Z(n32084) );
  XNOR U33405 ( .A(n32085), .B(n32084), .Z(n32086) );
  XNOR U33406 ( .A(n32087), .B(n32086), .Z(n32092) );
  XOR U33407 ( .A(n32093), .B(n32092), .Z(n32071) );
  NANDN U33408 ( .A(n32048), .B(n32047), .Z(n32052) );
  NANDN U33409 ( .A(n32050), .B(n32049), .Z(n32051) );
  AND U33410 ( .A(n32052), .B(n32051), .Z(n32070) );
  XNOR U33411 ( .A(n32071), .B(n32070), .Z(n32072) );
  NANDN U33412 ( .A(n32054), .B(n32053), .Z(n32058) );
  NAND U33413 ( .A(n32056), .B(n32055), .Z(n32057) );
  NAND U33414 ( .A(n32058), .B(n32057), .Z(n32073) );
  XNOR U33415 ( .A(n32072), .B(n32073), .Z(n32064) );
  XNOR U33416 ( .A(n32065), .B(n32064), .Z(n32066) );
  XNOR U33417 ( .A(n32067), .B(n32066), .Z(n32096) );
  XNOR U33418 ( .A(sreg[1772]), .B(n32096), .Z(n32098) );
  NANDN U33419 ( .A(sreg[1771]), .B(n32059), .Z(n32063) );
  NAND U33420 ( .A(n32061), .B(n32060), .Z(n32062) );
  NAND U33421 ( .A(n32063), .B(n32062), .Z(n32097) );
  XNOR U33422 ( .A(n32098), .B(n32097), .Z(c[1772]) );
  NANDN U33423 ( .A(n32065), .B(n32064), .Z(n32069) );
  NANDN U33424 ( .A(n32067), .B(n32066), .Z(n32068) );
  AND U33425 ( .A(n32069), .B(n32068), .Z(n32104) );
  NANDN U33426 ( .A(n32071), .B(n32070), .Z(n32075) );
  NANDN U33427 ( .A(n32073), .B(n32072), .Z(n32074) );
  AND U33428 ( .A(n32075), .B(n32074), .Z(n32102) );
  NAND U33429 ( .A(n42143), .B(n32076), .Z(n32078) );
  XNOR U33430 ( .A(a[751]), .B(n4179), .Z(n32113) );
  NAND U33431 ( .A(n42144), .B(n32113), .Z(n32077) );
  AND U33432 ( .A(n32078), .B(n32077), .Z(n32128) );
  XOR U33433 ( .A(a[755]), .B(n42012), .Z(n32116) );
  XNOR U33434 ( .A(n32128), .B(n32127), .Z(n32130) );
  AND U33435 ( .A(a[757]), .B(b[0]), .Z(n32080) );
  XNOR U33436 ( .A(n32080), .B(n4071), .Z(n32082) );
  NANDN U33437 ( .A(b[0]), .B(a[756]), .Z(n32081) );
  NAND U33438 ( .A(n32082), .B(n32081), .Z(n32124) );
  XOR U33439 ( .A(a[753]), .B(n42085), .Z(n32120) );
  AND U33440 ( .A(a[749]), .B(b[7]), .Z(n32121) );
  XNOR U33441 ( .A(n32122), .B(n32121), .Z(n32123) );
  XNOR U33442 ( .A(n32124), .B(n32123), .Z(n32129) );
  XOR U33443 ( .A(n32130), .B(n32129), .Z(n32108) );
  NANDN U33444 ( .A(n32085), .B(n32084), .Z(n32089) );
  NANDN U33445 ( .A(n32087), .B(n32086), .Z(n32088) );
  AND U33446 ( .A(n32089), .B(n32088), .Z(n32107) );
  XNOR U33447 ( .A(n32108), .B(n32107), .Z(n32109) );
  NANDN U33448 ( .A(n32091), .B(n32090), .Z(n32095) );
  NAND U33449 ( .A(n32093), .B(n32092), .Z(n32094) );
  NAND U33450 ( .A(n32095), .B(n32094), .Z(n32110) );
  XNOR U33451 ( .A(n32109), .B(n32110), .Z(n32101) );
  XNOR U33452 ( .A(n32102), .B(n32101), .Z(n32103) );
  XNOR U33453 ( .A(n32104), .B(n32103), .Z(n32133) );
  XNOR U33454 ( .A(sreg[1773]), .B(n32133), .Z(n32135) );
  NANDN U33455 ( .A(sreg[1772]), .B(n32096), .Z(n32100) );
  NAND U33456 ( .A(n32098), .B(n32097), .Z(n32099) );
  NAND U33457 ( .A(n32100), .B(n32099), .Z(n32134) );
  XNOR U33458 ( .A(n32135), .B(n32134), .Z(c[1773]) );
  NANDN U33459 ( .A(n32102), .B(n32101), .Z(n32106) );
  NANDN U33460 ( .A(n32104), .B(n32103), .Z(n32105) );
  AND U33461 ( .A(n32106), .B(n32105), .Z(n32141) );
  NANDN U33462 ( .A(n32108), .B(n32107), .Z(n32112) );
  NANDN U33463 ( .A(n32110), .B(n32109), .Z(n32111) );
  AND U33464 ( .A(n32112), .B(n32111), .Z(n32139) );
  NAND U33465 ( .A(n42143), .B(n32113), .Z(n32115) );
  XNOR U33466 ( .A(a[752]), .B(n4179), .Z(n32150) );
  NAND U33467 ( .A(n42144), .B(n32150), .Z(n32114) );
  AND U33468 ( .A(n32115), .B(n32114), .Z(n32165) );
  XOR U33469 ( .A(a[756]), .B(n42012), .Z(n32153) );
  XNOR U33470 ( .A(n32165), .B(n32164), .Z(n32167) );
  AND U33471 ( .A(a[758]), .B(b[0]), .Z(n32117) );
  XNOR U33472 ( .A(n32117), .B(n4071), .Z(n32119) );
  NANDN U33473 ( .A(b[0]), .B(a[757]), .Z(n32118) );
  NAND U33474 ( .A(n32119), .B(n32118), .Z(n32161) );
  XOR U33475 ( .A(a[754]), .B(n42085), .Z(n32157) );
  AND U33476 ( .A(a[750]), .B(b[7]), .Z(n32158) );
  XNOR U33477 ( .A(n32159), .B(n32158), .Z(n32160) );
  XNOR U33478 ( .A(n32161), .B(n32160), .Z(n32166) );
  XOR U33479 ( .A(n32167), .B(n32166), .Z(n32145) );
  NANDN U33480 ( .A(n32122), .B(n32121), .Z(n32126) );
  NANDN U33481 ( .A(n32124), .B(n32123), .Z(n32125) );
  AND U33482 ( .A(n32126), .B(n32125), .Z(n32144) );
  XNOR U33483 ( .A(n32145), .B(n32144), .Z(n32146) );
  NANDN U33484 ( .A(n32128), .B(n32127), .Z(n32132) );
  NAND U33485 ( .A(n32130), .B(n32129), .Z(n32131) );
  NAND U33486 ( .A(n32132), .B(n32131), .Z(n32147) );
  XNOR U33487 ( .A(n32146), .B(n32147), .Z(n32138) );
  XNOR U33488 ( .A(n32139), .B(n32138), .Z(n32140) );
  XNOR U33489 ( .A(n32141), .B(n32140), .Z(n32170) );
  XNOR U33490 ( .A(sreg[1774]), .B(n32170), .Z(n32172) );
  NANDN U33491 ( .A(sreg[1773]), .B(n32133), .Z(n32137) );
  NAND U33492 ( .A(n32135), .B(n32134), .Z(n32136) );
  NAND U33493 ( .A(n32137), .B(n32136), .Z(n32171) );
  XNOR U33494 ( .A(n32172), .B(n32171), .Z(c[1774]) );
  NANDN U33495 ( .A(n32139), .B(n32138), .Z(n32143) );
  NANDN U33496 ( .A(n32141), .B(n32140), .Z(n32142) );
  AND U33497 ( .A(n32143), .B(n32142), .Z(n32178) );
  NANDN U33498 ( .A(n32145), .B(n32144), .Z(n32149) );
  NANDN U33499 ( .A(n32147), .B(n32146), .Z(n32148) );
  AND U33500 ( .A(n32149), .B(n32148), .Z(n32176) );
  NAND U33501 ( .A(n42143), .B(n32150), .Z(n32152) );
  XNOR U33502 ( .A(a[753]), .B(n4179), .Z(n32187) );
  NAND U33503 ( .A(n42144), .B(n32187), .Z(n32151) );
  AND U33504 ( .A(n32152), .B(n32151), .Z(n32202) );
  XOR U33505 ( .A(a[757]), .B(n42012), .Z(n32190) );
  XNOR U33506 ( .A(n32202), .B(n32201), .Z(n32204) );
  AND U33507 ( .A(a[759]), .B(b[0]), .Z(n32154) );
  XNOR U33508 ( .A(n32154), .B(n4071), .Z(n32156) );
  NANDN U33509 ( .A(b[0]), .B(a[758]), .Z(n32155) );
  NAND U33510 ( .A(n32156), .B(n32155), .Z(n32198) );
  XOR U33511 ( .A(a[755]), .B(n42085), .Z(n32194) );
  AND U33512 ( .A(a[751]), .B(b[7]), .Z(n32195) );
  XNOR U33513 ( .A(n32196), .B(n32195), .Z(n32197) );
  XNOR U33514 ( .A(n32198), .B(n32197), .Z(n32203) );
  XOR U33515 ( .A(n32204), .B(n32203), .Z(n32182) );
  NANDN U33516 ( .A(n32159), .B(n32158), .Z(n32163) );
  NANDN U33517 ( .A(n32161), .B(n32160), .Z(n32162) );
  AND U33518 ( .A(n32163), .B(n32162), .Z(n32181) );
  XNOR U33519 ( .A(n32182), .B(n32181), .Z(n32183) );
  NANDN U33520 ( .A(n32165), .B(n32164), .Z(n32169) );
  NAND U33521 ( .A(n32167), .B(n32166), .Z(n32168) );
  NAND U33522 ( .A(n32169), .B(n32168), .Z(n32184) );
  XNOR U33523 ( .A(n32183), .B(n32184), .Z(n32175) );
  XNOR U33524 ( .A(n32176), .B(n32175), .Z(n32177) );
  XNOR U33525 ( .A(n32178), .B(n32177), .Z(n32207) );
  XNOR U33526 ( .A(sreg[1775]), .B(n32207), .Z(n32209) );
  NANDN U33527 ( .A(sreg[1774]), .B(n32170), .Z(n32174) );
  NAND U33528 ( .A(n32172), .B(n32171), .Z(n32173) );
  NAND U33529 ( .A(n32174), .B(n32173), .Z(n32208) );
  XNOR U33530 ( .A(n32209), .B(n32208), .Z(c[1775]) );
  NANDN U33531 ( .A(n32176), .B(n32175), .Z(n32180) );
  NANDN U33532 ( .A(n32178), .B(n32177), .Z(n32179) );
  AND U33533 ( .A(n32180), .B(n32179), .Z(n32215) );
  NANDN U33534 ( .A(n32182), .B(n32181), .Z(n32186) );
  NANDN U33535 ( .A(n32184), .B(n32183), .Z(n32185) );
  AND U33536 ( .A(n32186), .B(n32185), .Z(n32213) );
  NAND U33537 ( .A(n42143), .B(n32187), .Z(n32189) );
  XNOR U33538 ( .A(a[754]), .B(n4179), .Z(n32224) );
  NAND U33539 ( .A(n42144), .B(n32224), .Z(n32188) );
  AND U33540 ( .A(n32189), .B(n32188), .Z(n32239) );
  XOR U33541 ( .A(a[758]), .B(n42012), .Z(n32227) );
  XNOR U33542 ( .A(n32239), .B(n32238), .Z(n32241) );
  AND U33543 ( .A(a[760]), .B(b[0]), .Z(n32191) );
  XNOR U33544 ( .A(n32191), .B(n4071), .Z(n32193) );
  NANDN U33545 ( .A(b[0]), .B(a[759]), .Z(n32192) );
  NAND U33546 ( .A(n32193), .B(n32192), .Z(n32235) );
  XOR U33547 ( .A(a[756]), .B(n42085), .Z(n32231) );
  AND U33548 ( .A(a[752]), .B(b[7]), .Z(n32232) );
  XNOR U33549 ( .A(n32233), .B(n32232), .Z(n32234) );
  XNOR U33550 ( .A(n32235), .B(n32234), .Z(n32240) );
  XOR U33551 ( .A(n32241), .B(n32240), .Z(n32219) );
  NANDN U33552 ( .A(n32196), .B(n32195), .Z(n32200) );
  NANDN U33553 ( .A(n32198), .B(n32197), .Z(n32199) );
  AND U33554 ( .A(n32200), .B(n32199), .Z(n32218) );
  XNOR U33555 ( .A(n32219), .B(n32218), .Z(n32220) );
  NANDN U33556 ( .A(n32202), .B(n32201), .Z(n32206) );
  NAND U33557 ( .A(n32204), .B(n32203), .Z(n32205) );
  NAND U33558 ( .A(n32206), .B(n32205), .Z(n32221) );
  XNOR U33559 ( .A(n32220), .B(n32221), .Z(n32212) );
  XNOR U33560 ( .A(n32213), .B(n32212), .Z(n32214) );
  XNOR U33561 ( .A(n32215), .B(n32214), .Z(n32244) );
  XNOR U33562 ( .A(sreg[1776]), .B(n32244), .Z(n32246) );
  NANDN U33563 ( .A(sreg[1775]), .B(n32207), .Z(n32211) );
  NAND U33564 ( .A(n32209), .B(n32208), .Z(n32210) );
  NAND U33565 ( .A(n32211), .B(n32210), .Z(n32245) );
  XNOR U33566 ( .A(n32246), .B(n32245), .Z(c[1776]) );
  NANDN U33567 ( .A(n32213), .B(n32212), .Z(n32217) );
  NANDN U33568 ( .A(n32215), .B(n32214), .Z(n32216) );
  AND U33569 ( .A(n32217), .B(n32216), .Z(n32252) );
  NANDN U33570 ( .A(n32219), .B(n32218), .Z(n32223) );
  NANDN U33571 ( .A(n32221), .B(n32220), .Z(n32222) );
  AND U33572 ( .A(n32223), .B(n32222), .Z(n32250) );
  NAND U33573 ( .A(n42143), .B(n32224), .Z(n32226) );
  XNOR U33574 ( .A(a[755]), .B(n4179), .Z(n32261) );
  NAND U33575 ( .A(n42144), .B(n32261), .Z(n32225) );
  AND U33576 ( .A(n32226), .B(n32225), .Z(n32276) );
  XOR U33577 ( .A(a[759]), .B(n42012), .Z(n32264) );
  XNOR U33578 ( .A(n32276), .B(n32275), .Z(n32278) );
  AND U33579 ( .A(a[761]), .B(b[0]), .Z(n32228) );
  XNOR U33580 ( .A(n32228), .B(n4071), .Z(n32230) );
  NANDN U33581 ( .A(b[0]), .B(a[760]), .Z(n32229) );
  NAND U33582 ( .A(n32230), .B(n32229), .Z(n32272) );
  XOR U33583 ( .A(a[757]), .B(n42085), .Z(n32268) );
  AND U33584 ( .A(a[753]), .B(b[7]), .Z(n32269) );
  XNOR U33585 ( .A(n32270), .B(n32269), .Z(n32271) );
  XNOR U33586 ( .A(n32272), .B(n32271), .Z(n32277) );
  XOR U33587 ( .A(n32278), .B(n32277), .Z(n32256) );
  NANDN U33588 ( .A(n32233), .B(n32232), .Z(n32237) );
  NANDN U33589 ( .A(n32235), .B(n32234), .Z(n32236) );
  AND U33590 ( .A(n32237), .B(n32236), .Z(n32255) );
  XNOR U33591 ( .A(n32256), .B(n32255), .Z(n32257) );
  NANDN U33592 ( .A(n32239), .B(n32238), .Z(n32243) );
  NAND U33593 ( .A(n32241), .B(n32240), .Z(n32242) );
  NAND U33594 ( .A(n32243), .B(n32242), .Z(n32258) );
  XNOR U33595 ( .A(n32257), .B(n32258), .Z(n32249) );
  XNOR U33596 ( .A(n32250), .B(n32249), .Z(n32251) );
  XNOR U33597 ( .A(n32252), .B(n32251), .Z(n32281) );
  XNOR U33598 ( .A(sreg[1777]), .B(n32281), .Z(n32283) );
  NANDN U33599 ( .A(sreg[1776]), .B(n32244), .Z(n32248) );
  NAND U33600 ( .A(n32246), .B(n32245), .Z(n32247) );
  NAND U33601 ( .A(n32248), .B(n32247), .Z(n32282) );
  XNOR U33602 ( .A(n32283), .B(n32282), .Z(c[1777]) );
  NANDN U33603 ( .A(n32250), .B(n32249), .Z(n32254) );
  NANDN U33604 ( .A(n32252), .B(n32251), .Z(n32253) );
  AND U33605 ( .A(n32254), .B(n32253), .Z(n32289) );
  NANDN U33606 ( .A(n32256), .B(n32255), .Z(n32260) );
  NANDN U33607 ( .A(n32258), .B(n32257), .Z(n32259) );
  AND U33608 ( .A(n32260), .B(n32259), .Z(n32287) );
  NAND U33609 ( .A(n42143), .B(n32261), .Z(n32263) );
  XNOR U33610 ( .A(a[756]), .B(n4179), .Z(n32298) );
  NAND U33611 ( .A(n42144), .B(n32298), .Z(n32262) );
  AND U33612 ( .A(n32263), .B(n32262), .Z(n32313) );
  XOR U33613 ( .A(a[760]), .B(n42012), .Z(n32301) );
  XNOR U33614 ( .A(n32313), .B(n32312), .Z(n32315) );
  AND U33615 ( .A(a[762]), .B(b[0]), .Z(n32265) );
  XNOR U33616 ( .A(n32265), .B(n4071), .Z(n32267) );
  NANDN U33617 ( .A(b[0]), .B(a[761]), .Z(n32266) );
  NAND U33618 ( .A(n32267), .B(n32266), .Z(n32309) );
  XOR U33619 ( .A(a[758]), .B(n42085), .Z(n32302) );
  AND U33620 ( .A(a[754]), .B(b[7]), .Z(n32306) );
  XNOR U33621 ( .A(n32307), .B(n32306), .Z(n32308) );
  XNOR U33622 ( .A(n32309), .B(n32308), .Z(n32314) );
  XOR U33623 ( .A(n32315), .B(n32314), .Z(n32293) );
  NANDN U33624 ( .A(n32270), .B(n32269), .Z(n32274) );
  NANDN U33625 ( .A(n32272), .B(n32271), .Z(n32273) );
  AND U33626 ( .A(n32274), .B(n32273), .Z(n32292) );
  XNOR U33627 ( .A(n32293), .B(n32292), .Z(n32294) );
  NANDN U33628 ( .A(n32276), .B(n32275), .Z(n32280) );
  NAND U33629 ( .A(n32278), .B(n32277), .Z(n32279) );
  NAND U33630 ( .A(n32280), .B(n32279), .Z(n32295) );
  XNOR U33631 ( .A(n32294), .B(n32295), .Z(n32286) );
  XNOR U33632 ( .A(n32287), .B(n32286), .Z(n32288) );
  XNOR U33633 ( .A(n32289), .B(n32288), .Z(n32318) );
  XNOR U33634 ( .A(sreg[1778]), .B(n32318), .Z(n32320) );
  NANDN U33635 ( .A(sreg[1777]), .B(n32281), .Z(n32285) );
  NAND U33636 ( .A(n32283), .B(n32282), .Z(n32284) );
  NAND U33637 ( .A(n32285), .B(n32284), .Z(n32319) );
  XNOR U33638 ( .A(n32320), .B(n32319), .Z(c[1778]) );
  NANDN U33639 ( .A(n32287), .B(n32286), .Z(n32291) );
  NANDN U33640 ( .A(n32289), .B(n32288), .Z(n32290) );
  AND U33641 ( .A(n32291), .B(n32290), .Z(n32326) );
  NANDN U33642 ( .A(n32293), .B(n32292), .Z(n32297) );
  NANDN U33643 ( .A(n32295), .B(n32294), .Z(n32296) );
  AND U33644 ( .A(n32297), .B(n32296), .Z(n32324) );
  NAND U33645 ( .A(n42143), .B(n32298), .Z(n32300) );
  XNOR U33646 ( .A(a[757]), .B(n4180), .Z(n32335) );
  NAND U33647 ( .A(n42144), .B(n32335), .Z(n32299) );
  AND U33648 ( .A(n32300), .B(n32299), .Z(n32350) );
  XOR U33649 ( .A(a[761]), .B(n42012), .Z(n32338) );
  XNOR U33650 ( .A(n32350), .B(n32349), .Z(n32352) );
  XOR U33651 ( .A(a[759]), .B(n42085), .Z(n32339) );
  AND U33652 ( .A(a[755]), .B(b[7]), .Z(n32343) );
  XNOR U33653 ( .A(n32344), .B(n32343), .Z(n32345) );
  AND U33654 ( .A(a[763]), .B(b[0]), .Z(n32303) );
  XNOR U33655 ( .A(n32303), .B(n4071), .Z(n32305) );
  NANDN U33656 ( .A(b[0]), .B(a[762]), .Z(n32304) );
  NAND U33657 ( .A(n32305), .B(n32304), .Z(n32346) );
  XNOR U33658 ( .A(n32345), .B(n32346), .Z(n32351) );
  XOR U33659 ( .A(n32352), .B(n32351), .Z(n32330) );
  NANDN U33660 ( .A(n32307), .B(n32306), .Z(n32311) );
  NANDN U33661 ( .A(n32309), .B(n32308), .Z(n32310) );
  AND U33662 ( .A(n32311), .B(n32310), .Z(n32329) );
  XNOR U33663 ( .A(n32330), .B(n32329), .Z(n32331) );
  NANDN U33664 ( .A(n32313), .B(n32312), .Z(n32317) );
  NAND U33665 ( .A(n32315), .B(n32314), .Z(n32316) );
  NAND U33666 ( .A(n32317), .B(n32316), .Z(n32332) );
  XNOR U33667 ( .A(n32331), .B(n32332), .Z(n32323) );
  XNOR U33668 ( .A(n32324), .B(n32323), .Z(n32325) );
  XNOR U33669 ( .A(n32326), .B(n32325), .Z(n32355) );
  XNOR U33670 ( .A(sreg[1779]), .B(n32355), .Z(n32357) );
  NANDN U33671 ( .A(sreg[1778]), .B(n32318), .Z(n32322) );
  NAND U33672 ( .A(n32320), .B(n32319), .Z(n32321) );
  NAND U33673 ( .A(n32322), .B(n32321), .Z(n32356) );
  XNOR U33674 ( .A(n32357), .B(n32356), .Z(c[1779]) );
  NANDN U33675 ( .A(n32324), .B(n32323), .Z(n32328) );
  NANDN U33676 ( .A(n32326), .B(n32325), .Z(n32327) );
  AND U33677 ( .A(n32328), .B(n32327), .Z(n32363) );
  NANDN U33678 ( .A(n32330), .B(n32329), .Z(n32334) );
  NANDN U33679 ( .A(n32332), .B(n32331), .Z(n32333) );
  AND U33680 ( .A(n32334), .B(n32333), .Z(n32361) );
  NAND U33681 ( .A(n42143), .B(n32335), .Z(n32337) );
  XNOR U33682 ( .A(a[758]), .B(n4180), .Z(n32372) );
  NAND U33683 ( .A(n42144), .B(n32372), .Z(n32336) );
  AND U33684 ( .A(n32337), .B(n32336), .Z(n32387) );
  XOR U33685 ( .A(a[762]), .B(n42012), .Z(n32375) );
  XNOR U33686 ( .A(n32387), .B(n32386), .Z(n32389) );
  XOR U33687 ( .A(a[760]), .B(n42085), .Z(n32376) );
  AND U33688 ( .A(a[756]), .B(b[7]), .Z(n32380) );
  XNOR U33689 ( .A(n32381), .B(n32380), .Z(n32382) );
  AND U33690 ( .A(a[764]), .B(b[0]), .Z(n32340) );
  XNOR U33691 ( .A(n32340), .B(n4071), .Z(n32342) );
  NANDN U33692 ( .A(b[0]), .B(a[763]), .Z(n32341) );
  NAND U33693 ( .A(n32342), .B(n32341), .Z(n32383) );
  XNOR U33694 ( .A(n32382), .B(n32383), .Z(n32388) );
  XOR U33695 ( .A(n32389), .B(n32388), .Z(n32367) );
  NANDN U33696 ( .A(n32344), .B(n32343), .Z(n32348) );
  NANDN U33697 ( .A(n32346), .B(n32345), .Z(n32347) );
  AND U33698 ( .A(n32348), .B(n32347), .Z(n32366) );
  XNOR U33699 ( .A(n32367), .B(n32366), .Z(n32368) );
  NANDN U33700 ( .A(n32350), .B(n32349), .Z(n32354) );
  NAND U33701 ( .A(n32352), .B(n32351), .Z(n32353) );
  NAND U33702 ( .A(n32354), .B(n32353), .Z(n32369) );
  XNOR U33703 ( .A(n32368), .B(n32369), .Z(n32360) );
  XNOR U33704 ( .A(n32361), .B(n32360), .Z(n32362) );
  XNOR U33705 ( .A(n32363), .B(n32362), .Z(n32392) );
  XNOR U33706 ( .A(sreg[1780]), .B(n32392), .Z(n32394) );
  NANDN U33707 ( .A(sreg[1779]), .B(n32355), .Z(n32359) );
  NAND U33708 ( .A(n32357), .B(n32356), .Z(n32358) );
  NAND U33709 ( .A(n32359), .B(n32358), .Z(n32393) );
  XNOR U33710 ( .A(n32394), .B(n32393), .Z(c[1780]) );
  NANDN U33711 ( .A(n32361), .B(n32360), .Z(n32365) );
  NANDN U33712 ( .A(n32363), .B(n32362), .Z(n32364) );
  AND U33713 ( .A(n32365), .B(n32364), .Z(n32400) );
  NANDN U33714 ( .A(n32367), .B(n32366), .Z(n32371) );
  NANDN U33715 ( .A(n32369), .B(n32368), .Z(n32370) );
  AND U33716 ( .A(n32371), .B(n32370), .Z(n32398) );
  NAND U33717 ( .A(n42143), .B(n32372), .Z(n32374) );
  XNOR U33718 ( .A(a[759]), .B(n4180), .Z(n32409) );
  NAND U33719 ( .A(n42144), .B(n32409), .Z(n32373) );
  AND U33720 ( .A(n32374), .B(n32373), .Z(n32424) );
  XOR U33721 ( .A(a[763]), .B(n42012), .Z(n32412) );
  XNOR U33722 ( .A(n32424), .B(n32423), .Z(n32426) );
  XOR U33723 ( .A(a[761]), .B(n42085), .Z(n32416) );
  AND U33724 ( .A(a[757]), .B(b[7]), .Z(n32417) );
  XNOR U33725 ( .A(n32418), .B(n32417), .Z(n32419) );
  AND U33726 ( .A(a[765]), .B(b[0]), .Z(n32377) );
  XNOR U33727 ( .A(n32377), .B(n4071), .Z(n32379) );
  NANDN U33728 ( .A(b[0]), .B(a[764]), .Z(n32378) );
  NAND U33729 ( .A(n32379), .B(n32378), .Z(n32420) );
  XNOR U33730 ( .A(n32419), .B(n32420), .Z(n32425) );
  XOR U33731 ( .A(n32426), .B(n32425), .Z(n32404) );
  NANDN U33732 ( .A(n32381), .B(n32380), .Z(n32385) );
  NANDN U33733 ( .A(n32383), .B(n32382), .Z(n32384) );
  AND U33734 ( .A(n32385), .B(n32384), .Z(n32403) );
  XNOR U33735 ( .A(n32404), .B(n32403), .Z(n32405) );
  NANDN U33736 ( .A(n32387), .B(n32386), .Z(n32391) );
  NAND U33737 ( .A(n32389), .B(n32388), .Z(n32390) );
  NAND U33738 ( .A(n32391), .B(n32390), .Z(n32406) );
  XNOR U33739 ( .A(n32405), .B(n32406), .Z(n32397) );
  XNOR U33740 ( .A(n32398), .B(n32397), .Z(n32399) );
  XNOR U33741 ( .A(n32400), .B(n32399), .Z(n32429) );
  XNOR U33742 ( .A(sreg[1781]), .B(n32429), .Z(n32431) );
  NANDN U33743 ( .A(sreg[1780]), .B(n32392), .Z(n32396) );
  NAND U33744 ( .A(n32394), .B(n32393), .Z(n32395) );
  NAND U33745 ( .A(n32396), .B(n32395), .Z(n32430) );
  XNOR U33746 ( .A(n32431), .B(n32430), .Z(c[1781]) );
  NANDN U33747 ( .A(n32398), .B(n32397), .Z(n32402) );
  NANDN U33748 ( .A(n32400), .B(n32399), .Z(n32401) );
  AND U33749 ( .A(n32402), .B(n32401), .Z(n32437) );
  NANDN U33750 ( .A(n32404), .B(n32403), .Z(n32408) );
  NANDN U33751 ( .A(n32406), .B(n32405), .Z(n32407) );
  AND U33752 ( .A(n32408), .B(n32407), .Z(n32435) );
  NAND U33753 ( .A(n42143), .B(n32409), .Z(n32411) );
  XNOR U33754 ( .A(a[760]), .B(n4180), .Z(n32446) );
  NAND U33755 ( .A(n42144), .B(n32446), .Z(n32410) );
  AND U33756 ( .A(n32411), .B(n32410), .Z(n32461) );
  XOR U33757 ( .A(a[764]), .B(n42012), .Z(n32449) );
  XNOR U33758 ( .A(n32461), .B(n32460), .Z(n32463) );
  AND U33759 ( .A(a[766]), .B(b[0]), .Z(n32413) );
  XNOR U33760 ( .A(n32413), .B(n4071), .Z(n32415) );
  NANDN U33761 ( .A(b[0]), .B(a[765]), .Z(n32414) );
  NAND U33762 ( .A(n32415), .B(n32414), .Z(n32457) );
  XOR U33763 ( .A(a[762]), .B(n42085), .Z(n32453) );
  AND U33764 ( .A(a[758]), .B(b[7]), .Z(n32454) );
  XNOR U33765 ( .A(n32455), .B(n32454), .Z(n32456) );
  XNOR U33766 ( .A(n32457), .B(n32456), .Z(n32462) );
  XOR U33767 ( .A(n32463), .B(n32462), .Z(n32441) );
  NANDN U33768 ( .A(n32418), .B(n32417), .Z(n32422) );
  NANDN U33769 ( .A(n32420), .B(n32419), .Z(n32421) );
  AND U33770 ( .A(n32422), .B(n32421), .Z(n32440) );
  XNOR U33771 ( .A(n32441), .B(n32440), .Z(n32442) );
  NANDN U33772 ( .A(n32424), .B(n32423), .Z(n32428) );
  NAND U33773 ( .A(n32426), .B(n32425), .Z(n32427) );
  NAND U33774 ( .A(n32428), .B(n32427), .Z(n32443) );
  XNOR U33775 ( .A(n32442), .B(n32443), .Z(n32434) );
  XNOR U33776 ( .A(n32435), .B(n32434), .Z(n32436) );
  XNOR U33777 ( .A(n32437), .B(n32436), .Z(n32466) );
  XNOR U33778 ( .A(sreg[1782]), .B(n32466), .Z(n32468) );
  NANDN U33779 ( .A(sreg[1781]), .B(n32429), .Z(n32433) );
  NAND U33780 ( .A(n32431), .B(n32430), .Z(n32432) );
  NAND U33781 ( .A(n32433), .B(n32432), .Z(n32467) );
  XNOR U33782 ( .A(n32468), .B(n32467), .Z(c[1782]) );
  NANDN U33783 ( .A(n32435), .B(n32434), .Z(n32439) );
  NANDN U33784 ( .A(n32437), .B(n32436), .Z(n32438) );
  AND U33785 ( .A(n32439), .B(n32438), .Z(n32474) );
  NANDN U33786 ( .A(n32441), .B(n32440), .Z(n32445) );
  NANDN U33787 ( .A(n32443), .B(n32442), .Z(n32444) );
  AND U33788 ( .A(n32445), .B(n32444), .Z(n32472) );
  NAND U33789 ( .A(n42143), .B(n32446), .Z(n32448) );
  XNOR U33790 ( .A(a[761]), .B(n4180), .Z(n32483) );
  NAND U33791 ( .A(n42144), .B(n32483), .Z(n32447) );
  AND U33792 ( .A(n32448), .B(n32447), .Z(n32498) );
  XOR U33793 ( .A(a[765]), .B(n42012), .Z(n32486) );
  XNOR U33794 ( .A(n32498), .B(n32497), .Z(n32500) );
  AND U33795 ( .A(a[767]), .B(b[0]), .Z(n32450) );
  XNOR U33796 ( .A(n32450), .B(n4071), .Z(n32452) );
  NANDN U33797 ( .A(b[0]), .B(a[766]), .Z(n32451) );
  NAND U33798 ( .A(n32452), .B(n32451), .Z(n32494) );
  XOR U33799 ( .A(a[763]), .B(n42085), .Z(n32490) );
  AND U33800 ( .A(a[759]), .B(b[7]), .Z(n32491) );
  XNOR U33801 ( .A(n32492), .B(n32491), .Z(n32493) );
  XNOR U33802 ( .A(n32494), .B(n32493), .Z(n32499) );
  XOR U33803 ( .A(n32500), .B(n32499), .Z(n32478) );
  NANDN U33804 ( .A(n32455), .B(n32454), .Z(n32459) );
  NANDN U33805 ( .A(n32457), .B(n32456), .Z(n32458) );
  AND U33806 ( .A(n32459), .B(n32458), .Z(n32477) );
  XNOR U33807 ( .A(n32478), .B(n32477), .Z(n32479) );
  NANDN U33808 ( .A(n32461), .B(n32460), .Z(n32465) );
  NAND U33809 ( .A(n32463), .B(n32462), .Z(n32464) );
  NAND U33810 ( .A(n32465), .B(n32464), .Z(n32480) );
  XNOR U33811 ( .A(n32479), .B(n32480), .Z(n32471) );
  XNOR U33812 ( .A(n32472), .B(n32471), .Z(n32473) );
  XNOR U33813 ( .A(n32474), .B(n32473), .Z(n32503) );
  XNOR U33814 ( .A(sreg[1783]), .B(n32503), .Z(n32505) );
  NANDN U33815 ( .A(sreg[1782]), .B(n32466), .Z(n32470) );
  NAND U33816 ( .A(n32468), .B(n32467), .Z(n32469) );
  NAND U33817 ( .A(n32470), .B(n32469), .Z(n32504) );
  XNOR U33818 ( .A(n32505), .B(n32504), .Z(c[1783]) );
  NANDN U33819 ( .A(n32472), .B(n32471), .Z(n32476) );
  NANDN U33820 ( .A(n32474), .B(n32473), .Z(n32475) );
  AND U33821 ( .A(n32476), .B(n32475), .Z(n32511) );
  NANDN U33822 ( .A(n32478), .B(n32477), .Z(n32482) );
  NANDN U33823 ( .A(n32480), .B(n32479), .Z(n32481) );
  AND U33824 ( .A(n32482), .B(n32481), .Z(n32509) );
  NAND U33825 ( .A(n42143), .B(n32483), .Z(n32485) );
  XNOR U33826 ( .A(a[762]), .B(n4180), .Z(n32520) );
  NAND U33827 ( .A(n42144), .B(n32520), .Z(n32484) );
  AND U33828 ( .A(n32485), .B(n32484), .Z(n32535) );
  XOR U33829 ( .A(a[766]), .B(n42012), .Z(n32523) );
  XNOR U33830 ( .A(n32535), .B(n32534), .Z(n32537) );
  AND U33831 ( .A(a[768]), .B(b[0]), .Z(n32487) );
  XNOR U33832 ( .A(n32487), .B(n4071), .Z(n32489) );
  NANDN U33833 ( .A(b[0]), .B(a[767]), .Z(n32488) );
  NAND U33834 ( .A(n32489), .B(n32488), .Z(n32531) );
  XOR U33835 ( .A(a[764]), .B(n42085), .Z(n32527) );
  AND U33836 ( .A(a[760]), .B(b[7]), .Z(n32528) );
  XNOR U33837 ( .A(n32529), .B(n32528), .Z(n32530) );
  XNOR U33838 ( .A(n32531), .B(n32530), .Z(n32536) );
  XOR U33839 ( .A(n32537), .B(n32536), .Z(n32515) );
  NANDN U33840 ( .A(n32492), .B(n32491), .Z(n32496) );
  NANDN U33841 ( .A(n32494), .B(n32493), .Z(n32495) );
  AND U33842 ( .A(n32496), .B(n32495), .Z(n32514) );
  XNOR U33843 ( .A(n32515), .B(n32514), .Z(n32516) );
  NANDN U33844 ( .A(n32498), .B(n32497), .Z(n32502) );
  NAND U33845 ( .A(n32500), .B(n32499), .Z(n32501) );
  NAND U33846 ( .A(n32502), .B(n32501), .Z(n32517) );
  XNOR U33847 ( .A(n32516), .B(n32517), .Z(n32508) );
  XNOR U33848 ( .A(n32509), .B(n32508), .Z(n32510) );
  XNOR U33849 ( .A(n32511), .B(n32510), .Z(n32540) );
  XNOR U33850 ( .A(sreg[1784]), .B(n32540), .Z(n32542) );
  NANDN U33851 ( .A(sreg[1783]), .B(n32503), .Z(n32507) );
  NAND U33852 ( .A(n32505), .B(n32504), .Z(n32506) );
  NAND U33853 ( .A(n32507), .B(n32506), .Z(n32541) );
  XNOR U33854 ( .A(n32542), .B(n32541), .Z(c[1784]) );
  NANDN U33855 ( .A(n32509), .B(n32508), .Z(n32513) );
  NANDN U33856 ( .A(n32511), .B(n32510), .Z(n32512) );
  AND U33857 ( .A(n32513), .B(n32512), .Z(n32548) );
  NANDN U33858 ( .A(n32515), .B(n32514), .Z(n32519) );
  NANDN U33859 ( .A(n32517), .B(n32516), .Z(n32518) );
  AND U33860 ( .A(n32519), .B(n32518), .Z(n32546) );
  NAND U33861 ( .A(n42143), .B(n32520), .Z(n32522) );
  XNOR U33862 ( .A(a[763]), .B(n4180), .Z(n32557) );
  NAND U33863 ( .A(n42144), .B(n32557), .Z(n32521) );
  AND U33864 ( .A(n32522), .B(n32521), .Z(n32572) );
  XOR U33865 ( .A(a[767]), .B(n42012), .Z(n32560) );
  XNOR U33866 ( .A(n32572), .B(n32571), .Z(n32574) );
  NAND U33867 ( .A(a[769]), .B(b[0]), .Z(n32524) );
  XNOR U33868 ( .A(b[1]), .B(n32524), .Z(n32526) );
  NANDN U33869 ( .A(b[0]), .B(a[768]), .Z(n32525) );
  AND U33870 ( .A(n32526), .B(n32525), .Z(n32567) );
  XOR U33871 ( .A(a[765]), .B(n42085), .Z(n32564) );
  AND U33872 ( .A(a[761]), .B(b[7]), .Z(n32565) );
  XOR U33873 ( .A(n32566), .B(n32565), .Z(n32568) );
  XNOR U33874 ( .A(n32567), .B(n32568), .Z(n32573) );
  XOR U33875 ( .A(n32574), .B(n32573), .Z(n32552) );
  NANDN U33876 ( .A(n32529), .B(n32528), .Z(n32533) );
  NANDN U33877 ( .A(n32531), .B(n32530), .Z(n32532) );
  AND U33878 ( .A(n32533), .B(n32532), .Z(n32551) );
  XNOR U33879 ( .A(n32552), .B(n32551), .Z(n32553) );
  NANDN U33880 ( .A(n32535), .B(n32534), .Z(n32539) );
  NAND U33881 ( .A(n32537), .B(n32536), .Z(n32538) );
  NAND U33882 ( .A(n32539), .B(n32538), .Z(n32554) );
  XNOR U33883 ( .A(n32553), .B(n32554), .Z(n32545) );
  XNOR U33884 ( .A(n32546), .B(n32545), .Z(n32547) );
  XNOR U33885 ( .A(n32548), .B(n32547), .Z(n32577) );
  XNOR U33886 ( .A(sreg[1785]), .B(n32577), .Z(n32579) );
  NANDN U33887 ( .A(sreg[1784]), .B(n32540), .Z(n32544) );
  NAND U33888 ( .A(n32542), .B(n32541), .Z(n32543) );
  NAND U33889 ( .A(n32544), .B(n32543), .Z(n32578) );
  XNOR U33890 ( .A(n32579), .B(n32578), .Z(c[1785]) );
  NANDN U33891 ( .A(n32546), .B(n32545), .Z(n32550) );
  NANDN U33892 ( .A(n32548), .B(n32547), .Z(n32549) );
  AND U33893 ( .A(n32550), .B(n32549), .Z(n32585) );
  NANDN U33894 ( .A(n32552), .B(n32551), .Z(n32556) );
  NANDN U33895 ( .A(n32554), .B(n32553), .Z(n32555) );
  AND U33896 ( .A(n32556), .B(n32555), .Z(n32583) );
  NAND U33897 ( .A(n42143), .B(n32557), .Z(n32559) );
  XNOR U33898 ( .A(a[764]), .B(n4181), .Z(n32594) );
  NAND U33899 ( .A(n42144), .B(n32594), .Z(n32558) );
  AND U33900 ( .A(n32559), .B(n32558), .Z(n32609) );
  XOR U33901 ( .A(a[768]), .B(n42012), .Z(n32597) );
  XNOR U33902 ( .A(n32609), .B(n32608), .Z(n32611) );
  AND U33903 ( .A(a[770]), .B(b[0]), .Z(n32561) );
  XNOR U33904 ( .A(n32561), .B(n4071), .Z(n32563) );
  NANDN U33905 ( .A(b[0]), .B(a[769]), .Z(n32562) );
  NAND U33906 ( .A(n32563), .B(n32562), .Z(n32605) );
  XOR U33907 ( .A(a[766]), .B(n42085), .Z(n32598) );
  AND U33908 ( .A(a[762]), .B(b[7]), .Z(n32602) );
  XNOR U33909 ( .A(n32603), .B(n32602), .Z(n32604) );
  XNOR U33910 ( .A(n32605), .B(n32604), .Z(n32610) );
  XOR U33911 ( .A(n32611), .B(n32610), .Z(n32589) );
  NANDN U33912 ( .A(n32566), .B(n32565), .Z(n32570) );
  NANDN U33913 ( .A(n32568), .B(n32567), .Z(n32569) );
  AND U33914 ( .A(n32570), .B(n32569), .Z(n32588) );
  XNOR U33915 ( .A(n32589), .B(n32588), .Z(n32590) );
  NANDN U33916 ( .A(n32572), .B(n32571), .Z(n32576) );
  NAND U33917 ( .A(n32574), .B(n32573), .Z(n32575) );
  NAND U33918 ( .A(n32576), .B(n32575), .Z(n32591) );
  XNOR U33919 ( .A(n32590), .B(n32591), .Z(n32582) );
  XNOR U33920 ( .A(n32583), .B(n32582), .Z(n32584) );
  XNOR U33921 ( .A(n32585), .B(n32584), .Z(n32614) );
  XNOR U33922 ( .A(sreg[1786]), .B(n32614), .Z(n32616) );
  NANDN U33923 ( .A(sreg[1785]), .B(n32577), .Z(n32581) );
  NAND U33924 ( .A(n32579), .B(n32578), .Z(n32580) );
  NAND U33925 ( .A(n32581), .B(n32580), .Z(n32615) );
  XNOR U33926 ( .A(n32616), .B(n32615), .Z(c[1786]) );
  NANDN U33927 ( .A(n32583), .B(n32582), .Z(n32587) );
  NANDN U33928 ( .A(n32585), .B(n32584), .Z(n32586) );
  AND U33929 ( .A(n32587), .B(n32586), .Z(n32622) );
  NANDN U33930 ( .A(n32589), .B(n32588), .Z(n32593) );
  NANDN U33931 ( .A(n32591), .B(n32590), .Z(n32592) );
  AND U33932 ( .A(n32593), .B(n32592), .Z(n32620) );
  NAND U33933 ( .A(n42143), .B(n32594), .Z(n32596) );
  XNOR U33934 ( .A(a[765]), .B(n4181), .Z(n32631) );
  NAND U33935 ( .A(n42144), .B(n32631), .Z(n32595) );
  AND U33936 ( .A(n32596), .B(n32595), .Z(n32646) );
  XOR U33937 ( .A(a[769]), .B(n42012), .Z(n32634) );
  XNOR U33938 ( .A(n32646), .B(n32645), .Z(n32648) );
  XOR U33939 ( .A(a[767]), .B(n42085), .Z(n32635) );
  AND U33940 ( .A(a[763]), .B(b[7]), .Z(n32639) );
  XNOR U33941 ( .A(n32640), .B(n32639), .Z(n32641) );
  AND U33942 ( .A(a[771]), .B(b[0]), .Z(n32599) );
  XNOR U33943 ( .A(n32599), .B(n4071), .Z(n32601) );
  NANDN U33944 ( .A(b[0]), .B(a[770]), .Z(n32600) );
  NAND U33945 ( .A(n32601), .B(n32600), .Z(n32642) );
  XNOR U33946 ( .A(n32641), .B(n32642), .Z(n32647) );
  XOR U33947 ( .A(n32648), .B(n32647), .Z(n32626) );
  NANDN U33948 ( .A(n32603), .B(n32602), .Z(n32607) );
  NANDN U33949 ( .A(n32605), .B(n32604), .Z(n32606) );
  AND U33950 ( .A(n32607), .B(n32606), .Z(n32625) );
  XNOR U33951 ( .A(n32626), .B(n32625), .Z(n32627) );
  NANDN U33952 ( .A(n32609), .B(n32608), .Z(n32613) );
  NAND U33953 ( .A(n32611), .B(n32610), .Z(n32612) );
  NAND U33954 ( .A(n32613), .B(n32612), .Z(n32628) );
  XNOR U33955 ( .A(n32627), .B(n32628), .Z(n32619) );
  XNOR U33956 ( .A(n32620), .B(n32619), .Z(n32621) );
  XNOR U33957 ( .A(n32622), .B(n32621), .Z(n32651) );
  XNOR U33958 ( .A(sreg[1787]), .B(n32651), .Z(n32653) );
  NANDN U33959 ( .A(sreg[1786]), .B(n32614), .Z(n32618) );
  NAND U33960 ( .A(n32616), .B(n32615), .Z(n32617) );
  NAND U33961 ( .A(n32618), .B(n32617), .Z(n32652) );
  XNOR U33962 ( .A(n32653), .B(n32652), .Z(c[1787]) );
  NANDN U33963 ( .A(n32620), .B(n32619), .Z(n32624) );
  NANDN U33964 ( .A(n32622), .B(n32621), .Z(n32623) );
  AND U33965 ( .A(n32624), .B(n32623), .Z(n32659) );
  NANDN U33966 ( .A(n32626), .B(n32625), .Z(n32630) );
  NANDN U33967 ( .A(n32628), .B(n32627), .Z(n32629) );
  AND U33968 ( .A(n32630), .B(n32629), .Z(n32657) );
  NAND U33969 ( .A(n42143), .B(n32631), .Z(n32633) );
  XNOR U33970 ( .A(a[766]), .B(n4181), .Z(n32668) );
  NAND U33971 ( .A(n42144), .B(n32668), .Z(n32632) );
  AND U33972 ( .A(n32633), .B(n32632), .Z(n32683) );
  XOR U33973 ( .A(a[770]), .B(n42012), .Z(n32671) );
  XNOR U33974 ( .A(n32683), .B(n32682), .Z(n32685) );
  XOR U33975 ( .A(a[768]), .B(n42085), .Z(n32672) );
  AND U33976 ( .A(a[764]), .B(b[7]), .Z(n32676) );
  XNOR U33977 ( .A(n32677), .B(n32676), .Z(n32678) );
  AND U33978 ( .A(a[772]), .B(b[0]), .Z(n32636) );
  XNOR U33979 ( .A(n32636), .B(n4071), .Z(n32638) );
  NANDN U33980 ( .A(b[0]), .B(a[771]), .Z(n32637) );
  NAND U33981 ( .A(n32638), .B(n32637), .Z(n32679) );
  XNOR U33982 ( .A(n32678), .B(n32679), .Z(n32684) );
  XOR U33983 ( .A(n32685), .B(n32684), .Z(n32663) );
  NANDN U33984 ( .A(n32640), .B(n32639), .Z(n32644) );
  NANDN U33985 ( .A(n32642), .B(n32641), .Z(n32643) );
  AND U33986 ( .A(n32644), .B(n32643), .Z(n32662) );
  XNOR U33987 ( .A(n32663), .B(n32662), .Z(n32664) );
  NANDN U33988 ( .A(n32646), .B(n32645), .Z(n32650) );
  NAND U33989 ( .A(n32648), .B(n32647), .Z(n32649) );
  NAND U33990 ( .A(n32650), .B(n32649), .Z(n32665) );
  XNOR U33991 ( .A(n32664), .B(n32665), .Z(n32656) );
  XNOR U33992 ( .A(n32657), .B(n32656), .Z(n32658) );
  XNOR U33993 ( .A(n32659), .B(n32658), .Z(n32688) );
  XNOR U33994 ( .A(sreg[1788]), .B(n32688), .Z(n32690) );
  NANDN U33995 ( .A(sreg[1787]), .B(n32651), .Z(n32655) );
  NAND U33996 ( .A(n32653), .B(n32652), .Z(n32654) );
  NAND U33997 ( .A(n32655), .B(n32654), .Z(n32689) );
  XNOR U33998 ( .A(n32690), .B(n32689), .Z(c[1788]) );
  NANDN U33999 ( .A(n32657), .B(n32656), .Z(n32661) );
  NANDN U34000 ( .A(n32659), .B(n32658), .Z(n32660) );
  AND U34001 ( .A(n32661), .B(n32660), .Z(n32696) );
  NANDN U34002 ( .A(n32663), .B(n32662), .Z(n32667) );
  NANDN U34003 ( .A(n32665), .B(n32664), .Z(n32666) );
  AND U34004 ( .A(n32667), .B(n32666), .Z(n32694) );
  NAND U34005 ( .A(n42143), .B(n32668), .Z(n32670) );
  XNOR U34006 ( .A(a[767]), .B(n4181), .Z(n32705) );
  NAND U34007 ( .A(n42144), .B(n32705), .Z(n32669) );
  AND U34008 ( .A(n32670), .B(n32669), .Z(n32720) );
  XOR U34009 ( .A(a[771]), .B(n42012), .Z(n32708) );
  XNOR U34010 ( .A(n32720), .B(n32719), .Z(n32722) );
  XOR U34011 ( .A(a[769]), .B(n42085), .Z(n32709) );
  AND U34012 ( .A(a[765]), .B(b[7]), .Z(n32713) );
  XNOR U34013 ( .A(n32714), .B(n32713), .Z(n32715) );
  AND U34014 ( .A(a[773]), .B(b[0]), .Z(n32673) );
  XNOR U34015 ( .A(n32673), .B(n4071), .Z(n32675) );
  NANDN U34016 ( .A(b[0]), .B(a[772]), .Z(n32674) );
  NAND U34017 ( .A(n32675), .B(n32674), .Z(n32716) );
  XNOR U34018 ( .A(n32715), .B(n32716), .Z(n32721) );
  XOR U34019 ( .A(n32722), .B(n32721), .Z(n32700) );
  NANDN U34020 ( .A(n32677), .B(n32676), .Z(n32681) );
  NANDN U34021 ( .A(n32679), .B(n32678), .Z(n32680) );
  AND U34022 ( .A(n32681), .B(n32680), .Z(n32699) );
  XNOR U34023 ( .A(n32700), .B(n32699), .Z(n32701) );
  NANDN U34024 ( .A(n32683), .B(n32682), .Z(n32687) );
  NAND U34025 ( .A(n32685), .B(n32684), .Z(n32686) );
  NAND U34026 ( .A(n32687), .B(n32686), .Z(n32702) );
  XNOR U34027 ( .A(n32701), .B(n32702), .Z(n32693) );
  XNOR U34028 ( .A(n32694), .B(n32693), .Z(n32695) );
  XNOR U34029 ( .A(n32696), .B(n32695), .Z(n32725) );
  XNOR U34030 ( .A(sreg[1789]), .B(n32725), .Z(n32727) );
  NANDN U34031 ( .A(sreg[1788]), .B(n32688), .Z(n32692) );
  NAND U34032 ( .A(n32690), .B(n32689), .Z(n32691) );
  NAND U34033 ( .A(n32692), .B(n32691), .Z(n32726) );
  XNOR U34034 ( .A(n32727), .B(n32726), .Z(c[1789]) );
  NANDN U34035 ( .A(n32694), .B(n32693), .Z(n32698) );
  NANDN U34036 ( .A(n32696), .B(n32695), .Z(n32697) );
  AND U34037 ( .A(n32698), .B(n32697), .Z(n32733) );
  NANDN U34038 ( .A(n32700), .B(n32699), .Z(n32704) );
  NANDN U34039 ( .A(n32702), .B(n32701), .Z(n32703) );
  AND U34040 ( .A(n32704), .B(n32703), .Z(n32731) );
  NAND U34041 ( .A(n42143), .B(n32705), .Z(n32707) );
  XNOR U34042 ( .A(a[768]), .B(n4181), .Z(n32742) );
  NAND U34043 ( .A(n42144), .B(n32742), .Z(n32706) );
  AND U34044 ( .A(n32707), .B(n32706), .Z(n32757) );
  XOR U34045 ( .A(a[772]), .B(n42012), .Z(n32745) );
  XNOR U34046 ( .A(n32757), .B(n32756), .Z(n32759) );
  XOR U34047 ( .A(a[770]), .B(n42085), .Z(n32746) );
  AND U34048 ( .A(a[766]), .B(b[7]), .Z(n32750) );
  XNOR U34049 ( .A(n32751), .B(n32750), .Z(n32752) );
  AND U34050 ( .A(a[774]), .B(b[0]), .Z(n32710) );
  XNOR U34051 ( .A(n32710), .B(n4071), .Z(n32712) );
  NANDN U34052 ( .A(b[0]), .B(a[773]), .Z(n32711) );
  NAND U34053 ( .A(n32712), .B(n32711), .Z(n32753) );
  XNOR U34054 ( .A(n32752), .B(n32753), .Z(n32758) );
  XOR U34055 ( .A(n32759), .B(n32758), .Z(n32737) );
  NANDN U34056 ( .A(n32714), .B(n32713), .Z(n32718) );
  NANDN U34057 ( .A(n32716), .B(n32715), .Z(n32717) );
  AND U34058 ( .A(n32718), .B(n32717), .Z(n32736) );
  XNOR U34059 ( .A(n32737), .B(n32736), .Z(n32738) );
  NANDN U34060 ( .A(n32720), .B(n32719), .Z(n32724) );
  NAND U34061 ( .A(n32722), .B(n32721), .Z(n32723) );
  NAND U34062 ( .A(n32724), .B(n32723), .Z(n32739) );
  XNOR U34063 ( .A(n32738), .B(n32739), .Z(n32730) );
  XNOR U34064 ( .A(n32731), .B(n32730), .Z(n32732) );
  XNOR U34065 ( .A(n32733), .B(n32732), .Z(n32762) );
  XNOR U34066 ( .A(sreg[1790]), .B(n32762), .Z(n32764) );
  NANDN U34067 ( .A(sreg[1789]), .B(n32725), .Z(n32729) );
  NAND U34068 ( .A(n32727), .B(n32726), .Z(n32728) );
  NAND U34069 ( .A(n32729), .B(n32728), .Z(n32763) );
  XNOR U34070 ( .A(n32764), .B(n32763), .Z(c[1790]) );
  NANDN U34071 ( .A(n32731), .B(n32730), .Z(n32735) );
  NANDN U34072 ( .A(n32733), .B(n32732), .Z(n32734) );
  AND U34073 ( .A(n32735), .B(n32734), .Z(n32770) );
  NANDN U34074 ( .A(n32737), .B(n32736), .Z(n32741) );
  NANDN U34075 ( .A(n32739), .B(n32738), .Z(n32740) );
  AND U34076 ( .A(n32741), .B(n32740), .Z(n32768) );
  NAND U34077 ( .A(n42143), .B(n32742), .Z(n32744) );
  XNOR U34078 ( .A(a[769]), .B(n4181), .Z(n32779) );
  NAND U34079 ( .A(n42144), .B(n32779), .Z(n32743) );
  AND U34080 ( .A(n32744), .B(n32743), .Z(n32794) );
  XOR U34081 ( .A(a[773]), .B(n42012), .Z(n32782) );
  XNOR U34082 ( .A(n32794), .B(n32793), .Z(n32796) );
  XOR U34083 ( .A(a[771]), .B(n42085), .Z(n32783) );
  AND U34084 ( .A(a[767]), .B(b[7]), .Z(n32787) );
  XNOR U34085 ( .A(n32788), .B(n32787), .Z(n32789) );
  AND U34086 ( .A(a[775]), .B(b[0]), .Z(n32747) );
  XNOR U34087 ( .A(n32747), .B(n4071), .Z(n32749) );
  NANDN U34088 ( .A(b[0]), .B(a[774]), .Z(n32748) );
  NAND U34089 ( .A(n32749), .B(n32748), .Z(n32790) );
  XNOR U34090 ( .A(n32789), .B(n32790), .Z(n32795) );
  XOR U34091 ( .A(n32796), .B(n32795), .Z(n32774) );
  NANDN U34092 ( .A(n32751), .B(n32750), .Z(n32755) );
  NANDN U34093 ( .A(n32753), .B(n32752), .Z(n32754) );
  AND U34094 ( .A(n32755), .B(n32754), .Z(n32773) );
  XNOR U34095 ( .A(n32774), .B(n32773), .Z(n32775) );
  NANDN U34096 ( .A(n32757), .B(n32756), .Z(n32761) );
  NAND U34097 ( .A(n32759), .B(n32758), .Z(n32760) );
  NAND U34098 ( .A(n32761), .B(n32760), .Z(n32776) );
  XNOR U34099 ( .A(n32775), .B(n32776), .Z(n32767) );
  XNOR U34100 ( .A(n32768), .B(n32767), .Z(n32769) );
  XNOR U34101 ( .A(n32770), .B(n32769), .Z(n32799) );
  XNOR U34102 ( .A(sreg[1791]), .B(n32799), .Z(n32801) );
  NANDN U34103 ( .A(sreg[1790]), .B(n32762), .Z(n32766) );
  NAND U34104 ( .A(n32764), .B(n32763), .Z(n32765) );
  NAND U34105 ( .A(n32766), .B(n32765), .Z(n32800) );
  XNOR U34106 ( .A(n32801), .B(n32800), .Z(c[1791]) );
  NANDN U34107 ( .A(n32768), .B(n32767), .Z(n32772) );
  NANDN U34108 ( .A(n32770), .B(n32769), .Z(n32771) );
  AND U34109 ( .A(n32772), .B(n32771), .Z(n32807) );
  NANDN U34110 ( .A(n32774), .B(n32773), .Z(n32778) );
  NANDN U34111 ( .A(n32776), .B(n32775), .Z(n32777) );
  AND U34112 ( .A(n32778), .B(n32777), .Z(n32805) );
  NAND U34113 ( .A(n42143), .B(n32779), .Z(n32781) );
  XNOR U34114 ( .A(a[770]), .B(n4181), .Z(n32816) );
  NAND U34115 ( .A(n42144), .B(n32816), .Z(n32780) );
  AND U34116 ( .A(n32781), .B(n32780), .Z(n32831) );
  XOR U34117 ( .A(a[774]), .B(n42012), .Z(n32819) );
  XNOR U34118 ( .A(n32831), .B(n32830), .Z(n32833) );
  XOR U34119 ( .A(a[772]), .B(n42085), .Z(n32820) );
  AND U34120 ( .A(a[768]), .B(b[7]), .Z(n32824) );
  XNOR U34121 ( .A(n32825), .B(n32824), .Z(n32826) );
  AND U34122 ( .A(a[776]), .B(b[0]), .Z(n32784) );
  XNOR U34123 ( .A(n32784), .B(n4071), .Z(n32786) );
  NANDN U34124 ( .A(b[0]), .B(a[775]), .Z(n32785) );
  NAND U34125 ( .A(n32786), .B(n32785), .Z(n32827) );
  XNOR U34126 ( .A(n32826), .B(n32827), .Z(n32832) );
  XOR U34127 ( .A(n32833), .B(n32832), .Z(n32811) );
  NANDN U34128 ( .A(n32788), .B(n32787), .Z(n32792) );
  NANDN U34129 ( .A(n32790), .B(n32789), .Z(n32791) );
  AND U34130 ( .A(n32792), .B(n32791), .Z(n32810) );
  XNOR U34131 ( .A(n32811), .B(n32810), .Z(n32812) );
  NANDN U34132 ( .A(n32794), .B(n32793), .Z(n32798) );
  NAND U34133 ( .A(n32796), .B(n32795), .Z(n32797) );
  NAND U34134 ( .A(n32798), .B(n32797), .Z(n32813) );
  XNOR U34135 ( .A(n32812), .B(n32813), .Z(n32804) );
  XNOR U34136 ( .A(n32805), .B(n32804), .Z(n32806) );
  XNOR U34137 ( .A(n32807), .B(n32806), .Z(n32836) );
  XNOR U34138 ( .A(sreg[1792]), .B(n32836), .Z(n32838) );
  NANDN U34139 ( .A(sreg[1791]), .B(n32799), .Z(n32803) );
  NAND U34140 ( .A(n32801), .B(n32800), .Z(n32802) );
  NAND U34141 ( .A(n32803), .B(n32802), .Z(n32837) );
  XNOR U34142 ( .A(n32838), .B(n32837), .Z(c[1792]) );
  NANDN U34143 ( .A(n32805), .B(n32804), .Z(n32809) );
  NANDN U34144 ( .A(n32807), .B(n32806), .Z(n32808) );
  AND U34145 ( .A(n32809), .B(n32808), .Z(n32844) );
  NANDN U34146 ( .A(n32811), .B(n32810), .Z(n32815) );
  NANDN U34147 ( .A(n32813), .B(n32812), .Z(n32814) );
  AND U34148 ( .A(n32815), .B(n32814), .Z(n32842) );
  NAND U34149 ( .A(n42143), .B(n32816), .Z(n32818) );
  XNOR U34150 ( .A(a[771]), .B(n4182), .Z(n32853) );
  NAND U34151 ( .A(n42144), .B(n32853), .Z(n32817) );
  AND U34152 ( .A(n32818), .B(n32817), .Z(n32868) );
  XOR U34153 ( .A(a[775]), .B(n42012), .Z(n32856) );
  XNOR U34154 ( .A(n32868), .B(n32867), .Z(n32870) );
  XOR U34155 ( .A(a[773]), .B(n42085), .Z(n32857) );
  AND U34156 ( .A(a[769]), .B(b[7]), .Z(n32861) );
  XNOR U34157 ( .A(n32862), .B(n32861), .Z(n32863) );
  AND U34158 ( .A(a[777]), .B(b[0]), .Z(n32821) );
  XNOR U34159 ( .A(n32821), .B(n4071), .Z(n32823) );
  NANDN U34160 ( .A(b[0]), .B(a[776]), .Z(n32822) );
  NAND U34161 ( .A(n32823), .B(n32822), .Z(n32864) );
  XNOR U34162 ( .A(n32863), .B(n32864), .Z(n32869) );
  XOR U34163 ( .A(n32870), .B(n32869), .Z(n32848) );
  NANDN U34164 ( .A(n32825), .B(n32824), .Z(n32829) );
  NANDN U34165 ( .A(n32827), .B(n32826), .Z(n32828) );
  AND U34166 ( .A(n32829), .B(n32828), .Z(n32847) );
  XNOR U34167 ( .A(n32848), .B(n32847), .Z(n32849) );
  NANDN U34168 ( .A(n32831), .B(n32830), .Z(n32835) );
  NAND U34169 ( .A(n32833), .B(n32832), .Z(n32834) );
  NAND U34170 ( .A(n32835), .B(n32834), .Z(n32850) );
  XNOR U34171 ( .A(n32849), .B(n32850), .Z(n32841) );
  XNOR U34172 ( .A(n32842), .B(n32841), .Z(n32843) );
  XNOR U34173 ( .A(n32844), .B(n32843), .Z(n32873) );
  XNOR U34174 ( .A(sreg[1793]), .B(n32873), .Z(n32875) );
  NANDN U34175 ( .A(sreg[1792]), .B(n32836), .Z(n32840) );
  NAND U34176 ( .A(n32838), .B(n32837), .Z(n32839) );
  NAND U34177 ( .A(n32840), .B(n32839), .Z(n32874) );
  XNOR U34178 ( .A(n32875), .B(n32874), .Z(c[1793]) );
  NANDN U34179 ( .A(n32842), .B(n32841), .Z(n32846) );
  NANDN U34180 ( .A(n32844), .B(n32843), .Z(n32845) );
  AND U34181 ( .A(n32846), .B(n32845), .Z(n32881) );
  NANDN U34182 ( .A(n32848), .B(n32847), .Z(n32852) );
  NANDN U34183 ( .A(n32850), .B(n32849), .Z(n32851) );
  AND U34184 ( .A(n32852), .B(n32851), .Z(n32879) );
  NAND U34185 ( .A(n42143), .B(n32853), .Z(n32855) );
  XNOR U34186 ( .A(a[772]), .B(n4182), .Z(n32890) );
  NAND U34187 ( .A(n42144), .B(n32890), .Z(n32854) );
  AND U34188 ( .A(n32855), .B(n32854), .Z(n32905) );
  XOR U34189 ( .A(a[776]), .B(n42012), .Z(n32893) );
  XNOR U34190 ( .A(n32905), .B(n32904), .Z(n32907) );
  XOR U34191 ( .A(a[774]), .B(n42085), .Z(n32897) );
  AND U34192 ( .A(a[770]), .B(b[7]), .Z(n32898) );
  XNOR U34193 ( .A(n32899), .B(n32898), .Z(n32900) );
  AND U34194 ( .A(a[778]), .B(b[0]), .Z(n32858) );
  XNOR U34195 ( .A(n32858), .B(n4071), .Z(n32860) );
  NANDN U34196 ( .A(b[0]), .B(a[777]), .Z(n32859) );
  NAND U34197 ( .A(n32860), .B(n32859), .Z(n32901) );
  XNOR U34198 ( .A(n32900), .B(n32901), .Z(n32906) );
  XOR U34199 ( .A(n32907), .B(n32906), .Z(n32885) );
  NANDN U34200 ( .A(n32862), .B(n32861), .Z(n32866) );
  NANDN U34201 ( .A(n32864), .B(n32863), .Z(n32865) );
  AND U34202 ( .A(n32866), .B(n32865), .Z(n32884) );
  XNOR U34203 ( .A(n32885), .B(n32884), .Z(n32886) );
  NANDN U34204 ( .A(n32868), .B(n32867), .Z(n32872) );
  NAND U34205 ( .A(n32870), .B(n32869), .Z(n32871) );
  NAND U34206 ( .A(n32872), .B(n32871), .Z(n32887) );
  XNOR U34207 ( .A(n32886), .B(n32887), .Z(n32878) );
  XNOR U34208 ( .A(n32879), .B(n32878), .Z(n32880) );
  XNOR U34209 ( .A(n32881), .B(n32880), .Z(n32910) );
  XNOR U34210 ( .A(sreg[1794]), .B(n32910), .Z(n32912) );
  NANDN U34211 ( .A(sreg[1793]), .B(n32873), .Z(n32877) );
  NAND U34212 ( .A(n32875), .B(n32874), .Z(n32876) );
  NAND U34213 ( .A(n32877), .B(n32876), .Z(n32911) );
  XNOR U34214 ( .A(n32912), .B(n32911), .Z(c[1794]) );
  NANDN U34215 ( .A(n32879), .B(n32878), .Z(n32883) );
  NANDN U34216 ( .A(n32881), .B(n32880), .Z(n32882) );
  AND U34217 ( .A(n32883), .B(n32882), .Z(n32918) );
  NANDN U34218 ( .A(n32885), .B(n32884), .Z(n32889) );
  NANDN U34219 ( .A(n32887), .B(n32886), .Z(n32888) );
  AND U34220 ( .A(n32889), .B(n32888), .Z(n32916) );
  NAND U34221 ( .A(n42143), .B(n32890), .Z(n32892) );
  XNOR U34222 ( .A(a[773]), .B(n4182), .Z(n32927) );
  NAND U34223 ( .A(n42144), .B(n32927), .Z(n32891) );
  AND U34224 ( .A(n32892), .B(n32891), .Z(n32942) );
  XOR U34225 ( .A(a[777]), .B(n42012), .Z(n32930) );
  XNOR U34226 ( .A(n32942), .B(n32941), .Z(n32944) );
  AND U34227 ( .A(a[779]), .B(b[0]), .Z(n32894) );
  XNOR U34228 ( .A(n32894), .B(n4071), .Z(n32896) );
  NANDN U34229 ( .A(b[0]), .B(a[778]), .Z(n32895) );
  NAND U34230 ( .A(n32896), .B(n32895), .Z(n32938) );
  XOR U34231 ( .A(a[775]), .B(n42085), .Z(n32934) );
  AND U34232 ( .A(a[771]), .B(b[7]), .Z(n32935) );
  XNOR U34233 ( .A(n32936), .B(n32935), .Z(n32937) );
  XNOR U34234 ( .A(n32938), .B(n32937), .Z(n32943) );
  XOR U34235 ( .A(n32944), .B(n32943), .Z(n32922) );
  NANDN U34236 ( .A(n32899), .B(n32898), .Z(n32903) );
  NANDN U34237 ( .A(n32901), .B(n32900), .Z(n32902) );
  AND U34238 ( .A(n32903), .B(n32902), .Z(n32921) );
  XNOR U34239 ( .A(n32922), .B(n32921), .Z(n32923) );
  NANDN U34240 ( .A(n32905), .B(n32904), .Z(n32909) );
  NAND U34241 ( .A(n32907), .B(n32906), .Z(n32908) );
  NAND U34242 ( .A(n32909), .B(n32908), .Z(n32924) );
  XNOR U34243 ( .A(n32923), .B(n32924), .Z(n32915) );
  XNOR U34244 ( .A(n32916), .B(n32915), .Z(n32917) );
  XNOR U34245 ( .A(n32918), .B(n32917), .Z(n32947) );
  XNOR U34246 ( .A(sreg[1795]), .B(n32947), .Z(n32949) );
  NANDN U34247 ( .A(sreg[1794]), .B(n32910), .Z(n32914) );
  NAND U34248 ( .A(n32912), .B(n32911), .Z(n32913) );
  NAND U34249 ( .A(n32914), .B(n32913), .Z(n32948) );
  XNOR U34250 ( .A(n32949), .B(n32948), .Z(c[1795]) );
  NANDN U34251 ( .A(n32916), .B(n32915), .Z(n32920) );
  NANDN U34252 ( .A(n32918), .B(n32917), .Z(n32919) );
  AND U34253 ( .A(n32920), .B(n32919), .Z(n32955) );
  NANDN U34254 ( .A(n32922), .B(n32921), .Z(n32926) );
  NANDN U34255 ( .A(n32924), .B(n32923), .Z(n32925) );
  AND U34256 ( .A(n32926), .B(n32925), .Z(n32953) );
  NAND U34257 ( .A(n42143), .B(n32927), .Z(n32929) );
  XNOR U34258 ( .A(a[774]), .B(n4182), .Z(n32964) );
  NAND U34259 ( .A(n42144), .B(n32964), .Z(n32928) );
  AND U34260 ( .A(n32929), .B(n32928), .Z(n32979) );
  XOR U34261 ( .A(a[778]), .B(n42012), .Z(n32967) );
  XNOR U34262 ( .A(n32979), .B(n32978), .Z(n32981) );
  AND U34263 ( .A(a[780]), .B(b[0]), .Z(n32931) );
  XNOR U34264 ( .A(n32931), .B(n4071), .Z(n32933) );
  NANDN U34265 ( .A(b[0]), .B(a[779]), .Z(n32932) );
  NAND U34266 ( .A(n32933), .B(n32932), .Z(n32975) );
  XOR U34267 ( .A(a[776]), .B(n42085), .Z(n32971) );
  AND U34268 ( .A(a[772]), .B(b[7]), .Z(n32972) );
  XNOR U34269 ( .A(n32973), .B(n32972), .Z(n32974) );
  XNOR U34270 ( .A(n32975), .B(n32974), .Z(n32980) );
  XOR U34271 ( .A(n32981), .B(n32980), .Z(n32959) );
  NANDN U34272 ( .A(n32936), .B(n32935), .Z(n32940) );
  NANDN U34273 ( .A(n32938), .B(n32937), .Z(n32939) );
  AND U34274 ( .A(n32940), .B(n32939), .Z(n32958) );
  XNOR U34275 ( .A(n32959), .B(n32958), .Z(n32960) );
  NANDN U34276 ( .A(n32942), .B(n32941), .Z(n32946) );
  NAND U34277 ( .A(n32944), .B(n32943), .Z(n32945) );
  NAND U34278 ( .A(n32946), .B(n32945), .Z(n32961) );
  XNOR U34279 ( .A(n32960), .B(n32961), .Z(n32952) );
  XNOR U34280 ( .A(n32953), .B(n32952), .Z(n32954) );
  XNOR U34281 ( .A(n32955), .B(n32954), .Z(n32984) );
  XNOR U34282 ( .A(sreg[1796]), .B(n32984), .Z(n32986) );
  NANDN U34283 ( .A(sreg[1795]), .B(n32947), .Z(n32951) );
  NAND U34284 ( .A(n32949), .B(n32948), .Z(n32950) );
  NAND U34285 ( .A(n32951), .B(n32950), .Z(n32985) );
  XNOR U34286 ( .A(n32986), .B(n32985), .Z(c[1796]) );
  NANDN U34287 ( .A(n32953), .B(n32952), .Z(n32957) );
  NANDN U34288 ( .A(n32955), .B(n32954), .Z(n32956) );
  AND U34289 ( .A(n32957), .B(n32956), .Z(n32992) );
  NANDN U34290 ( .A(n32959), .B(n32958), .Z(n32963) );
  NANDN U34291 ( .A(n32961), .B(n32960), .Z(n32962) );
  AND U34292 ( .A(n32963), .B(n32962), .Z(n32990) );
  NAND U34293 ( .A(n42143), .B(n32964), .Z(n32966) );
  XNOR U34294 ( .A(a[775]), .B(n4182), .Z(n33001) );
  NAND U34295 ( .A(n42144), .B(n33001), .Z(n32965) );
  AND U34296 ( .A(n32966), .B(n32965), .Z(n33016) );
  XOR U34297 ( .A(a[779]), .B(n42012), .Z(n33004) );
  XNOR U34298 ( .A(n33016), .B(n33015), .Z(n33018) );
  AND U34299 ( .A(a[781]), .B(b[0]), .Z(n32968) );
  XNOR U34300 ( .A(n32968), .B(n4071), .Z(n32970) );
  NANDN U34301 ( .A(b[0]), .B(a[780]), .Z(n32969) );
  NAND U34302 ( .A(n32970), .B(n32969), .Z(n33012) );
  XOR U34303 ( .A(a[777]), .B(n42085), .Z(n33008) );
  AND U34304 ( .A(a[773]), .B(b[7]), .Z(n33009) );
  XNOR U34305 ( .A(n33010), .B(n33009), .Z(n33011) );
  XNOR U34306 ( .A(n33012), .B(n33011), .Z(n33017) );
  XOR U34307 ( .A(n33018), .B(n33017), .Z(n32996) );
  NANDN U34308 ( .A(n32973), .B(n32972), .Z(n32977) );
  NANDN U34309 ( .A(n32975), .B(n32974), .Z(n32976) );
  AND U34310 ( .A(n32977), .B(n32976), .Z(n32995) );
  XNOR U34311 ( .A(n32996), .B(n32995), .Z(n32997) );
  NANDN U34312 ( .A(n32979), .B(n32978), .Z(n32983) );
  NAND U34313 ( .A(n32981), .B(n32980), .Z(n32982) );
  NAND U34314 ( .A(n32983), .B(n32982), .Z(n32998) );
  XNOR U34315 ( .A(n32997), .B(n32998), .Z(n32989) );
  XNOR U34316 ( .A(n32990), .B(n32989), .Z(n32991) );
  XNOR U34317 ( .A(n32992), .B(n32991), .Z(n33021) );
  XNOR U34318 ( .A(sreg[1797]), .B(n33021), .Z(n33023) );
  NANDN U34319 ( .A(sreg[1796]), .B(n32984), .Z(n32988) );
  NAND U34320 ( .A(n32986), .B(n32985), .Z(n32987) );
  NAND U34321 ( .A(n32988), .B(n32987), .Z(n33022) );
  XNOR U34322 ( .A(n33023), .B(n33022), .Z(c[1797]) );
  NANDN U34323 ( .A(n32990), .B(n32989), .Z(n32994) );
  NANDN U34324 ( .A(n32992), .B(n32991), .Z(n32993) );
  AND U34325 ( .A(n32994), .B(n32993), .Z(n33029) );
  NANDN U34326 ( .A(n32996), .B(n32995), .Z(n33000) );
  NANDN U34327 ( .A(n32998), .B(n32997), .Z(n32999) );
  AND U34328 ( .A(n33000), .B(n32999), .Z(n33027) );
  NAND U34329 ( .A(n42143), .B(n33001), .Z(n33003) );
  XNOR U34330 ( .A(a[776]), .B(n4182), .Z(n33038) );
  NAND U34331 ( .A(n42144), .B(n33038), .Z(n33002) );
  AND U34332 ( .A(n33003), .B(n33002), .Z(n33053) );
  XOR U34333 ( .A(a[780]), .B(n42012), .Z(n33041) );
  XNOR U34334 ( .A(n33053), .B(n33052), .Z(n33055) );
  AND U34335 ( .A(a[782]), .B(b[0]), .Z(n33005) );
  XNOR U34336 ( .A(n33005), .B(n4071), .Z(n33007) );
  NANDN U34337 ( .A(b[0]), .B(a[781]), .Z(n33006) );
  NAND U34338 ( .A(n33007), .B(n33006), .Z(n33049) );
  XOR U34339 ( .A(a[778]), .B(n42085), .Z(n33045) );
  AND U34340 ( .A(a[774]), .B(b[7]), .Z(n33046) );
  XNOR U34341 ( .A(n33047), .B(n33046), .Z(n33048) );
  XNOR U34342 ( .A(n33049), .B(n33048), .Z(n33054) );
  XOR U34343 ( .A(n33055), .B(n33054), .Z(n33033) );
  NANDN U34344 ( .A(n33010), .B(n33009), .Z(n33014) );
  NANDN U34345 ( .A(n33012), .B(n33011), .Z(n33013) );
  AND U34346 ( .A(n33014), .B(n33013), .Z(n33032) );
  XNOR U34347 ( .A(n33033), .B(n33032), .Z(n33034) );
  NANDN U34348 ( .A(n33016), .B(n33015), .Z(n33020) );
  NAND U34349 ( .A(n33018), .B(n33017), .Z(n33019) );
  NAND U34350 ( .A(n33020), .B(n33019), .Z(n33035) );
  XNOR U34351 ( .A(n33034), .B(n33035), .Z(n33026) );
  XNOR U34352 ( .A(n33027), .B(n33026), .Z(n33028) );
  XNOR U34353 ( .A(n33029), .B(n33028), .Z(n33058) );
  XNOR U34354 ( .A(sreg[1798]), .B(n33058), .Z(n33060) );
  NANDN U34355 ( .A(sreg[1797]), .B(n33021), .Z(n33025) );
  NAND U34356 ( .A(n33023), .B(n33022), .Z(n33024) );
  NAND U34357 ( .A(n33025), .B(n33024), .Z(n33059) );
  XNOR U34358 ( .A(n33060), .B(n33059), .Z(c[1798]) );
  NANDN U34359 ( .A(n33027), .B(n33026), .Z(n33031) );
  NANDN U34360 ( .A(n33029), .B(n33028), .Z(n33030) );
  AND U34361 ( .A(n33031), .B(n33030), .Z(n33066) );
  NANDN U34362 ( .A(n33033), .B(n33032), .Z(n33037) );
  NANDN U34363 ( .A(n33035), .B(n33034), .Z(n33036) );
  AND U34364 ( .A(n33037), .B(n33036), .Z(n33064) );
  NAND U34365 ( .A(n42143), .B(n33038), .Z(n33040) );
  XNOR U34366 ( .A(a[777]), .B(n4182), .Z(n33075) );
  NAND U34367 ( .A(n42144), .B(n33075), .Z(n33039) );
  AND U34368 ( .A(n33040), .B(n33039), .Z(n33090) );
  XOR U34369 ( .A(a[781]), .B(n42012), .Z(n33078) );
  XNOR U34370 ( .A(n33090), .B(n33089), .Z(n33092) );
  AND U34371 ( .A(a[783]), .B(b[0]), .Z(n33042) );
  XNOR U34372 ( .A(n33042), .B(n4071), .Z(n33044) );
  NANDN U34373 ( .A(b[0]), .B(a[782]), .Z(n33043) );
  NAND U34374 ( .A(n33044), .B(n33043), .Z(n33086) );
  XOR U34375 ( .A(a[779]), .B(n42085), .Z(n33082) );
  AND U34376 ( .A(a[775]), .B(b[7]), .Z(n33083) );
  XNOR U34377 ( .A(n33084), .B(n33083), .Z(n33085) );
  XNOR U34378 ( .A(n33086), .B(n33085), .Z(n33091) );
  XOR U34379 ( .A(n33092), .B(n33091), .Z(n33070) );
  NANDN U34380 ( .A(n33047), .B(n33046), .Z(n33051) );
  NANDN U34381 ( .A(n33049), .B(n33048), .Z(n33050) );
  AND U34382 ( .A(n33051), .B(n33050), .Z(n33069) );
  XNOR U34383 ( .A(n33070), .B(n33069), .Z(n33071) );
  NANDN U34384 ( .A(n33053), .B(n33052), .Z(n33057) );
  NAND U34385 ( .A(n33055), .B(n33054), .Z(n33056) );
  NAND U34386 ( .A(n33057), .B(n33056), .Z(n33072) );
  XNOR U34387 ( .A(n33071), .B(n33072), .Z(n33063) );
  XNOR U34388 ( .A(n33064), .B(n33063), .Z(n33065) );
  XNOR U34389 ( .A(n33066), .B(n33065), .Z(n33095) );
  XNOR U34390 ( .A(sreg[1799]), .B(n33095), .Z(n33097) );
  NANDN U34391 ( .A(sreg[1798]), .B(n33058), .Z(n33062) );
  NAND U34392 ( .A(n33060), .B(n33059), .Z(n33061) );
  NAND U34393 ( .A(n33062), .B(n33061), .Z(n33096) );
  XNOR U34394 ( .A(n33097), .B(n33096), .Z(c[1799]) );
  NANDN U34395 ( .A(n33064), .B(n33063), .Z(n33068) );
  NANDN U34396 ( .A(n33066), .B(n33065), .Z(n33067) );
  AND U34397 ( .A(n33068), .B(n33067), .Z(n33103) );
  NANDN U34398 ( .A(n33070), .B(n33069), .Z(n33074) );
  NANDN U34399 ( .A(n33072), .B(n33071), .Z(n33073) );
  AND U34400 ( .A(n33074), .B(n33073), .Z(n33101) );
  NAND U34401 ( .A(n42143), .B(n33075), .Z(n33077) );
  XNOR U34402 ( .A(a[778]), .B(n4183), .Z(n33112) );
  NAND U34403 ( .A(n42144), .B(n33112), .Z(n33076) );
  AND U34404 ( .A(n33077), .B(n33076), .Z(n33127) );
  XOR U34405 ( .A(a[782]), .B(n42012), .Z(n33115) );
  XNOR U34406 ( .A(n33127), .B(n33126), .Z(n33129) );
  AND U34407 ( .A(a[784]), .B(b[0]), .Z(n33079) );
  XNOR U34408 ( .A(n33079), .B(n4071), .Z(n33081) );
  NANDN U34409 ( .A(b[0]), .B(a[783]), .Z(n33080) );
  NAND U34410 ( .A(n33081), .B(n33080), .Z(n33123) );
  XOR U34411 ( .A(a[780]), .B(n42085), .Z(n33116) );
  AND U34412 ( .A(a[776]), .B(b[7]), .Z(n33120) );
  XNOR U34413 ( .A(n33121), .B(n33120), .Z(n33122) );
  XNOR U34414 ( .A(n33123), .B(n33122), .Z(n33128) );
  XOR U34415 ( .A(n33129), .B(n33128), .Z(n33107) );
  NANDN U34416 ( .A(n33084), .B(n33083), .Z(n33088) );
  NANDN U34417 ( .A(n33086), .B(n33085), .Z(n33087) );
  AND U34418 ( .A(n33088), .B(n33087), .Z(n33106) );
  XNOR U34419 ( .A(n33107), .B(n33106), .Z(n33108) );
  NANDN U34420 ( .A(n33090), .B(n33089), .Z(n33094) );
  NAND U34421 ( .A(n33092), .B(n33091), .Z(n33093) );
  NAND U34422 ( .A(n33094), .B(n33093), .Z(n33109) );
  XNOR U34423 ( .A(n33108), .B(n33109), .Z(n33100) );
  XNOR U34424 ( .A(n33101), .B(n33100), .Z(n33102) );
  XNOR U34425 ( .A(n33103), .B(n33102), .Z(n33132) );
  XNOR U34426 ( .A(sreg[1800]), .B(n33132), .Z(n33134) );
  NANDN U34427 ( .A(sreg[1799]), .B(n33095), .Z(n33099) );
  NAND U34428 ( .A(n33097), .B(n33096), .Z(n33098) );
  NAND U34429 ( .A(n33099), .B(n33098), .Z(n33133) );
  XNOR U34430 ( .A(n33134), .B(n33133), .Z(c[1800]) );
  NANDN U34431 ( .A(n33101), .B(n33100), .Z(n33105) );
  NANDN U34432 ( .A(n33103), .B(n33102), .Z(n33104) );
  AND U34433 ( .A(n33105), .B(n33104), .Z(n33140) );
  NANDN U34434 ( .A(n33107), .B(n33106), .Z(n33111) );
  NANDN U34435 ( .A(n33109), .B(n33108), .Z(n33110) );
  AND U34436 ( .A(n33111), .B(n33110), .Z(n33138) );
  NAND U34437 ( .A(n42143), .B(n33112), .Z(n33114) );
  XNOR U34438 ( .A(a[779]), .B(n4183), .Z(n33149) );
  NAND U34439 ( .A(n42144), .B(n33149), .Z(n33113) );
  AND U34440 ( .A(n33114), .B(n33113), .Z(n33164) );
  XOR U34441 ( .A(a[783]), .B(n42012), .Z(n33152) );
  XNOR U34442 ( .A(n33164), .B(n33163), .Z(n33166) );
  XOR U34443 ( .A(a[781]), .B(n42085), .Z(n33156) );
  AND U34444 ( .A(a[777]), .B(b[7]), .Z(n33157) );
  XNOR U34445 ( .A(n33158), .B(n33157), .Z(n33159) );
  AND U34446 ( .A(a[785]), .B(b[0]), .Z(n33117) );
  XNOR U34447 ( .A(n33117), .B(n4071), .Z(n33119) );
  NANDN U34448 ( .A(b[0]), .B(a[784]), .Z(n33118) );
  NAND U34449 ( .A(n33119), .B(n33118), .Z(n33160) );
  XNOR U34450 ( .A(n33159), .B(n33160), .Z(n33165) );
  XOR U34451 ( .A(n33166), .B(n33165), .Z(n33144) );
  NANDN U34452 ( .A(n33121), .B(n33120), .Z(n33125) );
  NANDN U34453 ( .A(n33123), .B(n33122), .Z(n33124) );
  AND U34454 ( .A(n33125), .B(n33124), .Z(n33143) );
  XNOR U34455 ( .A(n33144), .B(n33143), .Z(n33145) );
  NANDN U34456 ( .A(n33127), .B(n33126), .Z(n33131) );
  NAND U34457 ( .A(n33129), .B(n33128), .Z(n33130) );
  NAND U34458 ( .A(n33131), .B(n33130), .Z(n33146) );
  XNOR U34459 ( .A(n33145), .B(n33146), .Z(n33137) );
  XNOR U34460 ( .A(n33138), .B(n33137), .Z(n33139) );
  XNOR U34461 ( .A(n33140), .B(n33139), .Z(n33169) );
  XNOR U34462 ( .A(sreg[1801]), .B(n33169), .Z(n33171) );
  NANDN U34463 ( .A(sreg[1800]), .B(n33132), .Z(n33136) );
  NAND U34464 ( .A(n33134), .B(n33133), .Z(n33135) );
  NAND U34465 ( .A(n33136), .B(n33135), .Z(n33170) );
  XNOR U34466 ( .A(n33171), .B(n33170), .Z(c[1801]) );
  NANDN U34467 ( .A(n33138), .B(n33137), .Z(n33142) );
  NANDN U34468 ( .A(n33140), .B(n33139), .Z(n33141) );
  AND U34469 ( .A(n33142), .B(n33141), .Z(n33177) );
  NANDN U34470 ( .A(n33144), .B(n33143), .Z(n33148) );
  NANDN U34471 ( .A(n33146), .B(n33145), .Z(n33147) );
  AND U34472 ( .A(n33148), .B(n33147), .Z(n33175) );
  NAND U34473 ( .A(n42143), .B(n33149), .Z(n33151) );
  XNOR U34474 ( .A(a[780]), .B(n4183), .Z(n33186) );
  NAND U34475 ( .A(n42144), .B(n33186), .Z(n33150) );
  AND U34476 ( .A(n33151), .B(n33150), .Z(n33201) );
  XOR U34477 ( .A(a[784]), .B(n42012), .Z(n33189) );
  XNOR U34478 ( .A(n33201), .B(n33200), .Z(n33203) );
  AND U34479 ( .A(a[786]), .B(b[0]), .Z(n33153) );
  XNOR U34480 ( .A(n33153), .B(n4071), .Z(n33155) );
  NANDN U34481 ( .A(b[0]), .B(a[785]), .Z(n33154) );
  NAND U34482 ( .A(n33155), .B(n33154), .Z(n33197) );
  XOR U34483 ( .A(a[782]), .B(n42085), .Z(n33190) );
  AND U34484 ( .A(a[778]), .B(b[7]), .Z(n33194) );
  XNOR U34485 ( .A(n33195), .B(n33194), .Z(n33196) );
  XNOR U34486 ( .A(n33197), .B(n33196), .Z(n33202) );
  XOR U34487 ( .A(n33203), .B(n33202), .Z(n33181) );
  NANDN U34488 ( .A(n33158), .B(n33157), .Z(n33162) );
  NANDN U34489 ( .A(n33160), .B(n33159), .Z(n33161) );
  AND U34490 ( .A(n33162), .B(n33161), .Z(n33180) );
  XNOR U34491 ( .A(n33181), .B(n33180), .Z(n33182) );
  NANDN U34492 ( .A(n33164), .B(n33163), .Z(n33168) );
  NAND U34493 ( .A(n33166), .B(n33165), .Z(n33167) );
  NAND U34494 ( .A(n33168), .B(n33167), .Z(n33183) );
  XNOR U34495 ( .A(n33182), .B(n33183), .Z(n33174) );
  XNOR U34496 ( .A(n33175), .B(n33174), .Z(n33176) );
  XNOR U34497 ( .A(n33177), .B(n33176), .Z(n33206) );
  XNOR U34498 ( .A(sreg[1802]), .B(n33206), .Z(n33208) );
  NANDN U34499 ( .A(sreg[1801]), .B(n33169), .Z(n33173) );
  NAND U34500 ( .A(n33171), .B(n33170), .Z(n33172) );
  NAND U34501 ( .A(n33173), .B(n33172), .Z(n33207) );
  XNOR U34502 ( .A(n33208), .B(n33207), .Z(c[1802]) );
  NANDN U34503 ( .A(n33175), .B(n33174), .Z(n33179) );
  NANDN U34504 ( .A(n33177), .B(n33176), .Z(n33178) );
  AND U34505 ( .A(n33179), .B(n33178), .Z(n33214) );
  NANDN U34506 ( .A(n33181), .B(n33180), .Z(n33185) );
  NANDN U34507 ( .A(n33183), .B(n33182), .Z(n33184) );
  AND U34508 ( .A(n33185), .B(n33184), .Z(n33212) );
  NAND U34509 ( .A(n42143), .B(n33186), .Z(n33188) );
  XNOR U34510 ( .A(a[781]), .B(n4183), .Z(n33223) );
  NAND U34511 ( .A(n42144), .B(n33223), .Z(n33187) );
  AND U34512 ( .A(n33188), .B(n33187), .Z(n33238) );
  XOR U34513 ( .A(a[785]), .B(n42012), .Z(n33226) );
  XNOR U34514 ( .A(n33238), .B(n33237), .Z(n33240) );
  XOR U34515 ( .A(a[783]), .B(n42085), .Z(n33227) );
  AND U34516 ( .A(a[779]), .B(b[7]), .Z(n33231) );
  XNOR U34517 ( .A(n33232), .B(n33231), .Z(n33233) );
  AND U34518 ( .A(a[787]), .B(b[0]), .Z(n33191) );
  XNOR U34519 ( .A(n33191), .B(n4071), .Z(n33193) );
  NANDN U34520 ( .A(b[0]), .B(a[786]), .Z(n33192) );
  NAND U34521 ( .A(n33193), .B(n33192), .Z(n33234) );
  XNOR U34522 ( .A(n33233), .B(n33234), .Z(n33239) );
  XOR U34523 ( .A(n33240), .B(n33239), .Z(n33218) );
  NANDN U34524 ( .A(n33195), .B(n33194), .Z(n33199) );
  NANDN U34525 ( .A(n33197), .B(n33196), .Z(n33198) );
  AND U34526 ( .A(n33199), .B(n33198), .Z(n33217) );
  XNOR U34527 ( .A(n33218), .B(n33217), .Z(n33219) );
  NANDN U34528 ( .A(n33201), .B(n33200), .Z(n33205) );
  NAND U34529 ( .A(n33203), .B(n33202), .Z(n33204) );
  NAND U34530 ( .A(n33205), .B(n33204), .Z(n33220) );
  XNOR U34531 ( .A(n33219), .B(n33220), .Z(n33211) );
  XNOR U34532 ( .A(n33212), .B(n33211), .Z(n33213) );
  XNOR U34533 ( .A(n33214), .B(n33213), .Z(n33243) );
  XNOR U34534 ( .A(sreg[1803]), .B(n33243), .Z(n33245) );
  NANDN U34535 ( .A(sreg[1802]), .B(n33206), .Z(n33210) );
  NAND U34536 ( .A(n33208), .B(n33207), .Z(n33209) );
  NAND U34537 ( .A(n33210), .B(n33209), .Z(n33244) );
  XNOR U34538 ( .A(n33245), .B(n33244), .Z(c[1803]) );
  NANDN U34539 ( .A(n33212), .B(n33211), .Z(n33216) );
  NANDN U34540 ( .A(n33214), .B(n33213), .Z(n33215) );
  AND U34541 ( .A(n33216), .B(n33215), .Z(n33251) );
  NANDN U34542 ( .A(n33218), .B(n33217), .Z(n33222) );
  NANDN U34543 ( .A(n33220), .B(n33219), .Z(n33221) );
  AND U34544 ( .A(n33222), .B(n33221), .Z(n33249) );
  NAND U34545 ( .A(n42143), .B(n33223), .Z(n33225) );
  XNOR U34546 ( .A(a[782]), .B(n4183), .Z(n33260) );
  NAND U34547 ( .A(n42144), .B(n33260), .Z(n33224) );
  AND U34548 ( .A(n33225), .B(n33224), .Z(n33275) );
  XOR U34549 ( .A(a[786]), .B(n42012), .Z(n33263) );
  XNOR U34550 ( .A(n33275), .B(n33274), .Z(n33277) );
  XOR U34551 ( .A(a[784]), .B(n42085), .Z(n33267) );
  AND U34552 ( .A(a[780]), .B(b[7]), .Z(n33268) );
  XNOR U34553 ( .A(n33269), .B(n33268), .Z(n33270) );
  AND U34554 ( .A(a[788]), .B(b[0]), .Z(n33228) );
  XNOR U34555 ( .A(n33228), .B(n4071), .Z(n33230) );
  NANDN U34556 ( .A(b[0]), .B(a[787]), .Z(n33229) );
  NAND U34557 ( .A(n33230), .B(n33229), .Z(n33271) );
  XNOR U34558 ( .A(n33270), .B(n33271), .Z(n33276) );
  XOR U34559 ( .A(n33277), .B(n33276), .Z(n33255) );
  NANDN U34560 ( .A(n33232), .B(n33231), .Z(n33236) );
  NANDN U34561 ( .A(n33234), .B(n33233), .Z(n33235) );
  AND U34562 ( .A(n33236), .B(n33235), .Z(n33254) );
  XNOR U34563 ( .A(n33255), .B(n33254), .Z(n33256) );
  NANDN U34564 ( .A(n33238), .B(n33237), .Z(n33242) );
  NAND U34565 ( .A(n33240), .B(n33239), .Z(n33241) );
  NAND U34566 ( .A(n33242), .B(n33241), .Z(n33257) );
  XNOR U34567 ( .A(n33256), .B(n33257), .Z(n33248) );
  XNOR U34568 ( .A(n33249), .B(n33248), .Z(n33250) );
  XNOR U34569 ( .A(n33251), .B(n33250), .Z(n33280) );
  XNOR U34570 ( .A(sreg[1804]), .B(n33280), .Z(n33282) );
  NANDN U34571 ( .A(sreg[1803]), .B(n33243), .Z(n33247) );
  NAND U34572 ( .A(n33245), .B(n33244), .Z(n33246) );
  NAND U34573 ( .A(n33247), .B(n33246), .Z(n33281) );
  XNOR U34574 ( .A(n33282), .B(n33281), .Z(c[1804]) );
  NANDN U34575 ( .A(n33249), .B(n33248), .Z(n33253) );
  NANDN U34576 ( .A(n33251), .B(n33250), .Z(n33252) );
  AND U34577 ( .A(n33253), .B(n33252), .Z(n33288) );
  NANDN U34578 ( .A(n33255), .B(n33254), .Z(n33259) );
  NANDN U34579 ( .A(n33257), .B(n33256), .Z(n33258) );
  AND U34580 ( .A(n33259), .B(n33258), .Z(n33286) );
  NAND U34581 ( .A(n42143), .B(n33260), .Z(n33262) );
  XNOR U34582 ( .A(a[783]), .B(n4183), .Z(n33297) );
  NAND U34583 ( .A(n42144), .B(n33297), .Z(n33261) );
  AND U34584 ( .A(n33262), .B(n33261), .Z(n33312) );
  XOR U34585 ( .A(a[787]), .B(n42012), .Z(n33300) );
  XNOR U34586 ( .A(n33312), .B(n33311), .Z(n33314) );
  AND U34587 ( .A(a[789]), .B(b[0]), .Z(n33264) );
  XNOR U34588 ( .A(n33264), .B(n4071), .Z(n33266) );
  NANDN U34589 ( .A(b[0]), .B(a[788]), .Z(n33265) );
  NAND U34590 ( .A(n33266), .B(n33265), .Z(n33308) );
  XOR U34591 ( .A(a[785]), .B(n42085), .Z(n33301) );
  AND U34592 ( .A(a[781]), .B(b[7]), .Z(n33305) );
  XNOR U34593 ( .A(n33306), .B(n33305), .Z(n33307) );
  XNOR U34594 ( .A(n33308), .B(n33307), .Z(n33313) );
  XOR U34595 ( .A(n33314), .B(n33313), .Z(n33292) );
  NANDN U34596 ( .A(n33269), .B(n33268), .Z(n33273) );
  NANDN U34597 ( .A(n33271), .B(n33270), .Z(n33272) );
  AND U34598 ( .A(n33273), .B(n33272), .Z(n33291) );
  XNOR U34599 ( .A(n33292), .B(n33291), .Z(n33293) );
  NANDN U34600 ( .A(n33275), .B(n33274), .Z(n33279) );
  NAND U34601 ( .A(n33277), .B(n33276), .Z(n33278) );
  NAND U34602 ( .A(n33279), .B(n33278), .Z(n33294) );
  XNOR U34603 ( .A(n33293), .B(n33294), .Z(n33285) );
  XNOR U34604 ( .A(n33286), .B(n33285), .Z(n33287) );
  XNOR U34605 ( .A(n33288), .B(n33287), .Z(n33317) );
  XNOR U34606 ( .A(sreg[1805]), .B(n33317), .Z(n33319) );
  NANDN U34607 ( .A(sreg[1804]), .B(n33280), .Z(n33284) );
  NAND U34608 ( .A(n33282), .B(n33281), .Z(n33283) );
  NAND U34609 ( .A(n33284), .B(n33283), .Z(n33318) );
  XNOR U34610 ( .A(n33319), .B(n33318), .Z(c[1805]) );
  NANDN U34611 ( .A(n33286), .B(n33285), .Z(n33290) );
  NANDN U34612 ( .A(n33288), .B(n33287), .Z(n33289) );
  AND U34613 ( .A(n33290), .B(n33289), .Z(n33325) );
  NANDN U34614 ( .A(n33292), .B(n33291), .Z(n33296) );
  NANDN U34615 ( .A(n33294), .B(n33293), .Z(n33295) );
  AND U34616 ( .A(n33296), .B(n33295), .Z(n33323) );
  NAND U34617 ( .A(n42143), .B(n33297), .Z(n33299) );
  XNOR U34618 ( .A(a[784]), .B(n4183), .Z(n33334) );
  NAND U34619 ( .A(n42144), .B(n33334), .Z(n33298) );
  AND U34620 ( .A(n33299), .B(n33298), .Z(n33349) );
  XOR U34621 ( .A(a[788]), .B(n42012), .Z(n33337) );
  XNOR U34622 ( .A(n33349), .B(n33348), .Z(n33351) );
  XOR U34623 ( .A(a[786]), .B(n42085), .Z(n33341) );
  AND U34624 ( .A(a[782]), .B(b[7]), .Z(n33342) );
  XNOR U34625 ( .A(n33343), .B(n33342), .Z(n33344) );
  AND U34626 ( .A(a[790]), .B(b[0]), .Z(n33302) );
  XNOR U34627 ( .A(n33302), .B(n4071), .Z(n33304) );
  NANDN U34628 ( .A(b[0]), .B(a[789]), .Z(n33303) );
  NAND U34629 ( .A(n33304), .B(n33303), .Z(n33345) );
  XNOR U34630 ( .A(n33344), .B(n33345), .Z(n33350) );
  XOR U34631 ( .A(n33351), .B(n33350), .Z(n33329) );
  NANDN U34632 ( .A(n33306), .B(n33305), .Z(n33310) );
  NANDN U34633 ( .A(n33308), .B(n33307), .Z(n33309) );
  AND U34634 ( .A(n33310), .B(n33309), .Z(n33328) );
  XNOR U34635 ( .A(n33329), .B(n33328), .Z(n33330) );
  NANDN U34636 ( .A(n33312), .B(n33311), .Z(n33316) );
  NAND U34637 ( .A(n33314), .B(n33313), .Z(n33315) );
  NAND U34638 ( .A(n33316), .B(n33315), .Z(n33331) );
  XNOR U34639 ( .A(n33330), .B(n33331), .Z(n33322) );
  XNOR U34640 ( .A(n33323), .B(n33322), .Z(n33324) );
  XNOR U34641 ( .A(n33325), .B(n33324), .Z(n33354) );
  XNOR U34642 ( .A(sreg[1806]), .B(n33354), .Z(n33356) );
  NANDN U34643 ( .A(sreg[1805]), .B(n33317), .Z(n33321) );
  NAND U34644 ( .A(n33319), .B(n33318), .Z(n33320) );
  NAND U34645 ( .A(n33321), .B(n33320), .Z(n33355) );
  XNOR U34646 ( .A(n33356), .B(n33355), .Z(c[1806]) );
  NANDN U34647 ( .A(n33323), .B(n33322), .Z(n33327) );
  NANDN U34648 ( .A(n33325), .B(n33324), .Z(n33326) );
  AND U34649 ( .A(n33327), .B(n33326), .Z(n33362) );
  NANDN U34650 ( .A(n33329), .B(n33328), .Z(n33333) );
  NANDN U34651 ( .A(n33331), .B(n33330), .Z(n33332) );
  AND U34652 ( .A(n33333), .B(n33332), .Z(n33360) );
  NAND U34653 ( .A(n42143), .B(n33334), .Z(n33336) );
  XNOR U34654 ( .A(a[785]), .B(n4184), .Z(n33371) );
  NAND U34655 ( .A(n42144), .B(n33371), .Z(n33335) );
  AND U34656 ( .A(n33336), .B(n33335), .Z(n33386) );
  XOR U34657 ( .A(a[789]), .B(n42012), .Z(n33374) );
  XNOR U34658 ( .A(n33386), .B(n33385), .Z(n33388) );
  AND U34659 ( .A(a[791]), .B(b[0]), .Z(n33338) );
  XNOR U34660 ( .A(n33338), .B(n4071), .Z(n33340) );
  NANDN U34661 ( .A(b[0]), .B(a[790]), .Z(n33339) );
  NAND U34662 ( .A(n33340), .B(n33339), .Z(n33382) );
  XOR U34663 ( .A(a[787]), .B(n42085), .Z(n33378) );
  AND U34664 ( .A(a[783]), .B(b[7]), .Z(n33379) );
  XNOR U34665 ( .A(n33380), .B(n33379), .Z(n33381) );
  XNOR U34666 ( .A(n33382), .B(n33381), .Z(n33387) );
  XOR U34667 ( .A(n33388), .B(n33387), .Z(n33366) );
  NANDN U34668 ( .A(n33343), .B(n33342), .Z(n33347) );
  NANDN U34669 ( .A(n33345), .B(n33344), .Z(n33346) );
  AND U34670 ( .A(n33347), .B(n33346), .Z(n33365) );
  XNOR U34671 ( .A(n33366), .B(n33365), .Z(n33367) );
  NANDN U34672 ( .A(n33349), .B(n33348), .Z(n33353) );
  NAND U34673 ( .A(n33351), .B(n33350), .Z(n33352) );
  NAND U34674 ( .A(n33353), .B(n33352), .Z(n33368) );
  XNOR U34675 ( .A(n33367), .B(n33368), .Z(n33359) );
  XNOR U34676 ( .A(n33360), .B(n33359), .Z(n33361) );
  XNOR U34677 ( .A(n33362), .B(n33361), .Z(n33391) );
  XNOR U34678 ( .A(sreg[1807]), .B(n33391), .Z(n33393) );
  NANDN U34679 ( .A(sreg[1806]), .B(n33354), .Z(n33358) );
  NAND U34680 ( .A(n33356), .B(n33355), .Z(n33357) );
  NAND U34681 ( .A(n33358), .B(n33357), .Z(n33392) );
  XNOR U34682 ( .A(n33393), .B(n33392), .Z(c[1807]) );
  NANDN U34683 ( .A(n33360), .B(n33359), .Z(n33364) );
  NANDN U34684 ( .A(n33362), .B(n33361), .Z(n33363) );
  AND U34685 ( .A(n33364), .B(n33363), .Z(n33399) );
  NANDN U34686 ( .A(n33366), .B(n33365), .Z(n33370) );
  NANDN U34687 ( .A(n33368), .B(n33367), .Z(n33369) );
  AND U34688 ( .A(n33370), .B(n33369), .Z(n33397) );
  NAND U34689 ( .A(n42143), .B(n33371), .Z(n33373) );
  XNOR U34690 ( .A(a[786]), .B(n4184), .Z(n33408) );
  NAND U34691 ( .A(n42144), .B(n33408), .Z(n33372) );
  AND U34692 ( .A(n33373), .B(n33372), .Z(n33423) );
  XOR U34693 ( .A(a[790]), .B(n42012), .Z(n33411) );
  XNOR U34694 ( .A(n33423), .B(n33422), .Z(n33425) );
  AND U34695 ( .A(a[792]), .B(b[0]), .Z(n33375) );
  XNOR U34696 ( .A(n33375), .B(n4071), .Z(n33377) );
  NANDN U34697 ( .A(b[0]), .B(a[791]), .Z(n33376) );
  NAND U34698 ( .A(n33377), .B(n33376), .Z(n33419) );
  XOR U34699 ( .A(a[788]), .B(n42085), .Z(n33415) );
  AND U34700 ( .A(a[784]), .B(b[7]), .Z(n33416) );
  XNOR U34701 ( .A(n33417), .B(n33416), .Z(n33418) );
  XNOR U34702 ( .A(n33419), .B(n33418), .Z(n33424) );
  XOR U34703 ( .A(n33425), .B(n33424), .Z(n33403) );
  NANDN U34704 ( .A(n33380), .B(n33379), .Z(n33384) );
  NANDN U34705 ( .A(n33382), .B(n33381), .Z(n33383) );
  AND U34706 ( .A(n33384), .B(n33383), .Z(n33402) );
  XNOR U34707 ( .A(n33403), .B(n33402), .Z(n33404) );
  NANDN U34708 ( .A(n33386), .B(n33385), .Z(n33390) );
  NAND U34709 ( .A(n33388), .B(n33387), .Z(n33389) );
  NAND U34710 ( .A(n33390), .B(n33389), .Z(n33405) );
  XNOR U34711 ( .A(n33404), .B(n33405), .Z(n33396) );
  XNOR U34712 ( .A(n33397), .B(n33396), .Z(n33398) );
  XNOR U34713 ( .A(n33399), .B(n33398), .Z(n33428) );
  XNOR U34714 ( .A(sreg[1808]), .B(n33428), .Z(n33430) );
  NANDN U34715 ( .A(sreg[1807]), .B(n33391), .Z(n33395) );
  NAND U34716 ( .A(n33393), .B(n33392), .Z(n33394) );
  NAND U34717 ( .A(n33395), .B(n33394), .Z(n33429) );
  XNOR U34718 ( .A(n33430), .B(n33429), .Z(c[1808]) );
  NANDN U34719 ( .A(n33397), .B(n33396), .Z(n33401) );
  NANDN U34720 ( .A(n33399), .B(n33398), .Z(n33400) );
  AND U34721 ( .A(n33401), .B(n33400), .Z(n33436) );
  NANDN U34722 ( .A(n33403), .B(n33402), .Z(n33407) );
  NANDN U34723 ( .A(n33405), .B(n33404), .Z(n33406) );
  AND U34724 ( .A(n33407), .B(n33406), .Z(n33434) );
  NAND U34725 ( .A(n42143), .B(n33408), .Z(n33410) );
  XNOR U34726 ( .A(a[787]), .B(n4184), .Z(n33445) );
  NAND U34727 ( .A(n42144), .B(n33445), .Z(n33409) );
  AND U34728 ( .A(n33410), .B(n33409), .Z(n33460) );
  XOR U34729 ( .A(a[791]), .B(n42012), .Z(n33448) );
  XNOR U34730 ( .A(n33460), .B(n33459), .Z(n33462) );
  AND U34731 ( .A(a[793]), .B(b[0]), .Z(n33412) );
  XNOR U34732 ( .A(n33412), .B(n4071), .Z(n33414) );
  NANDN U34733 ( .A(b[0]), .B(a[792]), .Z(n33413) );
  NAND U34734 ( .A(n33414), .B(n33413), .Z(n33456) );
  XOR U34735 ( .A(a[789]), .B(n42085), .Z(n33449) );
  AND U34736 ( .A(a[785]), .B(b[7]), .Z(n33453) );
  XNOR U34737 ( .A(n33454), .B(n33453), .Z(n33455) );
  XNOR U34738 ( .A(n33456), .B(n33455), .Z(n33461) );
  XOR U34739 ( .A(n33462), .B(n33461), .Z(n33440) );
  NANDN U34740 ( .A(n33417), .B(n33416), .Z(n33421) );
  NANDN U34741 ( .A(n33419), .B(n33418), .Z(n33420) );
  AND U34742 ( .A(n33421), .B(n33420), .Z(n33439) );
  XNOR U34743 ( .A(n33440), .B(n33439), .Z(n33441) );
  NANDN U34744 ( .A(n33423), .B(n33422), .Z(n33427) );
  NAND U34745 ( .A(n33425), .B(n33424), .Z(n33426) );
  NAND U34746 ( .A(n33427), .B(n33426), .Z(n33442) );
  XNOR U34747 ( .A(n33441), .B(n33442), .Z(n33433) );
  XNOR U34748 ( .A(n33434), .B(n33433), .Z(n33435) );
  XNOR U34749 ( .A(n33436), .B(n33435), .Z(n33465) );
  XNOR U34750 ( .A(sreg[1809]), .B(n33465), .Z(n33467) );
  NANDN U34751 ( .A(sreg[1808]), .B(n33428), .Z(n33432) );
  NAND U34752 ( .A(n33430), .B(n33429), .Z(n33431) );
  NAND U34753 ( .A(n33432), .B(n33431), .Z(n33466) );
  XNOR U34754 ( .A(n33467), .B(n33466), .Z(c[1809]) );
  NANDN U34755 ( .A(n33434), .B(n33433), .Z(n33438) );
  NANDN U34756 ( .A(n33436), .B(n33435), .Z(n33437) );
  AND U34757 ( .A(n33438), .B(n33437), .Z(n33473) );
  NANDN U34758 ( .A(n33440), .B(n33439), .Z(n33444) );
  NANDN U34759 ( .A(n33442), .B(n33441), .Z(n33443) );
  AND U34760 ( .A(n33444), .B(n33443), .Z(n33471) );
  NAND U34761 ( .A(n42143), .B(n33445), .Z(n33447) );
  XNOR U34762 ( .A(a[788]), .B(n4184), .Z(n33482) );
  NAND U34763 ( .A(n42144), .B(n33482), .Z(n33446) );
  AND U34764 ( .A(n33447), .B(n33446), .Z(n33497) );
  XOR U34765 ( .A(a[792]), .B(n42012), .Z(n33485) );
  XNOR U34766 ( .A(n33497), .B(n33496), .Z(n33499) );
  XOR U34767 ( .A(a[790]), .B(n42085), .Z(n33489) );
  AND U34768 ( .A(a[786]), .B(b[7]), .Z(n33490) );
  XNOR U34769 ( .A(n33491), .B(n33490), .Z(n33492) );
  AND U34770 ( .A(a[794]), .B(b[0]), .Z(n33450) );
  XNOR U34771 ( .A(n33450), .B(n4071), .Z(n33452) );
  NANDN U34772 ( .A(b[0]), .B(a[793]), .Z(n33451) );
  NAND U34773 ( .A(n33452), .B(n33451), .Z(n33493) );
  XNOR U34774 ( .A(n33492), .B(n33493), .Z(n33498) );
  XOR U34775 ( .A(n33499), .B(n33498), .Z(n33477) );
  NANDN U34776 ( .A(n33454), .B(n33453), .Z(n33458) );
  NANDN U34777 ( .A(n33456), .B(n33455), .Z(n33457) );
  AND U34778 ( .A(n33458), .B(n33457), .Z(n33476) );
  XNOR U34779 ( .A(n33477), .B(n33476), .Z(n33478) );
  NANDN U34780 ( .A(n33460), .B(n33459), .Z(n33464) );
  NAND U34781 ( .A(n33462), .B(n33461), .Z(n33463) );
  NAND U34782 ( .A(n33464), .B(n33463), .Z(n33479) );
  XNOR U34783 ( .A(n33478), .B(n33479), .Z(n33470) );
  XNOR U34784 ( .A(n33471), .B(n33470), .Z(n33472) );
  XNOR U34785 ( .A(n33473), .B(n33472), .Z(n33502) );
  XNOR U34786 ( .A(sreg[1810]), .B(n33502), .Z(n33504) );
  NANDN U34787 ( .A(sreg[1809]), .B(n33465), .Z(n33469) );
  NAND U34788 ( .A(n33467), .B(n33466), .Z(n33468) );
  NAND U34789 ( .A(n33469), .B(n33468), .Z(n33503) );
  XNOR U34790 ( .A(n33504), .B(n33503), .Z(c[1810]) );
  NANDN U34791 ( .A(n33471), .B(n33470), .Z(n33475) );
  NANDN U34792 ( .A(n33473), .B(n33472), .Z(n33474) );
  AND U34793 ( .A(n33475), .B(n33474), .Z(n33510) );
  NANDN U34794 ( .A(n33477), .B(n33476), .Z(n33481) );
  NANDN U34795 ( .A(n33479), .B(n33478), .Z(n33480) );
  AND U34796 ( .A(n33481), .B(n33480), .Z(n33508) );
  NAND U34797 ( .A(n42143), .B(n33482), .Z(n33484) );
  XNOR U34798 ( .A(a[789]), .B(n4184), .Z(n33519) );
  NAND U34799 ( .A(n42144), .B(n33519), .Z(n33483) );
  AND U34800 ( .A(n33484), .B(n33483), .Z(n33534) );
  XOR U34801 ( .A(a[793]), .B(n42012), .Z(n33522) );
  XNOR U34802 ( .A(n33534), .B(n33533), .Z(n33536) );
  AND U34803 ( .A(a[795]), .B(b[0]), .Z(n33486) );
  XNOR U34804 ( .A(n33486), .B(n4071), .Z(n33488) );
  NANDN U34805 ( .A(b[0]), .B(a[794]), .Z(n33487) );
  NAND U34806 ( .A(n33488), .B(n33487), .Z(n33530) );
  XOR U34807 ( .A(a[791]), .B(n42085), .Z(n33523) );
  AND U34808 ( .A(a[787]), .B(b[7]), .Z(n33527) );
  XNOR U34809 ( .A(n33528), .B(n33527), .Z(n33529) );
  XNOR U34810 ( .A(n33530), .B(n33529), .Z(n33535) );
  XOR U34811 ( .A(n33536), .B(n33535), .Z(n33514) );
  NANDN U34812 ( .A(n33491), .B(n33490), .Z(n33495) );
  NANDN U34813 ( .A(n33493), .B(n33492), .Z(n33494) );
  AND U34814 ( .A(n33495), .B(n33494), .Z(n33513) );
  XNOR U34815 ( .A(n33514), .B(n33513), .Z(n33515) );
  NANDN U34816 ( .A(n33497), .B(n33496), .Z(n33501) );
  NAND U34817 ( .A(n33499), .B(n33498), .Z(n33500) );
  NAND U34818 ( .A(n33501), .B(n33500), .Z(n33516) );
  XNOR U34819 ( .A(n33515), .B(n33516), .Z(n33507) );
  XNOR U34820 ( .A(n33508), .B(n33507), .Z(n33509) );
  XNOR U34821 ( .A(n33510), .B(n33509), .Z(n33539) );
  XNOR U34822 ( .A(sreg[1811]), .B(n33539), .Z(n33541) );
  NANDN U34823 ( .A(sreg[1810]), .B(n33502), .Z(n33506) );
  NAND U34824 ( .A(n33504), .B(n33503), .Z(n33505) );
  NAND U34825 ( .A(n33506), .B(n33505), .Z(n33540) );
  XNOR U34826 ( .A(n33541), .B(n33540), .Z(c[1811]) );
  NANDN U34827 ( .A(n33508), .B(n33507), .Z(n33512) );
  NANDN U34828 ( .A(n33510), .B(n33509), .Z(n33511) );
  AND U34829 ( .A(n33512), .B(n33511), .Z(n33547) );
  NANDN U34830 ( .A(n33514), .B(n33513), .Z(n33518) );
  NANDN U34831 ( .A(n33516), .B(n33515), .Z(n33517) );
  AND U34832 ( .A(n33518), .B(n33517), .Z(n33545) );
  NAND U34833 ( .A(n42143), .B(n33519), .Z(n33521) );
  XNOR U34834 ( .A(a[790]), .B(n4184), .Z(n33556) );
  NAND U34835 ( .A(n42144), .B(n33556), .Z(n33520) );
  AND U34836 ( .A(n33521), .B(n33520), .Z(n33571) );
  XOR U34837 ( .A(a[794]), .B(n42012), .Z(n33559) );
  XNOR U34838 ( .A(n33571), .B(n33570), .Z(n33573) );
  XOR U34839 ( .A(a[792]), .B(n42085), .Z(n33563) );
  AND U34840 ( .A(a[788]), .B(b[7]), .Z(n33564) );
  XNOR U34841 ( .A(n33565), .B(n33564), .Z(n33566) );
  AND U34842 ( .A(a[796]), .B(b[0]), .Z(n33524) );
  XNOR U34843 ( .A(n33524), .B(n4071), .Z(n33526) );
  NANDN U34844 ( .A(b[0]), .B(a[795]), .Z(n33525) );
  NAND U34845 ( .A(n33526), .B(n33525), .Z(n33567) );
  XNOR U34846 ( .A(n33566), .B(n33567), .Z(n33572) );
  XOR U34847 ( .A(n33573), .B(n33572), .Z(n33551) );
  NANDN U34848 ( .A(n33528), .B(n33527), .Z(n33532) );
  NANDN U34849 ( .A(n33530), .B(n33529), .Z(n33531) );
  AND U34850 ( .A(n33532), .B(n33531), .Z(n33550) );
  XNOR U34851 ( .A(n33551), .B(n33550), .Z(n33552) );
  NANDN U34852 ( .A(n33534), .B(n33533), .Z(n33538) );
  NAND U34853 ( .A(n33536), .B(n33535), .Z(n33537) );
  NAND U34854 ( .A(n33538), .B(n33537), .Z(n33553) );
  XNOR U34855 ( .A(n33552), .B(n33553), .Z(n33544) );
  XNOR U34856 ( .A(n33545), .B(n33544), .Z(n33546) );
  XNOR U34857 ( .A(n33547), .B(n33546), .Z(n33576) );
  XNOR U34858 ( .A(sreg[1812]), .B(n33576), .Z(n33578) );
  NANDN U34859 ( .A(sreg[1811]), .B(n33539), .Z(n33543) );
  NAND U34860 ( .A(n33541), .B(n33540), .Z(n33542) );
  NAND U34861 ( .A(n33543), .B(n33542), .Z(n33577) );
  XNOR U34862 ( .A(n33578), .B(n33577), .Z(c[1812]) );
  NANDN U34863 ( .A(n33545), .B(n33544), .Z(n33549) );
  NANDN U34864 ( .A(n33547), .B(n33546), .Z(n33548) );
  AND U34865 ( .A(n33549), .B(n33548), .Z(n33584) );
  NANDN U34866 ( .A(n33551), .B(n33550), .Z(n33555) );
  NANDN U34867 ( .A(n33553), .B(n33552), .Z(n33554) );
  AND U34868 ( .A(n33555), .B(n33554), .Z(n33582) );
  NAND U34869 ( .A(n42143), .B(n33556), .Z(n33558) );
  XNOR U34870 ( .A(a[791]), .B(n4184), .Z(n33593) );
  NAND U34871 ( .A(n42144), .B(n33593), .Z(n33557) );
  AND U34872 ( .A(n33558), .B(n33557), .Z(n33608) );
  XOR U34873 ( .A(a[795]), .B(n42012), .Z(n33596) );
  XNOR U34874 ( .A(n33608), .B(n33607), .Z(n33610) );
  AND U34875 ( .A(a[797]), .B(b[0]), .Z(n33560) );
  XNOR U34876 ( .A(n33560), .B(n4071), .Z(n33562) );
  NANDN U34877 ( .A(b[0]), .B(a[796]), .Z(n33561) );
  NAND U34878 ( .A(n33562), .B(n33561), .Z(n33604) );
  XOR U34879 ( .A(a[793]), .B(n42085), .Z(n33600) );
  AND U34880 ( .A(a[789]), .B(b[7]), .Z(n33601) );
  XNOR U34881 ( .A(n33602), .B(n33601), .Z(n33603) );
  XNOR U34882 ( .A(n33604), .B(n33603), .Z(n33609) );
  XOR U34883 ( .A(n33610), .B(n33609), .Z(n33588) );
  NANDN U34884 ( .A(n33565), .B(n33564), .Z(n33569) );
  NANDN U34885 ( .A(n33567), .B(n33566), .Z(n33568) );
  AND U34886 ( .A(n33569), .B(n33568), .Z(n33587) );
  XNOR U34887 ( .A(n33588), .B(n33587), .Z(n33589) );
  NANDN U34888 ( .A(n33571), .B(n33570), .Z(n33575) );
  NAND U34889 ( .A(n33573), .B(n33572), .Z(n33574) );
  NAND U34890 ( .A(n33575), .B(n33574), .Z(n33590) );
  XNOR U34891 ( .A(n33589), .B(n33590), .Z(n33581) );
  XNOR U34892 ( .A(n33582), .B(n33581), .Z(n33583) );
  XNOR U34893 ( .A(n33584), .B(n33583), .Z(n33613) );
  XNOR U34894 ( .A(sreg[1813]), .B(n33613), .Z(n33615) );
  NANDN U34895 ( .A(sreg[1812]), .B(n33576), .Z(n33580) );
  NAND U34896 ( .A(n33578), .B(n33577), .Z(n33579) );
  NAND U34897 ( .A(n33580), .B(n33579), .Z(n33614) );
  XNOR U34898 ( .A(n33615), .B(n33614), .Z(c[1813]) );
  NANDN U34899 ( .A(n33582), .B(n33581), .Z(n33586) );
  NANDN U34900 ( .A(n33584), .B(n33583), .Z(n33585) );
  AND U34901 ( .A(n33586), .B(n33585), .Z(n33621) );
  NANDN U34902 ( .A(n33588), .B(n33587), .Z(n33592) );
  NANDN U34903 ( .A(n33590), .B(n33589), .Z(n33591) );
  AND U34904 ( .A(n33592), .B(n33591), .Z(n33619) );
  NAND U34905 ( .A(n42143), .B(n33593), .Z(n33595) );
  XNOR U34906 ( .A(a[792]), .B(n4185), .Z(n33630) );
  NAND U34907 ( .A(n42144), .B(n33630), .Z(n33594) );
  AND U34908 ( .A(n33595), .B(n33594), .Z(n33645) );
  XOR U34909 ( .A(a[796]), .B(n42012), .Z(n33633) );
  XNOR U34910 ( .A(n33645), .B(n33644), .Z(n33647) );
  AND U34911 ( .A(a[798]), .B(b[0]), .Z(n33597) );
  XNOR U34912 ( .A(n33597), .B(n4071), .Z(n33599) );
  NANDN U34913 ( .A(b[0]), .B(a[797]), .Z(n33598) );
  NAND U34914 ( .A(n33599), .B(n33598), .Z(n33641) );
  XOR U34915 ( .A(a[794]), .B(n42085), .Z(n33634) );
  AND U34916 ( .A(a[790]), .B(b[7]), .Z(n33638) );
  XNOR U34917 ( .A(n33639), .B(n33638), .Z(n33640) );
  XNOR U34918 ( .A(n33641), .B(n33640), .Z(n33646) );
  XOR U34919 ( .A(n33647), .B(n33646), .Z(n33625) );
  NANDN U34920 ( .A(n33602), .B(n33601), .Z(n33606) );
  NANDN U34921 ( .A(n33604), .B(n33603), .Z(n33605) );
  AND U34922 ( .A(n33606), .B(n33605), .Z(n33624) );
  XNOR U34923 ( .A(n33625), .B(n33624), .Z(n33626) );
  NANDN U34924 ( .A(n33608), .B(n33607), .Z(n33612) );
  NAND U34925 ( .A(n33610), .B(n33609), .Z(n33611) );
  NAND U34926 ( .A(n33612), .B(n33611), .Z(n33627) );
  XNOR U34927 ( .A(n33626), .B(n33627), .Z(n33618) );
  XNOR U34928 ( .A(n33619), .B(n33618), .Z(n33620) );
  XNOR U34929 ( .A(n33621), .B(n33620), .Z(n33650) );
  XNOR U34930 ( .A(sreg[1814]), .B(n33650), .Z(n33652) );
  NANDN U34931 ( .A(sreg[1813]), .B(n33613), .Z(n33617) );
  NAND U34932 ( .A(n33615), .B(n33614), .Z(n33616) );
  NAND U34933 ( .A(n33617), .B(n33616), .Z(n33651) );
  XNOR U34934 ( .A(n33652), .B(n33651), .Z(c[1814]) );
  NANDN U34935 ( .A(n33619), .B(n33618), .Z(n33623) );
  NANDN U34936 ( .A(n33621), .B(n33620), .Z(n33622) );
  AND U34937 ( .A(n33623), .B(n33622), .Z(n33658) );
  NANDN U34938 ( .A(n33625), .B(n33624), .Z(n33629) );
  NANDN U34939 ( .A(n33627), .B(n33626), .Z(n33628) );
  AND U34940 ( .A(n33629), .B(n33628), .Z(n33656) );
  NAND U34941 ( .A(n42143), .B(n33630), .Z(n33632) );
  XNOR U34942 ( .A(a[793]), .B(n4185), .Z(n33667) );
  NAND U34943 ( .A(n42144), .B(n33667), .Z(n33631) );
  AND U34944 ( .A(n33632), .B(n33631), .Z(n33682) );
  XOR U34945 ( .A(a[797]), .B(n42012), .Z(n33670) );
  XNOR U34946 ( .A(n33682), .B(n33681), .Z(n33684) );
  XOR U34947 ( .A(a[795]), .B(n42085), .Z(n33674) );
  AND U34948 ( .A(a[791]), .B(b[7]), .Z(n33675) );
  XNOR U34949 ( .A(n33676), .B(n33675), .Z(n33677) );
  AND U34950 ( .A(a[799]), .B(b[0]), .Z(n33635) );
  XNOR U34951 ( .A(n33635), .B(n4071), .Z(n33637) );
  NANDN U34952 ( .A(b[0]), .B(a[798]), .Z(n33636) );
  NAND U34953 ( .A(n33637), .B(n33636), .Z(n33678) );
  XNOR U34954 ( .A(n33677), .B(n33678), .Z(n33683) );
  XOR U34955 ( .A(n33684), .B(n33683), .Z(n33662) );
  NANDN U34956 ( .A(n33639), .B(n33638), .Z(n33643) );
  NANDN U34957 ( .A(n33641), .B(n33640), .Z(n33642) );
  AND U34958 ( .A(n33643), .B(n33642), .Z(n33661) );
  XNOR U34959 ( .A(n33662), .B(n33661), .Z(n33663) );
  NANDN U34960 ( .A(n33645), .B(n33644), .Z(n33649) );
  NAND U34961 ( .A(n33647), .B(n33646), .Z(n33648) );
  NAND U34962 ( .A(n33649), .B(n33648), .Z(n33664) );
  XNOR U34963 ( .A(n33663), .B(n33664), .Z(n33655) );
  XNOR U34964 ( .A(n33656), .B(n33655), .Z(n33657) );
  XNOR U34965 ( .A(n33658), .B(n33657), .Z(n33687) );
  XNOR U34966 ( .A(sreg[1815]), .B(n33687), .Z(n33689) );
  NANDN U34967 ( .A(sreg[1814]), .B(n33650), .Z(n33654) );
  NAND U34968 ( .A(n33652), .B(n33651), .Z(n33653) );
  NAND U34969 ( .A(n33654), .B(n33653), .Z(n33688) );
  XNOR U34970 ( .A(n33689), .B(n33688), .Z(c[1815]) );
  NANDN U34971 ( .A(n33656), .B(n33655), .Z(n33660) );
  NANDN U34972 ( .A(n33658), .B(n33657), .Z(n33659) );
  AND U34973 ( .A(n33660), .B(n33659), .Z(n33695) );
  NANDN U34974 ( .A(n33662), .B(n33661), .Z(n33666) );
  NANDN U34975 ( .A(n33664), .B(n33663), .Z(n33665) );
  AND U34976 ( .A(n33666), .B(n33665), .Z(n33693) );
  NAND U34977 ( .A(n42143), .B(n33667), .Z(n33669) );
  XNOR U34978 ( .A(a[794]), .B(n4185), .Z(n33704) );
  NAND U34979 ( .A(n42144), .B(n33704), .Z(n33668) );
  AND U34980 ( .A(n33669), .B(n33668), .Z(n33719) );
  XOR U34981 ( .A(a[798]), .B(n42012), .Z(n33707) );
  XNOR U34982 ( .A(n33719), .B(n33718), .Z(n33721) );
  AND U34983 ( .A(a[800]), .B(b[0]), .Z(n33671) );
  XNOR U34984 ( .A(n33671), .B(n4071), .Z(n33673) );
  NANDN U34985 ( .A(b[0]), .B(a[799]), .Z(n33672) );
  NAND U34986 ( .A(n33673), .B(n33672), .Z(n33715) );
  XOR U34987 ( .A(a[796]), .B(n42085), .Z(n33711) );
  AND U34988 ( .A(a[792]), .B(b[7]), .Z(n33712) );
  XNOR U34989 ( .A(n33713), .B(n33712), .Z(n33714) );
  XNOR U34990 ( .A(n33715), .B(n33714), .Z(n33720) );
  XOR U34991 ( .A(n33721), .B(n33720), .Z(n33699) );
  NANDN U34992 ( .A(n33676), .B(n33675), .Z(n33680) );
  NANDN U34993 ( .A(n33678), .B(n33677), .Z(n33679) );
  AND U34994 ( .A(n33680), .B(n33679), .Z(n33698) );
  XNOR U34995 ( .A(n33699), .B(n33698), .Z(n33700) );
  NANDN U34996 ( .A(n33682), .B(n33681), .Z(n33686) );
  NAND U34997 ( .A(n33684), .B(n33683), .Z(n33685) );
  NAND U34998 ( .A(n33686), .B(n33685), .Z(n33701) );
  XNOR U34999 ( .A(n33700), .B(n33701), .Z(n33692) );
  XNOR U35000 ( .A(n33693), .B(n33692), .Z(n33694) );
  XNOR U35001 ( .A(n33695), .B(n33694), .Z(n33724) );
  XNOR U35002 ( .A(sreg[1816]), .B(n33724), .Z(n33726) );
  NANDN U35003 ( .A(sreg[1815]), .B(n33687), .Z(n33691) );
  NAND U35004 ( .A(n33689), .B(n33688), .Z(n33690) );
  NAND U35005 ( .A(n33691), .B(n33690), .Z(n33725) );
  XNOR U35006 ( .A(n33726), .B(n33725), .Z(c[1816]) );
  NANDN U35007 ( .A(n33693), .B(n33692), .Z(n33697) );
  NANDN U35008 ( .A(n33695), .B(n33694), .Z(n33696) );
  AND U35009 ( .A(n33697), .B(n33696), .Z(n33732) );
  NANDN U35010 ( .A(n33699), .B(n33698), .Z(n33703) );
  NANDN U35011 ( .A(n33701), .B(n33700), .Z(n33702) );
  AND U35012 ( .A(n33703), .B(n33702), .Z(n33730) );
  NAND U35013 ( .A(n42143), .B(n33704), .Z(n33706) );
  XNOR U35014 ( .A(a[795]), .B(n4185), .Z(n33741) );
  NAND U35015 ( .A(n42144), .B(n33741), .Z(n33705) );
  AND U35016 ( .A(n33706), .B(n33705), .Z(n33756) );
  XOR U35017 ( .A(a[799]), .B(n42012), .Z(n33744) );
  XNOR U35018 ( .A(n33756), .B(n33755), .Z(n33758) );
  AND U35019 ( .A(a[801]), .B(b[0]), .Z(n33708) );
  XNOR U35020 ( .A(n33708), .B(n4071), .Z(n33710) );
  NANDN U35021 ( .A(b[0]), .B(a[800]), .Z(n33709) );
  NAND U35022 ( .A(n33710), .B(n33709), .Z(n33752) );
  XOR U35023 ( .A(a[797]), .B(n42085), .Z(n33748) );
  AND U35024 ( .A(a[793]), .B(b[7]), .Z(n33749) );
  XNOR U35025 ( .A(n33750), .B(n33749), .Z(n33751) );
  XNOR U35026 ( .A(n33752), .B(n33751), .Z(n33757) );
  XOR U35027 ( .A(n33758), .B(n33757), .Z(n33736) );
  NANDN U35028 ( .A(n33713), .B(n33712), .Z(n33717) );
  NANDN U35029 ( .A(n33715), .B(n33714), .Z(n33716) );
  AND U35030 ( .A(n33717), .B(n33716), .Z(n33735) );
  XNOR U35031 ( .A(n33736), .B(n33735), .Z(n33737) );
  NANDN U35032 ( .A(n33719), .B(n33718), .Z(n33723) );
  NAND U35033 ( .A(n33721), .B(n33720), .Z(n33722) );
  NAND U35034 ( .A(n33723), .B(n33722), .Z(n33738) );
  XNOR U35035 ( .A(n33737), .B(n33738), .Z(n33729) );
  XNOR U35036 ( .A(n33730), .B(n33729), .Z(n33731) );
  XNOR U35037 ( .A(n33732), .B(n33731), .Z(n33761) );
  XNOR U35038 ( .A(sreg[1817]), .B(n33761), .Z(n33763) );
  NANDN U35039 ( .A(sreg[1816]), .B(n33724), .Z(n33728) );
  NAND U35040 ( .A(n33726), .B(n33725), .Z(n33727) );
  NAND U35041 ( .A(n33728), .B(n33727), .Z(n33762) );
  XNOR U35042 ( .A(n33763), .B(n33762), .Z(c[1817]) );
  NANDN U35043 ( .A(n33730), .B(n33729), .Z(n33734) );
  NANDN U35044 ( .A(n33732), .B(n33731), .Z(n33733) );
  AND U35045 ( .A(n33734), .B(n33733), .Z(n33769) );
  NANDN U35046 ( .A(n33736), .B(n33735), .Z(n33740) );
  NANDN U35047 ( .A(n33738), .B(n33737), .Z(n33739) );
  AND U35048 ( .A(n33740), .B(n33739), .Z(n33767) );
  NAND U35049 ( .A(n42143), .B(n33741), .Z(n33743) );
  XNOR U35050 ( .A(a[796]), .B(n4185), .Z(n33778) );
  NAND U35051 ( .A(n42144), .B(n33778), .Z(n33742) );
  AND U35052 ( .A(n33743), .B(n33742), .Z(n33793) );
  XOR U35053 ( .A(a[800]), .B(n42012), .Z(n33781) );
  XNOR U35054 ( .A(n33793), .B(n33792), .Z(n33795) );
  AND U35055 ( .A(a[802]), .B(b[0]), .Z(n33745) );
  XNOR U35056 ( .A(n33745), .B(n4071), .Z(n33747) );
  NANDN U35057 ( .A(b[0]), .B(a[801]), .Z(n33746) );
  NAND U35058 ( .A(n33747), .B(n33746), .Z(n33789) );
  XOR U35059 ( .A(a[798]), .B(n42085), .Z(n33782) );
  AND U35060 ( .A(a[794]), .B(b[7]), .Z(n33786) );
  XNOR U35061 ( .A(n33787), .B(n33786), .Z(n33788) );
  XNOR U35062 ( .A(n33789), .B(n33788), .Z(n33794) );
  XOR U35063 ( .A(n33795), .B(n33794), .Z(n33773) );
  NANDN U35064 ( .A(n33750), .B(n33749), .Z(n33754) );
  NANDN U35065 ( .A(n33752), .B(n33751), .Z(n33753) );
  AND U35066 ( .A(n33754), .B(n33753), .Z(n33772) );
  XNOR U35067 ( .A(n33773), .B(n33772), .Z(n33774) );
  NANDN U35068 ( .A(n33756), .B(n33755), .Z(n33760) );
  NAND U35069 ( .A(n33758), .B(n33757), .Z(n33759) );
  NAND U35070 ( .A(n33760), .B(n33759), .Z(n33775) );
  XNOR U35071 ( .A(n33774), .B(n33775), .Z(n33766) );
  XNOR U35072 ( .A(n33767), .B(n33766), .Z(n33768) );
  XNOR U35073 ( .A(n33769), .B(n33768), .Z(n33798) );
  XNOR U35074 ( .A(sreg[1818]), .B(n33798), .Z(n33800) );
  NANDN U35075 ( .A(sreg[1817]), .B(n33761), .Z(n33765) );
  NAND U35076 ( .A(n33763), .B(n33762), .Z(n33764) );
  NAND U35077 ( .A(n33765), .B(n33764), .Z(n33799) );
  XNOR U35078 ( .A(n33800), .B(n33799), .Z(c[1818]) );
  NANDN U35079 ( .A(n33767), .B(n33766), .Z(n33771) );
  NANDN U35080 ( .A(n33769), .B(n33768), .Z(n33770) );
  AND U35081 ( .A(n33771), .B(n33770), .Z(n33806) );
  NANDN U35082 ( .A(n33773), .B(n33772), .Z(n33777) );
  NANDN U35083 ( .A(n33775), .B(n33774), .Z(n33776) );
  AND U35084 ( .A(n33777), .B(n33776), .Z(n33804) );
  NAND U35085 ( .A(n42143), .B(n33778), .Z(n33780) );
  XNOR U35086 ( .A(a[797]), .B(n4185), .Z(n33815) );
  NAND U35087 ( .A(n42144), .B(n33815), .Z(n33779) );
  AND U35088 ( .A(n33780), .B(n33779), .Z(n33830) );
  XOR U35089 ( .A(a[801]), .B(n42012), .Z(n33818) );
  XNOR U35090 ( .A(n33830), .B(n33829), .Z(n33832) );
  XOR U35091 ( .A(a[799]), .B(n42085), .Z(n33822) );
  AND U35092 ( .A(a[795]), .B(b[7]), .Z(n33823) );
  XNOR U35093 ( .A(n33824), .B(n33823), .Z(n33825) );
  AND U35094 ( .A(a[803]), .B(b[0]), .Z(n33783) );
  XNOR U35095 ( .A(n33783), .B(n4071), .Z(n33785) );
  NANDN U35096 ( .A(b[0]), .B(a[802]), .Z(n33784) );
  NAND U35097 ( .A(n33785), .B(n33784), .Z(n33826) );
  XNOR U35098 ( .A(n33825), .B(n33826), .Z(n33831) );
  XOR U35099 ( .A(n33832), .B(n33831), .Z(n33810) );
  NANDN U35100 ( .A(n33787), .B(n33786), .Z(n33791) );
  NANDN U35101 ( .A(n33789), .B(n33788), .Z(n33790) );
  AND U35102 ( .A(n33791), .B(n33790), .Z(n33809) );
  XNOR U35103 ( .A(n33810), .B(n33809), .Z(n33811) );
  NANDN U35104 ( .A(n33793), .B(n33792), .Z(n33797) );
  NAND U35105 ( .A(n33795), .B(n33794), .Z(n33796) );
  NAND U35106 ( .A(n33797), .B(n33796), .Z(n33812) );
  XNOR U35107 ( .A(n33811), .B(n33812), .Z(n33803) );
  XNOR U35108 ( .A(n33804), .B(n33803), .Z(n33805) );
  XNOR U35109 ( .A(n33806), .B(n33805), .Z(n33835) );
  XNOR U35110 ( .A(sreg[1819]), .B(n33835), .Z(n33837) );
  NANDN U35111 ( .A(sreg[1818]), .B(n33798), .Z(n33802) );
  NAND U35112 ( .A(n33800), .B(n33799), .Z(n33801) );
  NAND U35113 ( .A(n33802), .B(n33801), .Z(n33836) );
  XNOR U35114 ( .A(n33837), .B(n33836), .Z(c[1819]) );
  NANDN U35115 ( .A(n33804), .B(n33803), .Z(n33808) );
  NANDN U35116 ( .A(n33806), .B(n33805), .Z(n33807) );
  AND U35117 ( .A(n33808), .B(n33807), .Z(n33843) );
  NANDN U35118 ( .A(n33810), .B(n33809), .Z(n33814) );
  NANDN U35119 ( .A(n33812), .B(n33811), .Z(n33813) );
  AND U35120 ( .A(n33814), .B(n33813), .Z(n33841) );
  NAND U35121 ( .A(n42143), .B(n33815), .Z(n33817) );
  XNOR U35122 ( .A(a[798]), .B(n4185), .Z(n33852) );
  NAND U35123 ( .A(n42144), .B(n33852), .Z(n33816) );
  AND U35124 ( .A(n33817), .B(n33816), .Z(n33867) );
  XOR U35125 ( .A(a[802]), .B(n42012), .Z(n33855) );
  XNOR U35126 ( .A(n33867), .B(n33866), .Z(n33869) );
  AND U35127 ( .A(a[804]), .B(b[0]), .Z(n33819) );
  XNOR U35128 ( .A(n33819), .B(n4071), .Z(n33821) );
  NANDN U35129 ( .A(b[0]), .B(a[803]), .Z(n33820) );
  NAND U35130 ( .A(n33821), .B(n33820), .Z(n33863) );
  XOR U35131 ( .A(a[800]), .B(n42085), .Z(n33859) );
  AND U35132 ( .A(a[796]), .B(b[7]), .Z(n33860) );
  XNOR U35133 ( .A(n33861), .B(n33860), .Z(n33862) );
  XNOR U35134 ( .A(n33863), .B(n33862), .Z(n33868) );
  XOR U35135 ( .A(n33869), .B(n33868), .Z(n33847) );
  NANDN U35136 ( .A(n33824), .B(n33823), .Z(n33828) );
  NANDN U35137 ( .A(n33826), .B(n33825), .Z(n33827) );
  AND U35138 ( .A(n33828), .B(n33827), .Z(n33846) );
  XNOR U35139 ( .A(n33847), .B(n33846), .Z(n33848) );
  NANDN U35140 ( .A(n33830), .B(n33829), .Z(n33834) );
  NAND U35141 ( .A(n33832), .B(n33831), .Z(n33833) );
  NAND U35142 ( .A(n33834), .B(n33833), .Z(n33849) );
  XNOR U35143 ( .A(n33848), .B(n33849), .Z(n33840) );
  XNOR U35144 ( .A(n33841), .B(n33840), .Z(n33842) );
  XNOR U35145 ( .A(n33843), .B(n33842), .Z(n33872) );
  XNOR U35146 ( .A(sreg[1820]), .B(n33872), .Z(n33874) );
  NANDN U35147 ( .A(sreg[1819]), .B(n33835), .Z(n33839) );
  NAND U35148 ( .A(n33837), .B(n33836), .Z(n33838) );
  NAND U35149 ( .A(n33839), .B(n33838), .Z(n33873) );
  XNOR U35150 ( .A(n33874), .B(n33873), .Z(c[1820]) );
  NANDN U35151 ( .A(n33841), .B(n33840), .Z(n33845) );
  NANDN U35152 ( .A(n33843), .B(n33842), .Z(n33844) );
  AND U35153 ( .A(n33845), .B(n33844), .Z(n33880) );
  NANDN U35154 ( .A(n33847), .B(n33846), .Z(n33851) );
  NANDN U35155 ( .A(n33849), .B(n33848), .Z(n33850) );
  AND U35156 ( .A(n33851), .B(n33850), .Z(n33878) );
  NAND U35157 ( .A(n42143), .B(n33852), .Z(n33854) );
  XNOR U35158 ( .A(a[799]), .B(n4186), .Z(n33889) );
  NAND U35159 ( .A(n42144), .B(n33889), .Z(n33853) );
  AND U35160 ( .A(n33854), .B(n33853), .Z(n33904) );
  XOR U35161 ( .A(a[803]), .B(n42012), .Z(n33892) );
  XNOR U35162 ( .A(n33904), .B(n33903), .Z(n33906) );
  AND U35163 ( .A(a[805]), .B(b[0]), .Z(n33856) );
  XNOR U35164 ( .A(n33856), .B(n4071), .Z(n33858) );
  NANDN U35165 ( .A(b[0]), .B(a[804]), .Z(n33857) );
  NAND U35166 ( .A(n33858), .B(n33857), .Z(n33900) );
  XOR U35167 ( .A(a[801]), .B(n42085), .Z(n33893) );
  AND U35168 ( .A(a[797]), .B(b[7]), .Z(n33897) );
  XNOR U35169 ( .A(n33898), .B(n33897), .Z(n33899) );
  XNOR U35170 ( .A(n33900), .B(n33899), .Z(n33905) );
  XOR U35171 ( .A(n33906), .B(n33905), .Z(n33884) );
  NANDN U35172 ( .A(n33861), .B(n33860), .Z(n33865) );
  NANDN U35173 ( .A(n33863), .B(n33862), .Z(n33864) );
  AND U35174 ( .A(n33865), .B(n33864), .Z(n33883) );
  XNOR U35175 ( .A(n33884), .B(n33883), .Z(n33885) );
  NANDN U35176 ( .A(n33867), .B(n33866), .Z(n33871) );
  NAND U35177 ( .A(n33869), .B(n33868), .Z(n33870) );
  NAND U35178 ( .A(n33871), .B(n33870), .Z(n33886) );
  XNOR U35179 ( .A(n33885), .B(n33886), .Z(n33877) );
  XNOR U35180 ( .A(n33878), .B(n33877), .Z(n33879) );
  XNOR U35181 ( .A(n33880), .B(n33879), .Z(n33909) );
  XNOR U35182 ( .A(sreg[1821]), .B(n33909), .Z(n33911) );
  NANDN U35183 ( .A(sreg[1820]), .B(n33872), .Z(n33876) );
  NAND U35184 ( .A(n33874), .B(n33873), .Z(n33875) );
  NAND U35185 ( .A(n33876), .B(n33875), .Z(n33910) );
  XNOR U35186 ( .A(n33911), .B(n33910), .Z(c[1821]) );
  NANDN U35187 ( .A(n33878), .B(n33877), .Z(n33882) );
  NANDN U35188 ( .A(n33880), .B(n33879), .Z(n33881) );
  AND U35189 ( .A(n33882), .B(n33881), .Z(n33917) );
  NANDN U35190 ( .A(n33884), .B(n33883), .Z(n33888) );
  NANDN U35191 ( .A(n33886), .B(n33885), .Z(n33887) );
  AND U35192 ( .A(n33888), .B(n33887), .Z(n33915) );
  NAND U35193 ( .A(n42143), .B(n33889), .Z(n33891) );
  XNOR U35194 ( .A(a[800]), .B(n4186), .Z(n33926) );
  NAND U35195 ( .A(n42144), .B(n33926), .Z(n33890) );
  AND U35196 ( .A(n33891), .B(n33890), .Z(n33941) );
  XOR U35197 ( .A(a[804]), .B(n42012), .Z(n33929) );
  XNOR U35198 ( .A(n33941), .B(n33940), .Z(n33943) );
  XOR U35199 ( .A(a[802]), .B(n42085), .Z(n33933) );
  AND U35200 ( .A(a[798]), .B(b[7]), .Z(n33934) );
  XNOR U35201 ( .A(n33935), .B(n33934), .Z(n33936) );
  AND U35202 ( .A(a[806]), .B(b[0]), .Z(n33894) );
  XNOR U35203 ( .A(n33894), .B(n4071), .Z(n33896) );
  NANDN U35204 ( .A(b[0]), .B(a[805]), .Z(n33895) );
  NAND U35205 ( .A(n33896), .B(n33895), .Z(n33937) );
  XNOR U35206 ( .A(n33936), .B(n33937), .Z(n33942) );
  XOR U35207 ( .A(n33943), .B(n33942), .Z(n33921) );
  NANDN U35208 ( .A(n33898), .B(n33897), .Z(n33902) );
  NANDN U35209 ( .A(n33900), .B(n33899), .Z(n33901) );
  AND U35210 ( .A(n33902), .B(n33901), .Z(n33920) );
  XNOR U35211 ( .A(n33921), .B(n33920), .Z(n33922) );
  NANDN U35212 ( .A(n33904), .B(n33903), .Z(n33908) );
  NAND U35213 ( .A(n33906), .B(n33905), .Z(n33907) );
  NAND U35214 ( .A(n33908), .B(n33907), .Z(n33923) );
  XNOR U35215 ( .A(n33922), .B(n33923), .Z(n33914) );
  XNOR U35216 ( .A(n33915), .B(n33914), .Z(n33916) );
  XNOR U35217 ( .A(n33917), .B(n33916), .Z(n33946) );
  XNOR U35218 ( .A(sreg[1822]), .B(n33946), .Z(n33948) );
  NANDN U35219 ( .A(sreg[1821]), .B(n33909), .Z(n33913) );
  NAND U35220 ( .A(n33911), .B(n33910), .Z(n33912) );
  NAND U35221 ( .A(n33913), .B(n33912), .Z(n33947) );
  XNOR U35222 ( .A(n33948), .B(n33947), .Z(c[1822]) );
  NANDN U35223 ( .A(n33915), .B(n33914), .Z(n33919) );
  NANDN U35224 ( .A(n33917), .B(n33916), .Z(n33918) );
  AND U35225 ( .A(n33919), .B(n33918), .Z(n33954) );
  NANDN U35226 ( .A(n33921), .B(n33920), .Z(n33925) );
  NANDN U35227 ( .A(n33923), .B(n33922), .Z(n33924) );
  AND U35228 ( .A(n33925), .B(n33924), .Z(n33952) );
  NAND U35229 ( .A(n42143), .B(n33926), .Z(n33928) );
  XNOR U35230 ( .A(a[801]), .B(n4186), .Z(n33963) );
  NAND U35231 ( .A(n42144), .B(n33963), .Z(n33927) );
  AND U35232 ( .A(n33928), .B(n33927), .Z(n33978) );
  XOR U35233 ( .A(a[805]), .B(n42012), .Z(n33966) );
  XNOR U35234 ( .A(n33978), .B(n33977), .Z(n33980) );
  AND U35235 ( .A(a[807]), .B(b[0]), .Z(n33930) );
  XNOR U35236 ( .A(n33930), .B(n4071), .Z(n33932) );
  NANDN U35237 ( .A(b[0]), .B(a[806]), .Z(n33931) );
  NAND U35238 ( .A(n33932), .B(n33931), .Z(n33974) );
  XOR U35239 ( .A(a[803]), .B(n42085), .Z(n33967) );
  AND U35240 ( .A(a[799]), .B(b[7]), .Z(n33971) );
  XNOR U35241 ( .A(n33972), .B(n33971), .Z(n33973) );
  XNOR U35242 ( .A(n33974), .B(n33973), .Z(n33979) );
  XOR U35243 ( .A(n33980), .B(n33979), .Z(n33958) );
  NANDN U35244 ( .A(n33935), .B(n33934), .Z(n33939) );
  NANDN U35245 ( .A(n33937), .B(n33936), .Z(n33938) );
  AND U35246 ( .A(n33939), .B(n33938), .Z(n33957) );
  XNOR U35247 ( .A(n33958), .B(n33957), .Z(n33959) );
  NANDN U35248 ( .A(n33941), .B(n33940), .Z(n33945) );
  NAND U35249 ( .A(n33943), .B(n33942), .Z(n33944) );
  NAND U35250 ( .A(n33945), .B(n33944), .Z(n33960) );
  XNOR U35251 ( .A(n33959), .B(n33960), .Z(n33951) );
  XNOR U35252 ( .A(n33952), .B(n33951), .Z(n33953) );
  XNOR U35253 ( .A(n33954), .B(n33953), .Z(n33983) );
  XNOR U35254 ( .A(sreg[1823]), .B(n33983), .Z(n33985) );
  NANDN U35255 ( .A(sreg[1822]), .B(n33946), .Z(n33950) );
  NAND U35256 ( .A(n33948), .B(n33947), .Z(n33949) );
  NAND U35257 ( .A(n33950), .B(n33949), .Z(n33984) );
  XNOR U35258 ( .A(n33985), .B(n33984), .Z(c[1823]) );
  NANDN U35259 ( .A(n33952), .B(n33951), .Z(n33956) );
  NANDN U35260 ( .A(n33954), .B(n33953), .Z(n33955) );
  AND U35261 ( .A(n33956), .B(n33955), .Z(n33991) );
  NANDN U35262 ( .A(n33958), .B(n33957), .Z(n33962) );
  NANDN U35263 ( .A(n33960), .B(n33959), .Z(n33961) );
  AND U35264 ( .A(n33962), .B(n33961), .Z(n33989) );
  NAND U35265 ( .A(n42143), .B(n33963), .Z(n33965) );
  XNOR U35266 ( .A(a[802]), .B(n4186), .Z(n34000) );
  NAND U35267 ( .A(n42144), .B(n34000), .Z(n33964) );
  AND U35268 ( .A(n33965), .B(n33964), .Z(n34015) );
  XOR U35269 ( .A(a[806]), .B(n42012), .Z(n34003) );
  XNOR U35270 ( .A(n34015), .B(n34014), .Z(n34017) );
  XOR U35271 ( .A(a[804]), .B(n42085), .Z(n34007) );
  AND U35272 ( .A(a[800]), .B(b[7]), .Z(n34008) );
  XNOR U35273 ( .A(n34009), .B(n34008), .Z(n34010) );
  AND U35274 ( .A(a[808]), .B(b[0]), .Z(n33968) );
  XNOR U35275 ( .A(n33968), .B(n4071), .Z(n33970) );
  NANDN U35276 ( .A(b[0]), .B(a[807]), .Z(n33969) );
  NAND U35277 ( .A(n33970), .B(n33969), .Z(n34011) );
  XNOR U35278 ( .A(n34010), .B(n34011), .Z(n34016) );
  XOR U35279 ( .A(n34017), .B(n34016), .Z(n33995) );
  NANDN U35280 ( .A(n33972), .B(n33971), .Z(n33976) );
  NANDN U35281 ( .A(n33974), .B(n33973), .Z(n33975) );
  AND U35282 ( .A(n33976), .B(n33975), .Z(n33994) );
  XNOR U35283 ( .A(n33995), .B(n33994), .Z(n33996) );
  NANDN U35284 ( .A(n33978), .B(n33977), .Z(n33982) );
  NAND U35285 ( .A(n33980), .B(n33979), .Z(n33981) );
  NAND U35286 ( .A(n33982), .B(n33981), .Z(n33997) );
  XNOR U35287 ( .A(n33996), .B(n33997), .Z(n33988) );
  XNOR U35288 ( .A(n33989), .B(n33988), .Z(n33990) );
  XNOR U35289 ( .A(n33991), .B(n33990), .Z(n34020) );
  XNOR U35290 ( .A(sreg[1824]), .B(n34020), .Z(n34022) );
  NANDN U35291 ( .A(sreg[1823]), .B(n33983), .Z(n33987) );
  NAND U35292 ( .A(n33985), .B(n33984), .Z(n33986) );
  NAND U35293 ( .A(n33987), .B(n33986), .Z(n34021) );
  XNOR U35294 ( .A(n34022), .B(n34021), .Z(c[1824]) );
  NANDN U35295 ( .A(n33989), .B(n33988), .Z(n33993) );
  NANDN U35296 ( .A(n33991), .B(n33990), .Z(n33992) );
  AND U35297 ( .A(n33993), .B(n33992), .Z(n34028) );
  NANDN U35298 ( .A(n33995), .B(n33994), .Z(n33999) );
  NANDN U35299 ( .A(n33997), .B(n33996), .Z(n33998) );
  AND U35300 ( .A(n33999), .B(n33998), .Z(n34026) );
  NAND U35301 ( .A(n42143), .B(n34000), .Z(n34002) );
  XNOR U35302 ( .A(a[803]), .B(n4186), .Z(n34037) );
  NAND U35303 ( .A(n42144), .B(n34037), .Z(n34001) );
  AND U35304 ( .A(n34002), .B(n34001), .Z(n34052) );
  XOR U35305 ( .A(a[807]), .B(n42012), .Z(n34040) );
  XNOR U35306 ( .A(n34052), .B(n34051), .Z(n34054) );
  AND U35307 ( .A(a[809]), .B(b[0]), .Z(n34004) );
  XNOR U35308 ( .A(n34004), .B(n4071), .Z(n34006) );
  NANDN U35309 ( .A(b[0]), .B(a[808]), .Z(n34005) );
  NAND U35310 ( .A(n34006), .B(n34005), .Z(n34048) );
  XOR U35311 ( .A(a[805]), .B(n42085), .Z(n34044) );
  AND U35312 ( .A(a[801]), .B(b[7]), .Z(n34045) );
  XNOR U35313 ( .A(n34046), .B(n34045), .Z(n34047) );
  XNOR U35314 ( .A(n34048), .B(n34047), .Z(n34053) );
  XOR U35315 ( .A(n34054), .B(n34053), .Z(n34032) );
  NANDN U35316 ( .A(n34009), .B(n34008), .Z(n34013) );
  NANDN U35317 ( .A(n34011), .B(n34010), .Z(n34012) );
  AND U35318 ( .A(n34013), .B(n34012), .Z(n34031) );
  XNOR U35319 ( .A(n34032), .B(n34031), .Z(n34033) );
  NANDN U35320 ( .A(n34015), .B(n34014), .Z(n34019) );
  NAND U35321 ( .A(n34017), .B(n34016), .Z(n34018) );
  NAND U35322 ( .A(n34019), .B(n34018), .Z(n34034) );
  XNOR U35323 ( .A(n34033), .B(n34034), .Z(n34025) );
  XNOR U35324 ( .A(n34026), .B(n34025), .Z(n34027) );
  XNOR U35325 ( .A(n34028), .B(n34027), .Z(n34057) );
  XNOR U35326 ( .A(sreg[1825]), .B(n34057), .Z(n34059) );
  NANDN U35327 ( .A(sreg[1824]), .B(n34020), .Z(n34024) );
  NAND U35328 ( .A(n34022), .B(n34021), .Z(n34023) );
  NAND U35329 ( .A(n34024), .B(n34023), .Z(n34058) );
  XNOR U35330 ( .A(n34059), .B(n34058), .Z(c[1825]) );
  NANDN U35331 ( .A(n34026), .B(n34025), .Z(n34030) );
  NANDN U35332 ( .A(n34028), .B(n34027), .Z(n34029) );
  AND U35333 ( .A(n34030), .B(n34029), .Z(n34065) );
  NANDN U35334 ( .A(n34032), .B(n34031), .Z(n34036) );
  NANDN U35335 ( .A(n34034), .B(n34033), .Z(n34035) );
  AND U35336 ( .A(n34036), .B(n34035), .Z(n34063) );
  NAND U35337 ( .A(n42143), .B(n34037), .Z(n34039) );
  XNOR U35338 ( .A(a[804]), .B(n4186), .Z(n34074) );
  NAND U35339 ( .A(n42144), .B(n34074), .Z(n34038) );
  AND U35340 ( .A(n34039), .B(n34038), .Z(n34089) );
  XOR U35341 ( .A(a[808]), .B(n42012), .Z(n34077) );
  XNOR U35342 ( .A(n34089), .B(n34088), .Z(n34091) );
  AND U35343 ( .A(a[810]), .B(b[0]), .Z(n34041) );
  XNOR U35344 ( .A(n34041), .B(n4071), .Z(n34043) );
  NANDN U35345 ( .A(b[0]), .B(a[809]), .Z(n34042) );
  NAND U35346 ( .A(n34043), .B(n34042), .Z(n34085) );
  XOR U35347 ( .A(a[806]), .B(n42085), .Z(n34078) );
  AND U35348 ( .A(a[802]), .B(b[7]), .Z(n34082) );
  XNOR U35349 ( .A(n34083), .B(n34082), .Z(n34084) );
  XNOR U35350 ( .A(n34085), .B(n34084), .Z(n34090) );
  XOR U35351 ( .A(n34091), .B(n34090), .Z(n34069) );
  NANDN U35352 ( .A(n34046), .B(n34045), .Z(n34050) );
  NANDN U35353 ( .A(n34048), .B(n34047), .Z(n34049) );
  AND U35354 ( .A(n34050), .B(n34049), .Z(n34068) );
  XNOR U35355 ( .A(n34069), .B(n34068), .Z(n34070) );
  NANDN U35356 ( .A(n34052), .B(n34051), .Z(n34056) );
  NAND U35357 ( .A(n34054), .B(n34053), .Z(n34055) );
  NAND U35358 ( .A(n34056), .B(n34055), .Z(n34071) );
  XNOR U35359 ( .A(n34070), .B(n34071), .Z(n34062) );
  XNOR U35360 ( .A(n34063), .B(n34062), .Z(n34064) );
  XNOR U35361 ( .A(n34065), .B(n34064), .Z(n34094) );
  XNOR U35362 ( .A(sreg[1826]), .B(n34094), .Z(n34096) );
  NANDN U35363 ( .A(sreg[1825]), .B(n34057), .Z(n34061) );
  NAND U35364 ( .A(n34059), .B(n34058), .Z(n34060) );
  NAND U35365 ( .A(n34061), .B(n34060), .Z(n34095) );
  XNOR U35366 ( .A(n34096), .B(n34095), .Z(c[1826]) );
  NANDN U35367 ( .A(n34063), .B(n34062), .Z(n34067) );
  NANDN U35368 ( .A(n34065), .B(n34064), .Z(n34066) );
  AND U35369 ( .A(n34067), .B(n34066), .Z(n34102) );
  NANDN U35370 ( .A(n34069), .B(n34068), .Z(n34073) );
  NANDN U35371 ( .A(n34071), .B(n34070), .Z(n34072) );
  AND U35372 ( .A(n34073), .B(n34072), .Z(n34100) );
  NAND U35373 ( .A(n42143), .B(n34074), .Z(n34076) );
  XNOR U35374 ( .A(a[805]), .B(n4186), .Z(n34111) );
  NAND U35375 ( .A(n42144), .B(n34111), .Z(n34075) );
  AND U35376 ( .A(n34076), .B(n34075), .Z(n34126) );
  XOR U35377 ( .A(a[809]), .B(n42012), .Z(n34114) );
  XNOR U35378 ( .A(n34126), .B(n34125), .Z(n34128) );
  XOR U35379 ( .A(a[807]), .B(n42085), .Z(n34115) );
  AND U35380 ( .A(a[803]), .B(b[7]), .Z(n34119) );
  XNOR U35381 ( .A(n34120), .B(n34119), .Z(n34121) );
  AND U35382 ( .A(a[811]), .B(b[0]), .Z(n34079) );
  XNOR U35383 ( .A(n34079), .B(n4071), .Z(n34081) );
  NANDN U35384 ( .A(b[0]), .B(a[810]), .Z(n34080) );
  NAND U35385 ( .A(n34081), .B(n34080), .Z(n34122) );
  XNOR U35386 ( .A(n34121), .B(n34122), .Z(n34127) );
  XOR U35387 ( .A(n34128), .B(n34127), .Z(n34106) );
  NANDN U35388 ( .A(n34083), .B(n34082), .Z(n34087) );
  NANDN U35389 ( .A(n34085), .B(n34084), .Z(n34086) );
  AND U35390 ( .A(n34087), .B(n34086), .Z(n34105) );
  XNOR U35391 ( .A(n34106), .B(n34105), .Z(n34107) );
  NANDN U35392 ( .A(n34089), .B(n34088), .Z(n34093) );
  NAND U35393 ( .A(n34091), .B(n34090), .Z(n34092) );
  NAND U35394 ( .A(n34093), .B(n34092), .Z(n34108) );
  XNOR U35395 ( .A(n34107), .B(n34108), .Z(n34099) );
  XNOR U35396 ( .A(n34100), .B(n34099), .Z(n34101) );
  XNOR U35397 ( .A(n34102), .B(n34101), .Z(n34131) );
  XNOR U35398 ( .A(sreg[1827]), .B(n34131), .Z(n34133) );
  NANDN U35399 ( .A(sreg[1826]), .B(n34094), .Z(n34098) );
  NAND U35400 ( .A(n34096), .B(n34095), .Z(n34097) );
  NAND U35401 ( .A(n34098), .B(n34097), .Z(n34132) );
  XNOR U35402 ( .A(n34133), .B(n34132), .Z(c[1827]) );
  NANDN U35403 ( .A(n34100), .B(n34099), .Z(n34104) );
  NANDN U35404 ( .A(n34102), .B(n34101), .Z(n34103) );
  AND U35405 ( .A(n34104), .B(n34103), .Z(n34139) );
  NANDN U35406 ( .A(n34106), .B(n34105), .Z(n34110) );
  NANDN U35407 ( .A(n34108), .B(n34107), .Z(n34109) );
  AND U35408 ( .A(n34110), .B(n34109), .Z(n34137) );
  NAND U35409 ( .A(n42143), .B(n34111), .Z(n34113) );
  XNOR U35410 ( .A(a[806]), .B(n4187), .Z(n34148) );
  NAND U35411 ( .A(n42144), .B(n34148), .Z(n34112) );
  AND U35412 ( .A(n34113), .B(n34112), .Z(n34163) );
  XOR U35413 ( .A(a[810]), .B(n42012), .Z(n34151) );
  XNOR U35414 ( .A(n34163), .B(n34162), .Z(n34165) );
  XOR U35415 ( .A(a[808]), .B(n42085), .Z(n34155) );
  AND U35416 ( .A(a[804]), .B(b[7]), .Z(n34156) );
  XNOR U35417 ( .A(n34157), .B(n34156), .Z(n34158) );
  AND U35418 ( .A(a[812]), .B(b[0]), .Z(n34116) );
  XNOR U35419 ( .A(n34116), .B(n4071), .Z(n34118) );
  NANDN U35420 ( .A(b[0]), .B(a[811]), .Z(n34117) );
  NAND U35421 ( .A(n34118), .B(n34117), .Z(n34159) );
  XNOR U35422 ( .A(n34158), .B(n34159), .Z(n34164) );
  XOR U35423 ( .A(n34165), .B(n34164), .Z(n34143) );
  NANDN U35424 ( .A(n34120), .B(n34119), .Z(n34124) );
  NANDN U35425 ( .A(n34122), .B(n34121), .Z(n34123) );
  AND U35426 ( .A(n34124), .B(n34123), .Z(n34142) );
  XNOR U35427 ( .A(n34143), .B(n34142), .Z(n34144) );
  NANDN U35428 ( .A(n34126), .B(n34125), .Z(n34130) );
  NAND U35429 ( .A(n34128), .B(n34127), .Z(n34129) );
  NAND U35430 ( .A(n34130), .B(n34129), .Z(n34145) );
  XNOR U35431 ( .A(n34144), .B(n34145), .Z(n34136) );
  XNOR U35432 ( .A(n34137), .B(n34136), .Z(n34138) );
  XNOR U35433 ( .A(n34139), .B(n34138), .Z(n34168) );
  XNOR U35434 ( .A(sreg[1828]), .B(n34168), .Z(n34170) );
  NANDN U35435 ( .A(sreg[1827]), .B(n34131), .Z(n34135) );
  NAND U35436 ( .A(n34133), .B(n34132), .Z(n34134) );
  NAND U35437 ( .A(n34135), .B(n34134), .Z(n34169) );
  XNOR U35438 ( .A(n34170), .B(n34169), .Z(c[1828]) );
  NANDN U35439 ( .A(n34137), .B(n34136), .Z(n34141) );
  NANDN U35440 ( .A(n34139), .B(n34138), .Z(n34140) );
  AND U35441 ( .A(n34141), .B(n34140), .Z(n34176) );
  NANDN U35442 ( .A(n34143), .B(n34142), .Z(n34147) );
  NANDN U35443 ( .A(n34145), .B(n34144), .Z(n34146) );
  AND U35444 ( .A(n34147), .B(n34146), .Z(n34174) );
  NAND U35445 ( .A(n42143), .B(n34148), .Z(n34150) );
  XNOR U35446 ( .A(a[807]), .B(n4187), .Z(n34185) );
  NAND U35447 ( .A(n42144), .B(n34185), .Z(n34149) );
  AND U35448 ( .A(n34150), .B(n34149), .Z(n34200) );
  XOR U35449 ( .A(a[811]), .B(n42012), .Z(n34188) );
  XNOR U35450 ( .A(n34200), .B(n34199), .Z(n34202) );
  AND U35451 ( .A(a[813]), .B(b[0]), .Z(n34152) );
  XNOR U35452 ( .A(n34152), .B(n4071), .Z(n34154) );
  NANDN U35453 ( .A(b[0]), .B(a[812]), .Z(n34153) );
  NAND U35454 ( .A(n34154), .B(n34153), .Z(n34196) );
  XOR U35455 ( .A(a[809]), .B(n42085), .Z(n34189) );
  AND U35456 ( .A(a[805]), .B(b[7]), .Z(n34193) );
  XNOR U35457 ( .A(n34194), .B(n34193), .Z(n34195) );
  XNOR U35458 ( .A(n34196), .B(n34195), .Z(n34201) );
  XOR U35459 ( .A(n34202), .B(n34201), .Z(n34180) );
  NANDN U35460 ( .A(n34157), .B(n34156), .Z(n34161) );
  NANDN U35461 ( .A(n34159), .B(n34158), .Z(n34160) );
  AND U35462 ( .A(n34161), .B(n34160), .Z(n34179) );
  XNOR U35463 ( .A(n34180), .B(n34179), .Z(n34181) );
  NANDN U35464 ( .A(n34163), .B(n34162), .Z(n34167) );
  NAND U35465 ( .A(n34165), .B(n34164), .Z(n34166) );
  NAND U35466 ( .A(n34167), .B(n34166), .Z(n34182) );
  XNOR U35467 ( .A(n34181), .B(n34182), .Z(n34173) );
  XNOR U35468 ( .A(n34174), .B(n34173), .Z(n34175) );
  XNOR U35469 ( .A(n34176), .B(n34175), .Z(n34205) );
  XNOR U35470 ( .A(sreg[1829]), .B(n34205), .Z(n34207) );
  NANDN U35471 ( .A(sreg[1828]), .B(n34168), .Z(n34172) );
  NAND U35472 ( .A(n34170), .B(n34169), .Z(n34171) );
  NAND U35473 ( .A(n34172), .B(n34171), .Z(n34206) );
  XNOR U35474 ( .A(n34207), .B(n34206), .Z(c[1829]) );
  NANDN U35475 ( .A(n34174), .B(n34173), .Z(n34178) );
  NANDN U35476 ( .A(n34176), .B(n34175), .Z(n34177) );
  AND U35477 ( .A(n34178), .B(n34177), .Z(n34213) );
  NANDN U35478 ( .A(n34180), .B(n34179), .Z(n34184) );
  NANDN U35479 ( .A(n34182), .B(n34181), .Z(n34183) );
  AND U35480 ( .A(n34184), .B(n34183), .Z(n34211) );
  NAND U35481 ( .A(n42143), .B(n34185), .Z(n34187) );
  XNOR U35482 ( .A(a[808]), .B(n4187), .Z(n34222) );
  NAND U35483 ( .A(n42144), .B(n34222), .Z(n34186) );
  AND U35484 ( .A(n34187), .B(n34186), .Z(n34237) );
  XOR U35485 ( .A(a[812]), .B(n42012), .Z(n34225) );
  XNOR U35486 ( .A(n34237), .B(n34236), .Z(n34239) );
  XOR U35487 ( .A(a[810]), .B(n42085), .Z(n34229) );
  AND U35488 ( .A(a[806]), .B(b[7]), .Z(n34230) );
  XNOR U35489 ( .A(n34231), .B(n34230), .Z(n34232) );
  AND U35490 ( .A(a[814]), .B(b[0]), .Z(n34190) );
  XNOR U35491 ( .A(n34190), .B(n4071), .Z(n34192) );
  NANDN U35492 ( .A(b[0]), .B(a[813]), .Z(n34191) );
  NAND U35493 ( .A(n34192), .B(n34191), .Z(n34233) );
  XNOR U35494 ( .A(n34232), .B(n34233), .Z(n34238) );
  XOR U35495 ( .A(n34239), .B(n34238), .Z(n34217) );
  NANDN U35496 ( .A(n34194), .B(n34193), .Z(n34198) );
  NANDN U35497 ( .A(n34196), .B(n34195), .Z(n34197) );
  AND U35498 ( .A(n34198), .B(n34197), .Z(n34216) );
  XNOR U35499 ( .A(n34217), .B(n34216), .Z(n34218) );
  NANDN U35500 ( .A(n34200), .B(n34199), .Z(n34204) );
  NAND U35501 ( .A(n34202), .B(n34201), .Z(n34203) );
  NAND U35502 ( .A(n34204), .B(n34203), .Z(n34219) );
  XNOR U35503 ( .A(n34218), .B(n34219), .Z(n34210) );
  XNOR U35504 ( .A(n34211), .B(n34210), .Z(n34212) );
  XNOR U35505 ( .A(n34213), .B(n34212), .Z(n34242) );
  XNOR U35506 ( .A(sreg[1830]), .B(n34242), .Z(n34244) );
  NANDN U35507 ( .A(sreg[1829]), .B(n34205), .Z(n34209) );
  NAND U35508 ( .A(n34207), .B(n34206), .Z(n34208) );
  NAND U35509 ( .A(n34209), .B(n34208), .Z(n34243) );
  XNOR U35510 ( .A(n34244), .B(n34243), .Z(c[1830]) );
  NANDN U35511 ( .A(n34211), .B(n34210), .Z(n34215) );
  NANDN U35512 ( .A(n34213), .B(n34212), .Z(n34214) );
  AND U35513 ( .A(n34215), .B(n34214), .Z(n34250) );
  NANDN U35514 ( .A(n34217), .B(n34216), .Z(n34221) );
  NANDN U35515 ( .A(n34219), .B(n34218), .Z(n34220) );
  AND U35516 ( .A(n34221), .B(n34220), .Z(n34248) );
  NAND U35517 ( .A(n42143), .B(n34222), .Z(n34224) );
  XNOR U35518 ( .A(a[809]), .B(n4187), .Z(n34259) );
  NAND U35519 ( .A(n42144), .B(n34259), .Z(n34223) );
  AND U35520 ( .A(n34224), .B(n34223), .Z(n34274) );
  XOR U35521 ( .A(a[813]), .B(n42012), .Z(n34262) );
  XNOR U35522 ( .A(n34274), .B(n34273), .Z(n34276) );
  AND U35523 ( .A(a[815]), .B(b[0]), .Z(n34226) );
  XNOR U35524 ( .A(n34226), .B(n4071), .Z(n34228) );
  NANDN U35525 ( .A(b[0]), .B(a[814]), .Z(n34227) );
  NAND U35526 ( .A(n34228), .B(n34227), .Z(n34270) );
  XOR U35527 ( .A(a[811]), .B(n42085), .Z(n34266) );
  AND U35528 ( .A(a[807]), .B(b[7]), .Z(n34267) );
  XNOR U35529 ( .A(n34268), .B(n34267), .Z(n34269) );
  XNOR U35530 ( .A(n34270), .B(n34269), .Z(n34275) );
  XOR U35531 ( .A(n34276), .B(n34275), .Z(n34254) );
  NANDN U35532 ( .A(n34231), .B(n34230), .Z(n34235) );
  NANDN U35533 ( .A(n34233), .B(n34232), .Z(n34234) );
  AND U35534 ( .A(n34235), .B(n34234), .Z(n34253) );
  XNOR U35535 ( .A(n34254), .B(n34253), .Z(n34255) );
  NANDN U35536 ( .A(n34237), .B(n34236), .Z(n34241) );
  NAND U35537 ( .A(n34239), .B(n34238), .Z(n34240) );
  NAND U35538 ( .A(n34241), .B(n34240), .Z(n34256) );
  XNOR U35539 ( .A(n34255), .B(n34256), .Z(n34247) );
  XNOR U35540 ( .A(n34248), .B(n34247), .Z(n34249) );
  XNOR U35541 ( .A(n34250), .B(n34249), .Z(n34279) );
  XNOR U35542 ( .A(sreg[1831]), .B(n34279), .Z(n34281) );
  NANDN U35543 ( .A(sreg[1830]), .B(n34242), .Z(n34246) );
  NAND U35544 ( .A(n34244), .B(n34243), .Z(n34245) );
  NAND U35545 ( .A(n34246), .B(n34245), .Z(n34280) );
  XNOR U35546 ( .A(n34281), .B(n34280), .Z(c[1831]) );
  NANDN U35547 ( .A(n34248), .B(n34247), .Z(n34252) );
  NANDN U35548 ( .A(n34250), .B(n34249), .Z(n34251) );
  AND U35549 ( .A(n34252), .B(n34251), .Z(n34287) );
  NANDN U35550 ( .A(n34254), .B(n34253), .Z(n34258) );
  NANDN U35551 ( .A(n34256), .B(n34255), .Z(n34257) );
  AND U35552 ( .A(n34258), .B(n34257), .Z(n34285) );
  NAND U35553 ( .A(n42143), .B(n34259), .Z(n34261) );
  XNOR U35554 ( .A(a[810]), .B(n4187), .Z(n34296) );
  NAND U35555 ( .A(n42144), .B(n34296), .Z(n34260) );
  AND U35556 ( .A(n34261), .B(n34260), .Z(n34311) );
  XOR U35557 ( .A(a[814]), .B(n42012), .Z(n34299) );
  XNOR U35558 ( .A(n34311), .B(n34310), .Z(n34313) );
  AND U35559 ( .A(a[816]), .B(b[0]), .Z(n34263) );
  XNOR U35560 ( .A(n34263), .B(n4071), .Z(n34265) );
  NANDN U35561 ( .A(b[0]), .B(a[815]), .Z(n34264) );
  NAND U35562 ( .A(n34265), .B(n34264), .Z(n34307) );
  XOR U35563 ( .A(a[812]), .B(n42085), .Z(n34300) );
  AND U35564 ( .A(a[808]), .B(b[7]), .Z(n34304) );
  XNOR U35565 ( .A(n34305), .B(n34304), .Z(n34306) );
  XNOR U35566 ( .A(n34307), .B(n34306), .Z(n34312) );
  XOR U35567 ( .A(n34313), .B(n34312), .Z(n34291) );
  NANDN U35568 ( .A(n34268), .B(n34267), .Z(n34272) );
  NANDN U35569 ( .A(n34270), .B(n34269), .Z(n34271) );
  AND U35570 ( .A(n34272), .B(n34271), .Z(n34290) );
  XNOR U35571 ( .A(n34291), .B(n34290), .Z(n34292) );
  NANDN U35572 ( .A(n34274), .B(n34273), .Z(n34278) );
  NAND U35573 ( .A(n34276), .B(n34275), .Z(n34277) );
  NAND U35574 ( .A(n34278), .B(n34277), .Z(n34293) );
  XNOR U35575 ( .A(n34292), .B(n34293), .Z(n34284) );
  XNOR U35576 ( .A(n34285), .B(n34284), .Z(n34286) );
  XNOR U35577 ( .A(n34287), .B(n34286), .Z(n34316) );
  XNOR U35578 ( .A(sreg[1832]), .B(n34316), .Z(n34318) );
  NANDN U35579 ( .A(sreg[1831]), .B(n34279), .Z(n34283) );
  NAND U35580 ( .A(n34281), .B(n34280), .Z(n34282) );
  NAND U35581 ( .A(n34283), .B(n34282), .Z(n34317) );
  XNOR U35582 ( .A(n34318), .B(n34317), .Z(c[1832]) );
  NANDN U35583 ( .A(n34285), .B(n34284), .Z(n34289) );
  NANDN U35584 ( .A(n34287), .B(n34286), .Z(n34288) );
  AND U35585 ( .A(n34289), .B(n34288), .Z(n34324) );
  NANDN U35586 ( .A(n34291), .B(n34290), .Z(n34295) );
  NANDN U35587 ( .A(n34293), .B(n34292), .Z(n34294) );
  AND U35588 ( .A(n34295), .B(n34294), .Z(n34322) );
  NAND U35589 ( .A(n42143), .B(n34296), .Z(n34298) );
  XNOR U35590 ( .A(a[811]), .B(n4187), .Z(n34333) );
  NAND U35591 ( .A(n42144), .B(n34333), .Z(n34297) );
  AND U35592 ( .A(n34298), .B(n34297), .Z(n34348) );
  XOR U35593 ( .A(a[815]), .B(n42012), .Z(n34336) );
  XNOR U35594 ( .A(n34348), .B(n34347), .Z(n34350) );
  XOR U35595 ( .A(a[813]), .B(n42085), .Z(n34340) );
  AND U35596 ( .A(a[809]), .B(b[7]), .Z(n34341) );
  XNOR U35597 ( .A(n34342), .B(n34341), .Z(n34343) );
  AND U35598 ( .A(a[817]), .B(b[0]), .Z(n34301) );
  XNOR U35599 ( .A(n34301), .B(n4071), .Z(n34303) );
  NANDN U35600 ( .A(b[0]), .B(a[816]), .Z(n34302) );
  NAND U35601 ( .A(n34303), .B(n34302), .Z(n34344) );
  XNOR U35602 ( .A(n34343), .B(n34344), .Z(n34349) );
  XOR U35603 ( .A(n34350), .B(n34349), .Z(n34328) );
  NANDN U35604 ( .A(n34305), .B(n34304), .Z(n34309) );
  NANDN U35605 ( .A(n34307), .B(n34306), .Z(n34308) );
  AND U35606 ( .A(n34309), .B(n34308), .Z(n34327) );
  XNOR U35607 ( .A(n34328), .B(n34327), .Z(n34329) );
  NANDN U35608 ( .A(n34311), .B(n34310), .Z(n34315) );
  NAND U35609 ( .A(n34313), .B(n34312), .Z(n34314) );
  NAND U35610 ( .A(n34315), .B(n34314), .Z(n34330) );
  XNOR U35611 ( .A(n34329), .B(n34330), .Z(n34321) );
  XNOR U35612 ( .A(n34322), .B(n34321), .Z(n34323) );
  XNOR U35613 ( .A(n34324), .B(n34323), .Z(n34353) );
  XNOR U35614 ( .A(sreg[1833]), .B(n34353), .Z(n34355) );
  NANDN U35615 ( .A(sreg[1832]), .B(n34316), .Z(n34320) );
  NAND U35616 ( .A(n34318), .B(n34317), .Z(n34319) );
  NAND U35617 ( .A(n34320), .B(n34319), .Z(n34354) );
  XNOR U35618 ( .A(n34355), .B(n34354), .Z(c[1833]) );
  NANDN U35619 ( .A(n34322), .B(n34321), .Z(n34326) );
  NANDN U35620 ( .A(n34324), .B(n34323), .Z(n34325) );
  AND U35621 ( .A(n34326), .B(n34325), .Z(n34361) );
  NANDN U35622 ( .A(n34328), .B(n34327), .Z(n34332) );
  NANDN U35623 ( .A(n34330), .B(n34329), .Z(n34331) );
  AND U35624 ( .A(n34332), .B(n34331), .Z(n34359) );
  NAND U35625 ( .A(n42143), .B(n34333), .Z(n34335) );
  XNOR U35626 ( .A(a[812]), .B(n4187), .Z(n34370) );
  NAND U35627 ( .A(n42144), .B(n34370), .Z(n34334) );
  AND U35628 ( .A(n34335), .B(n34334), .Z(n34385) );
  XOR U35629 ( .A(a[816]), .B(n42012), .Z(n34373) );
  XNOR U35630 ( .A(n34385), .B(n34384), .Z(n34387) );
  AND U35631 ( .A(a[818]), .B(b[0]), .Z(n34337) );
  XNOR U35632 ( .A(n34337), .B(n4071), .Z(n34339) );
  NANDN U35633 ( .A(b[0]), .B(a[817]), .Z(n34338) );
  NAND U35634 ( .A(n34339), .B(n34338), .Z(n34381) );
  XOR U35635 ( .A(a[814]), .B(n42085), .Z(n34374) );
  AND U35636 ( .A(a[810]), .B(b[7]), .Z(n34378) );
  XNOR U35637 ( .A(n34379), .B(n34378), .Z(n34380) );
  XNOR U35638 ( .A(n34381), .B(n34380), .Z(n34386) );
  XOR U35639 ( .A(n34387), .B(n34386), .Z(n34365) );
  NANDN U35640 ( .A(n34342), .B(n34341), .Z(n34346) );
  NANDN U35641 ( .A(n34344), .B(n34343), .Z(n34345) );
  AND U35642 ( .A(n34346), .B(n34345), .Z(n34364) );
  XNOR U35643 ( .A(n34365), .B(n34364), .Z(n34366) );
  NANDN U35644 ( .A(n34348), .B(n34347), .Z(n34352) );
  NAND U35645 ( .A(n34350), .B(n34349), .Z(n34351) );
  NAND U35646 ( .A(n34352), .B(n34351), .Z(n34367) );
  XNOR U35647 ( .A(n34366), .B(n34367), .Z(n34358) );
  XNOR U35648 ( .A(n34359), .B(n34358), .Z(n34360) );
  XNOR U35649 ( .A(n34361), .B(n34360), .Z(n34390) );
  XNOR U35650 ( .A(sreg[1834]), .B(n34390), .Z(n34392) );
  NANDN U35651 ( .A(sreg[1833]), .B(n34353), .Z(n34357) );
  NAND U35652 ( .A(n34355), .B(n34354), .Z(n34356) );
  NAND U35653 ( .A(n34357), .B(n34356), .Z(n34391) );
  XNOR U35654 ( .A(n34392), .B(n34391), .Z(c[1834]) );
  NANDN U35655 ( .A(n34359), .B(n34358), .Z(n34363) );
  NANDN U35656 ( .A(n34361), .B(n34360), .Z(n34362) );
  AND U35657 ( .A(n34363), .B(n34362), .Z(n34398) );
  NANDN U35658 ( .A(n34365), .B(n34364), .Z(n34369) );
  NANDN U35659 ( .A(n34367), .B(n34366), .Z(n34368) );
  AND U35660 ( .A(n34369), .B(n34368), .Z(n34396) );
  NAND U35661 ( .A(n42143), .B(n34370), .Z(n34372) );
  XNOR U35662 ( .A(a[813]), .B(n4188), .Z(n34407) );
  NAND U35663 ( .A(n42144), .B(n34407), .Z(n34371) );
  AND U35664 ( .A(n34372), .B(n34371), .Z(n34422) );
  XOR U35665 ( .A(a[817]), .B(n42012), .Z(n34410) );
  XNOR U35666 ( .A(n34422), .B(n34421), .Z(n34424) );
  XOR U35667 ( .A(a[815]), .B(n42085), .Z(n34411) );
  AND U35668 ( .A(a[811]), .B(b[7]), .Z(n34415) );
  XNOR U35669 ( .A(n34416), .B(n34415), .Z(n34417) );
  AND U35670 ( .A(a[819]), .B(b[0]), .Z(n34375) );
  XNOR U35671 ( .A(n34375), .B(n4071), .Z(n34377) );
  NANDN U35672 ( .A(b[0]), .B(a[818]), .Z(n34376) );
  NAND U35673 ( .A(n34377), .B(n34376), .Z(n34418) );
  XNOR U35674 ( .A(n34417), .B(n34418), .Z(n34423) );
  XOR U35675 ( .A(n34424), .B(n34423), .Z(n34402) );
  NANDN U35676 ( .A(n34379), .B(n34378), .Z(n34383) );
  NANDN U35677 ( .A(n34381), .B(n34380), .Z(n34382) );
  AND U35678 ( .A(n34383), .B(n34382), .Z(n34401) );
  XNOR U35679 ( .A(n34402), .B(n34401), .Z(n34403) );
  NANDN U35680 ( .A(n34385), .B(n34384), .Z(n34389) );
  NAND U35681 ( .A(n34387), .B(n34386), .Z(n34388) );
  NAND U35682 ( .A(n34389), .B(n34388), .Z(n34404) );
  XNOR U35683 ( .A(n34403), .B(n34404), .Z(n34395) );
  XNOR U35684 ( .A(n34396), .B(n34395), .Z(n34397) );
  XNOR U35685 ( .A(n34398), .B(n34397), .Z(n34427) );
  XNOR U35686 ( .A(sreg[1835]), .B(n34427), .Z(n34429) );
  NANDN U35687 ( .A(sreg[1834]), .B(n34390), .Z(n34394) );
  NAND U35688 ( .A(n34392), .B(n34391), .Z(n34393) );
  NAND U35689 ( .A(n34394), .B(n34393), .Z(n34428) );
  XNOR U35690 ( .A(n34429), .B(n34428), .Z(c[1835]) );
  NANDN U35691 ( .A(n34396), .B(n34395), .Z(n34400) );
  NANDN U35692 ( .A(n34398), .B(n34397), .Z(n34399) );
  AND U35693 ( .A(n34400), .B(n34399), .Z(n34435) );
  NANDN U35694 ( .A(n34402), .B(n34401), .Z(n34406) );
  NANDN U35695 ( .A(n34404), .B(n34403), .Z(n34405) );
  AND U35696 ( .A(n34406), .B(n34405), .Z(n34433) );
  NAND U35697 ( .A(n42143), .B(n34407), .Z(n34409) );
  XNOR U35698 ( .A(a[814]), .B(n4188), .Z(n34444) );
  NAND U35699 ( .A(n42144), .B(n34444), .Z(n34408) );
  AND U35700 ( .A(n34409), .B(n34408), .Z(n34459) );
  XOR U35701 ( .A(a[818]), .B(n42012), .Z(n34447) );
  XNOR U35702 ( .A(n34459), .B(n34458), .Z(n34461) );
  XOR U35703 ( .A(a[816]), .B(n42085), .Z(n34448) );
  AND U35704 ( .A(a[812]), .B(b[7]), .Z(n34452) );
  XNOR U35705 ( .A(n34453), .B(n34452), .Z(n34454) );
  AND U35706 ( .A(a[820]), .B(b[0]), .Z(n34412) );
  XNOR U35707 ( .A(n34412), .B(n4071), .Z(n34414) );
  NANDN U35708 ( .A(b[0]), .B(a[819]), .Z(n34413) );
  NAND U35709 ( .A(n34414), .B(n34413), .Z(n34455) );
  XNOR U35710 ( .A(n34454), .B(n34455), .Z(n34460) );
  XOR U35711 ( .A(n34461), .B(n34460), .Z(n34439) );
  NANDN U35712 ( .A(n34416), .B(n34415), .Z(n34420) );
  NANDN U35713 ( .A(n34418), .B(n34417), .Z(n34419) );
  AND U35714 ( .A(n34420), .B(n34419), .Z(n34438) );
  XNOR U35715 ( .A(n34439), .B(n34438), .Z(n34440) );
  NANDN U35716 ( .A(n34422), .B(n34421), .Z(n34426) );
  NAND U35717 ( .A(n34424), .B(n34423), .Z(n34425) );
  NAND U35718 ( .A(n34426), .B(n34425), .Z(n34441) );
  XNOR U35719 ( .A(n34440), .B(n34441), .Z(n34432) );
  XNOR U35720 ( .A(n34433), .B(n34432), .Z(n34434) );
  XNOR U35721 ( .A(n34435), .B(n34434), .Z(n34464) );
  XNOR U35722 ( .A(sreg[1836]), .B(n34464), .Z(n34466) );
  NANDN U35723 ( .A(sreg[1835]), .B(n34427), .Z(n34431) );
  NAND U35724 ( .A(n34429), .B(n34428), .Z(n34430) );
  NAND U35725 ( .A(n34431), .B(n34430), .Z(n34465) );
  XNOR U35726 ( .A(n34466), .B(n34465), .Z(c[1836]) );
  NANDN U35727 ( .A(n34433), .B(n34432), .Z(n34437) );
  NANDN U35728 ( .A(n34435), .B(n34434), .Z(n34436) );
  AND U35729 ( .A(n34437), .B(n34436), .Z(n34472) );
  NANDN U35730 ( .A(n34439), .B(n34438), .Z(n34443) );
  NANDN U35731 ( .A(n34441), .B(n34440), .Z(n34442) );
  AND U35732 ( .A(n34443), .B(n34442), .Z(n34470) );
  NAND U35733 ( .A(n42143), .B(n34444), .Z(n34446) );
  XNOR U35734 ( .A(a[815]), .B(n4188), .Z(n34481) );
  NAND U35735 ( .A(n42144), .B(n34481), .Z(n34445) );
  AND U35736 ( .A(n34446), .B(n34445), .Z(n34496) );
  XOR U35737 ( .A(a[819]), .B(n42012), .Z(n34484) );
  XNOR U35738 ( .A(n34496), .B(n34495), .Z(n34498) );
  XOR U35739 ( .A(a[817]), .B(n42085), .Z(n34485) );
  AND U35740 ( .A(a[813]), .B(b[7]), .Z(n34489) );
  XNOR U35741 ( .A(n34490), .B(n34489), .Z(n34491) );
  AND U35742 ( .A(a[821]), .B(b[0]), .Z(n34449) );
  XNOR U35743 ( .A(n34449), .B(n4071), .Z(n34451) );
  NANDN U35744 ( .A(b[0]), .B(a[820]), .Z(n34450) );
  NAND U35745 ( .A(n34451), .B(n34450), .Z(n34492) );
  XNOR U35746 ( .A(n34491), .B(n34492), .Z(n34497) );
  XOR U35747 ( .A(n34498), .B(n34497), .Z(n34476) );
  NANDN U35748 ( .A(n34453), .B(n34452), .Z(n34457) );
  NANDN U35749 ( .A(n34455), .B(n34454), .Z(n34456) );
  AND U35750 ( .A(n34457), .B(n34456), .Z(n34475) );
  XNOR U35751 ( .A(n34476), .B(n34475), .Z(n34477) );
  NANDN U35752 ( .A(n34459), .B(n34458), .Z(n34463) );
  NAND U35753 ( .A(n34461), .B(n34460), .Z(n34462) );
  NAND U35754 ( .A(n34463), .B(n34462), .Z(n34478) );
  XNOR U35755 ( .A(n34477), .B(n34478), .Z(n34469) );
  XNOR U35756 ( .A(n34470), .B(n34469), .Z(n34471) );
  XNOR U35757 ( .A(n34472), .B(n34471), .Z(n34501) );
  XNOR U35758 ( .A(sreg[1837]), .B(n34501), .Z(n34503) );
  NANDN U35759 ( .A(sreg[1836]), .B(n34464), .Z(n34468) );
  NAND U35760 ( .A(n34466), .B(n34465), .Z(n34467) );
  NAND U35761 ( .A(n34468), .B(n34467), .Z(n34502) );
  XNOR U35762 ( .A(n34503), .B(n34502), .Z(c[1837]) );
  NANDN U35763 ( .A(n34470), .B(n34469), .Z(n34474) );
  NANDN U35764 ( .A(n34472), .B(n34471), .Z(n34473) );
  AND U35765 ( .A(n34474), .B(n34473), .Z(n34509) );
  NANDN U35766 ( .A(n34476), .B(n34475), .Z(n34480) );
  NANDN U35767 ( .A(n34478), .B(n34477), .Z(n34479) );
  AND U35768 ( .A(n34480), .B(n34479), .Z(n34507) );
  NAND U35769 ( .A(n42143), .B(n34481), .Z(n34483) );
  XNOR U35770 ( .A(a[816]), .B(n4188), .Z(n34518) );
  NAND U35771 ( .A(n42144), .B(n34518), .Z(n34482) );
  AND U35772 ( .A(n34483), .B(n34482), .Z(n34533) );
  XOR U35773 ( .A(a[820]), .B(n42012), .Z(n34521) );
  XNOR U35774 ( .A(n34533), .B(n34532), .Z(n34535) );
  XOR U35775 ( .A(a[818]), .B(n42085), .Z(n34525) );
  AND U35776 ( .A(a[814]), .B(b[7]), .Z(n34526) );
  XNOR U35777 ( .A(n34527), .B(n34526), .Z(n34528) );
  AND U35778 ( .A(a[822]), .B(b[0]), .Z(n34486) );
  XNOR U35779 ( .A(n34486), .B(n4071), .Z(n34488) );
  NANDN U35780 ( .A(b[0]), .B(a[821]), .Z(n34487) );
  NAND U35781 ( .A(n34488), .B(n34487), .Z(n34529) );
  XNOR U35782 ( .A(n34528), .B(n34529), .Z(n34534) );
  XOR U35783 ( .A(n34535), .B(n34534), .Z(n34513) );
  NANDN U35784 ( .A(n34490), .B(n34489), .Z(n34494) );
  NANDN U35785 ( .A(n34492), .B(n34491), .Z(n34493) );
  AND U35786 ( .A(n34494), .B(n34493), .Z(n34512) );
  XNOR U35787 ( .A(n34513), .B(n34512), .Z(n34514) );
  NANDN U35788 ( .A(n34496), .B(n34495), .Z(n34500) );
  NAND U35789 ( .A(n34498), .B(n34497), .Z(n34499) );
  NAND U35790 ( .A(n34500), .B(n34499), .Z(n34515) );
  XNOR U35791 ( .A(n34514), .B(n34515), .Z(n34506) );
  XNOR U35792 ( .A(n34507), .B(n34506), .Z(n34508) );
  XNOR U35793 ( .A(n34509), .B(n34508), .Z(n34538) );
  XNOR U35794 ( .A(sreg[1838]), .B(n34538), .Z(n34540) );
  NANDN U35795 ( .A(sreg[1837]), .B(n34501), .Z(n34505) );
  NAND U35796 ( .A(n34503), .B(n34502), .Z(n34504) );
  NAND U35797 ( .A(n34505), .B(n34504), .Z(n34539) );
  XNOR U35798 ( .A(n34540), .B(n34539), .Z(c[1838]) );
  NANDN U35799 ( .A(n34507), .B(n34506), .Z(n34511) );
  NANDN U35800 ( .A(n34509), .B(n34508), .Z(n34510) );
  AND U35801 ( .A(n34511), .B(n34510), .Z(n34546) );
  NANDN U35802 ( .A(n34513), .B(n34512), .Z(n34517) );
  NANDN U35803 ( .A(n34515), .B(n34514), .Z(n34516) );
  AND U35804 ( .A(n34517), .B(n34516), .Z(n34544) );
  NAND U35805 ( .A(n42143), .B(n34518), .Z(n34520) );
  XNOR U35806 ( .A(a[817]), .B(n4188), .Z(n34555) );
  NAND U35807 ( .A(n42144), .B(n34555), .Z(n34519) );
  AND U35808 ( .A(n34520), .B(n34519), .Z(n34570) );
  XOR U35809 ( .A(a[821]), .B(n42012), .Z(n34558) );
  XNOR U35810 ( .A(n34570), .B(n34569), .Z(n34572) );
  AND U35811 ( .A(a[823]), .B(b[0]), .Z(n34522) );
  XNOR U35812 ( .A(n34522), .B(n4071), .Z(n34524) );
  NANDN U35813 ( .A(b[0]), .B(a[822]), .Z(n34523) );
  NAND U35814 ( .A(n34524), .B(n34523), .Z(n34566) );
  XOR U35815 ( .A(a[819]), .B(n42085), .Z(n34562) );
  AND U35816 ( .A(a[815]), .B(b[7]), .Z(n34563) );
  XNOR U35817 ( .A(n34564), .B(n34563), .Z(n34565) );
  XNOR U35818 ( .A(n34566), .B(n34565), .Z(n34571) );
  XOR U35819 ( .A(n34572), .B(n34571), .Z(n34550) );
  NANDN U35820 ( .A(n34527), .B(n34526), .Z(n34531) );
  NANDN U35821 ( .A(n34529), .B(n34528), .Z(n34530) );
  AND U35822 ( .A(n34531), .B(n34530), .Z(n34549) );
  XNOR U35823 ( .A(n34550), .B(n34549), .Z(n34551) );
  NANDN U35824 ( .A(n34533), .B(n34532), .Z(n34537) );
  NAND U35825 ( .A(n34535), .B(n34534), .Z(n34536) );
  NAND U35826 ( .A(n34537), .B(n34536), .Z(n34552) );
  XNOR U35827 ( .A(n34551), .B(n34552), .Z(n34543) );
  XNOR U35828 ( .A(n34544), .B(n34543), .Z(n34545) );
  XNOR U35829 ( .A(n34546), .B(n34545), .Z(n34575) );
  XNOR U35830 ( .A(sreg[1839]), .B(n34575), .Z(n34577) );
  NANDN U35831 ( .A(sreg[1838]), .B(n34538), .Z(n34542) );
  NAND U35832 ( .A(n34540), .B(n34539), .Z(n34541) );
  NAND U35833 ( .A(n34542), .B(n34541), .Z(n34576) );
  XNOR U35834 ( .A(n34577), .B(n34576), .Z(c[1839]) );
  NANDN U35835 ( .A(n34544), .B(n34543), .Z(n34548) );
  NANDN U35836 ( .A(n34546), .B(n34545), .Z(n34547) );
  AND U35837 ( .A(n34548), .B(n34547), .Z(n34583) );
  NANDN U35838 ( .A(n34550), .B(n34549), .Z(n34554) );
  NANDN U35839 ( .A(n34552), .B(n34551), .Z(n34553) );
  AND U35840 ( .A(n34554), .B(n34553), .Z(n34581) );
  NAND U35841 ( .A(n42143), .B(n34555), .Z(n34557) );
  XNOR U35842 ( .A(a[818]), .B(n4188), .Z(n34592) );
  NAND U35843 ( .A(n42144), .B(n34592), .Z(n34556) );
  AND U35844 ( .A(n34557), .B(n34556), .Z(n34607) );
  XOR U35845 ( .A(a[822]), .B(n42012), .Z(n34595) );
  XNOR U35846 ( .A(n34607), .B(n34606), .Z(n34609) );
  AND U35847 ( .A(a[824]), .B(b[0]), .Z(n34559) );
  XNOR U35848 ( .A(n34559), .B(n4071), .Z(n34561) );
  NANDN U35849 ( .A(b[0]), .B(a[823]), .Z(n34560) );
  NAND U35850 ( .A(n34561), .B(n34560), .Z(n34603) );
  XOR U35851 ( .A(a[820]), .B(n42085), .Z(n34596) );
  AND U35852 ( .A(a[816]), .B(b[7]), .Z(n34600) );
  XNOR U35853 ( .A(n34601), .B(n34600), .Z(n34602) );
  XNOR U35854 ( .A(n34603), .B(n34602), .Z(n34608) );
  XOR U35855 ( .A(n34609), .B(n34608), .Z(n34587) );
  NANDN U35856 ( .A(n34564), .B(n34563), .Z(n34568) );
  NANDN U35857 ( .A(n34566), .B(n34565), .Z(n34567) );
  AND U35858 ( .A(n34568), .B(n34567), .Z(n34586) );
  XNOR U35859 ( .A(n34587), .B(n34586), .Z(n34588) );
  NANDN U35860 ( .A(n34570), .B(n34569), .Z(n34574) );
  NAND U35861 ( .A(n34572), .B(n34571), .Z(n34573) );
  NAND U35862 ( .A(n34574), .B(n34573), .Z(n34589) );
  XNOR U35863 ( .A(n34588), .B(n34589), .Z(n34580) );
  XNOR U35864 ( .A(n34581), .B(n34580), .Z(n34582) );
  XNOR U35865 ( .A(n34583), .B(n34582), .Z(n34612) );
  XNOR U35866 ( .A(sreg[1840]), .B(n34612), .Z(n34614) );
  NANDN U35867 ( .A(sreg[1839]), .B(n34575), .Z(n34579) );
  NAND U35868 ( .A(n34577), .B(n34576), .Z(n34578) );
  NAND U35869 ( .A(n34579), .B(n34578), .Z(n34613) );
  XNOR U35870 ( .A(n34614), .B(n34613), .Z(c[1840]) );
  NANDN U35871 ( .A(n34581), .B(n34580), .Z(n34585) );
  NANDN U35872 ( .A(n34583), .B(n34582), .Z(n34584) );
  AND U35873 ( .A(n34585), .B(n34584), .Z(n34620) );
  NANDN U35874 ( .A(n34587), .B(n34586), .Z(n34591) );
  NANDN U35875 ( .A(n34589), .B(n34588), .Z(n34590) );
  AND U35876 ( .A(n34591), .B(n34590), .Z(n34618) );
  NAND U35877 ( .A(n42143), .B(n34592), .Z(n34594) );
  XNOR U35878 ( .A(a[819]), .B(n4188), .Z(n34629) );
  NAND U35879 ( .A(n42144), .B(n34629), .Z(n34593) );
  AND U35880 ( .A(n34594), .B(n34593), .Z(n34644) );
  XOR U35881 ( .A(a[823]), .B(n42012), .Z(n34632) );
  XNOR U35882 ( .A(n34644), .B(n34643), .Z(n34646) );
  XOR U35883 ( .A(a[821]), .B(n42085), .Z(n34636) );
  AND U35884 ( .A(a[817]), .B(b[7]), .Z(n34637) );
  XNOR U35885 ( .A(n34638), .B(n34637), .Z(n34639) );
  AND U35886 ( .A(a[825]), .B(b[0]), .Z(n34597) );
  XNOR U35887 ( .A(n34597), .B(n4071), .Z(n34599) );
  NANDN U35888 ( .A(b[0]), .B(a[824]), .Z(n34598) );
  NAND U35889 ( .A(n34599), .B(n34598), .Z(n34640) );
  XNOR U35890 ( .A(n34639), .B(n34640), .Z(n34645) );
  XOR U35891 ( .A(n34646), .B(n34645), .Z(n34624) );
  NANDN U35892 ( .A(n34601), .B(n34600), .Z(n34605) );
  NANDN U35893 ( .A(n34603), .B(n34602), .Z(n34604) );
  AND U35894 ( .A(n34605), .B(n34604), .Z(n34623) );
  XNOR U35895 ( .A(n34624), .B(n34623), .Z(n34625) );
  NANDN U35896 ( .A(n34607), .B(n34606), .Z(n34611) );
  NAND U35897 ( .A(n34609), .B(n34608), .Z(n34610) );
  NAND U35898 ( .A(n34611), .B(n34610), .Z(n34626) );
  XNOR U35899 ( .A(n34625), .B(n34626), .Z(n34617) );
  XNOR U35900 ( .A(n34618), .B(n34617), .Z(n34619) );
  XNOR U35901 ( .A(n34620), .B(n34619), .Z(n34649) );
  XNOR U35902 ( .A(sreg[1841]), .B(n34649), .Z(n34651) );
  NANDN U35903 ( .A(sreg[1840]), .B(n34612), .Z(n34616) );
  NAND U35904 ( .A(n34614), .B(n34613), .Z(n34615) );
  NAND U35905 ( .A(n34616), .B(n34615), .Z(n34650) );
  XNOR U35906 ( .A(n34651), .B(n34650), .Z(c[1841]) );
  NANDN U35907 ( .A(n34618), .B(n34617), .Z(n34622) );
  NANDN U35908 ( .A(n34620), .B(n34619), .Z(n34621) );
  AND U35909 ( .A(n34622), .B(n34621), .Z(n34657) );
  NANDN U35910 ( .A(n34624), .B(n34623), .Z(n34628) );
  NANDN U35911 ( .A(n34626), .B(n34625), .Z(n34627) );
  AND U35912 ( .A(n34628), .B(n34627), .Z(n34655) );
  NAND U35913 ( .A(n42143), .B(n34629), .Z(n34631) );
  XNOR U35914 ( .A(a[820]), .B(n4189), .Z(n34666) );
  NAND U35915 ( .A(n42144), .B(n34666), .Z(n34630) );
  AND U35916 ( .A(n34631), .B(n34630), .Z(n34681) );
  XOR U35917 ( .A(a[824]), .B(n42012), .Z(n34669) );
  XNOR U35918 ( .A(n34681), .B(n34680), .Z(n34683) );
  AND U35919 ( .A(a[826]), .B(b[0]), .Z(n34633) );
  XNOR U35920 ( .A(n34633), .B(n4071), .Z(n34635) );
  NANDN U35921 ( .A(b[0]), .B(a[825]), .Z(n34634) );
  NAND U35922 ( .A(n34635), .B(n34634), .Z(n34677) );
  XOR U35923 ( .A(a[822]), .B(n42085), .Z(n34670) );
  AND U35924 ( .A(a[818]), .B(b[7]), .Z(n34674) );
  XNOR U35925 ( .A(n34675), .B(n34674), .Z(n34676) );
  XNOR U35926 ( .A(n34677), .B(n34676), .Z(n34682) );
  XOR U35927 ( .A(n34683), .B(n34682), .Z(n34661) );
  NANDN U35928 ( .A(n34638), .B(n34637), .Z(n34642) );
  NANDN U35929 ( .A(n34640), .B(n34639), .Z(n34641) );
  AND U35930 ( .A(n34642), .B(n34641), .Z(n34660) );
  XNOR U35931 ( .A(n34661), .B(n34660), .Z(n34662) );
  NANDN U35932 ( .A(n34644), .B(n34643), .Z(n34648) );
  NAND U35933 ( .A(n34646), .B(n34645), .Z(n34647) );
  NAND U35934 ( .A(n34648), .B(n34647), .Z(n34663) );
  XNOR U35935 ( .A(n34662), .B(n34663), .Z(n34654) );
  XNOR U35936 ( .A(n34655), .B(n34654), .Z(n34656) );
  XNOR U35937 ( .A(n34657), .B(n34656), .Z(n34686) );
  XNOR U35938 ( .A(sreg[1842]), .B(n34686), .Z(n34688) );
  NANDN U35939 ( .A(sreg[1841]), .B(n34649), .Z(n34653) );
  NAND U35940 ( .A(n34651), .B(n34650), .Z(n34652) );
  NAND U35941 ( .A(n34653), .B(n34652), .Z(n34687) );
  XNOR U35942 ( .A(n34688), .B(n34687), .Z(c[1842]) );
  NANDN U35943 ( .A(n34655), .B(n34654), .Z(n34659) );
  NANDN U35944 ( .A(n34657), .B(n34656), .Z(n34658) );
  AND U35945 ( .A(n34659), .B(n34658), .Z(n34694) );
  NANDN U35946 ( .A(n34661), .B(n34660), .Z(n34665) );
  NANDN U35947 ( .A(n34663), .B(n34662), .Z(n34664) );
  AND U35948 ( .A(n34665), .B(n34664), .Z(n34692) );
  NAND U35949 ( .A(n42143), .B(n34666), .Z(n34668) );
  XNOR U35950 ( .A(a[821]), .B(n4189), .Z(n34703) );
  NAND U35951 ( .A(n42144), .B(n34703), .Z(n34667) );
  AND U35952 ( .A(n34668), .B(n34667), .Z(n34718) );
  XOR U35953 ( .A(a[825]), .B(n42012), .Z(n34706) );
  XNOR U35954 ( .A(n34718), .B(n34717), .Z(n34720) );
  XOR U35955 ( .A(a[823]), .B(n42085), .Z(n34707) );
  AND U35956 ( .A(a[819]), .B(b[7]), .Z(n34711) );
  XNOR U35957 ( .A(n34712), .B(n34711), .Z(n34713) );
  AND U35958 ( .A(a[827]), .B(b[0]), .Z(n34671) );
  XNOR U35959 ( .A(n34671), .B(n4071), .Z(n34673) );
  NANDN U35960 ( .A(b[0]), .B(a[826]), .Z(n34672) );
  NAND U35961 ( .A(n34673), .B(n34672), .Z(n34714) );
  XNOR U35962 ( .A(n34713), .B(n34714), .Z(n34719) );
  XOR U35963 ( .A(n34720), .B(n34719), .Z(n34698) );
  NANDN U35964 ( .A(n34675), .B(n34674), .Z(n34679) );
  NANDN U35965 ( .A(n34677), .B(n34676), .Z(n34678) );
  AND U35966 ( .A(n34679), .B(n34678), .Z(n34697) );
  XNOR U35967 ( .A(n34698), .B(n34697), .Z(n34699) );
  NANDN U35968 ( .A(n34681), .B(n34680), .Z(n34685) );
  NAND U35969 ( .A(n34683), .B(n34682), .Z(n34684) );
  NAND U35970 ( .A(n34685), .B(n34684), .Z(n34700) );
  XNOR U35971 ( .A(n34699), .B(n34700), .Z(n34691) );
  XNOR U35972 ( .A(n34692), .B(n34691), .Z(n34693) );
  XNOR U35973 ( .A(n34694), .B(n34693), .Z(n34723) );
  XNOR U35974 ( .A(sreg[1843]), .B(n34723), .Z(n34725) );
  NANDN U35975 ( .A(sreg[1842]), .B(n34686), .Z(n34690) );
  NAND U35976 ( .A(n34688), .B(n34687), .Z(n34689) );
  NAND U35977 ( .A(n34690), .B(n34689), .Z(n34724) );
  XNOR U35978 ( .A(n34725), .B(n34724), .Z(c[1843]) );
  NANDN U35979 ( .A(n34692), .B(n34691), .Z(n34696) );
  NANDN U35980 ( .A(n34694), .B(n34693), .Z(n34695) );
  AND U35981 ( .A(n34696), .B(n34695), .Z(n34731) );
  NANDN U35982 ( .A(n34698), .B(n34697), .Z(n34702) );
  NANDN U35983 ( .A(n34700), .B(n34699), .Z(n34701) );
  AND U35984 ( .A(n34702), .B(n34701), .Z(n34729) );
  NAND U35985 ( .A(n42143), .B(n34703), .Z(n34705) );
  XNOR U35986 ( .A(a[822]), .B(n4189), .Z(n34740) );
  NAND U35987 ( .A(n42144), .B(n34740), .Z(n34704) );
  AND U35988 ( .A(n34705), .B(n34704), .Z(n34755) );
  XOR U35989 ( .A(a[826]), .B(n42012), .Z(n34743) );
  XNOR U35990 ( .A(n34755), .B(n34754), .Z(n34757) );
  XOR U35991 ( .A(a[824]), .B(n42085), .Z(n34744) );
  AND U35992 ( .A(a[820]), .B(b[7]), .Z(n34748) );
  XNOR U35993 ( .A(n34749), .B(n34748), .Z(n34750) );
  AND U35994 ( .A(a[828]), .B(b[0]), .Z(n34708) );
  XNOR U35995 ( .A(n34708), .B(n4071), .Z(n34710) );
  NANDN U35996 ( .A(b[0]), .B(a[827]), .Z(n34709) );
  NAND U35997 ( .A(n34710), .B(n34709), .Z(n34751) );
  XNOR U35998 ( .A(n34750), .B(n34751), .Z(n34756) );
  XOR U35999 ( .A(n34757), .B(n34756), .Z(n34735) );
  NANDN U36000 ( .A(n34712), .B(n34711), .Z(n34716) );
  NANDN U36001 ( .A(n34714), .B(n34713), .Z(n34715) );
  AND U36002 ( .A(n34716), .B(n34715), .Z(n34734) );
  XNOR U36003 ( .A(n34735), .B(n34734), .Z(n34736) );
  NANDN U36004 ( .A(n34718), .B(n34717), .Z(n34722) );
  NAND U36005 ( .A(n34720), .B(n34719), .Z(n34721) );
  NAND U36006 ( .A(n34722), .B(n34721), .Z(n34737) );
  XNOR U36007 ( .A(n34736), .B(n34737), .Z(n34728) );
  XNOR U36008 ( .A(n34729), .B(n34728), .Z(n34730) );
  XNOR U36009 ( .A(n34731), .B(n34730), .Z(n34760) );
  XNOR U36010 ( .A(sreg[1844]), .B(n34760), .Z(n34762) );
  NANDN U36011 ( .A(sreg[1843]), .B(n34723), .Z(n34727) );
  NAND U36012 ( .A(n34725), .B(n34724), .Z(n34726) );
  NAND U36013 ( .A(n34727), .B(n34726), .Z(n34761) );
  XNOR U36014 ( .A(n34762), .B(n34761), .Z(c[1844]) );
  NANDN U36015 ( .A(n34729), .B(n34728), .Z(n34733) );
  NANDN U36016 ( .A(n34731), .B(n34730), .Z(n34732) );
  AND U36017 ( .A(n34733), .B(n34732), .Z(n34768) );
  NANDN U36018 ( .A(n34735), .B(n34734), .Z(n34739) );
  NANDN U36019 ( .A(n34737), .B(n34736), .Z(n34738) );
  AND U36020 ( .A(n34739), .B(n34738), .Z(n34766) );
  NAND U36021 ( .A(n42143), .B(n34740), .Z(n34742) );
  XNOR U36022 ( .A(a[823]), .B(n4189), .Z(n34777) );
  NAND U36023 ( .A(n42144), .B(n34777), .Z(n34741) );
  AND U36024 ( .A(n34742), .B(n34741), .Z(n34792) );
  XOR U36025 ( .A(a[827]), .B(n42012), .Z(n34780) );
  XNOR U36026 ( .A(n34792), .B(n34791), .Z(n34794) );
  XOR U36027 ( .A(a[825]), .B(n42085), .Z(n34781) );
  AND U36028 ( .A(a[821]), .B(b[7]), .Z(n34785) );
  XNOR U36029 ( .A(n34786), .B(n34785), .Z(n34787) );
  AND U36030 ( .A(a[829]), .B(b[0]), .Z(n34745) );
  XNOR U36031 ( .A(n34745), .B(n4071), .Z(n34747) );
  NANDN U36032 ( .A(b[0]), .B(a[828]), .Z(n34746) );
  NAND U36033 ( .A(n34747), .B(n34746), .Z(n34788) );
  XNOR U36034 ( .A(n34787), .B(n34788), .Z(n34793) );
  XOR U36035 ( .A(n34794), .B(n34793), .Z(n34772) );
  NANDN U36036 ( .A(n34749), .B(n34748), .Z(n34753) );
  NANDN U36037 ( .A(n34751), .B(n34750), .Z(n34752) );
  AND U36038 ( .A(n34753), .B(n34752), .Z(n34771) );
  XNOR U36039 ( .A(n34772), .B(n34771), .Z(n34773) );
  NANDN U36040 ( .A(n34755), .B(n34754), .Z(n34759) );
  NAND U36041 ( .A(n34757), .B(n34756), .Z(n34758) );
  NAND U36042 ( .A(n34759), .B(n34758), .Z(n34774) );
  XNOR U36043 ( .A(n34773), .B(n34774), .Z(n34765) );
  XNOR U36044 ( .A(n34766), .B(n34765), .Z(n34767) );
  XNOR U36045 ( .A(n34768), .B(n34767), .Z(n34797) );
  XNOR U36046 ( .A(sreg[1845]), .B(n34797), .Z(n34799) );
  NANDN U36047 ( .A(sreg[1844]), .B(n34760), .Z(n34764) );
  NAND U36048 ( .A(n34762), .B(n34761), .Z(n34763) );
  NAND U36049 ( .A(n34764), .B(n34763), .Z(n34798) );
  XNOR U36050 ( .A(n34799), .B(n34798), .Z(c[1845]) );
  NANDN U36051 ( .A(n34766), .B(n34765), .Z(n34770) );
  NANDN U36052 ( .A(n34768), .B(n34767), .Z(n34769) );
  AND U36053 ( .A(n34770), .B(n34769), .Z(n34805) );
  NANDN U36054 ( .A(n34772), .B(n34771), .Z(n34776) );
  NANDN U36055 ( .A(n34774), .B(n34773), .Z(n34775) );
  AND U36056 ( .A(n34776), .B(n34775), .Z(n34803) );
  NAND U36057 ( .A(n42143), .B(n34777), .Z(n34779) );
  XNOR U36058 ( .A(a[824]), .B(n4189), .Z(n34814) );
  NAND U36059 ( .A(n42144), .B(n34814), .Z(n34778) );
  AND U36060 ( .A(n34779), .B(n34778), .Z(n34829) );
  XOR U36061 ( .A(a[828]), .B(n42012), .Z(n34817) );
  XNOR U36062 ( .A(n34829), .B(n34828), .Z(n34831) );
  XOR U36063 ( .A(a[826]), .B(n42085), .Z(n34818) );
  AND U36064 ( .A(a[822]), .B(b[7]), .Z(n34822) );
  XNOR U36065 ( .A(n34823), .B(n34822), .Z(n34824) );
  AND U36066 ( .A(a[830]), .B(b[0]), .Z(n34782) );
  XNOR U36067 ( .A(n34782), .B(n4071), .Z(n34784) );
  NANDN U36068 ( .A(b[0]), .B(a[829]), .Z(n34783) );
  NAND U36069 ( .A(n34784), .B(n34783), .Z(n34825) );
  XNOR U36070 ( .A(n34824), .B(n34825), .Z(n34830) );
  XOR U36071 ( .A(n34831), .B(n34830), .Z(n34809) );
  NANDN U36072 ( .A(n34786), .B(n34785), .Z(n34790) );
  NANDN U36073 ( .A(n34788), .B(n34787), .Z(n34789) );
  AND U36074 ( .A(n34790), .B(n34789), .Z(n34808) );
  XNOR U36075 ( .A(n34809), .B(n34808), .Z(n34810) );
  NANDN U36076 ( .A(n34792), .B(n34791), .Z(n34796) );
  NAND U36077 ( .A(n34794), .B(n34793), .Z(n34795) );
  NAND U36078 ( .A(n34796), .B(n34795), .Z(n34811) );
  XNOR U36079 ( .A(n34810), .B(n34811), .Z(n34802) );
  XNOR U36080 ( .A(n34803), .B(n34802), .Z(n34804) );
  XNOR U36081 ( .A(n34805), .B(n34804), .Z(n34834) );
  XNOR U36082 ( .A(sreg[1846]), .B(n34834), .Z(n34836) );
  NANDN U36083 ( .A(sreg[1845]), .B(n34797), .Z(n34801) );
  NAND U36084 ( .A(n34799), .B(n34798), .Z(n34800) );
  NAND U36085 ( .A(n34801), .B(n34800), .Z(n34835) );
  XNOR U36086 ( .A(n34836), .B(n34835), .Z(c[1846]) );
  NANDN U36087 ( .A(n34803), .B(n34802), .Z(n34807) );
  NANDN U36088 ( .A(n34805), .B(n34804), .Z(n34806) );
  AND U36089 ( .A(n34807), .B(n34806), .Z(n34842) );
  NANDN U36090 ( .A(n34809), .B(n34808), .Z(n34813) );
  NANDN U36091 ( .A(n34811), .B(n34810), .Z(n34812) );
  AND U36092 ( .A(n34813), .B(n34812), .Z(n34840) );
  NAND U36093 ( .A(n42143), .B(n34814), .Z(n34816) );
  XNOR U36094 ( .A(a[825]), .B(n4189), .Z(n34851) );
  NAND U36095 ( .A(n42144), .B(n34851), .Z(n34815) );
  AND U36096 ( .A(n34816), .B(n34815), .Z(n34866) );
  XOR U36097 ( .A(a[829]), .B(n42012), .Z(n34854) );
  XNOR U36098 ( .A(n34866), .B(n34865), .Z(n34868) );
  XOR U36099 ( .A(a[827]), .B(n42085), .Z(n34855) );
  AND U36100 ( .A(a[823]), .B(b[7]), .Z(n34859) );
  XNOR U36101 ( .A(n34860), .B(n34859), .Z(n34861) );
  AND U36102 ( .A(a[831]), .B(b[0]), .Z(n34819) );
  XNOR U36103 ( .A(n34819), .B(n4071), .Z(n34821) );
  NANDN U36104 ( .A(b[0]), .B(a[830]), .Z(n34820) );
  NAND U36105 ( .A(n34821), .B(n34820), .Z(n34862) );
  XNOR U36106 ( .A(n34861), .B(n34862), .Z(n34867) );
  XOR U36107 ( .A(n34868), .B(n34867), .Z(n34846) );
  NANDN U36108 ( .A(n34823), .B(n34822), .Z(n34827) );
  NANDN U36109 ( .A(n34825), .B(n34824), .Z(n34826) );
  AND U36110 ( .A(n34827), .B(n34826), .Z(n34845) );
  XNOR U36111 ( .A(n34846), .B(n34845), .Z(n34847) );
  NANDN U36112 ( .A(n34829), .B(n34828), .Z(n34833) );
  NAND U36113 ( .A(n34831), .B(n34830), .Z(n34832) );
  NAND U36114 ( .A(n34833), .B(n34832), .Z(n34848) );
  XNOR U36115 ( .A(n34847), .B(n34848), .Z(n34839) );
  XNOR U36116 ( .A(n34840), .B(n34839), .Z(n34841) );
  XNOR U36117 ( .A(n34842), .B(n34841), .Z(n34871) );
  XNOR U36118 ( .A(sreg[1847]), .B(n34871), .Z(n34873) );
  NANDN U36119 ( .A(sreg[1846]), .B(n34834), .Z(n34838) );
  NAND U36120 ( .A(n34836), .B(n34835), .Z(n34837) );
  NAND U36121 ( .A(n34838), .B(n34837), .Z(n34872) );
  XNOR U36122 ( .A(n34873), .B(n34872), .Z(c[1847]) );
  NANDN U36123 ( .A(n34840), .B(n34839), .Z(n34844) );
  NANDN U36124 ( .A(n34842), .B(n34841), .Z(n34843) );
  AND U36125 ( .A(n34844), .B(n34843), .Z(n34879) );
  NANDN U36126 ( .A(n34846), .B(n34845), .Z(n34850) );
  NANDN U36127 ( .A(n34848), .B(n34847), .Z(n34849) );
  AND U36128 ( .A(n34850), .B(n34849), .Z(n34877) );
  NAND U36129 ( .A(n42143), .B(n34851), .Z(n34853) );
  XNOR U36130 ( .A(a[826]), .B(n4189), .Z(n34888) );
  NAND U36131 ( .A(n42144), .B(n34888), .Z(n34852) );
  AND U36132 ( .A(n34853), .B(n34852), .Z(n34903) );
  XOR U36133 ( .A(a[830]), .B(n42012), .Z(n34891) );
  XNOR U36134 ( .A(n34903), .B(n34902), .Z(n34905) );
  XOR U36135 ( .A(a[828]), .B(n42085), .Z(n34892) );
  AND U36136 ( .A(a[824]), .B(b[7]), .Z(n34896) );
  XNOR U36137 ( .A(n34897), .B(n34896), .Z(n34898) );
  AND U36138 ( .A(a[832]), .B(b[0]), .Z(n34856) );
  XNOR U36139 ( .A(n34856), .B(n4071), .Z(n34858) );
  NANDN U36140 ( .A(b[0]), .B(a[831]), .Z(n34857) );
  NAND U36141 ( .A(n34858), .B(n34857), .Z(n34899) );
  XNOR U36142 ( .A(n34898), .B(n34899), .Z(n34904) );
  XOR U36143 ( .A(n34905), .B(n34904), .Z(n34883) );
  NANDN U36144 ( .A(n34860), .B(n34859), .Z(n34864) );
  NANDN U36145 ( .A(n34862), .B(n34861), .Z(n34863) );
  AND U36146 ( .A(n34864), .B(n34863), .Z(n34882) );
  XNOR U36147 ( .A(n34883), .B(n34882), .Z(n34884) );
  NANDN U36148 ( .A(n34866), .B(n34865), .Z(n34870) );
  NAND U36149 ( .A(n34868), .B(n34867), .Z(n34869) );
  NAND U36150 ( .A(n34870), .B(n34869), .Z(n34885) );
  XNOR U36151 ( .A(n34884), .B(n34885), .Z(n34876) );
  XNOR U36152 ( .A(n34877), .B(n34876), .Z(n34878) );
  XNOR U36153 ( .A(n34879), .B(n34878), .Z(n34908) );
  XNOR U36154 ( .A(sreg[1848]), .B(n34908), .Z(n34910) );
  NANDN U36155 ( .A(sreg[1847]), .B(n34871), .Z(n34875) );
  NAND U36156 ( .A(n34873), .B(n34872), .Z(n34874) );
  NAND U36157 ( .A(n34875), .B(n34874), .Z(n34909) );
  XNOR U36158 ( .A(n34910), .B(n34909), .Z(c[1848]) );
  NANDN U36159 ( .A(n34877), .B(n34876), .Z(n34881) );
  NANDN U36160 ( .A(n34879), .B(n34878), .Z(n34880) );
  AND U36161 ( .A(n34881), .B(n34880), .Z(n34916) );
  NANDN U36162 ( .A(n34883), .B(n34882), .Z(n34887) );
  NANDN U36163 ( .A(n34885), .B(n34884), .Z(n34886) );
  AND U36164 ( .A(n34887), .B(n34886), .Z(n34914) );
  NAND U36165 ( .A(n42143), .B(n34888), .Z(n34890) );
  XNOR U36166 ( .A(a[827]), .B(n4190), .Z(n34925) );
  NAND U36167 ( .A(n42144), .B(n34925), .Z(n34889) );
  AND U36168 ( .A(n34890), .B(n34889), .Z(n34940) );
  XOR U36169 ( .A(a[831]), .B(n42012), .Z(n34928) );
  XNOR U36170 ( .A(n34940), .B(n34939), .Z(n34942) );
  XOR U36171 ( .A(a[829]), .B(n42085), .Z(n34929) );
  AND U36172 ( .A(a[825]), .B(b[7]), .Z(n34933) );
  XNOR U36173 ( .A(n34934), .B(n34933), .Z(n34935) );
  AND U36174 ( .A(a[833]), .B(b[0]), .Z(n34893) );
  XNOR U36175 ( .A(n34893), .B(n4071), .Z(n34895) );
  NANDN U36176 ( .A(b[0]), .B(a[832]), .Z(n34894) );
  NAND U36177 ( .A(n34895), .B(n34894), .Z(n34936) );
  XNOR U36178 ( .A(n34935), .B(n34936), .Z(n34941) );
  XOR U36179 ( .A(n34942), .B(n34941), .Z(n34920) );
  NANDN U36180 ( .A(n34897), .B(n34896), .Z(n34901) );
  NANDN U36181 ( .A(n34899), .B(n34898), .Z(n34900) );
  AND U36182 ( .A(n34901), .B(n34900), .Z(n34919) );
  XNOR U36183 ( .A(n34920), .B(n34919), .Z(n34921) );
  NANDN U36184 ( .A(n34903), .B(n34902), .Z(n34907) );
  NAND U36185 ( .A(n34905), .B(n34904), .Z(n34906) );
  NAND U36186 ( .A(n34907), .B(n34906), .Z(n34922) );
  XNOR U36187 ( .A(n34921), .B(n34922), .Z(n34913) );
  XNOR U36188 ( .A(n34914), .B(n34913), .Z(n34915) );
  XNOR U36189 ( .A(n34916), .B(n34915), .Z(n34945) );
  XNOR U36190 ( .A(sreg[1849]), .B(n34945), .Z(n34947) );
  NANDN U36191 ( .A(sreg[1848]), .B(n34908), .Z(n34912) );
  NAND U36192 ( .A(n34910), .B(n34909), .Z(n34911) );
  NAND U36193 ( .A(n34912), .B(n34911), .Z(n34946) );
  XNOR U36194 ( .A(n34947), .B(n34946), .Z(c[1849]) );
  NANDN U36195 ( .A(n34914), .B(n34913), .Z(n34918) );
  NANDN U36196 ( .A(n34916), .B(n34915), .Z(n34917) );
  AND U36197 ( .A(n34918), .B(n34917), .Z(n34953) );
  NANDN U36198 ( .A(n34920), .B(n34919), .Z(n34924) );
  NANDN U36199 ( .A(n34922), .B(n34921), .Z(n34923) );
  AND U36200 ( .A(n34924), .B(n34923), .Z(n34951) );
  NAND U36201 ( .A(n42143), .B(n34925), .Z(n34927) );
  XNOR U36202 ( .A(a[828]), .B(n4190), .Z(n34962) );
  NAND U36203 ( .A(n42144), .B(n34962), .Z(n34926) );
  AND U36204 ( .A(n34927), .B(n34926), .Z(n34977) );
  XOR U36205 ( .A(a[832]), .B(n42012), .Z(n34965) );
  XNOR U36206 ( .A(n34977), .B(n34976), .Z(n34979) );
  XOR U36207 ( .A(a[830]), .B(n42085), .Z(n34969) );
  AND U36208 ( .A(a[826]), .B(b[7]), .Z(n34970) );
  XNOR U36209 ( .A(n34971), .B(n34970), .Z(n34972) );
  AND U36210 ( .A(a[834]), .B(b[0]), .Z(n34930) );
  XNOR U36211 ( .A(n34930), .B(n4071), .Z(n34932) );
  NANDN U36212 ( .A(b[0]), .B(a[833]), .Z(n34931) );
  NAND U36213 ( .A(n34932), .B(n34931), .Z(n34973) );
  XNOR U36214 ( .A(n34972), .B(n34973), .Z(n34978) );
  XOR U36215 ( .A(n34979), .B(n34978), .Z(n34957) );
  NANDN U36216 ( .A(n34934), .B(n34933), .Z(n34938) );
  NANDN U36217 ( .A(n34936), .B(n34935), .Z(n34937) );
  AND U36218 ( .A(n34938), .B(n34937), .Z(n34956) );
  XNOR U36219 ( .A(n34957), .B(n34956), .Z(n34958) );
  NANDN U36220 ( .A(n34940), .B(n34939), .Z(n34944) );
  NAND U36221 ( .A(n34942), .B(n34941), .Z(n34943) );
  NAND U36222 ( .A(n34944), .B(n34943), .Z(n34959) );
  XNOR U36223 ( .A(n34958), .B(n34959), .Z(n34950) );
  XNOR U36224 ( .A(n34951), .B(n34950), .Z(n34952) );
  XNOR U36225 ( .A(n34953), .B(n34952), .Z(n34982) );
  XNOR U36226 ( .A(sreg[1850]), .B(n34982), .Z(n34984) );
  NANDN U36227 ( .A(sreg[1849]), .B(n34945), .Z(n34949) );
  NAND U36228 ( .A(n34947), .B(n34946), .Z(n34948) );
  NAND U36229 ( .A(n34949), .B(n34948), .Z(n34983) );
  XNOR U36230 ( .A(n34984), .B(n34983), .Z(c[1850]) );
  NANDN U36231 ( .A(n34951), .B(n34950), .Z(n34955) );
  NANDN U36232 ( .A(n34953), .B(n34952), .Z(n34954) );
  AND U36233 ( .A(n34955), .B(n34954), .Z(n34990) );
  NANDN U36234 ( .A(n34957), .B(n34956), .Z(n34961) );
  NANDN U36235 ( .A(n34959), .B(n34958), .Z(n34960) );
  AND U36236 ( .A(n34961), .B(n34960), .Z(n34988) );
  NAND U36237 ( .A(n42143), .B(n34962), .Z(n34964) );
  XNOR U36238 ( .A(a[829]), .B(n4190), .Z(n34999) );
  NAND U36239 ( .A(n42144), .B(n34999), .Z(n34963) );
  AND U36240 ( .A(n34964), .B(n34963), .Z(n35014) );
  XOR U36241 ( .A(a[833]), .B(n42012), .Z(n35002) );
  XNOR U36242 ( .A(n35014), .B(n35013), .Z(n35016) );
  AND U36243 ( .A(a[835]), .B(b[0]), .Z(n34966) );
  XNOR U36244 ( .A(n34966), .B(n4071), .Z(n34968) );
  NANDN U36245 ( .A(b[0]), .B(a[834]), .Z(n34967) );
  NAND U36246 ( .A(n34968), .B(n34967), .Z(n35010) );
  XOR U36247 ( .A(a[831]), .B(n42085), .Z(n35006) );
  AND U36248 ( .A(a[827]), .B(b[7]), .Z(n35007) );
  XNOR U36249 ( .A(n35008), .B(n35007), .Z(n35009) );
  XNOR U36250 ( .A(n35010), .B(n35009), .Z(n35015) );
  XOR U36251 ( .A(n35016), .B(n35015), .Z(n34994) );
  NANDN U36252 ( .A(n34971), .B(n34970), .Z(n34975) );
  NANDN U36253 ( .A(n34973), .B(n34972), .Z(n34974) );
  AND U36254 ( .A(n34975), .B(n34974), .Z(n34993) );
  XNOR U36255 ( .A(n34994), .B(n34993), .Z(n34995) );
  NANDN U36256 ( .A(n34977), .B(n34976), .Z(n34981) );
  NAND U36257 ( .A(n34979), .B(n34978), .Z(n34980) );
  NAND U36258 ( .A(n34981), .B(n34980), .Z(n34996) );
  XNOR U36259 ( .A(n34995), .B(n34996), .Z(n34987) );
  XNOR U36260 ( .A(n34988), .B(n34987), .Z(n34989) );
  XNOR U36261 ( .A(n34990), .B(n34989), .Z(n35019) );
  XNOR U36262 ( .A(sreg[1851]), .B(n35019), .Z(n35021) );
  NANDN U36263 ( .A(sreg[1850]), .B(n34982), .Z(n34986) );
  NAND U36264 ( .A(n34984), .B(n34983), .Z(n34985) );
  NAND U36265 ( .A(n34986), .B(n34985), .Z(n35020) );
  XNOR U36266 ( .A(n35021), .B(n35020), .Z(c[1851]) );
  NANDN U36267 ( .A(n34988), .B(n34987), .Z(n34992) );
  NANDN U36268 ( .A(n34990), .B(n34989), .Z(n34991) );
  AND U36269 ( .A(n34992), .B(n34991), .Z(n35027) );
  NANDN U36270 ( .A(n34994), .B(n34993), .Z(n34998) );
  NANDN U36271 ( .A(n34996), .B(n34995), .Z(n34997) );
  AND U36272 ( .A(n34998), .B(n34997), .Z(n35025) );
  NAND U36273 ( .A(n42143), .B(n34999), .Z(n35001) );
  XNOR U36274 ( .A(a[830]), .B(n4190), .Z(n35036) );
  NAND U36275 ( .A(n42144), .B(n35036), .Z(n35000) );
  AND U36276 ( .A(n35001), .B(n35000), .Z(n35051) );
  XOR U36277 ( .A(a[834]), .B(n42012), .Z(n35039) );
  XNOR U36278 ( .A(n35051), .B(n35050), .Z(n35053) );
  AND U36279 ( .A(a[836]), .B(b[0]), .Z(n35003) );
  XNOR U36280 ( .A(n35003), .B(n4071), .Z(n35005) );
  NANDN U36281 ( .A(b[0]), .B(a[835]), .Z(n35004) );
  NAND U36282 ( .A(n35005), .B(n35004), .Z(n35047) );
  XOR U36283 ( .A(a[832]), .B(n42085), .Z(n35043) );
  AND U36284 ( .A(a[828]), .B(b[7]), .Z(n35044) );
  XNOR U36285 ( .A(n35045), .B(n35044), .Z(n35046) );
  XNOR U36286 ( .A(n35047), .B(n35046), .Z(n35052) );
  XOR U36287 ( .A(n35053), .B(n35052), .Z(n35031) );
  NANDN U36288 ( .A(n35008), .B(n35007), .Z(n35012) );
  NANDN U36289 ( .A(n35010), .B(n35009), .Z(n35011) );
  AND U36290 ( .A(n35012), .B(n35011), .Z(n35030) );
  XNOR U36291 ( .A(n35031), .B(n35030), .Z(n35032) );
  NANDN U36292 ( .A(n35014), .B(n35013), .Z(n35018) );
  NAND U36293 ( .A(n35016), .B(n35015), .Z(n35017) );
  NAND U36294 ( .A(n35018), .B(n35017), .Z(n35033) );
  XNOR U36295 ( .A(n35032), .B(n35033), .Z(n35024) );
  XNOR U36296 ( .A(n35025), .B(n35024), .Z(n35026) );
  XNOR U36297 ( .A(n35027), .B(n35026), .Z(n35056) );
  XNOR U36298 ( .A(sreg[1852]), .B(n35056), .Z(n35058) );
  NANDN U36299 ( .A(sreg[1851]), .B(n35019), .Z(n35023) );
  NAND U36300 ( .A(n35021), .B(n35020), .Z(n35022) );
  NAND U36301 ( .A(n35023), .B(n35022), .Z(n35057) );
  XNOR U36302 ( .A(n35058), .B(n35057), .Z(c[1852]) );
  NANDN U36303 ( .A(n35025), .B(n35024), .Z(n35029) );
  NANDN U36304 ( .A(n35027), .B(n35026), .Z(n35028) );
  AND U36305 ( .A(n35029), .B(n35028), .Z(n35064) );
  NANDN U36306 ( .A(n35031), .B(n35030), .Z(n35035) );
  NANDN U36307 ( .A(n35033), .B(n35032), .Z(n35034) );
  AND U36308 ( .A(n35035), .B(n35034), .Z(n35062) );
  NAND U36309 ( .A(n42143), .B(n35036), .Z(n35038) );
  XNOR U36310 ( .A(a[831]), .B(n4190), .Z(n35073) );
  NAND U36311 ( .A(n42144), .B(n35073), .Z(n35037) );
  AND U36312 ( .A(n35038), .B(n35037), .Z(n35088) );
  XOR U36313 ( .A(a[835]), .B(n42012), .Z(n35076) );
  XNOR U36314 ( .A(n35088), .B(n35087), .Z(n35090) );
  AND U36315 ( .A(a[837]), .B(b[0]), .Z(n35040) );
  XNOR U36316 ( .A(n35040), .B(n4071), .Z(n35042) );
  NANDN U36317 ( .A(b[0]), .B(a[836]), .Z(n35041) );
  NAND U36318 ( .A(n35042), .B(n35041), .Z(n35084) );
  XOR U36319 ( .A(a[833]), .B(n42085), .Z(n35077) );
  AND U36320 ( .A(a[829]), .B(b[7]), .Z(n35081) );
  XNOR U36321 ( .A(n35082), .B(n35081), .Z(n35083) );
  XNOR U36322 ( .A(n35084), .B(n35083), .Z(n35089) );
  XOR U36323 ( .A(n35090), .B(n35089), .Z(n35068) );
  NANDN U36324 ( .A(n35045), .B(n35044), .Z(n35049) );
  NANDN U36325 ( .A(n35047), .B(n35046), .Z(n35048) );
  AND U36326 ( .A(n35049), .B(n35048), .Z(n35067) );
  XNOR U36327 ( .A(n35068), .B(n35067), .Z(n35069) );
  NANDN U36328 ( .A(n35051), .B(n35050), .Z(n35055) );
  NAND U36329 ( .A(n35053), .B(n35052), .Z(n35054) );
  NAND U36330 ( .A(n35055), .B(n35054), .Z(n35070) );
  XNOR U36331 ( .A(n35069), .B(n35070), .Z(n35061) );
  XNOR U36332 ( .A(n35062), .B(n35061), .Z(n35063) );
  XNOR U36333 ( .A(n35064), .B(n35063), .Z(n35093) );
  XNOR U36334 ( .A(sreg[1853]), .B(n35093), .Z(n35095) );
  NANDN U36335 ( .A(sreg[1852]), .B(n35056), .Z(n35060) );
  NAND U36336 ( .A(n35058), .B(n35057), .Z(n35059) );
  NAND U36337 ( .A(n35060), .B(n35059), .Z(n35094) );
  XNOR U36338 ( .A(n35095), .B(n35094), .Z(c[1853]) );
  NANDN U36339 ( .A(n35062), .B(n35061), .Z(n35066) );
  NANDN U36340 ( .A(n35064), .B(n35063), .Z(n35065) );
  AND U36341 ( .A(n35066), .B(n35065), .Z(n35101) );
  NANDN U36342 ( .A(n35068), .B(n35067), .Z(n35072) );
  NANDN U36343 ( .A(n35070), .B(n35069), .Z(n35071) );
  AND U36344 ( .A(n35072), .B(n35071), .Z(n35099) );
  NAND U36345 ( .A(n42143), .B(n35073), .Z(n35075) );
  XNOR U36346 ( .A(a[832]), .B(n4190), .Z(n35110) );
  NAND U36347 ( .A(n42144), .B(n35110), .Z(n35074) );
  AND U36348 ( .A(n35075), .B(n35074), .Z(n35125) );
  XOR U36349 ( .A(a[836]), .B(n42012), .Z(n35113) );
  XNOR U36350 ( .A(n35125), .B(n35124), .Z(n35127) );
  XOR U36351 ( .A(a[834]), .B(n42085), .Z(n35114) );
  AND U36352 ( .A(a[830]), .B(b[7]), .Z(n35118) );
  XNOR U36353 ( .A(n35119), .B(n35118), .Z(n35120) );
  AND U36354 ( .A(a[838]), .B(b[0]), .Z(n35078) );
  XNOR U36355 ( .A(n35078), .B(n4071), .Z(n35080) );
  NANDN U36356 ( .A(b[0]), .B(a[837]), .Z(n35079) );
  NAND U36357 ( .A(n35080), .B(n35079), .Z(n35121) );
  XNOR U36358 ( .A(n35120), .B(n35121), .Z(n35126) );
  XOR U36359 ( .A(n35127), .B(n35126), .Z(n35105) );
  NANDN U36360 ( .A(n35082), .B(n35081), .Z(n35086) );
  NANDN U36361 ( .A(n35084), .B(n35083), .Z(n35085) );
  AND U36362 ( .A(n35086), .B(n35085), .Z(n35104) );
  XNOR U36363 ( .A(n35105), .B(n35104), .Z(n35106) );
  NANDN U36364 ( .A(n35088), .B(n35087), .Z(n35092) );
  NAND U36365 ( .A(n35090), .B(n35089), .Z(n35091) );
  NAND U36366 ( .A(n35092), .B(n35091), .Z(n35107) );
  XNOR U36367 ( .A(n35106), .B(n35107), .Z(n35098) );
  XNOR U36368 ( .A(n35099), .B(n35098), .Z(n35100) );
  XNOR U36369 ( .A(n35101), .B(n35100), .Z(n35130) );
  XNOR U36370 ( .A(sreg[1854]), .B(n35130), .Z(n35132) );
  NANDN U36371 ( .A(sreg[1853]), .B(n35093), .Z(n35097) );
  NAND U36372 ( .A(n35095), .B(n35094), .Z(n35096) );
  NAND U36373 ( .A(n35097), .B(n35096), .Z(n35131) );
  XNOR U36374 ( .A(n35132), .B(n35131), .Z(c[1854]) );
  NANDN U36375 ( .A(n35099), .B(n35098), .Z(n35103) );
  NANDN U36376 ( .A(n35101), .B(n35100), .Z(n35102) );
  AND U36377 ( .A(n35103), .B(n35102), .Z(n35138) );
  NANDN U36378 ( .A(n35105), .B(n35104), .Z(n35109) );
  NANDN U36379 ( .A(n35107), .B(n35106), .Z(n35108) );
  AND U36380 ( .A(n35109), .B(n35108), .Z(n35136) );
  NAND U36381 ( .A(n42143), .B(n35110), .Z(n35112) );
  XNOR U36382 ( .A(a[833]), .B(n4190), .Z(n35147) );
  NAND U36383 ( .A(n42144), .B(n35147), .Z(n35111) );
  AND U36384 ( .A(n35112), .B(n35111), .Z(n35162) );
  XOR U36385 ( .A(a[837]), .B(n42012), .Z(n35150) );
  XNOR U36386 ( .A(n35162), .B(n35161), .Z(n35164) );
  XOR U36387 ( .A(a[835]), .B(n42085), .Z(n35154) );
  AND U36388 ( .A(a[831]), .B(b[7]), .Z(n35155) );
  XNOR U36389 ( .A(n35156), .B(n35155), .Z(n35157) );
  AND U36390 ( .A(a[839]), .B(b[0]), .Z(n35115) );
  XNOR U36391 ( .A(n35115), .B(n4071), .Z(n35117) );
  NANDN U36392 ( .A(b[0]), .B(a[838]), .Z(n35116) );
  NAND U36393 ( .A(n35117), .B(n35116), .Z(n35158) );
  XNOR U36394 ( .A(n35157), .B(n35158), .Z(n35163) );
  XOR U36395 ( .A(n35164), .B(n35163), .Z(n35142) );
  NANDN U36396 ( .A(n35119), .B(n35118), .Z(n35123) );
  NANDN U36397 ( .A(n35121), .B(n35120), .Z(n35122) );
  AND U36398 ( .A(n35123), .B(n35122), .Z(n35141) );
  XNOR U36399 ( .A(n35142), .B(n35141), .Z(n35143) );
  NANDN U36400 ( .A(n35125), .B(n35124), .Z(n35129) );
  NAND U36401 ( .A(n35127), .B(n35126), .Z(n35128) );
  NAND U36402 ( .A(n35129), .B(n35128), .Z(n35144) );
  XNOR U36403 ( .A(n35143), .B(n35144), .Z(n35135) );
  XNOR U36404 ( .A(n35136), .B(n35135), .Z(n35137) );
  XNOR U36405 ( .A(n35138), .B(n35137), .Z(n35167) );
  XNOR U36406 ( .A(sreg[1855]), .B(n35167), .Z(n35169) );
  NANDN U36407 ( .A(sreg[1854]), .B(n35130), .Z(n35134) );
  NAND U36408 ( .A(n35132), .B(n35131), .Z(n35133) );
  NAND U36409 ( .A(n35134), .B(n35133), .Z(n35168) );
  XNOR U36410 ( .A(n35169), .B(n35168), .Z(c[1855]) );
  NANDN U36411 ( .A(n35136), .B(n35135), .Z(n35140) );
  NANDN U36412 ( .A(n35138), .B(n35137), .Z(n35139) );
  AND U36413 ( .A(n35140), .B(n35139), .Z(n35175) );
  NANDN U36414 ( .A(n35142), .B(n35141), .Z(n35146) );
  NANDN U36415 ( .A(n35144), .B(n35143), .Z(n35145) );
  AND U36416 ( .A(n35146), .B(n35145), .Z(n35173) );
  NAND U36417 ( .A(n42143), .B(n35147), .Z(n35149) );
  XNOR U36418 ( .A(a[834]), .B(n4191), .Z(n35184) );
  NAND U36419 ( .A(n42144), .B(n35184), .Z(n35148) );
  AND U36420 ( .A(n35149), .B(n35148), .Z(n35199) );
  XOR U36421 ( .A(a[838]), .B(n42012), .Z(n35187) );
  XNOR U36422 ( .A(n35199), .B(n35198), .Z(n35201) );
  AND U36423 ( .A(a[840]), .B(b[0]), .Z(n35151) );
  XNOR U36424 ( .A(n35151), .B(n4071), .Z(n35153) );
  NANDN U36425 ( .A(b[0]), .B(a[839]), .Z(n35152) );
  NAND U36426 ( .A(n35153), .B(n35152), .Z(n35195) );
  XOR U36427 ( .A(a[836]), .B(n42085), .Z(n35191) );
  AND U36428 ( .A(a[832]), .B(b[7]), .Z(n35192) );
  XNOR U36429 ( .A(n35193), .B(n35192), .Z(n35194) );
  XNOR U36430 ( .A(n35195), .B(n35194), .Z(n35200) );
  XOR U36431 ( .A(n35201), .B(n35200), .Z(n35179) );
  NANDN U36432 ( .A(n35156), .B(n35155), .Z(n35160) );
  NANDN U36433 ( .A(n35158), .B(n35157), .Z(n35159) );
  AND U36434 ( .A(n35160), .B(n35159), .Z(n35178) );
  XNOR U36435 ( .A(n35179), .B(n35178), .Z(n35180) );
  NANDN U36436 ( .A(n35162), .B(n35161), .Z(n35166) );
  NAND U36437 ( .A(n35164), .B(n35163), .Z(n35165) );
  NAND U36438 ( .A(n35166), .B(n35165), .Z(n35181) );
  XNOR U36439 ( .A(n35180), .B(n35181), .Z(n35172) );
  XNOR U36440 ( .A(n35173), .B(n35172), .Z(n35174) );
  XNOR U36441 ( .A(n35175), .B(n35174), .Z(n35204) );
  XNOR U36442 ( .A(sreg[1856]), .B(n35204), .Z(n35206) );
  NANDN U36443 ( .A(sreg[1855]), .B(n35167), .Z(n35171) );
  NAND U36444 ( .A(n35169), .B(n35168), .Z(n35170) );
  NAND U36445 ( .A(n35171), .B(n35170), .Z(n35205) );
  XNOR U36446 ( .A(n35206), .B(n35205), .Z(c[1856]) );
  NANDN U36447 ( .A(n35173), .B(n35172), .Z(n35177) );
  NANDN U36448 ( .A(n35175), .B(n35174), .Z(n35176) );
  AND U36449 ( .A(n35177), .B(n35176), .Z(n35212) );
  NANDN U36450 ( .A(n35179), .B(n35178), .Z(n35183) );
  NANDN U36451 ( .A(n35181), .B(n35180), .Z(n35182) );
  AND U36452 ( .A(n35183), .B(n35182), .Z(n35210) );
  NAND U36453 ( .A(n42143), .B(n35184), .Z(n35186) );
  XNOR U36454 ( .A(a[835]), .B(n4191), .Z(n35221) );
  NAND U36455 ( .A(n42144), .B(n35221), .Z(n35185) );
  AND U36456 ( .A(n35186), .B(n35185), .Z(n35236) );
  XOR U36457 ( .A(a[839]), .B(n42012), .Z(n35224) );
  XNOR U36458 ( .A(n35236), .B(n35235), .Z(n35238) );
  AND U36459 ( .A(a[841]), .B(b[0]), .Z(n35188) );
  XNOR U36460 ( .A(n35188), .B(n4071), .Z(n35190) );
  NANDN U36461 ( .A(b[0]), .B(a[840]), .Z(n35189) );
  NAND U36462 ( .A(n35190), .B(n35189), .Z(n35232) );
  XOR U36463 ( .A(a[837]), .B(n42085), .Z(n35228) );
  AND U36464 ( .A(a[833]), .B(b[7]), .Z(n35229) );
  XNOR U36465 ( .A(n35230), .B(n35229), .Z(n35231) );
  XNOR U36466 ( .A(n35232), .B(n35231), .Z(n35237) );
  XOR U36467 ( .A(n35238), .B(n35237), .Z(n35216) );
  NANDN U36468 ( .A(n35193), .B(n35192), .Z(n35197) );
  NANDN U36469 ( .A(n35195), .B(n35194), .Z(n35196) );
  AND U36470 ( .A(n35197), .B(n35196), .Z(n35215) );
  XNOR U36471 ( .A(n35216), .B(n35215), .Z(n35217) );
  NANDN U36472 ( .A(n35199), .B(n35198), .Z(n35203) );
  NAND U36473 ( .A(n35201), .B(n35200), .Z(n35202) );
  NAND U36474 ( .A(n35203), .B(n35202), .Z(n35218) );
  XNOR U36475 ( .A(n35217), .B(n35218), .Z(n35209) );
  XNOR U36476 ( .A(n35210), .B(n35209), .Z(n35211) );
  XNOR U36477 ( .A(n35212), .B(n35211), .Z(n35241) );
  XNOR U36478 ( .A(sreg[1857]), .B(n35241), .Z(n35243) );
  NANDN U36479 ( .A(sreg[1856]), .B(n35204), .Z(n35208) );
  NAND U36480 ( .A(n35206), .B(n35205), .Z(n35207) );
  NAND U36481 ( .A(n35208), .B(n35207), .Z(n35242) );
  XNOR U36482 ( .A(n35243), .B(n35242), .Z(c[1857]) );
  NANDN U36483 ( .A(n35210), .B(n35209), .Z(n35214) );
  NANDN U36484 ( .A(n35212), .B(n35211), .Z(n35213) );
  AND U36485 ( .A(n35214), .B(n35213), .Z(n35249) );
  NANDN U36486 ( .A(n35216), .B(n35215), .Z(n35220) );
  NANDN U36487 ( .A(n35218), .B(n35217), .Z(n35219) );
  AND U36488 ( .A(n35220), .B(n35219), .Z(n35247) );
  NAND U36489 ( .A(n42143), .B(n35221), .Z(n35223) );
  XNOR U36490 ( .A(a[836]), .B(n4191), .Z(n35258) );
  NAND U36491 ( .A(n42144), .B(n35258), .Z(n35222) );
  AND U36492 ( .A(n35223), .B(n35222), .Z(n35273) );
  XOR U36493 ( .A(a[840]), .B(n42012), .Z(n35261) );
  XNOR U36494 ( .A(n35273), .B(n35272), .Z(n35275) );
  AND U36495 ( .A(a[842]), .B(b[0]), .Z(n35225) );
  XNOR U36496 ( .A(n35225), .B(n4071), .Z(n35227) );
  NANDN U36497 ( .A(b[0]), .B(a[841]), .Z(n35226) );
  NAND U36498 ( .A(n35227), .B(n35226), .Z(n35269) );
  XOR U36499 ( .A(a[838]), .B(n42085), .Z(n35265) );
  AND U36500 ( .A(a[834]), .B(b[7]), .Z(n35266) );
  XNOR U36501 ( .A(n35267), .B(n35266), .Z(n35268) );
  XNOR U36502 ( .A(n35269), .B(n35268), .Z(n35274) );
  XOR U36503 ( .A(n35275), .B(n35274), .Z(n35253) );
  NANDN U36504 ( .A(n35230), .B(n35229), .Z(n35234) );
  NANDN U36505 ( .A(n35232), .B(n35231), .Z(n35233) );
  AND U36506 ( .A(n35234), .B(n35233), .Z(n35252) );
  XNOR U36507 ( .A(n35253), .B(n35252), .Z(n35254) );
  NANDN U36508 ( .A(n35236), .B(n35235), .Z(n35240) );
  NAND U36509 ( .A(n35238), .B(n35237), .Z(n35239) );
  NAND U36510 ( .A(n35240), .B(n35239), .Z(n35255) );
  XNOR U36511 ( .A(n35254), .B(n35255), .Z(n35246) );
  XNOR U36512 ( .A(n35247), .B(n35246), .Z(n35248) );
  XNOR U36513 ( .A(n35249), .B(n35248), .Z(n35278) );
  XNOR U36514 ( .A(sreg[1858]), .B(n35278), .Z(n35280) );
  NANDN U36515 ( .A(sreg[1857]), .B(n35241), .Z(n35245) );
  NAND U36516 ( .A(n35243), .B(n35242), .Z(n35244) );
  NAND U36517 ( .A(n35245), .B(n35244), .Z(n35279) );
  XNOR U36518 ( .A(n35280), .B(n35279), .Z(c[1858]) );
  NANDN U36519 ( .A(n35247), .B(n35246), .Z(n35251) );
  NANDN U36520 ( .A(n35249), .B(n35248), .Z(n35250) );
  AND U36521 ( .A(n35251), .B(n35250), .Z(n35286) );
  NANDN U36522 ( .A(n35253), .B(n35252), .Z(n35257) );
  NANDN U36523 ( .A(n35255), .B(n35254), .Z(n35256) );
  AND U36524 ( .A(n35257), .B(n35256), .Z(n35284) );
  NAND U36525 ( .A(n42143), .B(n35258), .Z(n35260) );
  XNOR U36526 ( .A(a[837]), .B(n4191), .Z(n35295) );
  NAND U36527 ( .A(n42144), .B(n35295), .Z(n35259) );
  AND U36528 ( .A(n35260), .B(n35259), .Z(n35310) );
  XOR U36529 ( .A(a[841]), .B(n42012), .Z(n35298) );
  XNOR U36530 ( .A(n35310), .B(n35309), .Z(n35312) );
  AND U36531 ( .A(a[843]), .B(b[0]), .Z(n35262) );
  XNOR U36532 ( .A(n35262), .B(n4071), .Z(n35264) );
  NANDN U36533 ( .A(b[0]), .B(a[842]), .Z(n35263) );
  NAND U36534 ( .A(n35264), .B(n35263), .Z(n35306) );
  XOR U36535 ( .A(a[839]), .B(n42085), .Z(n35299) );
  AND U36536 ( .A(a[835]), .B(b[7]), .Z(n35303) );
  XNOR U36537 ( .A(n35304), .B(n35303), .Z(n35305) );
  XNOR U36538 ( .A(n35306), .B(n35305), .Z(n35311) );
  XOR U36539 ( .A(n35312), .B(n35311), .Z(n35290) );
  NANDN U36540 ( .A(n35267), .B(n35266), .Z(n35271) );
  NANDN U36541 ( .A(n35269), .B(n35268), .Z(n35270) );
  AND U36542 ( .A(n35271), .B(n35270), .Z(n35289) );
  XNOR U36543 ( .A(n35290), .B(n35289), .Z(n35291) );
  NANDN U36544 ( .A(n35273), .B(n35272), .Z(n35277) );
  NAND U36545 ( .A(n35275), .B(n35274), .Z(n35276) );
  NAND U36546 ( .A(n35277), .B(n35276), .Z(n35292) );
  XNOR U36547 ( .A(n35291), .B(n35292), .Z(n35283) );
  XNOR U36548 ( .A(n35284), .B(n35283), .Z(n35285) );
  XNOR U36549 ( .A(n35286), .B(n35285), .Z(n35315) );
  XNOR U36550 ( .A(sreg[1859]), .B(n35315), .Z(n35317) );
  NANDN U36551 ( .A(sreg[1858]), .B(n35278), .Z(n35282) );
  NAND U36552 ( .A(n35280), .B(n35279), .Z(n35281) );
  NAND U36553 ( .A(n35282), .B(n35281), .Z(n35316) );
  XNOR U36554 ( .A(n35317), .B(n35316), .Z(c[1859]) );
  NANDN U36555 ( .A(n35284), .B(n35283), .Z(n35288) );
  NANDN U36556 ( .A(n35286), .B(n35285), .Z(n35287) );
  AND U36557 ( .A(n35288), .B(n35287), .Z(n35323) );
  NANDN U36558 ( .A(n35290), .B(n35289), .Z(n35294) );
  NANDN U36559 ( .A(n35292), .B(n35291), .Z(n35293) );
  AND U36560 ( .A(n35294), .B(n35293), .Z(n35321) );
  NAND U36561 ( .A(n42143), .B(n35295), .Z(n35297) );
  XNOR U36562 ( .A(a[838]), .B(n4191), .Z(n35332) );
  NAND U36563 ( .A(n42144), .B(n35332), .Z(n35296) );
  AND U36564 ( .A(n35297), .B(n35296), .Z(n35347) );
  XOR U36565 ( .A(a[842]), .B(n42012), .Z(n35335) );
  XNOR U36566 ( .A(n35347), .B(n35346), .Z(n35349) );
  XOR U36567 ( .A(a[840]), .B(n42085), .Z(n35336) );
  AND U36568 ( .A(a[836]), .B(b[7]), .Z(n35340) );
  XNOR U36569 ( .A(n35341), .B(n35340), .Z(n35342) );
  AND U36570 ( .A(a[844]), .B(b[0]), .Z(n35300) );
  XNOR U36571 ( .A(n35300), .B(n4071), .Z(n35302) );
  NANDN U36572 ( .A(b[0]), .B(a[843]), .Z(n35301) );
  NAND U36573 ( .A(n35302), .B(n35301), .Z(n35343) );
  XNOR U36574 ( .A(n35342), .B(n35343), .Z(n35348) );
  XOR U36575 ( .A(n35349), .B(n35348), .Z(n35327) );
  NANDN U36576 ( .A(n35304), .B(n35303), .Z(n35308) );
  NANDN U36577 ( .A(n35306), .B(n35305), .Z(n35307) );
  AND U36578 ( .A(n35308), .B(n35307), .Z(n35326) );
  XNOR U36579 ( .A(n35327), .B(n35326), .Z(n35328) );
  NANDN U36580 ( .A(n35310), .B(n35309), .Z(n35314) );
  NAND U36581 ( .A(n35312), .B(n35311), .Z(n35313) );
  NAND U36582 ( .A(n35314), .B(n35313), .Z(n35329) );
  XNOR U36583 ( .A(n35328), .B(n35329), .Z(n35320) );
  XNOR U36584 ( .A(n35321), .B(n35320), .Z(n35322) );
  XNOR U36585 ( .A(n35323), .B(n35322), .Z(n35352) );
  XNOR U36586 ( .A(sreg[1860]), .B(n35352), .Z(n35354) );
  NANDN U36587 ( .A(sreg[1859]), .B(n35315), .Z(n35319) );
  NAND U36588 ( .A(n35317), .B(n35316), .Z(n35318) );
  NAND U36589 ( .A(n35319), .B(n35318), .Z(n35353) );
  XNOR U36590 ( .A(n35354), .B(n35353), .Z(c[1860]) );
  NANDN U36591 ( .A(n35321), .B(n35320), .Z(n35325) );
  NANDN U36592 ( .A(n35323), .B(n35322), .Z(n35324) );
  AND U36593 ( .A(n35325), .B(n35324), .Z(n35360) );
  NANDN U36594 ( .A(n35327), .B(n35326), .Z(n35331) );
  NANDN U36595 ( .A(n35329), .B(n35328), .Z(n35330) );
  AND U36596 ( .A(n35331), .B(n35330), .Z(n35358) );
  NAND U36597 ( .A(n42143), .B(n35332), .Z(n35334) );
  XNOR U36598 ( .A(a[839]), .B(n4191), .Z(n35369) );
  NAND U36599 ( .A(n42144), .B(n35369), .Z(n35333) );
  AND U36600 ( .A(n35334), .B(n35333), .Z(n35384) );
  XOR U36601 ( .A(a[843]), .B(n42012), .Z(n35372) );
  XNOR U36602 ( .A(n35384), .B(n35383), .Z(n35386) );
  XOR U36603 ( .A(a[841]), .B(n42085), .Z(n35373) );
  AND U36604 ( .A(a[837]), .B(b[7]), .Z(n35377) );
  XNOR U36605 ( .A(n35378), .B(n35377), .Z(n35379) );
  AND U36606 ( .A(a[845]), .B(b[0]), .Z(n35337) );
  XNOR U36607 ( .A(n35337), .B(n4071), .Z(n35339) );
  NANDN U36608 ( .A(b[0]), .B(a[844]), .Z(n35338) );
  NAND U36609 ( .A(n35339), .B(n35338), .Z(n35380) );
  XNOR U36610 ( .A(n35379), .B(n35380), .Z(n35385) );
  XOR U36611 ( .A(n35386), .B(n35385), .Z(n35364) );
  NANDN U36612 ( .A(n35341), .B(n35340), .Z(n35345) );
  NANDN U36613 ( .A(n35343), .B(n35342), .Z(n35344) );
  AND U36614 ( .A(n35345), .B(n35344), .Z(n35363) );
  XNOR U36615 ( .A(n35364), .B(n35363), .Z(n35365) );
  NANDN U36616 ( .A(n35347), .B(n35346), .Z(n35351) );
  NAND U36617 ( .A(n35349), .B(n35348), .Z(n35350) );
  NAND U36618 ( .A(n35351), .B(n35350), .Z(n35366) );
  XNOR U36619 ( .A(n35365), .B(n35366), .Z(n35357) );
  XNOR U36620 ( .A(n35358), .B(n35357), .Z(n35359) );
  XNOR U36621 ( .A(n35360), .B(n35359), .Z(n35389) );
  XNOR U36622 ( .A(sreg[1861]), .B(n35389), .Z(n35391) );
  NANDN U36623 ( .A(sreg[1860]), .B(n35352), .Z(n35356) );
  NAND U36624 ( .A(n35354), .B(n35353), .Z(n35355) );
  NAND U36625 ( .A(n35356), .B(n35355), .Z(n35390) );
  XNOR U36626 ( .A(n35391), .B(n35390), .Z(c[1861]) );
  NANDN U36627 ( .A(n35358), .B(n35357), .Z(n35362) );
  NANDN U36628 ( .A(n35360), .B(n35359), .Z(n35361) );
  AND U36629 ( .A(n35362), .B(n35361), .Z(n35397) );
  NANDN U36630 ( .A(n35364), .B(n35363), .Z(n35368) );
  NANDN U36631 ( .A(n35366), .B(n35365), .Z(n35367) );
  AND U36632 ( .A(n35368), .B(n35367), .Z(n35395) );
  NAND U36633 ( .A(n42143), .B(n35369), .Z(n35371) );
  XNOR U36634 ( .A(a[840]), .B(n4191), .Z(n35406) );
  NAND U36635 ( .A(n42144), .B(n35406), .Z(n35370) );
  AND U36636 ( .A(n35371), .B(n35370), .Z(n35421) );
  XOR U36637 ( .A(a[844]), .B(n42012), .Z(n35409) );
  XNOR U36638 ( .A(n35421), .B(n35420), .Z(n35423) );
  XOR U36639 ( .A(a[842]), .B(n42085), .Z(n35410) );
  AND U36640 ( .A(a[838]), .B(b[7]), .Z(n35414) );
  XNOR U36641 ( .A(n35415), .B(n35414), .Z(n35416) );
  AND U36642 ( .A(a[846]), .B(b[0]), .Z(n35374) );
  XNOR U36643 ( .A(n35374), .B(n4071), .Z(n35376) );
  NANDN U36644 ( .A(b[0]), .B(a[845]), .Z(n35375) );
  NAND U36645 ( .A(n35376), .B(n35375), .Z(n35417) );
  XNOR U36646 ( .A(n35416), .B(n35417), .Z(n35422) );
  XOR U36647 ( .A(n35423), .B(n35422), .Z(n35401) );
  NANDN U36648 ( .A(n35378), .B(n35377), .Z(n35382) );
  NANDN U36649 ( .A(n35380), .B(n35379), .Z(n35381) );
  AND U36650 ( .A(n35382), .B(n35381), .Z(n35400) );
  XNOR U36651 ( .A(n35401), .B(n35400), .Z(n35402) );
  NANDN U36652 ( .A(n35384), .B(n35383), .Z(n35388) );
  NAND U36653 ( .A(n35386), .B(n35385), .Z(n35387) );
  NAND U36654 ( .A(n35388), .B(n35387), .Z(n35403) );
  XNOR U36655 ( .A(n35402), .B(n35403), .Z(n35394) );
  XNOR U36656 ( .A(n35395), .B(n35394), .Z(n35396) );
  XNOR U36657 ( .A(n35397), .B(n35396), .Z(n35426) );
  XNOR U36658 ( .A(sreg[1862]), .B(n35426), .Z(n35428) );
  NANDN U36659 ( .A(sreg[1861]), .B(n35389), .Z(n35393) );
  NAND U36660 ( .A(n35391), .B(n35390), .Z(n35392) );
  NAND U36661 ( .A(n35393), .B(n35392), .Z(n35427) );
  XNOR U36662 ( .A(n35428), .B(n35427), .Z(c[1862]) );
  NANDN U36663 ( .A(n35395), .B(n35394), .Z(n35399) );
  NANDN U36664 ( .A(n35397), .B(n35396), .Z(n35398) );
  AND U36665 ( .A(n35399), .B(n35398), .Z(n35434) );
  NANDN U36666 ( .A(n35401), .B(n35400), .Z(n35405) );
  NANDN U36667 ( .A(n35403), .B(n35402), .Z(n35404) );
  AND U36668 ( .A(n35405), .B(n35404), .Z(n35432) );
  NAND U36669 ( .A(n42143), .B(n35406), .Z(n35408) );
  XNOR U36670 ( .A(a[841]), .B(n4192), .Z(n35443) );
  NAND U36671 ( .A(n42144), .B(n35443), .Z(n35407) );
  AND U36672 ( .A(n35408), .B(n35407), .Z(n35458) );
  XOR U36673 ( .A(a[845]), .B(n42012), .Z(n35446) );
  XNOR U36674 ( .A(n35458), .B(n35457), .Z(n35460) );
  XOR U36675 ( .A(a[843]), .B(n42085), .Z(n35447) );
  AND U36676 ( .A(a[839]), .B(b[7]), .Z(n35451) );
  XNOR U36677 ( .A(n35452), .B(n35451), .Z(n35453) );
  AND U36678 ( .A(a[847]), .B(b[0]), .Z(n35411) );
  XNOR U36679 ( .A(n35411), .B(n4071), .Z(n35413) );
  NANDN U36680 ( .A(b[0]), .B(a[846]), .Z(n35412) );
  NAND U36681 ( .A(n35413), .B(n35412), .Z(n35454) );
  XNOR U36682 ( .A(n35453), .B(n35454), .Z(n35459) );
  XOR U36683 ( .A(n35460), .B(n35459), .Z(n35438) );
  NANDN U36684 ( .A(n35415), .B(n35414), .Z(n35419) );
  NANDN U36685 ( .A(n35417), .B(n35416), .Z(n35418) );
  AND U36686 ( .A(n35419), .B(n35418), .Z(n35437) );
  XNOR U36687 ( .A(n35438), .B(n35437), .Z(n35439) );
  NANDN U36688 ( .A(n35421), .B(n35420), .Z(n35425) );
  NAND U36689 ( .A(n35423), .B(n35422), .Z(n35424) );
  NAND U36690 ( .A(n35425), .B(n35424), .Z(n35440) );
  XNOR U36691 ( .A(n35439), .B(n35440), .Z(n35431) );
  XNOR U36692 ( .A(n35432), .B(n35431), .Z(n35433) );
  XNOR U36693 ( .A(n35434), .B(n35433), .Z(n35463) );
  XNOR U36694 ( .A(sreg[1863]), .B(n35463), .Z(n35465) );
  NANDN U36695 ( .A(sreg[1862]), .B(n35426), .Z(n35430) );
  NAND U36696 ( .A(n35428), .B(n35427), .Z(n35429) );
  NAND U36697 ( .A(n35430), .B(n35429), .Z(n35464) );
  XNOR U36698 ( .A(n35465), .B(n35464), .Z(c[1863]) );
  NANDN U36699 ( .A(n35432), .B(n35431), .Z(n35436) );
  NANDN U36700 ( .A(n35434), .B(n35433), .Z(n35435) );
  AND U36701 ( .A(n35436), .B(n35435), .Z(n35471) );
  NANDN U36702 ( .A(n35438), .B(n35437), .Z(n35442) );
  NANDN U36703 ( .A(n35440), .B(n35439), .Z(n35441) );
  AND U36704 ( .A(n35442), .B(n35441), .Z(n35469) );
  NAND U36705 ( .A(n42143), .B(n35443), .Z(n35445) );
  XNOR U36706 ( .A(a[842]), .B(n4192), .Z(n35480) );
  NAND U36707 ( .A(n42144), .B(n35480), .Z(n35444) );
  AND U36708 ( .A(n35445), .B(n35444), .Z(n35495) );
  XOR U36709 ( .A(a[846]), .B(n42012), .Z(n35483) );
  XNOR U36710 ( .A(n35495), .B(n35494), .Z(n35497) );
  XOR U36711 ( .A(a[844]), .B(n42085), .Z(n35484) );
  AND U36712 ( .A(a[840]), .B(b[7]), .Z(n35488) );
  XNOR U36713 ( .A(n35489), .B(n35488), .Z(n35490) );
  AND U36714 ( .A(a[848]), .B(b[0]), .Z(n35448) );
  XNOR U36715 ( .A(n35448), .B(n4071), .Z(n35450) );
  NANDN U36716 ( .A(b[0]), .B(a[847]), .Z(n35449) );
  NAND U36717 ( .A(n35450), .B(n35449), .Z(n35491) );
  XNOR U36718 ( .A(n35490), .B(n35491), .Z(n35496) );
  XOR U36719 ( .A(n35497), .B(n35496), .Z(n35475) );
  NANDN U36720 ( .A(n35452), .B(n35451), .Z(n35456) );
  NANDN U36721 ( .A(n35454), .B(n35453), .Z(n35455) );
  AND U36722 ( .A(n35456), .B(n35455), .Z(n35474) );
  XNOR U36723 ( .A(n35475), .B(n35474), .Z(n35476) );
  NANDN U36724 ( .A(n35458), .B(n35457), .Z(n35462) );
  NAND U36725 ( .A(n35460), .B(n35459), .Z(n35461) );
  NAND U36726 ( .A(n35462), .B(n35461), .Z(n35477) );
  XNOR U36727 ( .A(n35476), .B(n35477), .Z(n35468) );
  XNOR U36728 ( .A(n35469), .B(n35468), .Z(n35470) );
  XNOR U36729 ( .A(n35471), .B(n35470), .Z(n35500) );
  XNOR U36730 ( .A(sreg[1864]), .B(n35500), .Z(n35502) );
  NANDN U36731 ( .A(sreg[1863]), .B(n35463), .Z(n35467) );
  NAND U36732 ( .A(n35465), .B(n35464), .Z(n35466) );
  NAND U36733 ( .A(n35467), .B(n35466), .Z(n35501) );
  XNOR U36734 ( .A(n35502), .B(n35501), .Z(c[1864]) );
  NANDN U36735 ( .A(n35469), .B(n35468), .Z(n35473) );
  NANDN U36736 ( .A(n35471), .B(n35470), .Z(n35472) );
  AND U36737 ( .A(n35473), .B(n35472), .Z(n35508) );
  NANDN U36738 ( .A(n35475), .B(n35474), .Z(n35479) );
  NANDN U36739 ( .A(n35477), .B(n35476), .Z(n35478) );
  AND U36740 ( .A(n35479), .B(n35478), .Z(n35506) );
  NAND U36741 ( .A(n42143), .B(n35480), .Z(n35482) );
  XNOR U36742 ( .A(a[843]), .B(n4192), .Z(n35517) );
  NAND U36743 ( .A(n42144), .B(n35517), .Z(n35481) );
  AND U36744 ( .A(n35482), .B(n35481), .Z(n35532) );
  XOR U36745 ( .A(a[847]), .B(n42012), .Z(n35520) );
  XNOR U36746 ( .A(n35532), .B(n35531), .Z(n35534) );
  XOR U36747 ( .A(a[845]), .B(n42085), .Z(n35521) );
  AND U36748 ( .A(a[841]), .B(b[7]), .Z(n35525) );
  XNOR U36749 ( .A(n35526), .B(n35525), .Z(n35527) );
  AND U36750 ( .A(a[849]), .B(b[0]), .Z(n35485) );
  XNOR U36751 ( .A(n35485), .B(n4071), .Z(n35487) );
  NANDN U36752 ( .A(b[0]), .B(a[848]), .Z(n35486) );
  NAND U36753 ( .A(n35487), .B(n35486), .Z(n35528) );
  XNOR U36754 ( .A(n35527), .B(n35528), .Z(n35533) );
  XOR U36755 ( .A(n35534), .B(n35533), .Z(n35512) );
  NANDN U36756 ( .A(n35489), .B(n35488), .Z(n35493) );
  NANDN U36757 ( .A(n35491), .B(n35490), .Z(n35492) );
  AND U36758 ( .A(n35493), .B(n35492), .Z(n35511) );
  XNOR U36759 ( .A(n35512), .B(n35511), .Z(n35513) );
  NANDN U36760 ( .A(n35495), .B(n35494), .Z(n35499) );
  NAND U36761 ( .A(n35497), .B(n35496), .Z(n35498) );
  NAND U36762 ( .A(n35499), .B(n35498), .Z(n35514) );
  XNOR U36763 ( .A(n35513), .B(n35514), .Z(n35505) );
  XNOR U36764 ( .A(n35506), .B(n35505), .Z(n35507) );
  XNOR U36765 ( .A(n35508), .B(n35507), .Z(n35537) );
  XNOR U36766 ( .A(sreg[1865]), .B(n35537), .Z(n35539) );
  NANDN U36767 ( .A(sreg[1864]), .B(n35500), .Z(n35504) );
  NAND U36768 ( .A(n35502), .B(n35501), .Z(n35503) );
  NAND U36769 ( .A(n35504), .B(n35503), .Z(n35538) );
  XNOR U36770 ( .A(n35539), .B(n35538), .Z(c[1865]) );
  NANDN U36771 ( .A(n35506), .B(n35505), .Z(n35510) );
  NANDN U36772 ( .A(n35508), .B(n35507), .Z(n35509) );
  AND U36773 ( .A(n35510), .B(n35509), .Z(n35545) );
  NANDN U36774 ( .A(n35512), .B(n35511), .Z(n35516) );
  NANDN U36775 ( .A(n35514), .B(n35513), .Z(n35515) );
  AND U36776 ( .A(n35516), .B(n35515), .Z(n35543) );
  NAND U36777 ( .A(n42143), .B(n35517), .Z(n35519) );
  XNOR U36778 ( .A(a[844]), .B(n4192), .Z(n35554) );
  NAND U36779 ( .A(n42144), .B(n35554), .Z(n35518) );
  AND U36780 ( .A(n35519), .B(n35518), .Z(n35569) );
  XOR U36781 ( .A(a[848]), .B(n42012), .Z(n35557) );
  XNOR U36782 ( .A(n35569), .B(n35568), .Z(n35571) );
  XOR U36783 ( .A(a[846]), .B(n42085), .Z(n35558) );
  AND U36784 ( .A(a[842]), .B(b[7]), .Z(n35562) );
  XNOR U36785 ( .A(n35563), .B(n35562), .Z(n35564) );
  AND U36786 ( .A(a[850]), .B(b[0]), .Z(n35522) );
  XNOR U36787 ( .A(n35522), .B(n4071), .Z(n35524) );
  NANDN U36788 ( .A(b[0]), .B(a[849]), .Z(n35523) );
  NAND U36789 ( .A(n35524), .B(n35523), .Z(n35565) );
  XNOR U36790 ( .A(n35564), .B(n35565), .Z(n35570) );
  XOR U36791 ( .A(n35571), .B(n35570), .Z(n35549) );
  NANDN U36792 ( .A(n35526), .B(n35525), .Z(n35530) );
  NANDN U36793 ( .A(n35528), .B(n35527), .Z(n35529) );
  AND U36794 ( .A(n35530), .B(n35529), .Z(n35548) );
  XNOR U36795 ( .A(n35549), .B(n35548), .Z(n35550) );
  NANDN U36796 ( .A(n35532), .B(n35531), .Z(n35536) );
  NAND U36797 ( .A(n35534), .B(n35533), .Z(n35535) );
  NAND U36798 ( .A(n35536), .B(n35535), .Z(n35551) );
  XNOR U36799 ( .A(n35550), .B(n35551), .Z(n35542) );
  XNOR U36800 ( .A(n35543), .B(n35542), .Z(n35544) );
  XNOR U36801 ( .A(n35545), .B(n35544), .Z(n35574) );
  XNOR U36802 ( .A(sreg[1866]), .B(n35574), .Z(n35576) );
  NANDN U36803 ( .A(sreg[1865]), .B(n35537), .Z(n35541) );
  NAND U36804 ( .A(n35539), .B(n35538), .Z(n35540) );
  NAND U36805 ( .A(n35541), .B(n35540), .Z(n35575) );
  XNOR U36806 ( .A(n35576), .B(n35575), .Z(c[1866]) );
  NANDN U36807 ( .A(n35543), .B(n35542), .Z(n35547) );
  NANDN U36808 ( .A(n35545), .B(n35544), .Z(n35546) );
  AND U36809 ( .A(n35547), .B(n35546), .Z(n35582) );
  NANDN U36810 ( .A(n35549), .B(n35548), .Z(n35553) );
  NANDN U36811 ( .A(n35551), .B(n35550), .Z(n35552) );
  AND U36812 ( .A(n35553), .B(n35552), .Z(n35580) );
  NAND U36813 ( .A(n42143), .B(n35554), .Z(n35556) );
  XNOR U36814 ( .A(a[845]), .B(n4192), .Z(n35591) );
  NAND U36815 ( .A(n42144), .B(n35591), .Z(n35555) );
  AND U36816 ( .A(n35556), .B(n35555), .Z(n35606) );
  XOR U36817 ( .A(a[849]), .B(n42012), .Z(n35594) );
  XNOR U36818 ( .A(n35606), .B(n35605), .Z(n35608) );
  XOR U36819 ( .A(a[847]), .B(n42085), .Z(n35598) );
  AND U36820 ( .A(a[843]), .B(b[7]), .Z(n35599) );
  XNOR U36821 ( .A(n35600), .B(n35599), .Z(n35601) );
  AND U36822 ( .A(a[851]), .B(b[0]), .Z(n35559) );
  XNOR U36823 ( .A(n35559), .B(n4071), .Z(n35561) );
  NANDN U36824 ( .A(b[0]), .B(a[850]), .Z(n35560) );
  NAND U36825 ( .A(n35561), .B(n35560), .Z(n35602) );
  XNOR U36826 ( .A(n35601), .B(n35602), .Z(n35607) );
  XOR U36827 ( .A(n35608), .B(n35607), .Z(n35586) );
  NANDN U36828 ( .A(n35563), .B(n35562), .Z(n35567) );
  NANDN U36829 ( .A(n35565), .B(n35564), .Z(n35566) );
  AND U36830 ( .A(n35567), .B(n35566), .Z(n35585) );
  XNOR U36831 ( .A(n35586), .B(n35585), .Z(n35587) );
  NANDN U36832 ( .A(n35569), .B(n35568), .Z(n35573) );
  NAND U36833 ( .A(n35571), .B(n35570), .Z(n35572) );
  NAND U36834 ( .A(n35573), .B(n35572), .Z(n35588) );
  XNOR U36835 ( .A(n35587), .B(n35588), .Z(n35579) );
  XNOR U36836 ( .A(n35580), .B(n35579), .Z(n35581) );
  XNOR U36837 ( .A(n35582), .B(n35581), .Z(n35611) );
  XNOR U36838 ( .A(sreg[1867]), .B(n35611), .Z(n35613) );
  NANDN U36839 ( .A(sreg[1866]), .B(n35574), .Z(n35578) );
  NAND U36840 ( .A(n35576), .B(n35575), .Z(n35577) );
  NAND U36841 ( .A(n35578), .B(n35577), .Z(n35612) );
  XNOR U36842 ( .A(n35613), .B(n35612), .Z(c[1867]) );
  NANDN U36843 ( .A(n35580), .B(n35579), .Z(n35584) );
  NANDN U36844 ( .A(n35582), .B(n35581), .Z(n35583) );
  AND U36845 ( .A(n35584), .B(n35583), .Z(n35619) );
  NANDN U36846 ( .A(n35586), .B(n35585), .Z(n35590) );
  NANDN U36847 ( .A(n35588), .B(n35587), .Z(n35589) );
  AND U36848 ( .A(n35590), .B(n35589), .Z(n35617) );
  NAND U36849 ( .A(n42143), .B(n35591), .Z(n35593) );
  XNOR U36850 ( .A(a[846]), .B(n4192), .Z(n35628) );
  NAND U36851 ( .A(n42144), .B(n35628), .Z(n35592) );
  AND U36852 ( .A(n35593), .B(n35592), .Z(n35643) );
  XOR U36853 ( .A(a[850]), .B(n42012), .Z(n35631) );
  XNOR U36854 ( .A(n35643), .B(n35642), .Z(n35645) );
  AND U36855 ( .A(a[852]), .B(b[0]), .Z(n35595) );
  XNOR U36856 ( .A(n35595), .B(n4071), .Z(n35597) );
  NANDN U36857 ( .A(b[0]), .B(a[851]), .Z(n35596) );
  NAND U36858 ( .A(n35597), .B(n35596), .Z(n35639) );
  XOR U36859 ( .A(a[848]), .B(n42085), .Z(n35635) );
  AND U36860 ( .A(a[844]), .B(b[7]), .Z(n35636) );
  XNOR U36861 ( .A(n35637), .B(n35636), .Z(n35638) );
  XNOR U36862 ( .A(n35639), .B(n35638), .Z(n35644) );
  XOR U36863 ( .A(n35645), .B(n35644), .Z(n35623) );
  NANDN U36864 ( .A(n35600), .B(n35599), .Z(n35604) );
  NANDN U36865 ( .A(n35602), .B(n35601), .Z(n35603) );
  AND U36866 ( .A(n35604), .B(n35603), .Z(n35622) );
  XNOR U36867 ( .A(n35623), .B(n35622), .Z(n35624) );
  NANDN U36868 ( .A(n35606), .B(n35605), .Z(n35610) );
  NAND U36869 ( .A(n35608), .B(n35607), .Z(n35609) );
  NAND U36870 ( .A(n35610), .B(n35609), .Z(n35625) );
  XNOR U36871 ( .A(n35624), .B(n35625), .Z(n35616) );
  XNOR U36872 ( .A(n35617), .B(n35616), .Z(n35618) );
  XNOR U36873 ( .A(n35619), .B(n35618), .Z(n35648) );
  XNOR U36874 ( .A(sreg[1868]), .B(n35648), .Z(n35650) );
  NANDN U36875 ( .A(sreg[1867]), .B(n35611), .Z(n35615) );
  NAND U36876 ( .A(n35613), .B(n35612), .Z(n35614) );
  NAND U36877 ( .A(n35615), .B(n35614), .Z(n35649) );
  XNOR U36878 ( .A(n35650), .B(n35649), .Z(c[1868]) );
  NANDN U36879 ( .A(n35617), .B(n35616), .Z(n35621) );
  NANDN U36880 ( .A(n35619), .B(n35618), .Z(n35620) );
  AND U36881 ( .A(n35621), .B(n35620), .Z(n35656) );
  NANDN U36882 ( .A(n35623), .B(n35622), .Z(n35627) );
  NANDN U36883 ( .A(n35625), .B(n35624), .Z(n35626) );
  AND U36884 ( .A(n35627), .B(n35626), .Z(n35654) );
  NAND U36885 ( .A(n42143), .B(n35628), .Z(n35630) );
  XNOR U36886 ( .A(a[847]), .B(n4192), .Z(n35665) );
  NAND U36887 ( .A(n42144), .B(n35665), .Z(n35629) );
  AND U36888 ( .A(n35630), .B(n35629), .Z(n35680) );
  XOR U36889 ( .A(a[851]), .B(n42012), .Z(n35668) );
  XNOR U36890 ( .A(n35680), .B(n35679), .Z(n35682) );
  AND U36891 ( .A(a[853]), .B(b[0]), .Z(n35632) );
  XNOR U36892 ( .A(n35632), .B(n4071), .Z(n35634) );
  NANDN U36893 ( .A(b[0]), .B(a[852]), .Z(n35633) );
  NAND U36894 ( .A(n35634), .B(n35633), .Z(n35676) );
  XOR U36895 ( .A(a[849]), .B(n42085), .Z(n35669) );
  AND U36896 ( .A(a[845]), .B(b[7]), .Z(n35673) );
  XNOR U36897 ( .A(n35674), .B(n35673), .Z(n35675) );
  XNOR U36898 ( .A(n35676), .B(n35675), .Z(n35681) );
  XOR U36899 ( .A(n35682), .B(n35681), .Z(n35660) );
  NANDN U36900 ( .A(n35637), .B(n35636), .Z(n35641) );
  NANDN U36901 ( .A(n35639), .B(n35638), .Z(n35640) );
  AND U36902 ( .A(n35641), .B(n35640), .Z(n35659) );
  XNOR U36903 ( .A(n35660), .B(n35659), .Z(n35661) );
  NANDN U36904 ( .A(n35643), .B(n35642), .Z(n35647) );
  NAND U36905 ( .A(n35645), .B(n35644), .Z(n35646) );
  NAND U36906 ( .A(n35647), .B(n35646), .Z(n35662) );
  XNOR U36907 ( .A(n35661), .B(n35662), .Z(n35653) );
  XNOR U36908 ( .A(n35654), .B(n35653), .Z(n35655) );
  XNOR U36909 ( .A(n35656), .B(n35655), .Z(n35685) );
  XNOR U36910 ( .A(sreg[1869]), .B(n35685), .Z(n35687) );
  NANDN U36911 ( .A(sreg[1868]), .B(n35648), .Z(n35652) );
  NAND U36912 ( .A(n35650), .B(n35649), .Z(n35651) );
  NAND U36913 ( .A(n35652), .B(n35651), .Z(n35686) );
  XNOR U36914 ( .A(n35687), .B(n35686), .Z(c[1869]) );
  NANDN U36915 ( .A(n35654), .B(n35653), .Z(n35658) );
  NANDN U36916 ( .A(n35656), .B(n35655), .Z(n35657) );
  AND U36917 ( .A(n35658), .B(n35657), .Z(n35693) );
  NANDN U36918 ( .A(n35660), .B(n35659), .Z(n35664) );
  NANDN U36919 ( .A(n35662), .B(n35661), .Z(n35663) );
  AND U36920 ( .A(n35664), .B(n35663), .Z(n35691) );
  NAND U36921 ( .A(n42143), .B(n35665), .Z(n35667) );
  XNOR U36922 ( .A(a[848]), .B(n4193), .Z(n35702) );
  NAND U36923 ( .A(n42144), .B(n35702), .Z(n35666) );
  AND U36924 ( .A(n35667), .B(n35666), .Z(n35717) );
  XOR U36925 ( .A(a[852]), .B(n42012), .Z(n35705) );
  XNOR U36926 ( .A(n35717), .B(n35716), .Z(n35719) );
  XOR U36927 ( .A(a[850]), .B(n42085), .Z(n35706) );
  AND U36928 ( .A(a[846]), .B(b[7]), .Z(n35710) );
  XNOR U36929 ( .A(n35711), .B(n35710), .Z(n35712) );
  AND U36930 ( .A(a[854]), .B(b[0]), .Z(n35670) );
  XNOR U36931 ( .A(n35670), .B(n4071), .Z(n35672) );
  NANDN U36932 ( .A(b[0]), .B(a[853]), .Z(n35671) );
  NAND U36933 ( .A(n35672), .B(n35671), .Z(n35713) );
  XNOR U36934 ( .A(n35712), .B(n35713), .Z(n35718) );
  XOR U36935 ( .A(n35719), .B(n35718), .Z(n35697) );
  NANDN U36936 ( .A(n35674), .B(n35673), .Z(n35678) );
  NANDN U36937 ( .A(n35676), .B(n35675), .Z(n35677) );
  AND U36938 ( .A(n35678), .B(n35677), .Z(n35696) );
  XNOR U36939 ( .A(n35697), .B(n35696), .Z(n35698) );
  NANDN U36940 ( .A(n35680), .B(n35679), .Z(n35684) );
  NAND U36941 ( .A(n35682), .B(n35681), .Z(n35683) );
  NAND U36942 ( .A(n35684), .B(n35683), .Z(n35699) );
  XNOR U36943 ( .A(n35698), .B(n35699), .Z(n35690) );
  XNOR U36944 ( .A(n35691), .B(n35690), .Z(n35692) );
  XNOR U36945 ( .A(n35693), .B(n35692), .Z(n35722) );
  XNOR U36946 ( .A(sreg[1870]), .B(n35722), .Z(n35724) );
  NANDN U36947 ( .A(sreg[1869]), .B(n35685), .Z(n35689) );
  NAND U36948 ( .A(n35687), .B(n35686), .Z(n35688) );
  NAND U36949 ( .A(n35689), .B(n35688), .Z(n35723) );
  XNOR U36950 ( .A(n35724), .B(n35723), .Z(c[1870]) );
  NANDN U36951 ( .A(n35691), .B(n35690), .Z(n35695) );
  NANDN U36952 ( .A(n35693), .B(n35692), .Z(n35694) );
  AND U36953 ( .A(n35695), .B(n35694), .Z(n35730) );
  NANDN U36954 ( .A(n35697), .B(n35696), .Z(n35701) );
  NANDN U36955 ( .A(n35699), .B(n35698), .Z(n35700) );
  AND U36956 ( .A(n35701), .B(n35700), .Z(n35728) );
  NAND U36957 ( .A(n42143), .B(n35702), .Z(n35704) );
  XNOR U36958 ( .A(a[849]), .B(n4193), .Z(n35739) );
  NAND U36959 ( .A(n42144), .B(n35739), .Z(n35703) );
  AND U36960 ( .A(n35704), .B(n35703), .Z(n35754) );
  XOR U36961 ( .A(a[853]), .B(n42012), .Z(n35742) );
  XNOR U36962 ( .A(n35754), .B(n35753), .Z(n35756) );
  XOR U36963 ( .A(a[851]), .B(n42085), .Z(n35743) );
  AND U36964 ( .A(a[847]), .B(b[7]), .Z(n35747) );
  XNOR U36965 ( .A(n35748), .B(n35747), .Z(n35749) );
  AND U36966 ( .A(a[855]), .B(b[0]), .Z(n35707) );
  XNOR U36967 ( .A(n35707), .B(n4071), .Z(n35709) );
  NANDN U36968 ( .A(b[0]), .B(a[854]), .Z(n35708) );
  NAND U36969 ( .A(n35709), .B(n35708), .Z(n35750) );
  XNOR U36970 ( .A(n35749), .B(n35750), .Z(n35755) );
  XOR U36971 ( .A(n35756), .B(n35755), .Z(n35734) );
  NANDN U36972 ( .A(n35711), .B(n35710), .Z(n35715) );
  NANDN U36973 ( .A(n35713), .B(n35712), .Z(n35714) );
  AND U36974 ( .A(n35715), .B(n35714), .Z(n35733) );
  XNOR U36975 ( .A(n35734), .B(n35733), .Z(n35735) );
  NANDN U36976 ( .A(n35717), .B(n35716), .Z(n35721) );
  NAND U36977 ( .A(n35719), .B(n35718), .Z(n35720) );
  NAND U36978 ( .A(n35721), .B(n35720), .Z(n35736) );
  XNOR U36979 ( .A(n35735), .B(n35736), .Z(n35727) );
  XNOR U36980 ( .A(n35728), .B(n35727), .Z(n35729) );
  XNOR U36981 ( .A(n35730), .B(n35729), .Z(n35759) );
  XNOR U36982 ( .A(sreg[1871]), .B(n35759), .Z(n35761) );
  NANDN U36983 ( .A(sreg[1870]), .B(n35722), .Z(n35726) );
  NAND U36984 ( .A(n35724), .B(n35723), .Z(n35725) );
  NAND U36985 ( .A(n35726), .B(n35725), .Z(n35760) );
  XNOR U36986 ( .A(n35761), .B(n35760), .Z(c[1871]) );
  NANDN U36987 ( .A(n35728), .B(n35727), .Z(n35732) );
  NANDN U36988 ( .A(n35730), .B(n35729), .Z(n35731) );
  AND U36989 ( .A(n35732), .B(n35731), .Z(n35767) );
  NANDN U36990 ( .A(n35734), .B(n35733), .Z(n35738) );
  NANDN U36991 ( .A(n35736), .B(n35735), .Z(n35737) );
  AND U36992 ( .A(n35738), .B(n35737), .Z(n35765) );
  NAND U36993 ( .A(n42143), .B(n35739), .Z(n35741) );
  XNOR U36994 ( .A(a[850]), .B(n4193), .Z(n35776) );
  NAND U36995 ( .A(n42144), .B(n35776), .Z(n35740) );
  AND U36996 ( .A(n35741), .B(n35740), .Z(n35791) );
  XOR U36997 ( .A(a[854]), .B(n42012), .Z(n35779) );
  XNOR U36998 ( .A(n35791), .B(n35790), .Z(n35793) );
  XOR U36999 ( .A(a[852]), .B(n42085), .Z(n35780) );
  AND U37000 ( .A(a[848]), .B(b[7]), .Z(n35784) );
  XNOR U37001 ( .A(n35785), .B(n35784), .Z(n35786) );
  AND U37002 ( .A(a[856]), .B(b[0]), .Z(n35744) );
  XNOR U37003 ( .A(n35744), .B(n4071), .Z(n35746) );
  NANDN U37004 ( .A(b[0]), .B(a[855]), .Z(n35745) );
  NAND U37005 ( .A(n35746), .B(n35745), .Z(n35787) );
  XNOR U37006 ( .A(n35786), .B(n35787), .Z(n35792) );
  XOR U37007 ( .A(n35793), .B(n35792), .Z(n35771) );
  NANDN U37008 ( .A(n35748), .B(n35747), .Z(n35752) );
  NANDN U37009 ( .A(n35750), .B(n35749), .Z(n35751) );
  AND U37010 ( .A(n35752), .B(n35751), .Z(n35770) );
  XNOR U37011 ( .A(n35771), .B(n35770), .Z(n35772) );
  NANDN U37012 ( .A(n35754), .B(n35753), .Z(n35758) );
  NAND U37013 ( .A(n35756), .B(n35755), .Z(n35757) );
  NAND U37014 ( .A(n35758), .B(n35757), .Z(n35773) );
  XNOR U37015 ( .A(n35772), .B(n35773), .Z(n35764) );
  XNOR U37016 ( .A(n35765), .B(n35764), .Z(n35766) );
  XNOR U37017 ( .A(n35767), .B(n35766), .Z(n35796) );
  XNOR U37018 ( .A(sreg[1872]), .B(n35796), .Z(n35798) );
  NANDN U37019 ( .A(sreg[1871]), .B(n35759), .Z(n35763) );
  NAND U37020 ( .A(n35761), .B(n35760), .Z(n35762) );
  NAND U37021 ( .A(n35763), .B(n35762), .Z(n35797) );
  XNOR U37022 ( .A(n35798), .B(n35797), .Z(c[1872]) );
  NANDN U37023 ( .A(n35765), .B(n35764), .Z(n35769) );
  NANDN U37024 ( .A(n35767), .B(n35766), .Z(n35768) );
  AND U37025 ( .A(n35769), .B(n35768), .Z(n35804) );
  NANDN U37026 ( .A(n35771), .B(n35770), .Z(n35775) );
  NANDN U37027 ( .A(n35773), .B(n35772), .Z(n35774) );
  AND U37028 ( .A(n35775), .B(n35774), .Z(n35802) );
  NAND U37029 ( .A(n42143), .B(n35776), .Z(n35778) );
  XNOR U37030 ( .A(a[851]), .B(n4193), .Z(n35813) );
  NAND U37031 ( .A(n42144), .B(n35813), .Z(n35777) );
  AND U37032 ( .A(n35778), .B(n35777), .Z(n35828) );
  XOR U37033 ( .A(a[855]), .B(n42012), .Z(n35816) );
  XNOR U37034 ( .A(n35828), .B(n35827), .Z(n35830) );
  XOR U37035 ( .A(a[853]), .B(n42085), .Z(n35820) );
  AND U37036 ( .A(a[849]), .B(b[7]), .Z(n35821) );
  XNOR U37037 ( .A(n35822), .B(n35821), .Z(n35823) );
  AND U37038 ( .A(a[857]), .B(b[0]), .Z(n35781) );
  XNOR U37039 ( .A(n35781), .B(n4071), .Z(n35783) );
  NANDN U37040 ( .A(b[0]), .B(a[856]), .Z(n35782) );
  NAND U37041 ( .A(n35783), .B(n35782), .Z(n35824) );
  XNOR U37042 ( .A(n35823), .B(n35824), .Z(n35829) );
  XOR U37043 ( .A(n35830), .B(n35829), .Z(n35808) );
  NANDN U37044 ( .A(n35785), .B(n35784), .Z(n35789) );
  NANDN U37045 ( .A(n35787), .B(n35786), .Z(n35788) );
  AND U37046 ( .A(n35789), .B(n35788), .Z(n35807) );
  XNOR U37047 ( .A(n35808), .B(n35807), .Z(n35809) );
  NANDN U37048 ( .A(n35791), .B(n35790), .Z(n35795) );
  NAND U37049 ( .A(n35793), .B(n35792), .Z(n35794) );
  NAND U37050 ( .A(n35795), .B(n35794), .Z(n35810) );
  XNOR U37051 ( .A(n35809), .B(n35810), .Z(n35801) );
  XNOR U37052 ( .A(n35802), .B(n35801), .Z(n35803) );
  XNOR U37053 ( .A(n35804), .B(n35803), .Z(n35833) );
  XNOR U37054 ( .A(sreg[1873]), .B(n35833), .Z(n35835) );
  NANDN U37055 ( .A(sreg[1872]), .B(n35796), .Z(n35800) );
  NAND U37056 ( .A(n35798), .B(n35797), .Z(n35799) );
  NAND U37057 ( .A(n35800), .B(n35799), .Z(n35834) );
  XNOR U37058 ( .A(n35835), .B(n35834), .Z(c[1873]) );
  NANDN U37059 ( .A(n35802), .B(n35801), .Z(n35806) );
  NANDN U37060 ( .A(n35804), .B(n35803), .Z(n35805) );
  AND U37061 ( .A(n35806), .B(n35805), .Z(n35841) );
  NANDN U37062 ( .A(n35808), .B(n35807), .Z(n35812) );
  NANDN U37063 ( .A(n35810), .B(n35809), .Z(n35811) );
  AND U37064 ( .A(n35812), .B(n35811), .Z(n35839) );
  NAND U37065 ( .A(n42143), .B(n35813), .Z(n35815) );
  XNOR U37066 ( .A(a[852]), .B(n4193), .Z(n35850) );
  NAND U37067 ( .A(n42144), .B(n35850), .Z(n35814) );
  AND U37068 ( .A(n35815), .B(n35814), .Z(n35865) );
  XOR U37069 ( .A(a[856]), .B(n42012), .Z(n35853) );
  XNOR U37070 ( .A(n35865), .B(n35864), .Z(n35867) );
  AND U37071 ( .A(a[858]), .B(b[0]), .Z(n35817) );
  XNOR U37072 ( .A(n35817), .B(n4071), .Z(n35819) );
  NANDN U37073 ( .A(b[0]), .B(a[857]), .Z(n35818) );
  NAND U37074 ( .A(n35819), .B(n35818), .Z(n35861) );
  XOR U37075 ( .A(a[854]), .B(n42085), .Z(n35857) );
  AND U37076 ( .A(a[850]), .B(b[7]), .Z(n35858) );
  XNOR U37077 ( .A(n35859), .B(n35858), .Z(n35860) );
  XNOR U37078 ( .A(n35861), .B(n35860), .Z(n35866) );
  XOR U37079 ( .A(n35867), .B(n35866), .Z(n35845) );
  NANDN U37080 ( .A(n35822), .B(n35821), .Z(n35826) );
  NANDN U37081 ( .A(n35824), .B(n35823), .Z(n35825) );
  AND U37082 ( .A(n35826), .B(n35825), .Z(n35844) );
  XNOR U37083 ( .A(n35845), .B(n35844), .Z(n35846) );
  NANDN U37084 ( .A(n35828), .B(n35827), .Z(n35832) );
  NAND U37085 ( .A(n35830), .B(n35829), .Z(n35831) );
  NAND U37086 ( .A(n35832), .B(n35831), .Z(n35847) );
  XNOR U37087 ( .A(n35846), .B(n35847), .Z(n35838) );
  XNOR U37088 ( .A(n35839), .B(n35838), .Z(n35840) );
  XNOR U37089 ( .A(n35841), .B(n35840), .Z(n35870) );
  XNOR U37090 ( .A(sreg[1874]), .B(n35870), .Z(n35872) );
  NANDN U37091 ( .A(sreg[1873]), .B(n35833), .Z(n35837) );
  NAND U37092 ( .A(n35835), .B(n35834), .Z(n35836) );
  NAND U37093 ( .A(n35837), .B(n35836), .Z(n35871) );
  XNOR U37094 ( .A(n35872), .B(n35871), .Z(c[1874]) );
  NANDN U37095 ( .A(n35839), .B(n35838), .Z(n35843) );
  NANDN U37096 ( .A(n35841), .B(n35840), .Z(n35842) );
  AND U37097 ( .A(n35843), .B(n35842), .Z(n35878) );
  NANDN U37098 ( .A(n35845), .B(n35844), .Z(n35849) );
  NANDN U37099 ( .A(n35847), .B(n35846), .Z(n35848) );
  AND U37100 ( .A(n35849), .B(n35848), .Z(n35876) );
  NAND U37101 ( .A(n42143), .B(n35850), .Z(n35852) );
  XNOR U37102 ( .A(a[853]), .B(n4193), .Z(n35887) );
  NAND U37103 ( .A(n42144), .B(n35887), .Z(n35851) );
  AND U37104 ( .A(n35852), .B(n35851), .Z(n35902) );
  XOR U37105 ( .A(a[857]), .B(n42012), .Z(n35890) );
  XNOR U37106 ( .A(n35902), .B(n35901), .Z(n35904) );
  AND U37107 ( .A(a[859]), .B(b[0]), .Z(n35854) );
  XNOR U37108 ( .A(n35854), .B(n4071), .Z(n35856) );
  NANDN U37109 ( .A(b[0]), .B(a[858]), .Z(n35855) );
  NAND U37110 ( .A(n35856), .B(n35855), .Z(n35898) );
  XOR U37111 ( .A(a[855]), .B(n42085), .Z(n35894) );
  AND U37112 ( .A(a[851]), .B(b[7]), .Z(n35895) );
  XNOR U37113 ( .A(n35896), .B(n35895), .Z(n35897) );
  XNOR U37114 ( .A(n35898), .B(n35897), .Z(n35903) );
  XOR U37115 ( .A(n35904), .B(n35903), .Z(n35882) );
  NANDN U37116 ( .A(n35859), .B(n35858), .Z(n35863) );
  NANDN U37117 ( .A(n35861), .B(n35860), .Z(n35862) );
  AND U37118 ( .A(n35863), .B(n35862), .Z(n35881) );
  XNOR U37119 ( .A(n35882), .B(n35881), .Z(n35883) );
  NANDN U37120 ( .A(n35865), .B(n35864), .Z(n35869) );
  NAND U37121 ( .A(n35867), .B(n35866), .Z(n35868) );
  NAND U37122 ( .A(n35869), .B(n35868), .Z(n35884) );
  XNOR U37123 ( .A(n35883), .B(n35884), .Z(n35875) );
  XNOR U37124 ( .A(n35876), .B(n35875), .Z(n35877) );
  XNOR U37125 ( .A(n35878), .B(n35877), .Z(n35907) );
  XNOR U37126 ( .A(sreg[1875]), .B(n35907), .Z(n35909) );
  NANDN U37127 ( .A(sreg[1874]), .B(n35870), .Z(n35874) );
  NAND U37128 ( .A(n35872), .B(n35871), .Z(n35873) );
  NAND U37129 ( .A(n35874), .B(n35873), .Z(n35908) );
  XNOR U37130 ( .A(n35909), .B(n35908), .Z(c[1875]) );
  NANDN U37131 ( .A(n35876), .B(n35875), .Z(n35880) );
  NANDN U37132 ( .A(n35878), .B(n35877), .Z(n35879) );
  AND U37133 ( .A(n35880), .B(n35879), .Z(n35915) );
  NANDN U37134 ( .A(n35882), .B(n35881), .Z(n35886) );
  NANDN U37135 ( .A(n35884), .B(n35883), .Z(n35885) );
  AND U37136 ( .A(n35886), .B(n35885), .Z(n35913) );
  NAND U37137 ( .A(n42143), .B(n35887), .Z(n35889) );
  XNOR U37138 ( .A(a[854]), .B(n4193), .Z(n35924) );
  NAND U37139 ( .A(n42144), .B(n35924), .Z(n35888) );
  AND U37140 ( .A(n35889), .B(n35888), .Z(n35939) );
  XOR U37141 ( .A(a[858]), .B(n42012), .Z(n35927) );
  XNOR U37142 ( .A(n35939), .B(n35938), .Z(n35941) );
  AND U37143 ( .A(a[860]), .B(b[0]), .Z(n35891) );
  XNOR U37144 ( .A(n35891), .B(n4071), .Z(n35893) );
  NANDN U37145 ( .A(b[0]), .B(a[859]), .Z(n35892) );
  NAND U37146 ( .A(n35893), .B(n35892), .Z(n35935) );
  XOR U37147 ( .A(a[856]), .B(n42085), .Z(n35928) );
  AND U37148 ( .A(a[852]), .B(b[7]), .Z(n35932) );
  XNOR U37149 ( .A(n35933), .B(n35932), .Z(n35934) );
  XNOR U37150 ( .A(n35935), .B(n35934), .Z(n35940) );
  XOR U37151 ( .A(n35941), .B(n35940), .Z(n35919) );
  NANDN U37152 ( .A(n35896), .B(n35895), .Z(n35900) );
  NANDN U37153 ( .A(n35898), .B(n35897), .Z(n35899) );
  AND U37154 ( .A(n35900), .B(n35899), .Z(n35918) );
  XNOR U37155 ( .A(n35919), .B(n35918), .Z(n35920) );
  NANDN U37156 ( .A(n35902), .B(n35901), .Z(n35906) );
  NAND U37157 ( .A(n35904), .B(n35903), .Z(n35905) );
  NAND U37158 ( .A(n35906), .B(n35905), .Z(n35921) );
  XNOR U37159 ( .A(n35920), .B(n35921), .Z(n35912) );
  XNOR U37160 ( .A(n35913), .B(n35912), .Z(n35914) );
  XNOR U37161 ( .A(n35915), .B(n35914), .Z(n35944) );
  XNOR U37162 ( .A(sreg[1876]), .B(n35944), .Z(n35946) );
  NANDN U37163 ( .A(sreg[1875]), .B(n35907), .Z(n35911) );
  NAND U37164 ( .A(n35909), .B(n35908), .Z(n35910) );
  NAND U37165 ( .A(n35911), .B(n35910), .Z(n35945) );
  XNOR U37166 ( .A(n35946), .B(n35945), .Z(c[1876]) );
  NANDN U37167 ( .A(n35913), .B(n35912), .Z(n35917) );
  NANDN U37168 ( .A(n35915), .B(n35914), .Z(n35916) );
  AND U37169 ( .A(n35917), .B(n35916), .Z(n35952) );
  NANDN U37170 ( .A(n35919), .B(n35918), .Z(n35923) );
  NANDN U37171 ( .A(n35921), .B(n35920), .Z(n35922) );
  AND U37172 ( .A(n35923), .B(n35922), .Z(n35950) );
  NAND U37173 ( .A(n42143), .B(n35924), .Z(n35926) );
  XNOR U37174 ( .A(a[855]), .B(n4194), .Z(n35961) );
  NAND U37175 ( .A(n42144), .B(n35961), .Z(n35925) );
  AND U37176 ( .A(n35926), .B(n35925), .Z(n35976) );
  XOR U37177 ( .A(a[859]), .B(n42012), .Z(n35964) );
  XNOR U37178 ( .A(n35976), .B(n35975), .Z(n35978) );
  XOR U37179 ( .A(a[857]), .B(n42085), .Z(n35968) );
  AND U37180 ( .A(a[853]), .B(b[7]), .Z(n35969) );
  XNOR U37181 ( .A(n35970), .B(n35969), .Z(n35971) );
  AND U37182 ( .A(a[861]), .B(b[0]), .Z(n35929) );
  XNOR U37183 ( .A(n35929), .B(n4071), .Z(n35931) );
  NANDN U37184 ( .A(b[0]), .B(a[860]), .Z(n35930) );
  NAND U37185 ( .A(n35931), .B(n35930), .Z(n35972) );
  XNOR U37186 ( .A(n35971), .B(n35972), .Z(n35977) );
  XOR U37187 ( .A(n35978), .B(n35977), .Z(n35956) );
  NANDN U37188 ( .A(n35933), .B(n35932), .Z(n35937) );
  NANDN U37189 ( .A(n35935), .B(n35934), .Z(n35936) );
  AND U37190 ( .A(n35937), .B(n35936), .Z(n35955) );
  XNOR U37191 ( .A(n35956), .B(n35955), .Z(n35957) );
  NANDN U37192 ( .A(n35939), .B(n35938), .Z(n35943) );
  NAND U37193 ( .A(n35941), .B(n35940), .Z(n35942) );
  NAND U37194 ( .A(n35943), .B(n35942), .Z(n35958) );
  XNOR U37195 ( .A(n35957), .B(n35958), .Z(n35949) );
  XNOR U37196 ( .A(n35950), .B(n35949), .Z(n35951) );
  XNOR U37197 ( .A(n35952), .B(n35951), .Z(n35981) );
  XNOR U37198 ( .A(sreg[1877]), .B(n35981), .Z(n35983) );
  NANDN U37199 ( .A(sreg[1876]), .B(n35944), .Z(n35948) );
  NAND U37200 ( .A(n35946), .B(n35945), .Z(n35947) );
  NAND U37201 ( .A(n35948), .B(n35947), .Z(n35982) );
  XNOR U37202 ( .A(n35983), .B(n35982), .Z(c[1877]) );
  NANDN U37203 ( .A(n35950), .B(n35949), .Z(n35954) );
  NANDN U37204 ( .A(n35952), .B(n35951), .Z(n35953) );
  AND U37205 ( .A(n35954), .B(n35953), .Z(n35989) );
  NANDN U37206 ( .A(n35956), .B(n35955), .Z(n35960) );
  NANDN U37207 ( .A(n35958), .B(n35957), .Z(n35959) );
  AND U37208 ( .A(n35960), .B(n35959), .Z(n35987) );
  NAND U37209 ( .A(n42143), .B(n35961), .Z(n35963) );
  XNOR U37210 ( .A(a[856]), .B(n4194), .Z(n35998) );
  NAND U37211 ( .A(n42144), .B(n35998), .Z(n35962) );
  AND U37212 ( .A(n35963), .B(n35962), .Z(n36013) );
  XOR U37213 ( .A(a[860]), .B(n42012), .Z(n36001) );
  XNOR U37214 ( .A(n36013), .B(n36012), .Z(n36015) );
  AND U37215 ( .A(a[862]), .B(b[0]), .Z(n35965) );
  XNOR U37216 ( .A(n35965), .B(n4071), .Z(n35967) );
  NANDN U37217 ( .A(b[0]), .B(a[861]), .Z(n35966) );
  NAND U37218 ( .A(n35967), .B(n35966), .Z(n36009) );
  XOR U37219 ( .A(a[858]), .B(n42085), .Z(n36002) );
  AND U37220 ( .A(a[854]), .B(b[7]), .Z(n36006) );
  XNOR U37221 ( .A(n36007), .B(n36006), .Z(n36008) );
  XNOR U37222 ( .A(n36009), .B(n36008), .Z(n36014) );
  XOR U37223 ( .A(n36015), .B(n36014), .Z(n35993) );
  NANDN U37224 ( .A(n35970), .B(n35969), .Z(n35974) );
  NANDN U37225 ( .A(n35972), .B(n35971), .Z(n35973) );
  AND U37226 ( .A(n35974), .B(n35973), .Z(n35992) );
  XNOR U37227 ( .A(n35993), .B(n35992), .Z(n35994) );
  NANDN U37228 ( .A(n35976), .B(n35975), .Z(n35980) );
  NAND U37229 ( .A(n35978), .B(n35977), .Z(n35979) );
  NAND U37230 ( .A(n35980), .B(n35979), .Z(n35995) );
  XNOR U37231 ( .A(n35994), .B(n35995), .Z(n35986) );
  XNOR U37232 ( .A(n35987), .B(n35986), .Z(n35988) );
  XNOR U37233 ( .A(n35989), .B(n35988), .Z(n36018) );
  XNOR U37234 ( .A(sreg[1878]), .B(n36018), .Z(n36020) );
  NANDN U37235 ( .A(sreg[1877]), .B(n35981), .Z(n35985) );
  NAND U37236 ( .A(n35983), .B(n35982), .Z(n35984) );
  NAND U37237 ( .A(n35985), .B(n35984), .Z(n36019) );
  XNOR U37238 ( .A(n36020), .B(n36019), .Z(c[1878]) );
  NANDN U37239 ( .A(n35987), .B(n35986), .Z(n35991) );
  NANDN U37240 ( .A(n35989), .B(n35988), .Z(n35990) );
  AND U37241 ( .A(n35991), .B(n35990), .Z(n36026) );
  NANDN U37242 ( .A(n35993), .B(n35992), .Z(n35997) );
  NANDN U37243 ( .A(n35995), .B(n35994), .Z(n35996) );
  AND U37244 ( .A(n35997), .B(n35996), .Z(n36024) );
  NAND U37245 ( .A(n42143), .B(n35998), .Z(n36000) );
  XNOR U37246 ( .A(a[857]), .B(n4194), .Z(n36035) );
  NAND U37247 ( .A(n42144), .B(n36035), .Z(n35999) );
  AND U37248 ( .A(n36000), .B(n35999), .Z(n36050) );
  XOR U37249 ( .A(a[861]), .B(n42012), .Z(n36038) );
  XNOR U37250 ( .A(n36050), .B(n36049), .Z(n36052) );
  XOR U37251 ( .A(a[859]), .B(n42085), .Z(n36042) );
  AND U37252 ( .A(a[855]), .B(b[7]), .Z(n36043) );
  XNOR U37253 ( .A(n36044), .B(n36043), .Z(n36045) );
  AND U37254 ( .A(a[863]), .B(b[0]), .Z(n36003) );
  XNOR U37255 ( .A(n36003), .B(n4071), .Z(n36005) );
  NANDN U37256 ( .A(b[0]), .B(a[862]), .Z(n36004) );
  NAND U37257 ( .A(n36005), .B(n36004), .Z(n36046) );
  XNOR U37258 ( .A(n36045), .B(n36046), .Z(n36051) );
  XOR U37259 ( .A(n36052), .B(n36051), .Z(n36030) );
  NANDN U37260 ( .A(n36007), .B(n36006), .Z(n36011) );
  NANDN U37261 ( .A(n36009), .B(n36008), .Z(n36010) );
  AND U37262 ( .A(n36011), .B(n36010), .Z(n36029) );
  XNOR U37263 ( .A(n36030), .B(n36029), .Z(n36031) );
  NANDN U37264 ( .A(n36013), .B(n36012), .Z(n36017) );
  NAND U37265 ( .A(n36015), .B(n36014), .Z(n36016) );
  NAND U37266 ( .A(n36017), .B(n36016), .Z(n36032) );
  XNOR U37267 ( .A(n36031), .B(n36032), .Z(n36023) );
  XNOR U37268 ( .A(n36024), .B(n36023), .Z(n36025) );
  XNOR U37269 ( .A(n36026), .B(n36025), .Z(n36055) );
  XNOR U37270 ( .A(sreg[1879]), .B(n36055), .Z(n36057) );
  NANDN U37271 ( .A(sreg[1878]), .B(n36018), .Z(n36022) );
  NAND U37272 ( .A(n36020), .B(n36019), .Z(n36021) );
  NAND U37273 ( .A(n36022), .B(n36021), .Z(n36056) );
  XNOR U37274 ( .A(n36057), .B(n36056), .Z(c[1879]) );
  NANDN U37275 ( .A(n36024), .B(n36023), .Z(n36028) );
  NANDN U37276 ( .A(n36026), .B(n36025), .Z(n36027) );
  AND U37277 ( .A(n36028), .B(n36027), .Z(n36063) );
  NANDN U37278 ( .A(n36030), .B(n36029), .Z(n36034) );
  NANDN U37279 ( .A(n36032), .B(n36031), .Z(n36033) );
  AND U37280 ( .A(n36034), .B(n36033), .Z(n36061) );
  NAND U37281 ( .A(n42143), .B(n36035), .Z(n36037) );
  XNOR U37282 ( .A(a[858]), .B(n4194), .Z(n36072) );
  NAND U37283 ( .A(n42144), .B(n36072), .Z(n36036) );
  AND U37284 ( .A(n36037), .B(n36036), .Z(n36087) );
  XOR U37285 ( .A(a[862]), .B(n42012), .Z(n36075) );
  XNOR U37286 ( .A(n36087), .B(n36086), .Z(n36089) );
  AND U37287 ( .A(a[864]), .B(b[0]), .Z(n36039) );
  XNOR U37288 ( .A(n36039), .B(n4071), .Z(n36041) );
  NANDN U37289 ( .A(b[0]), .B(a[863]), .Z(n36040) );
  NAND U37290 ( .A(n36041), .B(n36040), .Z(n36083) );
  XOR U37291 ( .A(a[860]), .B(n42085), .Z(n36079) );
  AND U37292 ( .A(a[856]), .B(b[7]), .Z(n36080) );
  XNOR U37293 ( .A(n36081), .B(n36080), .Z(n36082) );
  XNOR U37294 ( .A(n36083), .B(n36082), .Z(n36088) );
  XOR U37295 ( .A(n36089), .B(n36088), .Z(n36067) );
  NANDN U37296 ( .A(n36044), .B(n36043), .Z(n36048) );
  NANDN U37297 ( .A(n36046), .B(n36045), .Z(n36047) );
  AND U37298 ( .A(n36048), .B(n36047), .Z(n36066) );
  XNOR U37299 ( .A(n36067), .B(n36066), .Z(n36068) );
  NANDN U37300 ( .A(n36050), .B(n36049), .Z(n36054) );
  NAND U37301 ( .A(n36052), .B(n36051), .Z(n36053) );
  NAND U37302 ( .A(n36054), .B(n36053), .Z(n36069) );
  XNOR U37303 ( .A(n36068), .B(n36069), .Z(n36060) );
  XNOR U37304 ( .A(n36061), .B(n36060), .Z(n36062) );
  XNOR U37305 ( .A(n36063), .B(n36062), .Z(n36092) );
  XNOR U37306 ( .A(sreg[1880]), .B(n36092), .Z(n36094) );
  NANDN U37307 ( .A(sreg[1879]), .B(n36055), .Z(n36059) );
  NAND U37308 ( .A(n36057), .B(n36056), .Z(n36058) );
  NAND U37309 ( .A(n36059), .B(n36058), .Z(n36093) );
  XNOR U37310 ( .A(n36094), .B(n36093), .Z(c[1880]) );
  NANDN U37311 ( .A(n36061), .B(n36060), .Z(n36065) );
  NANDN U37312 ( .A(n36063), .B(n36062), .Z(n36064) );
  AND U37313 ( .A(n36065), .B(n36064), .Z(n36100) );
  NANDN U37314 ( .A(n36067), .B(n36066), .Z(n36071) );
  NANDN U37315 ( .A(n36069), .B(n36068), .Z(n36070) );
  AND U37316 ( .A(n36071), .B(n36070), .Z(n36098) );
  NAND U37317 ( .A(n42143), .B(n36072), .Z(n36074) );
  XNOR U37318 ( .A(a[859]), .B(n4194), .Z(n36109) );
  NAND U37319 ( .A(n42144), .B(n36109), .Z(n36073) );
  AND U37320 ( .A(n36074), .B(n36073), .Z(n36124) );
  XOR U37321 ( .A(a[863]), .B(n42012), .Z(n36112) );
  XNOR U37322 ( .A(n36124), .B(n36123), .Z(n36126) );
  AND U37323 ( .A(a[865]), .B(b[0]), .Z(n36076) );
  XNOR U37324 ( .A(n36076), .B(n4071), .Z(n36078) );
  NANDN U37325 ( .A(b[0]), .B(a[864]), .Z(n36077) );
  NAND U37326 ( .A(n36078), .B(n36077), .Z(n36120) );
  XOR U37327 ( .A(a[861]), .B(n42085), .Z(n36113) );
  AND U37328 ( .A(a[857]), .B(b[7]), .Z(n36117) );
  XNOR U37329 ( .A(n36118), .B(n36117), .Z(n36119) );
  XNOR U37330 ( .A(n36120), .B(n36119), .Z(n36125) );
  XOR U37331 ( .A(n36126), .B(n36125), .Z(n36104) );
  NANDN U37332 ( .A(n36081), .B(n36080), .Z(n36085) );
  NANDN U37333 ( .A(n36083), .B(n36082), .Z(n36084) );
  AND U37334 ( .A(n36085), .B(n36084), .Z(n36103) );
  XNOR U37335 ( .A(n36104), .B(n36103), .Z(n36105) );
  NANDN U37336 ( .A(n36087), .B(n36086), .Z(n36091) );
  NAND U37337 ( .A(n36089), .B(n36088), .Z(n36090) );
  NAND U37338 ( .A(n36091), .B(n36090), .Z(n36106) );
  XNOR U37339 ( .A(n36105), .B(n36106), .Z(n36097) );
  XNOR U37340 ( .A(n36098), .B(n36097), .Z(n36099) );
  XNOR U37341 ( .A(n36100), .B(n36099), .Z(n36129) );
  XNOR U37342 ( .A(sreg[1881]), .B(n36129), .Z(n36131) );
  NANDN U37343 ( .A(sreg[1880]), .B(n36092), .Z(n36096) );
  NAND U37344 ( .A(n36094), .B(n36093), .Z(n36095) );
  NAND U37345 ( .A(n36096), .B(n36095), .Z(n36130) );
  XNOR U37346 ( .A(n36131), .B(n36130), .Z(c[1881]) );
  NANDN U37347 ( .A(n36098), .B(n36097), .Z(n36102) );
  NANDN U37348 ( .A(n36100), .B(n36099), .Z(n36101) );
  AND U37349 ( .A(n36102), .B(n36101), .Z(n36137) );
  NANDN U37350 ( .A(n36104), .B(n36103), .Z(n36108) );
  NANDN U37351 ( .A(n36106), .B(n36105), .Z(n36107) );
  AND U37352 ( .A(n36108), .B(n36107), .Z(n36135) );
  NAND U37353 ( .A(n42143), .B(n36109), .Z(n36111) );
  XNOR U37354 ( .A(a[860]), .B(n4194), .Z(n36146) );
  NAND U37355 ( .A(n42144), .B(n36146), .Z(n36110) );
  AND U37356 ( .A(n36111), .B(n36110), .Z(n36161) );
  XOR U37357 ( .A(a[864]), .B(n42012), .Z(n36149) );
  XNOR U37358 ( .A(n36161), .B(n36160), .Z(n36163) );
  XOR U37359 ( .A(a[862]), .B(n42085), .Z(n36153) );
  AND U37360 ( .A(a[858]), .B(b[7]), .Z(n36154) );
  XNOR U37361 ( .A(n36155), .B(n36154), .Z(n36156) );
  AND U37362 ( .A(a[866]), .B(b[0]), .Z(n36114) );
  XNOR U37363 ( .A(n36114), .B(n4071), .Z(n36116) );
  NANDN U37364 ( .A(b[0]), .B(a[865]), .Z(n36115) );
  NAND U37365 ( .A(n36116), .B(n36115), .Z(n36157) );
  XNOR U37366 ( .A(n36156), .B(n36157), .Z(n36162) );
  XOR U37367 ( .A(n36163), .B(n36162), .Z(n36141) );
  NANDN U37368 ( .A(n36118), .B(n36117), .Z(n36122) );
  NANDN U37369 ( .A(n36120), .B(n36119), .Z(n36121) );
  AND U37370 ( .A(n36122), .B(n36121), .Z(n36140) );
  XNOR U37371 ( .A(n36141), .B(n36140), .Z(n36142) );
  NANDN U37372 ( .A(n36124), .B(n36123), .Z(n36128) );
  NAND U37373 ( .A(n36126), .B(n36125), .Z(n36127) );
  NAND U37374 ( .A(n36128), .B(n36127), .Z(n36143) );
  XNOR U37375 ( .A(n36142), .B(n36143), .Z(n36134) );
  XNOR U37376 ( .A(n36135), .B(n36134), .Z(n36136) );
  XNOR U37377 ( .A(n36137), .B(n36136), .Z(n36166) );
  XNOR U37378 ( .A(sreg[1882]), .B(n36166), .Z(n36168) );
  NANDN U37379 ( .A(sreg[1881]), .B(n36129), .Z(n36133) );
  NAND U37380 ( .A(n36131), .B(n36130), .Z(n36132) );
  NAND U37381 ( .A(n36133), .B(n36132), .Z(n36167) );
  XNOR U37382 ( .A(n36168), .B(n36167), .Z(c[1882]) );
  NANDN U37383 ( .A(n36135), .B(n36134), .Z(n36139) );
  NANDN U37384 ( .A(n36137), .B(n36136), .Z(n36138) );
  AND U37385 ( .A(n36139), .B(n36138), .Z(n36174) );
  NANDN U37386 ( .A(n36141), .B(n36140), .Z(n36145) );
  NANDN U37387 ( .A(n36143), .B(n36142), .Z(n36144) );
  AND U37388 ( .A(n36145), .B(n36144), .Z(n36172) );
  NAND U37389 ( .A(n42143), .B(n36146), .Z(n36148) );
  XNOR U37390 ( .A(a[861]), .B(n4194), .Z(n36183) );
  NAND U37391 ( .A(n42144), .B(n36183), .Z(n36147) );
  AND U37392 ( .A(n36148), .B(n36147), .Z(n36198) );
  XOR U37393 ( .A(a[865]), .B(n42012), .Z(n36186) );
  XNOR U37394 ( .A(n36198), .B(n36197), .Z(n36200) );
  AND U37395 ( .A(a[867]), .B(b[0]), .Z(n36150) );
  XNOR U37396 ( .A(n36150), .B(n4071), .Z(n36152) );
  NANDN U37397 ( .A(b[0]), .B(a[866]), .Z(n36151) );
  NAND U37398 ( .A(n36152), .B(n36151), .Z(n36194) );
  XOR U37399 ( .A(a[863]), .B(n42085), .Z(n36190) );
  AND U37400 ( .A(a[859]), .B(b[7]), .Z(n36191) );
  XNOR U37401 ( .A(n36192), .B(n36191), .Z(n36193) );
  XNOR U37402 ( .A(n36194), .B(n36193), .Z(n36199) );
  XOR U37403 ( .A(n36200), .B(n36199), .Z(n36178) );
  NANDN U37404 ( .A(n36155), .B(n36154), .Z(n36159) );
  NANDN U37405 ( .A(n36157), .B(n36156), .Z(n36158) );
  AND U37406 ( .A(n36159), .B(n36158), .Z(n36177) );
  XNOR U37407 ( .A(n36178), .B(n36177), .Z(n36179) );
  NANDN U37408 ( .A(n36161), .B(n36160), .Z(n36165) );
  NAND U37409 ( .A(n36163), .B(n36162), .Z(n36164) );
  NAND U37410 ( .A(n36165), .B(n36164), .Z(n36180) );
  XNOR U37411 ( .A(n36179), .B(n36180), .Z(n36171) );
  XNOR U37412 ( .A(n36172), .B(n36171), .Z(n36173) );
  XNOR U37413 ( .A(n36174), .B(n36173), .Z(n36203) );
  XNOR U37414 ( .A(sreg[1883]), .B(n36203), .Z(n36205) );
  NANDN U37415 ( .A(sreg[1882]), .B(n36166), .Z(n36170) );
  NAND U37416 ( .A(n36168), .B(n36167), .Z(n36169) );
  NAND U37417 ( .A(n36170), .B(n36169), .Z(n36204) );
  XNOR U37418 ( .A(n36205), .B(n36204), .Z(c[1883]) );
  NANDN U37419 ( .A(n36172), .B(n36171), .Z(n36176) );
  NANDN U37420 ( .A(n36174), .B(n36173), .Z(n36175) );
  AND U37421 ( .A(n36176), .B(n36175), .Z(n36211) );
  NANDN U37422 ( .A(n36178), .B(n36177), .Z(n36182) );
  NANDN U37423 ( .A(n36180), .B(n36179), .Z(n36181) );
  AND U37424 ( .A(n36182), .B(n36181), .Z(n36209) );
  NAND U37425 ( .A(n42143), .B(n36183), .Z(n36185) );
  XNOR U37426 ( .A(a[862]), .B(n4195), .Z(n36220) );
  NAND U37427 ( .A(n42144), .B(n36220), .Z(n36184) );
  AND U37428 ( .A(n36185), .B(n36184), .Z(n36235) );
  XOR U37429 ( .A(a[866]), .B(n42012), .Z(n36223) );
  XNOR U37430 ( .A(n36235), .B(n36234), .Z(n36237) );
  AND U37431 ( .A(a[868]), .B(b[0]), .Z(n36187) );
  XNOR U37432 ( .A(n36187), .B(n4071), .Z(n36189) );
  NANDN U37433 ( .A(b[0]), .B(a[867]), .Z(n36188) );
  NAND U37434 ( .A(n36189), .B(n36188), .Z(n36231) );
  XOR U37435 ( .A(a[864]), .B(n42085), .Z(n36224) );
  AND U37436 ( .A(a[860]), .B(b[7]), .Z(n36228) );
  XNOR U37437 ( .A(n36229), .B(n36228), .Z(n36230) );
  XNOR U37438 ( .A(n36231), .B(n36230), .Z(n36236) );
  XOR U37439 ( .A(n36237), .B(n36236), .Z(n36215) );
  NANDN U37440 ( .A(n36192), .B(n36191), .Z(n36196) );
  NANDN U37441 ( .A(n36194), .B(n36193), .Z(n36195) );
  AND U37442 ( .A(n36196), .B(n36195), .Z(n36214) );
  XNOR U37443 ( .A(n36215), .B(n36214), .Z(n36216) );
  NANDN U37444 ( .A(n36198), .B(n36197), .Z(n36202) );
  NAND U37445 ( .A(n36200), .B(n36199), .Z(n36201) );
  NAND U37446 ( .A(n36202), .B(n36201), .Z(n36217) );
  XNOR U37447 ( .A(n36216), .B(n36217), .Z(n36208) );
  XNOR U37448 ( .A(n36209), .B(n36208), .Z(n36210) );
  XNOR U37449 ( .A(n36211), .B(n36210), .Z(n36240) );
  XNOR U37450 ( .A(sreg[1884]), .B(n36240), .Z(n36242) );
  NANDN U37451 ( .A(sreg[1883]), .B(n36203), .Z(n36207) );
  NAND U37452 ( .A(n36205), .B(n36204), .Z(n36206) );
  NAND U37453 ( .A(n36207), .B(n36206), .Z(n36241) );
  XNOR U37454 ( .A(n36242), .B(n36241), .Z(c[1884]) );
  NANDN U37455 ( .A(n36209), .B(n36208), .Z(n36213) );
  NANDN U37456 ( .A(n36211), .B(n36210), .Z(n36212) );
  AND U37457 ( .A(n36213), .B(n36212), .Z(n36248) );
  NANDN U37458 ( .A(n36215), .B(n36214), .Z(n36219) );
  NANDN U37459 ( .A(n36217), .B(n36216), .Z(n36218) );
  AND U37460 ( .A(n36219), .B(n36218), .Z(n36246) );
  NAND U37461 ( .A(n42143), .B(n36220), .Z(n36222) );
  XNOR U37462 ( .A(a[863]), .B(n4195), .Z(n36257) );
  NAND U37463 ( .A(n42144), .B(n36257), .Z(n36221) );
  AND U37464 ( .A(n36222), .B(n36221), .Z(n36272) );
  XOR U37465 ( .A(a[867]), .B(n42012), .Z(n36260) );
  XNOR U37466 ( .A(n36272), .B(n36271), .Z(n36274) );
  XOR U37467 ( .A(a[865]), .B(n42085), .Z(n36261) );
  AND U37468 ( .A(a[861]), .B(b[7]), .Z(n36265) );
  XNOR U37469 ( .A(n36266), .B(n36265), .Z(n36267) );
  AND U37470 ( .A(a[869]), .B(b[0]), .Z(n36225) );
  XNOR U37471 ( .A(n36225), .B(n4071), .Z(n36227) );
  NANDN U37472 ( .A(b[0]), .B(a[868]), .Z(n36226) );
  NAND U37473 ( .A(n36227), .B(n36226), .Z(n36268) );
  XNOR U37474 ( .A(n36267), .B(n36268), .Z(n36273) );
  XOR U37475 ( .A(n36274), .B(n36273), .Z(n36252) );
  NANDN U37476 ( .A(n36229), .B(n36228), .Z(n36233) );
  NANDN U37477 ( .A(n36231), .B(n36230), .Z(n36232) );
  AND U37478 ( .A(n36233), .B(n36232), .Z(n36251) );
  XNOR U37479 ( .A(n36252), .B(n36251), .Z(n36253) );
  NANDN U37480 ( .A(n36235), .B(n36234), .Z(n36239) );
  NAND U37481 ( .A(n36237), .B(n36236), .Z(n36238) );
  NAND U37482 ( .A(n36239), .B(n36238), .Z(n36254) );
  XNOR U37483 ( .A(n36253), .B(n36254), .Z(n36245) );
  XNOR U37484 ( .A(n36246), .B(n36245), .Z(n36247) );
  XNOR U37485 ( .A(n36248), .B(n36247), .Z(n36277) );
  XNOR U37486 ( .A(sreg[1885]), .B(n36277), .Z(n36279) );
  NANDN U37487 ( .A(sreg[1884]), .B(n36240), .Z(n36244) );
  NAND U37488 ( .A(n36242), .B(n36241), .Z(n36243) );
  NAND U37489 ( .A(n36244), .B(n36243), .Z(n36278) );
  XNOR U37490 ( .A(n36279), .B(n36278), .Z(c[1885]) );
  NANDN U37491 ( .A(n36246), .B(n36245), .Z(n36250) );
  NANDN U37492 ( .A(n36248), .B(n36247), .Z(n36249) );
  AND U37493 ( .A(n36250), .B(n36249), .Z(n36289) );
  NANDN U37494 ( .A(n36252), .B(n36251), .Z(n36256) );
  NANDN U37495 ( .A(n36254), .B(n36253), .Z(n36255) );
  AND U37496 ( .A(n36256), .B(n36255), .Z(n36288) );
  NAND U37497 ( .A(n42143), .B(n36257), .Z(n36259) );
  XNOR U37498 ( .A(a[864]), .B(n4195), .Z(n36299) );
  NAND U37499 ( .A(n42144), .B(n36299), .Z(n36258) );
  AND U37500 ( .A(n36259), .B(n36258), .Z(n36314) );
  XOR U37501 ( .A(a[868]), .B(n42012), .Z(n36302) );
  XNOR U37502 ( .A(n36314), .B(n36313), .Z(n36316) );
  XOR U37503 ( .A(a[866]), .B(n42085), .Z(n36306) );
  AND U37504 ( .A(a[862]), .B(b[7]), .Z(n36307) );
  XNOR U37505 ( .A(n36308), .B(n36307), .Z(n36309) );
  AND U37506 ( .A(a[870]), .B(b[0]), .Z(n36262) );
  XNOR U37507 ( .A(n36262), .B(n4071), .Z(n36264) );
  NANDN U37508 ( .A(b[0]), .B(a[869]), .Z(n36263) );
  NAND U37509 ( .A(n36264), .B(n36263), .Z(n36310) );
  XNOR U37510 ( .A(n36309), .B(n36310), .Z(n36315) );
  XOR U37511 ( .A(n36316), .B(n36315), .Z(n36294) );
  NANDN U37512 ( .A(n36266), .B(n36265), .Z(n36270) );
  NANDN U37513 ( .A(n36268), .B(n36267), .Z(n36269) );
  AND U37514 ( .A(n36270), .B(n36269), .Z(n36293) );
  XNOR U37515 ( .A(n36294), .B(n36293), .Z(n36295) );
  NANDN U37516 ( .A(n36272), .B(n36271), .Z(n36276) );
  NAND U37517 ( .A(n36274), .B(n36273), .Z(n36275) );
  NAND U37518 ( .A(n36276), .B(n36275), .Z(n36296) );
  XNOR U37519 ( .A(n36295), .B(n36296), .Z(n36287) );
  XOR U37520 ( .A(n36288), .B(n36287), .Z(n36290) );
  XOR U37521 ( .A(n36289), .B(n36290), .Z(n36282) );
  XNOR U37522 ( .A(n36282), .B(sreg[1886]), .Z(n36284) );
  NANDN U37523 ( .A(sreg[1885]), .B(n36277), .Z(n36281) );
  NAND U37524 ( .A(n36279), .B(n36278), .Z(n36280) );
  AND U37525 ( .A(n36281), .B(n36280), .Z(n36283) );
  XOR U37526 ( .A(n36284), .B(n36283), .Z(c[1886]) );
  NANDN U37527 ( .A(n36282), .B(sreg[1886]), .Z(n36286) );
  NAND U37528 ( .A(n36284), .B(n36283), .Z(n36285) );
  AND U37529 ( .A(n36286), .B(n36285), .Z(n36353) );
  NANDN U37530 ( .A(n36288), .B(n36287), .Z(n36292) );
  OR U37531 ( .A(n36290), .B(n36289), .Z(n36291) );
  AND U37532 ( .A(n36292), .B(n36291), .Z(n36322) );
  NANDN U37533 ( .A(n36294), .B(n36293), .Z(n36298) );
  NANDN U37534 ( .A(n36296), .B(n36295), .Z(n36297) );
  AND U37535 ( .A(n36298), .B(n36297), .Z(n36320) );
  NAND U37536 ( .A(n42143), .B(n36299), .Z(n36301) );
  XNOR U37537 ( .A(a[865]), .B(n4195), .Z(n36331) );
  NAND U37538 ( .A(n42144), .B(n36331), .Z(n36300) );
  AND U37539 ( .A(n36301), .B(n36300), .Z(n36346) );
  XOR U37540 ( .A(a[869]), .B(n42012), .Z(n36334) );
  XNOR U37541 ( .A(n36346), .B(n36345), .Z(n36348) );
  AND U37542 ( .A(a[871]), .B(b[0]), .Z(n36303) );
  XNOR U37543 ( .A(n36303), .B(n4071), .Z(n36305) );
  NANDN U37544 ( .A(b[0]), .B(a[870]), .Z(n36304) );
  NAND U37545 ( .A(n36305), .B(n36304), .Z(n36342) );
  XOR U37546 ( .A(a[867]), .B(n42085), .Z(n36335) );
  AND U37547 ( .A(a[863]), .B(b[7]), .Z(n36339) );
  XNOR U37548 ( .A(n36340), .B(n36339), .Z(n36341) );
  XNOR U37549 ( .A(n36342), .B(n36341), .Z(n36347) );
  XOR U37550 ( .A(n36348), .B(n36347), .Z(n36326) );
  NANDN U37551 ( .A(n36308), .B(n36307), .Z(n36312) );
  NANDN U37552 ( .A(n36310), .B(n36309), .Z(n36311) );
  AND U37553 ( .A(n36312), .B(n36311), .Z(n36325) );
  XNOR U37554 ( .A(n36326), .B(n36325), .Z(n36327) );
  NANDN U37555 ( .A(n36314), .B(n36313), .Z(n36318) );
  NAND U37556 ( .A(n36316), .B(n36315), .Z(n36317) );
  NAND U37557 ( .A(n36318), .B(n36317), .Z(n36328) );
  XNOR U37558 ( .A(n36327), .B(n36328), .Z(n36319) );
  XNOR U37559 ( .A(n36320), .B(n36319), .Z(n36321) );
  XNOR U37560 ( .A(n36322), .B(n36321), .Z(n36351) );
  XNOR U37561 ( .A(sreg[1887]), .B(n36351), .Z(n36352) );
  XNOR U37562 ( .A(n36353), .B(n36352), .Z(c[1887]) );
  NANDN U37563 ( .A(n36320), .B(n36319), .Z(n36324) );
  NANDN U37564 ( .A(n36322), .B(n36321), .Z(n36323) );
  AND U37565 ( .A(n36324), .B(n36323), .Z(n36359) );
  NANDN U37566 ( .A(n36326), .B(n36325), .Z(n36330) );
  NANDN U37567 ( .A(n36328), .B(n36327), .Z(n36329) );
  AND U37568 ( .A(n36330), .B(n36329), .Z(n36357) );
  NAND U37569 ( .A(n42143), .B(n36331), .Z(n36333) );
  XNOR U37570 ( .A(a[866]), .B(n4195), .Z(n36368) );
  NAND U37571 ( .A(n42144), .B(n36368), .Z(n36332) );
  AND U37572 ( .A(n36333), .B(n36332), .Z(n36383) );
  XOR U37573 ( .A(a[870]), .B(n42012), .Z(n36371) );
  XNOR U37574 ( .A(n36383), .B(n36382), .Z(n36385) );
  XOR U37575 ( .A(a[868]), .B(n42085), .Z(n36372) );
  AND U37576 ( .A(a[864]), .B(b[7]), .Z(n36376) );
  XNOR U37577 ( .A(n36377), .B(n36376), .Z(n36378) );
  AND U37578 ( .A(a[872]), .B(b[0]), .Z(n36336) );
  XNOR U37579 ( .A(n36336), .B(n4071), .Z(n36338) );
  NANDN U37580 ( .A(b[0]), .B(a[871]), .Z(n36337) );
  NAND U37581 ( .A(n36338), .B(n36337), .Z(n36379) );
  XNOR U37582 ( .A(n36378), .B(n36379), .Z(n36384) );
  XOR U37583 ( .A(n36385), .B(n36384), .Z(n36363) );
  NANDN U37584 ( .A(n36340), .B(n36339), .Z(n36344) );
  NANDN U37585 ( .A(n36342), .B(n36341), .Z(n36343) );
  AND U37586 ( .A(n36344), .B(n36343), .Z(n36362) );
  XNOR U37587 ( .A(n36363), .B(n36362), .Z(n36364) );
  NANDN U37588 ( .A(n36346), .B(n36345), .Z(n36350) );
  NAND U37589 ( .A(n36348), .B(n36347), .Z(n36349) );
  NAND U37590 ( .A(n36350), .B(n36349), .Z(n36365) );
  XNOR U37591 ( .A(n36364), .B(n36365), .Z(n36356) );
  XNOR U37592 ( .A(n36357), .B(n36356), .Z(n36358) );
  XNOR U37593 ( .A(n36359), .B(n36358), .Z(n36388) );
  XNOR U37594 ( .A(sreg[1888]), .B(n36388), .Z(n36390) );
  NANDN U37595 ( .A(sreg[1887]), .B(n36351), .Z(n36355) );
  NAND U37596 ( .A(n36353), .B(n36352), .Z(n36354) );
  NAND U37597 ( .A(n36355), .B(n36354), .Z(n36389) );
  XNOR U37598 ( .A(n36390), .B(n36389), .Z(c[1888]) );
  NANDN U37599 ( .A(n36357), .B(n36356), .Z(n36361) );
  NANDN U37600 ( .A(n36359), .B(n36358), .Z(n36360) );
  AND U37601 ( .A(n36361), .B(n36360), .Z(n36396) );
  NANDN U37602 ( .A(n36363), .B(n36362), .Z(n36367) );
  NANDN U37603 ( .A(n36365), .B(n36364), .Z(n36366) );
  AND U37604 ( .A(n36367), .B(n36366), .Z(n36394) );
  NAND U37605 ( .A(n42143), .B(n36368), .Z(n36370) );
  XNOR U37606 ( .A(a[867]), .B(n4195), .Z(n36405) );
  NAND U37607 ( .A(n42144), .B(n36405), .Z(n36369) );
  AND U37608 ( .A(n36370), .B(n36369), .Z(n36420) );
  XOR U37609 ( .A(a[871]), .B(n42012), .Z(n36408) );
  XNOR U37610 ( .A(n36420), .B(n36419), .Z(n36422) );
  XOR U37611 ( .A(a[869]), .B(n42085), .Z(n36412) );
  AND U37612 ( .A(a[865]), .B(b[7]), .Z(n36413) );
  XNOR U37613 ( .A(n36414), .B(n36413), .Z(n36415) );
  AND U37614 ( .A(a[873]), .B(b[0]), .Z(n36373) );
  XNOR U37615 ( .A(n36373), .B(n4071), .Z(n36375) );
  NANDN U37616 ( .A(b[0]), .B(a[872]), .Z(n36374) );
  NAND U37617 ( .A(n36375), .B(n36374), .Z(n36416) );
  XNOR U37618 ( .A(n36415), .B(n36416), .Z(n36421) );
  XOR U37619 ( .A(n36422), .B(n36421), .Z(n36400) );
  NANDN U37620 ( .A(n36377), .B(n36376), .Z(n36381) );
  NANDN U37621 ( .A(n36379), .B(n36378), .Z(n36380) );
  AND U37622 ( .A(n36381), .B(n36380), .Z(n36399) );
  XNOR U37623 ( .A(n36400), .B(n36399), .Z(n36401) );
  NANDN U37624 ( .A(n36383), .B(n36382), .Z(n36387) );
  NAND U37625 ( .A(n36385), .B(n36384), .Z(n36386) );
  NAND U37626 ( .A(n36387), .B(n36386), .Z(n36402) );
  XNOR U37627 ( .A(n36401), .B(n36402), .Z(n36393) );
  XNOR U37628 ( .A(n36394), .B(n36393), .Z(n36395) );
  XNOR U37629 ( .A(n36396), .B(n36395), .Z(n36425) );
  XNOR U37630 ( .A(sreg[1889]), .B(n36425), .Z(n36427) );
  NANDN U37631 ( .A(sreg[1888]), .B(n36388), .Z(n36392) );
  NAND U37632 ( .A(n36390), .B(n36389), .Z(n36391) );
  NAND U37633 ( .A(n36392), .B(n36391), .Z(n36426) );
  XNOR U37634 ( .A(n36427), .B(n36426), .Z(c[1889]) );
  NANDN U37635 ( .A(n36394), .B(n36393), .Z(n36398) );
  NANDN U37636 ( .A(n36396), .B(n36395), .Z(n36397) );
  AND U37637 ( .A(n36398), .B(n36397), .Z(n36433) );
  NANDN U37638 ( .A(n36400), .B(n36399), .Z(n36404) );
  NANDN U37639 ( .A(n36402), .B(n36401), .Z(n36403) );
  AND U37640 ( .A(n36404), .B(n36403), .Z(n36431) );
  NAND U37641 ( .A(n42143), .B(n36405), .Z(n36407) );
  XNOR U37642 ( .A(a[868]), .B(n4195), .Z(n36442) );
  NAND U37643 ( .A(n42144), .B(n36442), .Z(n36406) );
  AND U37644 ( .A(n36407), .B(n36406), .Z(n36457) );
  XOR U37645 ( .A(a[872]), .B(n42012), .Z(n36445) );
  XNOR U37646 ( .A(n36457), .B(n36456), .Z(n36459) );
  AND U37647 ( .A(a[874]), .B(b[0]), .Z(n36409) );
  XNOR U37648 ( .A(n36409), .B(n4071), .Z(n36411) );
  NANDN U37649 ( .A(b[0]), .B(a[873]), .Z(n36410) );
  NAND U37650 ( .A(n36411), .B(n36410), .Z(n36453) );
  XOR U37651 ( .A(a[870]), .B(n42085), .Z(n36449) );
  AND U37652 ( .A(a[866]), .B(b[7]), .Z(n36450) );
  XNOR U37653 ( .A(n36451), .B(n36450), .Z(n36452) );
  XNOR U37654 ( .A(n36453), .B(n36452), .Z(n36458) );
  XOR U37655 ( .A(n36459), .B(n36458), .Z(n36437) );
  NANDN U37656 ( .A(n36414), .B(n36413), .Z(n36418) );
  NANDN U37657 ( .A(n36416), .B(n36415), .Z(n36417) );
  AND U37658 ( .A(n36418), .B(n36417), .Z(n36436) );
  XNOR U37659 ( .A(n36437), .B(n36436), .Z(n36438) );
  NANDN U37660 ( .A(n36420), .B(n36419), .Z(n36424) );
  NAND U37661 ( .A(n36422), .B(n36421), .Z(n36423) );
  NAND U37662 ( .A(n36424), .B(n36423), .Z(n36439) );
  XNOR U37663 ( .A(n36438), .B(n36439), .Z(n36430) );
  XNOR U37664 ( .A(n36431), .B(n36430), .Z(n36432) );
  XNOR U37665 ( .A(n36433), .B(n36432), .Z(n36462) );
  XNOR U37666 ( .A(sreg[1890]), .B(n36462), .Z(n36464) );
  NANDN U37667 ( .A(sreg[1889]), .B(n36425), .Z(n36429) );
  NAND U37668 ( .A(n36427), .B(n36426), .Z(n36428) );
  NAND U37669 ( .A(n36429), .B(n36428), .Z(n36463) );
  XNOR U37670 ( .A(n36464), .B(n36463), .Z(c[1890]) );
  NANDN U37671 ( .A(n36431), .B(n36430), .Z(n36435) );
  NANDN U37672 ( .A(n36433), .B(n36432), .Z(n36434) );
  AND U37673 ( .A(n36435), .B(n36434), .Z(n36470) );
  NANDN U37674 ( .A(n36437), .B(n36436), .Z(n36441) );
  NANDN U37675 ( .A(n36439), .B(n36438), .Z(n36440) );
  AND U37676 ( .A(n36441), .B(n36440), .Z(n36468) );
  NAND U37677 ( .A(n42143), .B(n36442), .Z(n36444) );
  XNOR U37678 ( .A(a[869]), .B(n4196), .Z(n36479) );
  NAND U37679 ( .A(n42144), .B(n36479), .Z(n36443) );
  AND U37680 ( .A(n36444), .B(n36443), .Z(n36494) );
  XOR U37681 ( .A(a[873]), .B(n42012), .Z(n36482) );
  XNOR U37682 ( .A(n36494), .B(n36493), .Z(n36496) );
  AND U37683 ( .A(a[875]), .B(b[0]), .Z(n36446) );
  XNOR U37684 ( .A(n36446), .B(n4071), .Z(n36448) );
  NANDN U37685 ( .A(b[0]), .B(a[874]), .Z(n36447) );
  NAND U37686 ( .A(n36448), .B(n36447), .Z(n36490) );
  XOR U37687 ( .A(a[871]), .B(n42085), .Z(n36486) );
  AND U37688 ( .A(a[867]), .B(b[7]), .Z(n36487) );
  XNOR U37689 ( .A(n36488), .B(n36487), .Z(n36489) );
  XNOR U37690 ( .A(n36490), .B(n36489), .Z(n36495) );
  XOR U37691 ( .A(n36496), .B(n36495), .Z(n36474) );
  NANDN U37692 ( .A(n36451), .B(n36450), .Z(n36455) );
  NANDN U37693 ( .A(n36453), .B(n36452), .Z(n36454) );
  AND U37694 ( .A(n36455), .B(n36454), .Z(n36473) );
  XNOR U37695 ( .A(n36474), .B(n36473), .Z(n36475) );
  NANDN U37696 ( .A(n36457), .B(n36456), .Z(n36461) );
  NAND U37697 ( .A(n36459), .B(n36458), .Z(n36460) );
  NAND U37698 ( .A(n36461), .B(n36460), .Z(n36476) );
  XNOR U37699 ( .A(n36475), .B(n36476), .Z(n36467) );
  XNOR U37700 ( .A(n36468), .B(n36467), .Z(n36469) );
  XNOR U37701 ( .A(n36470), .B(n36469), .Z(n36499) );
  XNOR U37702 ( .A(sreg[1891]), .B(n36499), .Z(n36501) );
  NANDN U37703 ( .A(sreg[1890]), .B(n36462), .Z(n36466) );
  NAND U37704 ( .A(n36464), .B(n36463), .Z(n36465) );
  NAND U37705 ( .A(n36466), .B(n36465), .Z(n36500) );
  XNOR U37706 ( .A(n36501), .B(n36500), .Z(c[1891]) );
  NANDN U37707 ( .A(n36468), .B(n36467), .Z(n36472) );
  NANDN U37708 ( .A(n36470), .B(n36469), .Z(n36471) );
  AND U37709 ( .A(n36472), .B(n36471), .Z(n36507) );
  NANDN U37710 ( .A(n36474), .B(n36473), .Z(n36478) );
  NANDN U37711 ( .A(n36476), .B(n36475), .Z(n36477) );
  AND U37712 ( .A(n36478), .B(n36477), .Z(n36505) );
  NAND U37713 ( .A(n42143), .B(n36479), .Z(n36481) );
  XNOR U37714 ( .A(a[870]), .B(n4196), .Z(n36516) );
  NAND U37715 ( .A(n42144), .B(n36516), .Z(n36480) );
  AND U37716 ( .A(n36481), .B(n36480), .Z(n36531) );
  XOR U37717 ( .A(a[874]), .B(n42012), .Z(n36519) );
  XNOR U37718 ( .A(n36531), .B(n36530), .Z(n36533) );
  AND U37719 ( .A(a[876]), .B(b[0]), .Z(n36483) );
  XNOR U37720 ( .A(n36483), .B(n4071), .Z(n36485) );
  NANDN U37721 ( .A(b[0]), .B(a[875]), .Z(n36484) );
  NAND U37722 ( .A(n36485), .B(n36484), .Z(n36527) );
  XOR U37723 ( .A(a[872]), .B(n42085), .Z(n36523) );
  AND U37724 ( .A(a[868]), .B(b[7]), .Z(n36524) );
  XNOR U37725 ( .A(n36525), .B(n36524), .Z(n36526) );
  XNOR U37726 ( .A(n36527), .B(n36526), .Z(n36532) );
  XOR U37727 ( .A(n36533), .B(n36532), .Z(n36511) );
  NANDN U37728 ( .A(n36488), .B(n36487), .Z(n36492) );
  NANDN U37729 ( .A(n36490), .B(n36489), .Z(n36491) );
  AND U37730 ( .A(n36492), .B(n36491), .Z(n36510) );
  XNOR U37731 ( .A(n36511), .B(n36510), .Z(n36512) );
  NANDN U37732 ( .A(n36494), .B(n36493), .Z(n36498) );
  NAND U37733 ( .A(n36496), .B(n36495), .Z(n36497) );
  NAND U37734 ( .A(n36498), .B(n36497), .Z(n36513) );
  XNOR U37735 ( .A(n36512), .B(n36513), .Z(n36504) );
  XNOR U37736 ( .A(n36505), .B(n36504), .Z(n36506) );
  XNOR U37737 ( .A(n36507), .B(n36506), .Z(n36536) );
  XNOR U37738 ( .A(sreg[1892]), .B(n36536), .Z(n36538) );
  NANDN U37739 ( .A(sreg[1891]), .B(n36499), .Z(n36503) );
  NAND U37740 ( .A(n36501), .B(n36500), .Z(n36502) );
  NAND U37741 ( .A(n36503), .B(n36502), .Z(n36537) );
  XNOR U37742 ( .A(n36538), .B(n36537), .Z(c[1892]) );
  NANDN U37743 ( .A(n36505), .B(n36504), .Z(n36509) );
  NANDN U37744 ( .A(n36507), .B(n36506), .Z(n36508) );
  AND U37745 ( .A(n36509), .B(n36508), .Z(n36544) );
  NANDN U37746 ( .A(n36511), .B(n36510), .Z(n36515) );
  NANDN U37747 ( .A(n36513), .B(n36512), .Z(n36514) );
  AND U37748 ( .A(n36515), .B(n36514), .Z(n36542) );
  NAND U37749 ( .A(n42143), .B(n36516), .Z(n36518) );
  XNOR U37750 ( .A(a[871]), .B(n4196), .Z(n36553) );
  NAND U37751 ( .A(n42144), .B(n36553), .Z(n36517) );
  AND U37752 ( .A(n36518), .B(n36517), .Z(n36568) );
  XOR U37753 ( .A(a[875]), .B(n42012), .Z(n36556) );
  XNOR U37754 ( .A(n36568), .B(n36567), .Z(n36570) );
  AND U37755 ( .A(a[877]), .B(b[0]), .Z(n36520) );
  XNOR U37756 ( .A(n36520), .B(n4071), .Z(n36522) );
  NANDN U37757 ( .A(b[0]), .B(a[876]), .Z(n36521) );
  NAND U37758 ( .A(n36522), .B(n36521), .Z(n36564) );
  XOR U37759 ( .A(a[873]), .B(n42085), .Z(n36560) );
  AND U37760 ( .A(a[869]), .B(b[7]), .Z(n36561) );
  XNOR U37761 ( .A(n36562), .B(n36561), .Z(n36563) );
  XNOR U37762 ( .A(n36564), .B(n36563), .Z(n36569) );
  XOR U37763 ( .A(n36570), .B(n36569), .Z(n36548) );
  NANDN U37764 ( .A(n36525), .B(n36524), .Z(n36529) );
  NANDN U37765 ( .A(n36527), .B(n36526), .Z(n36528) );
  AND U37766 ( .A(n36529), .B(n36528), .Z(n36547) );
  XNOR U37767 ( .A(n36548), .B(n36547), .Z(n36549) );
  NANDN U37768 ( .A(n36531), .B(n36530), .Z(n36535) );
  NAND U37769 ( .A(n36533), .B(n36532), .Z(n36534) );
  NAND U37770 ( .A(n36535), .B(n36534), .Z(n36550) );
  XNOR U37771 ( .A(n36549), .B(n36550), .Z(n36541) );
  XNOR U37772 ( .A(n36542), .B(n36541), .Z(n36543) );
  XNOR U37773 ( .A(n36544), .B(n36543), .Z(n36573) );
  XNOR U37774 ( .A(sreg[1893]), .B(n36573), .Z(n36575) );
  NANDN U37775 ( .A(sreg[1892]), .B(n36536), .Z(n36540) );
  NAND U37776 ( .A(n36538), .B(n36537), .Z(n36539) );
  NAND U37777 ( .A(n36540), .B(n36539), .Z(n36574) );
  XNOR U37778 ( .A(n36575), .B(n36574), .Z(c[1893]) );
  NANDN U37779 ( .A(n36542), .B(n36541), .Z(n36546) );
  NANDN U37780 ( .A(n36544), .B(n36543), .Z(n36545) );
  AND U37781 ( .A(n36546), .B(n36545), .Z(n36581) );
  NANDN U37782 ( .A(n36548), .B(n36547), .Z(n36552) );
  NANDN U37783 ( .A(n36550), .B(n36549), .Z(n36551) );
  AND U37784 ( .A(n36552), .B(n36551), .Z(n36579) );
  NAND U37785 ( .A(n42143), .B(n36553), .Z(n36555) );
  XNOR U37786 ( .A(a[872]), .B(n4196), .Z(n36590) );
  NAND U37787 ( .A(n42144), .B(n36590), .Z(n36554) );
  AND U37788 ( .A(n36555), .B(n36554), .Z(n36605) );
  XOR U37789 ( .A(a[876]), .B(n42012), .Z(n36593) );
  XNOR U37790 ( .A(n36605), .B(n36604), .Z(n36607) );
  AND U37791 ( .A(a[878]), .B(b[0]), .Z(n36557) );
  XNOR U37792 ( .A(n36557), .B(n4071), .Z(n36559) );
  NANDN U37793 ( .A(b[0]), .B(a[877]), .Z(n36558) );
  NAND U37794 ( .A(n36559), .B(n36558), .Z(n36601) );
  XOR U37795 ( .A(a[874]), .B(n42085), .Z(n36597) );
  AND U37796 ( .A(a[870]), .B(b[7]), .Z(n36598) );
  XNOR U37797 ( .A(n36599), .B(n36598), .Z(n36600) );
  XNOR U37798 ( .A(n36601), .B(n36600), .Z(n36606) );
  XOR U37799 ( .A(n36607), .B(n36606), .Z(n36585) );
  NANDN U37800 ( .A(n36562), .B(n36561), .Z(n36566) );
  NANDN U37801 ( .A(n36564), .B(n36563), .Z(n36565) );
  AND U37802 ( .A(n36566), .B(n36565), .Z(n36584) );
  XNOR U37803 ( .A(n36585), .B(n36584), .Z(n36586) );
  NANDN U37804 ( .A(n36568), .B(n36567), .Z(n36572) );
  NAND U37805 ( .A(n36570), .B(n36569), .Z(n36571) );
  NAND U37806 ( .A(n36572), .B(n36571), .Z(n36587) );
  XNOR U37807 ( .A(n36586), .B(n36587), .Z(n36578) );
  XNOR U37808 ( .A(n36579), .B(n36578), .Z(n36580) );
  XNOR U37809 ( .A(n36581), .B(n36580), .Z(n36610) );
  XNOR U37810 ( .A(sreg[1894]), .B(n36610), .Z(n36612) );
  NANDN U37811 ( .A(sreg[1893]), .B(n36573), .Z(n36577) );
  NAND U37812 ( .A(n36575), .B(n36574), .Z(n36576) );
  NAND U37813 ( .A(n36577), .B(n36576), .Z(n36611) );
  XNOR U37814 ( .A(n36612), .B(n36611), .Z(c[1894]) );
  NANDN U37815 ( .A(n36579), .B(n36578), .Z(n36583) );
  NANDN U37816 ( .A(n36581), .B(n36580), .Z(n36582) );
  AND U37817 ( .A(n36583), .B(n36582), .Z(n36618) );
  NANDN U37818 ( .A(n36585), .B(n36584), .Z(n36589) );
  NANDN U37819 ( .A(n36587), .B(n36586), .Z(n36588) );
  AND U37820 ( .A(n36589), .B(n36588), .Z(n36616) );
  NAND U37821 ( .A(n42143), .B(n36590), .Z(n36592) );
  XNOR U37822 ( .A(a[873]), .B(n4196), .Z(n36627) );
  NAND U37823 ( .A(n42144), .B(n36627), .Z(n36591) );
  AND U37824 ( .A(n36592), .B(n36591), .Z(n36642) );
  XOR U37825 ( .A(a[877]), .B(n42012), .Z(n36630) );
  XNOR U37826 ( .A(n36642), .B(n36641), .Z(n36644) );
  AND U37827 ( .A(a[879]), .B(b[0]), .Z(n36594) );
  XNOR U37828 ( .A(n36594), .B(n4071), .Z(n36596) );
  NANDN U37829 ( .A(b[0]), .B(a[878]), .Z(n36595) );
  NAND U37830 ( .A(n36596), .B(n36595), .Z(n36638) );
  XOR U37831 ( .A(a[875]), .B(n42085), .Z(n36631) );
  AND U37832 ( .A(a[871]), .B(b[7]), .Z(n36635) );
  XNOR U37833 ( .A(n36636), .B(n36635), .Z(n36637) );
  XNOR U37834 ( .A(n36638), .B(n36637), .Z(n36643) );
  XOR U37835 ( .A(n36644), .B(n36643), .Z(n36622) );
  NANDN U37836 ( .A(n36599), .B(n36598), .Z(n36603) );
  NANDN U37837 ( .A(n36601), .B(n36600), .Z(n36602) );
  AND U37838 ( .A(n36603), .B(n36602), .Z(n36621) );
  XNOR U37839 ( .A(n36622), .B(n36621), .Z(n36623) );
  NANDN U37840 ( .A(n36605), .B(n36604), .Z(n36609) );
  NAND U37841 ( .A(n36607), .B(n36606), .Z(n36608) );
  NAND U37842 ( .A(n36609), .B(n36608), .Z(n36624) );
  XNOR U37843 ( .A(n36623), .B(n36624), .Z(n36615) );
  XNOR U37844 ( .A(n36616), .B(n36615), .Z(n36617) );
  XNOR U37845 ( .A(n36618), .B(n36617), .Z(n36647) );
  XNOR U37846 ( .A(sreg[1895]), .B(n36647), .Z(n36649) );
  NANDN U37847 ( .A(sreg[1894]), .B(n36610), .Z(n36614) );
  NAND U37848 ( .A(n36612), .B(n36611), .Z(n36613) );
  NAND U37849 ( .A(n36614), .B(n36613), .Z(n36648) );
  XNOR U37850 ( .A(n36649), .B(n36648), .Z(c[1895]) );
  NANDN U37851 ( .A(n36616), .B(n36615), .Z(n36620) );
  NANDN U37852 ( .A(n36618), .B(n36617), .Z(n36619) );
  AND U37853 ( .A(n36620), .B(n36619), .Z(n36655) );
  NANDN U37854 ( .A(n36622), .B(n36621), .Z(n36626) );
  NANDN U37855 ( .A(n36624), .B(n36623), .Z(n36625) );
  AND U37856 ( .A(n36626), .B(n36625), .Z(n36653) );
  NAND U37857 ( .A(n42143), .B(n36627), .Z(n36629) );
  XNOR U37858 ( .A(a[874]), .B(n4196), .Z(n36664) );
  NAND U37859 ( .A(n42144), .B(n36664), .Z(n36628) );
  AND U37860 ( .A(n36629), .B(n36628), .Z(n36679) );
  XOR U37861 ( .A(a[878]), .B(n42012), .Z(n36667) );
  XNOR U37862 ( .A(n36679), .B(n36678), .Z(n36681) );
  XOR U37863 ( .A(a[876]), .B(n42085), .Z(n36671) );
  AND U37864 ( .A(a[872]), .B(b[7]), .Z(n36672) );
  XNOR U37865 ( .A(n36673), .B(n36672), .Z(n36674) );
  AND U37866 ( .A(a[880]), .B(b[0]), .Z(n36632) );
  XNOR U37867 ( .A(n36632), .B(n4071), .Z(n36634) );
  NANDN U37868 ( .A(b[0]), .B(a[879]), .Z(n36633) );
  NAND U37869 ( .A(n36634), .B(n36633), .Z(n36675) );
  XNOR U37870 ( .A(n36674), .B(n36675), .Z(n36680) );
  XOR U37871 ( .A(n36681), .B(n36680), .Z(n36659) );
  NANDN U37872 ( .A(n36636), .B(n36635), .Z(n36640) );
  NANDN U37873 ( .A(n36638), .B(n36637), .Z(n36639) );
  AND U37874 ( .A(n36640), .B(n36639), .Z(n36658) );
  XNOR U37875 ( .A(n36659), .B(n36658), .Z(n36660) );
  NANDN U37876 ( .A(n36642), .B(n36641), .Z(n36646) );
  NAND U37877 ( .A(n36644), .B(n36643), .Z(n36645) );
  NAND U37878 ( .A(n36646), .B(n36645), .Z(n36661) );
  XNOR U37879 ( .A(n36660), .B(n36661), .Z(n36652) );
  XNOR U37880 ( .A(n36653), .B(n36652), .Z(n36654) );
  XNOR U37881 ( .A(n36655), .B(n36654), .Z(n36684) );
  XNOR U37882 ( .A(sreg[1896]), .B(n36684), .Z(n36686) );
  NANDN U37883 ( .A(sreg[1895]), .B(n36647), .Z(n36651) );
  NAND U37884 ( .A(n36649), .B(n36648), .Z(n36650) );
  NAND U37885 ( .A(n36651), .B(n36650), .Z(n36685) );
  XNOR U37886 ( .A(n36686), .B(n36685), .Z(c[1896]) );
  NANDN U37887 ( .A(n36653), .B(n36652), .Z(n36657) );
  NANDN U37888 ( .A(n36655), .B(n36654), .Z(n36656) );
  AND U37889 ( .A(n36657), .B(n36656), .Z(n36692) );
  NANDN U37890 ( .A(n36659), .B(n36658), .Z(n36663) );
  NANDN U37891 ( .A(n36661), .B(n36660), .Z(n36662) );
  AND U37892 ( .A(n36663), .B(n36662), .Z(n36690) );
  NAND U37893 ( .A(n42143), .B(n36664), .Z(n36666) );
  XNOR U37894 ( .A(a[875]), .B(n4196), .Z(n36701) );
  NAND U37895 ( .A(n42144), .B(n36701), .Z(n36665) );
  AND U37896 ( .A(n36666), .B(n36665), .Z(n36716) );
  XOR U37897 ( .A(a[879]), .B(n42012), .Z(n36704) );
  XNOR U37898 ( .A(n36716), .B(n36715), .Z(n36718) );
  AND U37899 ( .A(a[881]), .B(b[0]), .Z(n36668) );
  XNOR U37900 ( .A(n36668), .B(n4071), .Z(n36670) );
  NANDN U37901 ( .A(b[0]), .B(a[880]), .Z(n36669) );
  NAND U37902 ( .A(n36670), .B(n36669), .Z(n36712) );
  XOR U37903 ( .A(a[877]), .B(n42085), .Z(n36708) );
  AND U37904 ( .A(a[873]), .B(b[7]), .Z(n36709) );
  XNOR U37905 ( .A(n36710), .B(n36709), .Z(n36711) );
  XNOR U37906 ( .A(n36712), .B(n36711), .Z(n36717) );
  XOR U37907 ( .A(n36718), .B(n36717), .Z(n36696) );
  NANDN U37908 ( .A(n36673), .B(n36672), .Z(n36677) );
  NANDN U37909 ( .A(n36675), .B(n36674), .Z(n36676) );
  AND U37910 ( .A(n36677), .B(n36676), .Z(n36695) );
  XNOR U37911 ( .A(n36696), .B(n36695), .Z(n36697) );
  NANDN U37912 ( .A(n36679), .B(n36678), .Z(n36683) );
  NAND U37913 ( .A(n36681), .B(n36680), .Z(n36682) );
  NAND U37914 ( .A(n36683), .B(n36682), .Z(n36698) );
  XNOR U37915 ( .A(n36697), .B(n36698), .Z(n36689) );
  XNOR U37916 ( .A(n36690), .B(n36689), .Z(n36691) );
  XNOR U37917 ( .A(n36692), .B(n36691), .Z(n36721) );
  XNOR U37918 ( .A(sreg[1897]), .B(n36721), .Z(n36723) );
  NANDN U37919 ( .A(sreg[1896]), .B(n36684), .Z(n36688) );
  NAND U37920 ( .A(n36686), .B(n36685), .Z(n36687) );
  NAND U37921 ( .A(n36688), .B(n36687), .Z(n36722) );
  XNOR U37922 ( .A(n36723), .B(n36722), .Z(c[1897]) );
  NANDN U37923 ( .A(n36690), .B(n36689), .Z(n36694) );
  NANDN U37924 ( .A(n36692), .B(n36691), .Z(n36693) );
  AND U37925 ( .A(n36694), .B(n36693), .Z(n36729) );
  NANDN U37926 ( .A(n36696), .B(n36695), .Z(n36700) );
  NANDN U37927 ( .A(n36698), .B(n36697), .Z(n36699) );
  AND U37928 ( .A(n36700), .B(n36699), .Z(n36727) );
  NAND U37929 ( .A(n42143), .B(n36701), .Z(n36703) );
  XNOR U37930 ( .A(a[876]), .B(n4197), .Z(n36738) );
  NAND U37931 ( .A(n42144), .B(n36738), .Z(n36702) );
  AND U37932 ( .A(n36703), .B(n36702), .Z(n36753) );
  XOR U37933 ( .A(a[880]), .B(n42012), .Z(n36741) );
  XNOR U37934 ( .A(n36753), .B(n36752), .Z(n36755) );
  AND U37935 ( .A(a[882]), .B(b[0]), .Z(n36705) );
  XNOR U37936 ( .A(n36705), .B(n4071), .Z(n36707) );
  NANDN U37937 ( .A(b[0]), .B(a[881]), .Z(n36706) );
  NAND U37938 ( .A(n36707), .B(n36706), .Z(n36749) );
  XOR U37939 ( .A(a[878]), .B(n42085), .Z(n36742) );
  AND U37940 ( .A(a[874]), .B(b[7]), .Z(n36746) );
  XNOR U37941 ( .A(n36747), .B(n36746), .Z(n36748) );
  XNOR U37942 ( .A(n36749), .B(n36748), .Z(n36754) );
  XOR U37943 ( .A(n36755), .B(n36754), .Z(n36733) );
  NANDN U37944 ( .A(n36710), .B(n36709), .Z(n36714) );
  NANDN U37945 ( .A(n36712), .B(n36711), .Z(n36713) );
  AND U37946 ( .A(n36714), .B(n36713), .Z(n36732) );
  XNOR U37947 ( .A(n36733), .B(n36732), .Z(n36734) );
  NANDN U37948 ( .A(n36716), .B(n36715), .Z(n36720) );
  NAND U37949 ( .A(n36718), .B(n36717), .Z(n36719) );
  NAND U37950 ( .A(n36720), .B(n36719), .Z(n36735) );
  XNOR U37951 ( .A(n36734), .B(n36735), .Z(n36726) );
  XNOR U37952 ( .A(n36727), .B(n36726), .Z(n36728) );
  XNOR U37953 ( .A(n36729), .B(n36728), .Z(n36758) );
  XNOR U37954 ( .A(sreg[1898]), .B(n36758), .Z(n36760) );
  NANDN U37955 ( .A(sreg[1897]), .B(n36721), .Z(n36725) );
  NAND U37956 ( .A(n36723), .B(n36722), .Z(n36724) );
  NAND U37957 ( .A(n36725), .B(n36724), .Z(n36759) );
  XNOR U37958 ( .A(n36760), .B(n36759), .Z(c[1898]) );
  NANDN U37959 ( .A(n36727), .B(n36726), .Z(n36731) );
  NANDN U37960 ( .A(n36729), .B(n36728), .Z(n36730) );
  AND U37961 ( .A(n36731), .B(n36730), .Z(n36766) );
  NANDN U37962 ( .A(n36733), .B(n36732), .Z(n36737) );
  NANDN U37963 ( .A(n36735), .B(n36734), .Z(n36736) );
  AND U37964 ( .A(n36737), .B(n36736), .Z(n36764) );
  NAND U37965 ( .A(n42143), .B(n36738), .Z(n36740) );
  XNOR U37966 ( .A(a[877]), .B(n4197), .Z(n36775) );
  NAND U37967 ( .A(n42144), .B(n36775), .Z(n36739) );
  AND U37968 ( .A(n36740), .B(n36739), .Z(n36790) );
  XOR U37969 ( .A(a[881]), .B(n42012), .Z(n36778) );
  XNOR U37970 ( .A(n36790), .B(n36789), .Z(n36792) );
  XOR U37971 ( .A(a[879]), .B(n42085), .Z(n36782) );
  AND U37972 ( .A(a[875]), .B(b[7]), .Z(n36783) );
  XNOR U37973 ( .A(n36784), .B(n36783), .Z(n36785) );
  AND U37974 ( .A(a[883]), .B(b[0]), .Z(n36743) );
  XNOR U37975 ( .A(n36743), .B(n4071), .Z(n36745) );
  NANDN U37976 ( .A(b[0]), .B(a[882]), .Z(n36744) );
  NAND U37977 ( .A(n36745), .B(n36744), .Z(n36786) );
  XNOR U37978 ( .A(n36785), .B(n36786), .Z(n36791) );
  XOR U37979 ( .A(n36792), .B(n36791), .Z(n36770) );
  NANDN U37980 ( .A(n36747), .B(n36746), .Z(n36751) );
  NANDN U37981 ( .A(n36749), .B(n36748), .Z(n36750) );
  AND U37982 ( .A(n36751), .B(n36750), .Z(n36769) );
  XNOR U37983 ( .A(n36770), .B(n36769), .Z(n36771) );
  NANDN U37984 ( .A(n36753), .B(n36752), .Z(n36757) );
  NAND U37985 ( .A(n36755), .B(n36754), .Z(n36756) );
  NAND U37986 ( .A(n36757), .B(n36756), .Z(n36772) );
  XNOR U37987 ( .A(n36771), .B(n36772), .Z(n36763) );
  XNOR U37988 ( .A(n36764), .B(n36763), .Z(n36765) );
  XNOR U37989 ( .A(n36766), .B(n36765), .Z(n36795) );
  XNOR U37990 ( .A(sreg[1899]), .B(n36795), .Z(n36797) );
  NANDN U37991 ( .A(sreg[1898]), .B(n36758), .Z(n36762) );
  NAND U37992 ( .A(n36760), .B(n36759), .Z(n36761) );
  NAND U37993 ( .A(n36762), .B(n36761), .Z(n36796) );
  XNOR U37994 ( .A(n36797), .B(n36796), .Z(c[1899]) );
  NANDN U37995 ( .A(n36764), .B(n36763), .Z(n36768) );
  NANDN U37996 ( .A(n36766), .B(n36765), .Z(n36767) );
  AND U37997 ( .A(n36768), .B(n36767), .Z(n36803) );
  NANDN U37998 ( .A(n36770), .B(n36769), .Z(n36774) );
  NANDN U37999 ( .A(n36772), .B(n36771), .Z(n36773) );
  AND U38000 ( .A(n36774), .B(n36773), .Z(n36801) );
  NAND U38001 ( .A(n42143), .B(n36775), .Z(n36777) );
  XNOR U38002 ( .A(a[878]), .B(n4197), .Z(n36812) );
  NAND U38003 ( .A(n42144), .B(n36812), .Z(n36776) );
  AND U38004 ( .A(n36777), .B(n36776), .Z(n36827) );
  XOR U38005 ( .A(a[882]), .B(n42012), .Z(n36815) );
  XNOR U38006 ( .A(n36827), .B(n36826), .Z(n36829) );
  AND U38007 ( .A(a[884]), .B(b[0]), .Z(n36779) );
  XNOR U38008 ( .A(n36779), .B(n4071), .Z(n36781) );
  NANDN U38009 ( .A(b[0]), .B(a[883]), .Z(n36780) );
  NAND U38010 ( .A(n36781), .B(n36780), .Z(n36823) );
  XOR U38011 ( .A(a[880]), .B(n42085), .Z(n36816) );
  AND U38012 ( .A(a[876]), .B(b[7]), .Z(n36820) );
  XNOR U38013 ( .A(n36821), .B(n36820), .Z(n36822) );
  XNOR U38014 ( .A(n36823), .B(n36822), .Z(n36828) );
  XOR U38015 ( .A(n36829), .B(n36828), .Z(n36807) );
  NANDN U38016 ( .A(n36784), .B(n36783), .Z(n36788) );
  NANDN U38017 ( .A(n36786), .B(n36785), .Z(n36787) );
  AND U38018 ( .A(n36788), .B(n36787), .Z(n36806) );
  XNOR U38019 ( .A(n36807), .B(n36806), .Z(n36808) );
  NANDN U38020 ( .A(n36790), .B(n36789), .Z(n36794) );
  NAND U38021 ( .A(n36792), .B(n36791), .Z(n36793) );
  NAND U38022 ( .A(n36794), .B(n36793), .Z(n36809) );
  XNOR U38023 ( .A(n36808), .B(n36809), .Z(n36800) );
  XNOR U38024 ( .A(n36801), .B(n36800), .Z(n36802) );
  XNOR U38025 ( .A(n36803), .B(n36802), .Z(n36832) );
  XNOR U38026 ( .A(sreg[1900]), .B(n36832), .Z(n36834) );
  NANDN U38027 ( .A(sreg[1899]), .B(n36795), .Z(n36799) );
  NAND U38028 ( .A(n36797), .B(n36796), .Z(n36798) );
  NAND U38029 ( .A(n36799), .B(n36798), .Z(n36833) );
  XNOR U38030 ( .A(n36834), .B(n36833), .Z(c[1900]) );
  NANDN U38031 ( .A(n36801), .B(n36800), .Z(n36805) );
  NANDN U38032 ( .A(n36803), .B(n36802), .Z(n36804) );
  AND U38033 ( .A(n36805), .B(n36804), .Z(n36840) );
  NANDN U38034 ( .A(n36807), .B(n36806), .Z(n36811) );
  NANDN U38035 ( .A(n36809), .B(n36808), .Z(n36810) );
  AND U38036 ( .A(n36811), .B(n36810), .Z(n36838) );
  NAND U38037 ( .A(n42143), .B(n36812), .Z(n36814) );
  XNOR U38038 ( .A(a[879]), .B(n4197), .Z(n36849) );
  NAND U38039 ( .A(n42144), .B(n36849), .Z(n36813) );
  AND U38040 ( .A(n36814), .B(n36813), .Z(n36864) );
  XOR U38041 ( .A(a[883]), .B(n42012), .Z(n36852) );
  XNOR U38042 ( .A(n36864), .B(n36863), .Z(n36866) );
  XOR U38043 ( .A(a[881]), .B(n42085), .Z(n36856) );
  AND U38044 ( .A(a[877]), .B(b[7]), .Z(n36857) );
  XNOR U38045 ( .A(n36858), .B(n36857), .Z(n36859) );
  AND U38046 ( .A(a[885]), .B(b[0]), .Z(n36817) );
  XNOR U38047 ( .A(n36817), .B(n4071), .Z(n36819) );
  NANDN U38048 ( .A(b[0]), .B(a[884]), .Z(n36818) );
  NAND U38049 ( .A(n36819), .B(n36818), .Z(n36860) );
  XNOR U38050 ( .A(n36859), .B(n36860), .Z(n36865) );
  XOR U38051 ( .A(n36866), .B(n36865), .Z(n36844) );
  NANDN U38052 ( .A(n36821), .B(n36820), .Z(n36825) );
  NANDN U38053 ( .A(n36823), .B(n36822), .Z(n36824) );
  AND U38054 ( .A(n36825), .B(n36824), .Z(n36843) );
  XNOR U38055 ( .A(n36844), .B(n36843), .Z(n36845) );
  NANDN U38056 ( .A(n36827), .B(n36826), .Z(n36831) );
  NAND U38057 ( .A(n36829), .B(n36828), .Z(n36830) );
  NAND U38058 ( .A(n36831), .B(n36830), .Z(n36846) );
  XNOR U38059 ( .A(n36845), .B(n36846), .Z(n36837) );
  XNOR U38060 ( .A(n36838), .B(n36837), .Z(n36839) );
  XNOR U38061 ( .A(n36840), .B(n36839), .Z(n36869) );
  XNOR U38062 ( .A(sreg[1901]), .B(n36869), .Z(n36871) );
  NANDN U38063 ( .A(sreg[1900]), .B(n36832), .Z(n36836) );
  NAND U38064 ( .A(n36834), .B(n36833), .Z(n36835) );
  NAND U38065 ( .A(n36836), .B(n36835), .Z(n36870) );
  XNOR U38066 ( .A(n36871), .B(n36870), .Z(c[1901]) );
  NANDN U38067 ( .A(n36838), .B(n36837), .Z(n36842) );
  NANDN U38068 ( .A(n36840), .B(n36839), .Z(n36841) );
  AND U38069 ( .A(n36842), .B(n36841), .Z(n36877) );
  NANDN U38070 ( .A(n36844), .B(n36843), .Z(n36848) );
  NANDN U38071 ( .A(n36846), .B(n36845), .Z(n36847) );
  AND U38072 ( .A(n36848), .B(n36847), .Z(n36875) );
  NAND U38073 ( .A(n42143), .B(n36849), .Z(n36851) );
  XNOR U38074 ( .A(a[880]), .B(n4197), .Z(n36886) );
  NAND U38075 ( .A(n42144), .B(n36886), .Z(n36850) );
  AND U38076 ( .A(n36851), .B(n36850), .Z(n36901) );
  XOR U38077 ( .A(a[884]), .B(n42012), .Z(n36889) );
  XNOR U38078 ( .A(n36901), .B(n36900), .Z(n36903) );
  AND U38079 ( .A(a[886]), .B(b[0]), .Z(n36853) );
  XNOR U38080 ( .A(n36853), .B(n4071), .Z(n36855) );
  NANDN U38081 ( .A(b[0]), .B(a[885]), .Z(n36854) );
  NAND U38082 ( .A(n36855), .B(n36854), .Z(n36897) );
  XOR U38083 ( .A(a[882]), .B(n42085), .Z(n36893) );
  AND U38084 ( .A(a[878]), .B(b[7]), .Z(n36894) );
  XNOR U38085 ( .A(n36895), .B(n36894), .Z(n36896) );
  XNOR U38086 ( .A(n36897), .B(n36896), .Z(n36902) );
  XOR U38087 ( .A(n36903), .B(n36902), .Z(n36881) );
  NANDN U38088 ( .A(n36858), .B(n36857), .Z(n36862) );
  NANDN U38089 ( .A(n36860), .B(n36859), .Z(n36861) );
  AND U38090 ( .A(n36862), .B(n36861), .Z(n36880) );
  XNOR U38091 ( .A(n36881), .B(n36880), .Z(n36882) );
  NANDN U38092 ( .A(n36864), .B(n36863), .Z(n36868) );
  NAND U38093 ( .A(n36866), .B(n36865), .Z(n36867) );
  NAND U38094 ( .A(n36868), .B(n36867), .Z(n36883) );
  XNOR U38095 ( .A(n36882), .B(n36883), .Z(n36874) );
  XNOR U38096 ( .A(n36875), .B(n36874), .Z(n36876) );
  XNOR U38097 ( .A(n36877), .B(n36876), .Z(n36906) );
  XNOR U38098 ( .A(sreg[1902]), .B(n36906), .Z(n36908) );
  NANDN U38099 ( .A(sreg[1901]), .B(n36869), .Z(n36873) );
  NAND U38100 ( .A(n36871), .B(n36870), .Z(n36872) );
  NAND U38101 ( .A(n36873), .B(n36872), .Z(n36907) );
  XNOR U38102 ( .A(n36908), .B(n36907), .Z(c[1902]) );
  NANDN U38103 ( .A(n36875), .B(n36874), .Z(n36879) );
  NANDN U38104 ( .A(n36877), .B(n36876), .Z(n36878) );
  AND U38105 ( .A(n36879), .B(n36878), .Z(n36914) );
  NANDN U38106 ( .A(n36881), .B(n36880), .Z(n36885) );
  NANDN U38107 ( .A(n36883), .B(n36882), .Z(n36884) );
  AND U38108 ( .A(n36885), .B(n36884), .Z(n36912) );
  NAND U38109 ( .A(n42143), .B(n36886), .Z(n36888) );
  XNOR U38110 ( .A(a[881]), .B(n4197), .Z(n36923) );
  NAND U38111 ( .A(n42144), .B(n36923), .Z(n36887) );
  AND U38112 ( .A(n36888), .B(n36887), .Z(n36938) );
  XOR U38113 ( .A(a[885]), .B(n42012), .Z(n36926) );
  XNOR U38114 ( .A(n36938), .B(n36937), .Z(n36940) );
  AND U38115 ( .A(a[887]), .B(b[0]), .Z(n36890) );
  XNOR U38116 ( .A(n36890), .B(n4071), .Z(n36892) );
  NANDN U38117 ( .A(b[0]), .B(a[886]), .Z(n36891) );
  NAND U38118 ( .A(n36892), .B(n36891), .Z(n36934) );
  XOR U38119 ( .A(a[883]), .B(n42085), .Z(n36927) );
  AND U38120 ( .A(a[879]), .B(b[7]), .Z(n36931) );
  XNOR U38121 ( .A(n36932), .B(n36931), .Z(n36933) );
  XNOR U38122 ( .A(n36934), .B(n36933), .Z(n36939) );
  XOR U38123 ( .A(n36940), .B(n36939), .Z(n36918) );
  NANDN U38124 ( .A(n36895), .B(n36894), .Z(n36899) );
  NANDN U38125 ( .A(n36897), .B(n36896), .Z(n36898) );
  AND U38126 ( .A(n36899), .B(n36898), .Z(n36917) );
  XNOR U38127 ( .A(n36918), .B(n36917), .Z(n36919) );
  NANDN U38128 ( .A(n36901), .B(n36900), .Z(n36905) );
  NAND U38129 ( .A(n36903), .B(n36902), .Z(n36904) );
  NAND U38130 ( .A(n36905), .B(n36904), .Z(n36920) );
  XNOR U38131 ( .A(n36919), .B(n36920), .Z(n36911) );
  XNOR U38132 ( .A(n36912), .B(n36911), .Z(n36913) );
  XNOR U38133 ( .A(n36914), .B(n36913), .Z(n36943) );
  XNOR U38134 ( .A(sreg[1903]), .B(n36943), .Z(n36945) );
  NANDN U38135 ( .A(sreg[1902]), .B(n36906), .Z(n36910) );
  NAND U38136 ( .A(n36908), .B(n36907), .Z(n36909) );
  NAND U38137 ( .A(n36910), .B(n36909), .Z(n36944) );
  XNOR U38138 ( .A(n36945), .B(n36944), .Z(c[1903]) );
  NANDN U38139 ( .A(n36912), .B(n36911), .Z(n36916) );
  NANDN U38140 ( .A(n36914), .B(n36913), .Z(n36915) );
  AND U38141 ( .A(n36916), .B(n36915), .Z(n36951) );
  NANDN U38142 ( .A(n36918), .B(n36917), .Z(n36922) );
  NANDN U38143 ( .A(n36920), .B(n36919), .Z(n36921) );
  AND U38144 ( .A(n36922), .B(n36921), .Z(n36949) );
  NAND U38145 ( .A(n42143), .B(n36923), .Z(n36925) );
  XNOR U38146 ( .A(a[882]), .B(n4197), .Z(n36960) );
  NAND U38147 ( .A(n42144), .B(n36960), .Z(n36924) );
  AND U38148 ( .A(n36925), .B(n36924), .Z(n36975) );
  XOR U38149 ( .A(a[886]), .B(n42012), .Z(n36963) );
  XNOR U38150 ( .A(n36975), .B(n36974), .Z(n36977) );
  XOR U38151 ( .A(a[884]), .B(n42085), .Z(n36967) );
  AND U38152 ( .A(a[880]), .B(b[7]), .Z(n36968) );
  XNOR U38153 ( .A(n36969), .B(n36968), .Z(n36970) );
  AND U38154 ( .A(a[888]), .B(b[0]), .Z(n36928) );
  XNOR U38155 ( .A(n36928), .B(n4071), .Z(n36930) );
  NANDN U38156 ( .A(b[0]), .B(a[887]), .Z(n36929) );
  NAND U38157 ( .A(n36930), .B(n36929), .Z(n36971) );
  XNOR U38158 ( .A(n36970), .B(n36971), .Z(n36976) );
  XOR U38159 ( .A(n36977), .B(n36976), .Z(n36955) );
  NANDN U38160 ( .A(n36932), .B(n36931), .Z(n36936) );
  NANDN U38161 ( .A(n36934), .B(n36933), .Z(n36935) );
  AND U38162 ( .A(n36936), .B(n36935), .Z(n36954) );
  XNOR U38163 ( .A(n36955), .B(n36954), .Z(n36956) );
  NANDN U38164 ( .A(n36938), .B(n36937), .Z(n36942) );
  NAND U38165 ( .A(n36940), .B(n36939), .Z(n36941) );
  NAND U38166 ( .A(n36942), .B(n36941), .Z(n36957) );
  XNOR U38167 ( .A(n36956), .B(n36957), .Z(n36948) );
  XNOR U38168 ( .A(n36949), .B(n36948), .Z(n36950) );
  XNOR U38169 ( .A(n36951), .B(n36950), .Z(n36980) );
  XNOR U38170 ( .A(sreg[1904]), .B(n36980), .Z(n36982) );
  NANDN U38171 ( .A(sreg[1903]), .B(n36943), .Z(n36947) );
  NAND U38172 ( .A(n36945), .B(n36944), .Z(n36946) );
  NAND U38173 ( .A(n36947), .B(n36946), .Z(n36981) );
  XNOR U38174 ( .A(n36982), .B(n36981), .Z(c[1904]) );
  NANDN U38175 ( .A(n36949), .B(n36948), .Z(n36953) );
  NANDN U38176 ( .A(n36951), .B(n36950), .Z(n36952) );
  AND U38177 ( .A(n36953), .B(n36952), .Z(n36988) );
  NANDN U38178 ( .A(n36955), .B(n36954), .Z(n36959) );
  NANDN U38179 ( .A(n36957), .B(n36956), .Z(n36958) );
  AND U38180 ( .A(n36959), .B(n36958), .Z(n36986) );
  NAND U38181 ( .A(n42143), .B(n36960), .Z(n36962) );
  XNOR U38182 ( .A(a[883]), .B(n4198), .Z(n36997) );
  NAND U38183 ( .A(n42144), .B(n36997), .Z(n36961) );
  AND U38184 ( .A(n36962), .B(n36961), .Z(n37012) );
  XOR U38185 ( .A(a[887]), .B(n42012), .Z(n37000) );
  XNOR U38186 ( .A(n37012), .B(n37011), .Z(n37014) );
  AND U38187 ( .A(a[889]), .B(b[0]), .Z(n36964) );
  XNOR U38188 ( .A(n36964), .B(n4071), .Z(n36966) );
  NANDN U38189 ( .A(b[0]), .B(a[888]), .Z(n36965) );
  NAND U38190 ( .A(n36966), .B(n36965), .Z(n37008) );
  XOR U38191 ( .A(a[885]), .B(n42085), .Z(n37001) );
  AND U38192 ( .A(a[881]), .B(b[7]), .Z(n37005) );
  XNOR U38193 ( .A(n37006), .B(n37005), .Z(n37007) );
  XNOR U38194 ( .A(n37008), .B(n37007), .Z(n37013) );
  XOR U38195 ( .A(n37014), .B(n37013), .Z(n36992) );
  NANDN U38196 ( .A(n36969), .B(n36968), .Z(n36973) );
  NANDN U38197 ( .A(n36971), .B(n36970), .Z(n36972) );
  AND U38198 ( .A(n36973), .B(n36972), .Z(n36991) );
  XNOR U38199 ( .A(n36992), .B(n36991), .Z(n36993) );
  NANDN U38200 ( .A(n36975), .B(n36974), .Z(n36979) );
  NAND U38201 ( .A(n36977), .B(n36976), .Z(n36978) );
  NAND U38202 ( .A(n36979), .B(n36978), .Z(n36994) );
  XNOR U38203 ( .A(n36993), .B(n36994), .Z(n36985) );
  XNOR U38204 ( .A(n36986), .B(n36985), .Z(n36987) );
  XNOR U38205 ( .A(n36988), .B(n36987), .Z(n37017) );
  XNOR U38206 ( .A(sreg[1905]), .B(n37017), .Z(n37019) );
  NANDN U38207 ( .A(sreg[1904]), .B(n36980), .Z(n36984) );
  NAND U38208 ( .A(n36982), .B(n36981), .Z(n36983) );
  NAND U38209 ( .A(n36984), .B(n36983), .Z(n37018) );
  XNOR U38210 ( .A(n37019), .B(n37018), .Z(c[1905]) );
  NANDN U38211 ( .A(n36986), .B(n36985), .Z(n36990) );
  NANDN U38212 ( .A(n36988), .B(n36987), .Z(n36989) );
  AND U38213 ( .A(n36990), .B(n36989), .Z(n37025) );
  NANDN U38214 ( .A(n36992), .B(n36991), .Z(n36996) );
  NANDN U38215 ( .A(n36994), .B(n36993), .Z(n36995) );
  AND U38216 ( .A(n36996), .B(n36995), .Z(n37023) );
  NAND U38217 ( .A(n42143), .B(n36997), .Z(n36999) );
  XNOR U38218 ( .A(a[884]), .B(n4198), .Z(n37034) );
  NAND U38219 ( .A(n42144), .B(n37034), .Z(n36998) );
  AND U38220 ( .A(n36999), .B(n36998), .Z(n37049) );
  XOR U38221 ( .A(a[888]), .B(n42012), .Z(n37037) );
  XNOR U38222 ( .A(n37049), .B(n37048), .Z(n37051) );
  XOR U38223 ( .A(a[886]), .B(n42085), .Z(n37041) );
  AND U38224 ( .A(a[882]), .B(b[7]), .Z(n37042) );
  XNOR U38225 ( .A(n37043), .B(n37042), .Z(n37044) );
  AND U38226 ( .A(a[890]), .B(b[0]), .Z(n37002) );
  XNOR U38227 ( .A(n37002), .B(n4071), .Z(n37004) );
  NANDN U38228 ( .A(b[0]), .B(a[889]), .Z(n37003) );
  NAND U38229 ( .A(n37004), .B(n37003), .Z(n37045) );
  XNOR U38230 ( .A(n37044), .B(n37045), .Z(n37050) );
  XOR U38231 ( .A(n37051), .B(n37050), .Z(n37029) );
  NANDN U38232 ( .A(n37006), .B(n37005), .Z(n37010) );
  NANDN U38233 ( .A(n37008), .B(n37007), .Z(n37009) );
  AND U38234 ( .A(n37010), .B(n37009), .Z(n37028) );
  XNOR U38235 ( .A(n37029), .B(n37028), .Z(n37030) );
  NANDN U38236 ( .A(n37012), .B(n37011), .Z(n37016) );
  NAND U38237 ( .A(n37014), .B(n37013), .Z(n37015) );
  NAND U38238 ( .A(n37016), .B(n37015), .Z(n37031) );
  XNOR U38239 ( .A(n37030), .B(n37031), .Z(n37022) );
  XNOR U38240 ( .A(n37023), .B(n37022), .Z(n37024) );
  XNOR U38241 ( .A(n37025), .B(n37024), .Z(n37054) );
  XNOR U38242 ( .A(sreg[1906]), .B(n37054), .Z(n37056) );
  NANDN U38243 ( .A(sreg[1905]), .B(n37017), .Z(n37021) );
  NAND U38244 ( .A(n37019), .B(n37018), .Z(n37020) );
  NAND U38245 ( .A(n37021), .B(n37020), .Z(n37055) );
  XNOR U38246 ( .A(n37056), .B(n37055), .Z(c[1906]) );
  NANDN U38247 ( .A(n37023), .B(n37022), .Z(n37027) );
  NANDN U38248 ( .A(n37025), .B(n37024), .Z(n37026) );
  AND U38249 ( .A(n37027), .B(n37026), .Z(n37062) );
  NANDN U38250 ( .A(n37029), .B(n37028), .Z(n37033) );
  NANDN U38251 ( .A(n37031), .B(n37030), .Z(n37032) );
  AND U38252 ( .A(n37033), .B(n37032), .Z(n37060) );
  NAND U38253 ( .A(n42143), .B(n37034), .Z(n37036) );
  XNOR U38254 ( .A(a[885]), .B(n4198), .Z(n37071) );
  NAND U38255 ( .A(n42144), .B(n37071), .Z(n37035) );
  AND U38256 ( .A(n37036), .B(n37035), .Z(n37086) );
  XOR U38257 ( .A(a[889]), .B(n42012), .Z(n37074) );
  XNOR U38258 ( .A(n37086), .B(n37085), .Z(n37088) );
  AND U38259 ( .A(a[891]), .B(b[0]), .Z(n37038) );
  XNOR U38260 ( .A(n37038), .B(n4071), .Z(n37040) );
  NANDN U38261 ( .A(b[0]), .B(a[890]), .Z(n37039) );
  NAND U38262 ( .A(n37040), .B(n37039), .Z(n37082) );
  XOR U38263 ( .A(a[887]), .B(n42085), .Z(n37078) );
  AND U38264 ( .A(a[883]), .B(b[7]), .Z(n37079) );
  XNOR U38265 ( .A(n37080), .B(n37079), .Z(n37081) );
  XNOR U38266 ( .A(n37082), .B(n37081), .Z(n37087) );
  XOR U38267 ( .A(n37088), .B(n37087), .Z(n37066) );
  NANDN U38268 ( .A(n37043), .B(n37042), .Z(n37047) );
  NANDN U38269 ( .A(n37045), .B(n37044), .Z(n37046) );
  AND U38270 ( .A(n37047), .B(n37046), .Z(n37065) );
  XNOR U38271 ( .A(n37066), .B(n37065), .Z(n37067) );
  NANDN U38272 ( .A(n37049), .B(n37048), .Z(n37053) );
  NAND U38273 ( .A(n37051), .B(n37050), .Z(n37052) );
  NAND U38274 ( .A(n37053), .B(n37052), .Z(n37068) );
  XNOR U38275 ( .A(n37067), .B(n37068), .Z(n37059) );
  XNOR U38276 ( .A(n37060), .B(n37059), .Z(n37061) );
  XNOR U38277 ( .A(n37062), .B(n37061), .Z(n37091) );
  XNOR U38278 ( .A(sreg[1907]), .B(n37091), .Z(n37093) );
  NANDN U38279 ( .A(sreg[1906]), .B(n37054), .Z(n37058) );
  NAND U38280 ( .A(n37056), .B(n37055), .Z(n37057) );
  NAND U38281 ( .A(n37058), .B(n37057), .Z(n37092) );
  XNOR U38282 ( .A(n37093), .B(n37092), .Z(c[1907]) );
  NANDN U38283 ( .A(n37060), .B(n37059), .Z(n37064) );
  NANDN U38284 ( .A(n37062), .B(n37061), .Z(n37063) );
  AND U38285 ( .A(n37064), .B(n37063), .Z(n37099) );
  NANDN U38286 ( .A(n37066), .B(n37065), .Z(n37070) );
  NANDN U38287 ( .A(n37068), .B(n37067), .Z(n37069) );
  AND U38288 ( .A(n37070), .B(n37069), .Z(n37097) );
  NAND U38289 ( .A(n42143), .B(n37071), .Z(n37073) );
  XNOR U38290 ( .A(a[886]), .B(n4198), .Z(n37108) );
  NAND U38291 ( .A(n42144), .B(n37108), .Z(n37072) );
  AND U38292 ( .A(n37073), .B(n37072), .Z(n37123) );
  XOR U38293 ( .A(a[890]), .B(n42012), .Z(n37111) );
  XNOR U38294 ( .A(n37123), .B(n37122), .Z(n37125) );
  AND U38295 ( .A(a[892]), .B(b[0]), .Z(n37075) );
  XNOR U38296 ( .A(n37075), .B(n4071), .Z(n37077) );
  NANDN U38297 ( .A(b[0]), .B(a[891]), .Z(n37076) );
  NAND U38298 ( .A(n37077), .B(n37076), .Z(n37119) );
  XOR U38299 ( .A(a[888]), .B(n42085), .Z(n37112) );
  AND U38300 ( .A(a[884]), .B(b[7]), .Z(n37116) );
  XNOR U38301 ( .A(n37117), .B(n37116), .Z(n37118) );
  XNOR U38302 ( .A(n37119), .B(n37118), .Z(n37124) );
  XOR U38303 ( .A(n37125), .B(n37124), .Z(n37103) );
  NANDN U38304 ( .A(n37080), .B(n37079), .Z(n37084) );
  NANDN U38305 ( .A(n37082), .B(n37081), .Z(n37083) );
  AND U38306 ( .A(n37084), .B(n37083), .Z(n37102) );
  XNOR U38307 ( .A(n37103), .B(n37102), .Z(n37104) );
  NANDN U38308 ( .A(n37086), .B(n37085), .Z(n37090) );
  NAND U38309 ( .A(n37088), .B(n37087), .Z(n37089) );
  NAND U38310 ( .A(n37090), .B(n37089), .Z(n37105) );
  XNOR U38311 ( .A(n37104), .B(n37105), .Z(n37096) );
  XNOR U38312 ( .A(n37097), .B(n37096), .Z(n37098) );
  XNOR U38313 ( .A(n37099), .B(n37098), .Z(n37128) );
  XNOR U38314 ( .A(sreg[1908]), .B(n37128), .Z(n37130) );
  NANDN U38315 ( .A(sreg[1907]), .B(n37091), .Z(n37095) );
  NAND U38316 ( .A(n37093), .B(n37092), .Z(n37094) );
  NAND U38317 ( .A(n37095), .B(n37094), .Z(n37129) );
  XNOR U38318 ( .A(n37130), .B(n37129), .Z(c[1908]) );
  NANDN U38319 ( .A(n37097), .B(n37096), .Z(n37101) );
  NANDN U38320 ( .A(n37099), .B(n37098), .Z(n37100) );
  AND U38321 ( .A(n37101), .B(n37100), .Z(n37136) );
  NANDN U38322 ( .A(n37103), .B(n37102), .Z(n37107) );
  NANDN U38323 ( .A(n37105), .B(n37104), .Z(n37106) );
  AND U38324 ( .A(n37107), .B(n37106), .Z(n37134) );
  NAND U38325 ( .A(n42143), .B(n37108), .Z(n37110) );
  XNOR U38326 ( .A(a[887]), .B(n4198), .Z(n37145) );
  NAND U38327 ( .A(n42144), .B(n37145), .Z(n37109) );
  AND U38328 ( .A(n37110), .B(n37109), .Z(n37160) );
  XOR U38329 ( .A(a[891]), .B(n42012), .Z(n37148) );
  XNOR U38330 ( .A(n37160), .B(n37159), .Z(n37162) );
  XOR U38331 ( .A(a[889]), .B(n42085), .Z(n37152) );
  AND U38332 ( .A(a[885]), .B(b[7]), .Z(n37153) );
  XNOR U38333 ( .A(n37154), .B(n37153), .Z(n37155) );
  AND U38334 ( .A(a[893]), .B(b[0]), .Z(n37113) );
  XNOR U38335 ( .A(n37113), .B(n4071), .Z(n37115) );
  NANDN U38336 ( .A(b[0]), .B(a[892]), .Z(n37114) );
  NAND U38337 ( .A(n37115), .B(n37114), .Z(n37156) );
  XNOR U38338 ( .A(n37155), .B(n37156), .Z(n37161) );
  XOR U38339 ( .A(n37162), .B(n37161), .Z(n37140) );
  NANDN U38340 ( .A(n37117), .B(n37116), .Z(n37121) );
  NANDN U38341 ( .A(n37119), .B(n37118), .Z(n37120) );
  AND U38342 ( .A(n37121), .B(n37120), .Z(n37139) );
  XNOR U38343 ( .A(n37140), .B(n37139), .Z(n37141) );
  NANDN U38344 ( .A(n37123), .B(n37122), .Z(n37127) );
  NAND U38345 ( .A(n37125), .B(n37124), .Z(n37126) );
  NAND U38346 ( .A(n37127), .B(n37126), .Z(n37142) );
  XNOR U38347 ( .A(n37141), .B(n37142), .Z(n37133) );
  XNOR U38348 ( .A(n37134), .B(n37133), .Z(n37135) );
  XNOR U38349 ( .A(n37136), .B(n37135), .Z(n37165) );
  XNOR U38350 ( .A(sreg[1909]), .B(n37165), .Z(n37167) );
  NANDN U38351 ( .A(sreg[1908]), .B(n37128), .Z(n37132) );
  NAND U38352 ( .A(n37130), .B(n37129), .Z(n37131) );
  NAND U38353 ( .A(n37132), .B(n37131), .Z(n37166) );
  XNOR U38354 ( .A(n37167), .B(n37166), .Z(c[1909]) );
  NANDN U38355 ( .A(n37134), .B(n37133), .Z(n37138) );
  NANDN U38356 ( .A(n37136), .B(n37135), .Z(n37137) );
  AND U38357 ( .A(n37138), .B(n37137), .Z(n37173) );
  NANDN U38358 ( .A(n37140), .B(n37139), .Z(n37144) );
  NANDN U38359 ( .A(n37142), .B(n37141), .Z(n37143) );
  AND U38360 ( .A(n37144), .B(n37143), .Z(n37171) );
  NAND U38361 ( .A(n42143), .B(n37145), .Z(n37147) );
  XNOR U38362 ( .A(a[888]), .B(n4198), .Z(n37182) );
  NAND U38363 ( .A(n42144), .B(n37182), .Z(n37146) );
  AND U38364 ( .A(n37147), .B(n37146), .Z(n37197) );
  XOR U38365 ( .A(a[892]), .B(n42012), .Z(n37185) );
  XNOR U38366 ( .A(n37197), .B(n37196), .Z(n37199) );
  AND U38367 ( .A(a[894]), .B(b[0]), .Z(n37149) );
  XNOR U38368 ( .A(n37149), .B(n4071), .Z(n37151) );
  NANDN U38369 ( .A(b[0]), .B(a[893]), .Z(n37150) );
  NAND U38370 ( .A(n37151), .B(n37150), .Z(n37193) );
  XOR U38371 ( .A(a[890]), .B(n42085), .Z(n37189) );
  AND U38372 ( .A(a[886]), .B(b[7]), .Z(n37190) );
  XNOR U38373 ( .A(n37191), .B(n37190), .Z(n37192) );
  XNOR U38374 ( .A(n37193), .B(n37192), .Z(n37198) );
  XOR U38375 ( .A(n37199), .B(n37198), .Z(n37177) );
  NANDN U38376 ( .A(n37154), .B(n37153), .Z(n37158) );
  NANDN U38377 ( .A(n37156), .B(n37155), .Z(n37157) );
  AND U38378 ( .A(n37158), .B(n37157), .Z(n37176) );
  XNOR U38379 ( .A(n37177), .B(n37176), .Z(n37178) );
  NANDN U38380 ( .A(n37160), .B(n37159), .Z(n37164) );
  NAND U38381 ( .A(n37162), .B(n37161), .Z(n37163) );
  NAND U38382 ( .A(n37164), .B(n37163), .Z(n37179) );
  XNOR U38383 ( .A(n37178), .B(n37179), .Z(n37170) );
  XNOR U38384 ( .A(n37171), .B(n37170), .Z(n37172) );
  XNOR U38385 ( .A(n37173), .B(n37172), .Z(n37202) );
  XNOR U38386 ( .A(sreg[1910]), .B(n37202), .Z(n37204) );
  NANDN U38387 ( .A(sreg[1909]), .B(n37165), .Z(n37169) );
  NAND U38388 ( .A(n37167), .B(n37166), .Z(n37168) );
  NAND U38389 ( .A(n37169), .B(n37168), .Z(n37203) );
  XNOR U38390 ( .A(n37204), .B(n37203), .Z(c[1910]) );
  NANDN U38391 ( .A(n37171), .B(n37170), .Z(n37175) );
  NANDN U38392 ( .A(n37173), .B(n37172), .Z(n37174) );
  AND U38393 ( .A(n37175), .B(n37174), .Z(n37210) );
  NANDN U38394 ( .A(n37177), .B(n37176), .Z(n37181) );
  NANDN U38395 ( .A(n37179), .B(n37178), .Z(n37180) );
  AND U38396 ( .A(n37181), .B(n37180), .Z(n37208) );
  NAND U38397 ( .A(n42143), .B(n37182), .Z(n37184) );
  XNOR U38398 ( .A(a[889]), .B(n4198), .Z(n37219) );
  NAND U38399 ( .A(n42144), .B(n37219), .Z(n37183) );
  AND U38400 ( .A(n37184), .B(n37183), .Z(n37234) );
  XOR U38401 ( .A(a[893]), .B(n42012), .Z(n37222) );
  XNOR U38402 ( .A(n37234), .B(n37233), .Z(n37236) );
  AND U38403 ( .A(b[0]), .B(a[895]), .Z(n37186) );
  XOR U38404 ( .A(b[1]), .B(n37186), .Z(n37188) );
  NANDN U38405 ( .A(b[0]), .B(a[894]), .Z(n37187) );
  AND U38406 ( .A(n37188), .B(n37187), .Z(n37229) );
  XOR U38407 ( .A(a[891]), .B(n42085), .Z(n37226) );
  AND U38408 ( .A(a[887]), .B(b[7]), .Z(n37227) );
  XOR U38409 ( .A(n37228), .B(n37227), .Z(n37230) );
  XNOR U38410 ( .A(n37229), .B(n37230), .Z(n37235) );
  XOR U38411 ( .A(n37236), .B(n37235), .Z(n37214) );
  NANDN U38412 ( .A(n37191), .B(n37190), .Z(n37195) );
  NANDN U38413 ( .A(n37193), .B(n37192), .Z(n37194) );
  AND U38414 ( .A(n37195), .B(n37194), .Z(n37213) );
  XNOR U38415 ( .A(n37214), .B(n37213), .Z(n37215) );
  NANDN U38416 ( .A(n37197), .B(n37196), .Z(n37201) );
  NAND U38417 ( .A(n37199), .B(n37198), .Z(n37200) );
  NAND U38418 ( .A(n37201), .B(n37200), .Z(n37216) );
  XNOR U38419 ( .A(n37215), .B(n37216), .Z(n37207) );
  XNOR U38420 ( .A(n37208), .B(n37207), .Z(n37209) );
  XNOR U38421 ( .A(n37210), .B(n37209), .Z(n37239) );
  XNOR U38422 ( .A(sreg[1911]), .B(n37239), .Z(n37241) );
  NANDN U38423 ( .A(sreg[1910]), .B(n37202), .Z(n37206) );
  NAND U38424 ( .A(n37204), .B(n37203), .Z(n37205) );
  NAND U38425 ( .A(n37206), .B(n37205), .Z(n37240) );
  XNOR U38426 ( .A(n37241), .B(n37240), .Z(c[1911]) );
  NANDN U38427 ( .A(n37208), .B(n37207), .Z(n37212) );
  NANDN U38428 ( .A(n37210), .B(n37209), .Z(n37211) );
  AND U38429 ( .A(n37212), .B(n37211), .Z(n37247) );
  NANDN U38430 ( .A(n37214), .B(n37213), .Z(n37218) );
  NANDN U38431 ( .A(n37216), .B(n37215), .Z(n37217) );
  AND U38432 ( .A(n37218), .B(n37217), .Z(n37245) );
  NAND U38433 ( .A(n42143), .B(n37219), .Z(n37221) );
  XNOR U38434 ( .A(a[890]), .B(n4199), .Z(n37256) );
  NAND U38435 ( .A(n42144), .B(n37256), .Z(n37220) );
  AND U38436 ( .A(n37221), .B(n37220), .Z(n37271) );
  XOR U38437 ( .A(a[894]), .B(n42012), .Z(n37259) );
  XNOR U38438 ( .A(n37271), .B(n37270), .Z(n37273) );
  AND U38439 ( .A(a[896]), .B(b[0]), .Z(n37223) );
  XNOR U38440 ( .A(n37223), .B(n4071), .Z(n37225) );
  NANDN U38441 ( .A(b[0]), .B(a[895]), .Z(n37224) );
  NAND U38442 ( .A(n37225), .B(n37224), .Z(n37267) );
  XOR U38443 ( .A(a[892]), .B(n42085), .Z(n37263) );
  AND U38444 ( .A(a[888]), .B(b[7]), .Z(n37264) );
  XNOR U38445 ( .A(n37265), .B(n37264), .Z(n37266) );
  XNOR U38446 ( .A(n37267), .B(n37266), .Z(n37272) );
  XOR U38447 ( .A(n37273), .B(n37272), .Z(n37251) );
  NANDN U38448 ( .A(n37228), .B(n37227), .Z(n37232) );
  NANDN U38449 ( .A(n37230), .B(n37229), .Z(n37231) );
  AND U38450 ( .A(n37232), .B(n37231), .Z(n37250) );
  XNOR U38451 ( .A(n37251), .B(n37250), .Z(n37252) );
  NANDN U38452 ( .A(n37234), .B(n37233), .Z(n37238) );
  NAND U38453 ( .A(n37236), .B(n37235), .Z(n37237) );
  NAND U38454 ( .A(n37238), .B(n37237), .Z(n37253) );
  XNOR U38455 ( .A(n37252), .B(n37253), .Z(n37244) );
  XNOR U38456 ( .A(n37245), .B(n37244), .Z(n37246) );
  XNOR U38457 ( .A(n37247), .B(n37246), .Z(n37276) );
  XNOR U38458 ( .A(sreg[1912]), .B(n37276), .Z(n37278) );
  NANDN U38459 ( .A(sreg[1911]), .B(n37239), .Z(n37243) );
  NAND U38460 ( .A(n37241), .B(n37240), .Z(n37242) );
  NAND U38461 ( .A(n37243), .B(n37242), .Z(n37277) );
  XNOR U38462 ( .A(n37278), .B(n37277), .Z(c[1912]) );
  NANDN U38463 ( .A(n37245), .B(n37244), .Z(n37249) );
  NANDN U38464 ( .A(n37247), .B(n37246), .Z(n37248) );
  AND U38465 ( .A(n37249), .B(n37248), .Z(n37284) );
  NANDN U38466 ( .A(n37251), .B(n37250), .Z(n37255) );
  NANDN U38467 ( .A(n37253), .B(n37252), .Z(n37254) );
  AND U38468 ( .A(n37255), .B(n37254), .Z(n37282) );
  NAND U38469 ( .A(n42143), .B(n37256), .Z(n37258) );
  XNOR U38470 ( .A(a[891]), .B(n4199), .Z(n37293) );
  NAND U38471 ( .A(n42144), .B(n37293), .Z(n37257) );
  AND U38472 ( .A(n37258), .B(n37257), .Z(n37308) );
  XOR U38473 ( .A(a[895]), .B(n42012), .Z(n37296) );
  XNOR U38474 ( .A(n37308), .B(n37307), .Z(n37310) );
  AND U38475 ( .A(a[897]), .B(b[0]), .Z(n37260) );
  XNOR U38476 ( .A(n37260), .B(n4071), .Z(n37262) );
  NANDN U38477 ( .A(b[0]), .B(a[896]), .Z(n37261) );
  NAND U38478 ( .A(n37262), .B(n37261), .Z(n37304) );
  XOR U38479 ( .A(a[893]), .B(n42085), .Z(n37297) );
  AND U38480 ( .A(a[889]), .B(b[7]), .Z(n37301) );
  XNOR U38481 ( .A(n37302), .B(n37301), .Z(n37303) );
  XNOR U38482 ( .A(n37304), .B(n37303), .Z(n37309) );
  XOR U38483 ( .A(n37310), .B(n37309), .Z(n37288) );
  NANDN U38484 ( .A(n37265), .B(n37264), .Z(n37269) );
  NANDN U38485 ( .A(n37267), .B(n37266), .Z(n37268) );
  AND U38486 ( .A(n37269), .B(n37268), .Z(n37287) );
  XNOR U38487 ( .A(n37288), .B(n37287), .Z(n37289) );
  NANDN U38488 ( .A(n37271), .B(n37270), .Z(n37275) );
  NAND U38489 ( .A(n37273), .B(n37272), .Z(n37274) );
  NAND U38490 ( .A(n37275), .B(n37274), .Z(n37290) );
  XNOR U38491 ( .A(n37289), .B(n37290), .Z(n37281) );
  XNOR U38492 ( .A(n37282), .B(n37281), .Z(n37283) );
  XNOR U38493 ( .A(n37284), .B(n37283), .Z(n37313) );
  XNOR U38494 ( .A(sreg[1913]), .B(n37313), .Z(n37315) );
  NANDN U38495 ( .A(sreg[1912]), .B(n37276), .Z(n37280) );
  NAND U38496 ( .A(n37278), .B(n37277), .Z(n37279) );
  NAND U38497 ( .A(n37280), .B(n37279), .Z(n37314) );
  XNOR U38498 ( .A(n37315), .B(n37314), .Z(c[1913]) );
  NANDN U38499 ( .A(n37282), .B(n37281), .Z(n37286) );
  NANDN U38500 ( .A(n37284), .B(n37283), .Z(n37285) );
  AND U38501 ( .A(n37286), .B(n37285), .Z(n37321) );
  NANDN U38502 ( .A(n37288), .B(n37287), .Z(n37292) );
  NANDN U38503 ( .A(n37290), .B(n37289), .Z(n37291) );
  AND U38504 ( .A(n37292), .B(n37291), .Z(n37319) );
  NAND U38505 ( .A(n42143), .B(n37293), .Z(n37295) );
  XNOR U38506 ( .A(a[892]), .B(n4199), .Z(n37330) );
  NAND U38507 ( .A(n42144), .B(n37330), .Z(n37294) );
  AND U38508 ( .A(n37295), .B(n37294), .Z(n37345) );
  XOR U38509 ( .A(a[896]), .B(n42012), .Z(n37333) );
  XNOR U38510 ( .A(n37345), .B(n37344), .Z(n37347) );
  XOR U38511 ( .A(a[894]), .B(n42085), .Z(n37334) );
  AND U38512 ( .A(a[890]), .B(b[7]), .Z(n37338) );
  XNOR U38513 ( .A(n37339), .B(n37338), .Z(n37340) );
  AND U38514 ( .A(a[898]), .B(b[0]), .Z(n37298) );
  XNOR U38515 ( .A(n37298), .B(n4071), .Z(n37300) );
  NANDN U38516 ( .A(b[0]), .B(a[897]), .Z(n37299) );
  NAND U38517 ( .A(n37300), .B(n37299), .Z(n37341) );
  XNOR U38518 ( .A(n37340), .B(n37341), .Z(n37346) );
  XOR U38519 ( .A(n37347), .B(n37346), .Z(n37325) );
  NANDN U38520 ( .A(n37302), .B(n37301), .Z(n37306) );
  NANDN U38521 ( .A(n37304), .B(n37303), .Z(n37305) );
  AND U38522 ( .A(n37306), .B(n37305), .Z(n37324) );
  XNOR U38523 ( .A(n37325), .B(n37324), .Z(n37326) );
  NANDN U38524 ( .A(n37308), .B(n37307), .Z(n37312) );
  NAND U38525 ( .A(n37310), .B(n37309), .Z(n37311) );
  NAND U38526 ( .A(n37312), .B(n37311), .Z(n37327) );
  XNOR U38527 ( .A(n37326), .B(n37327), .Z(n37318) );
  XNOR U38528 ( .A(n37319), .B(n37318), .Z(n37320) );
  XNOR U38529 ( .A(n37321), .B(n37320), .Z(n37350) );
  XNOR U38530 ( .A(sreg[1914]), .B(n37350), .Z(n37352) );
  NANDN U38531 ( .A(sreg[1913]), .B(n37313), .Z(n37317) );
  NAND U38532 ( .A(n37315), .B(n37314), .Z(n37316) );
  NAND U38533 ( .A(n37317), .B(n37316), .Z(n37351) );
  XNOR U38534 ( .A(n37352), .B(n37351), .Z(c[1914]) );
  NANDN U38535 ( .A(n37319), .B(n37318), .Z(n37323) );
  NANDN U38536 ( .A(n37321), .B(n37320), .Z(n37322) );
  AND U38537 ( .A(n37323), .B(n37322), .Z(n37358) );
  NANDN U38538 ( .A(n37325), .B(n37324), .Z(n37329) );
  NANDN U38539 ( .A(n37327), .B(n37326), .Z(n37328) );
  AND U38540 ( .A(n37329), .B(n37328), .Z(n37356) );
  NAND U38541 ( .A(n42143), .B(n37330), .Z(n37332) );
  XNOR U38542 ( .A(a[893]), .B(n4199), .Z(n37367) );
  NAND U38543 ( .A(n42144), .B(n37367), .Z(n37331) );
  AND U38544 ( .A(n37332), .B(n37331), .Z(n37382) );
  XOR U38545 ( .A(a[897]), .B(n42012), .Z(n37370) );
  XNOR U38546 ( .A(n37382), .B(n37381), .Z(n37384) );
  XOR U38547 ( .A(a[895]), .B(n42085), .Z(n37371) );
  AND U38548 ( .A(a[891]), .B(b[7]), .Z(n37375) );
  XNOR U38549 ( .A(n37376), .B(n37375), .Z(n37377) );
  AND U38550 ( .A(a[899]), .B(b[0]), .Z(n37335) );
  XNOR U38551 ( .A(n37335), .B(n4071), .Z(n37337) );
  NANDN U38552 ( .A(b[0]), .B(a[898]), .Z(n37336) );
  NAND U38553 ( .A(n37337), .B(n37336), .Z(n37378) );
  XNOR U38554 ( .A(n37377), .B(n37378), .Z(n37383) );
  XOR U38555 ( .A(n37384), .B(n37383), .Z(n37362) );
  NANDN U38556 ( .A(n37339), .B(n37338), .Z(n37343) );
  NANDN U38557 ( .A(n37341), .B(n37340), .Z(n37342) );
  AND U38558 ( .A(n37343), .B(n37342), .Z(n37361) );
  XNOR U38559 ( .A(n37362), .B(n37361), .Z(n37363) );
  NANDN U38560 ( .A(n37345), .B(n37344), .Z(n37349) );
  NAND U38561 ( .A(n37347), .B(n37346), .Z(n37348) );
  NAND U38562 ( .A(n37349), .B(n37348), .Z(n37364) );
  XNOR U38563 ( .A(n37363), .B(n37364), .Z(n37355) );
  XNOR U38564 ( .A(n37356), .B(n37355), .Z(n37357) );
  XNOR U38565 ( .A(n37358), .B(n37357), .Z(n37387) );
  XNOR U38566 ( .A(sreg[1915]), .B(n37387), .Z(n37389) );
  NANDN U38567 ( .A(sreg[1914]), .B(n37350), .Z(n37354) );
  NAND U38568 ( .A(n37352), .B(n37351), .Z(n37353) );
  NAND U38569 ( .A(n37354), .B(n37353), .Z(n37388) );
  XNOR U38570 ( .A(n37389), .B(n37388), .Z(c[1915]) );
  NANDN U38571 ( .A(n37356), .B(n37355), .Z(n37360) );
  NANDN U38572 ( .A(n37358), .B(n37357), .Z(n37359) );
  AND U38573 ( .A(n37360), .B(n37359), .Z(n37395) );
  NANDN U38574 ( .A(n37362), .B(n37361), .Z(n37366) );
  NANDN U38575 ( .A(n37364), .B(n37363), .Z(n37365) );
  AND U38576 ( .A(n37366), .B(n37365), .Z(n37393) );
  NAND U38577 ( .A(n42143), .B(n37367), .Z(n37369) );
  XNOR U38578 ( .A(a[894]), .B(n4199), .Z(n37404) );
  NAND U38579 ( .A(n42144), .B(n37404), .Z(n37368) );
  AND U38580 ( .A(n37369), .B(n37368), .Z(n37419) );
  XOR U38581 ( .A(a[898]), .B(n42012), .Z(n37407) );
  XNOR U38582 ( .A(n37419), .B(n37418), .Z(n37421) );
  XOR U38583 ( .A(a[896]), .B(n42085), .Z(n37411) );
  AND U38584 ( .A(a[892]), .B(b[7]), .Z(n37412) );
  XNOR U38585 ( .A(n37413), .B(n37412), .Z(n37414) );
  AND U38586 ( .A(a[900]), .B(b[0]), .Z(n37372) );
  XNOR U38587 ( .A(n37372), .B(n4071), .Z(n37374) );
  NANDN U38588 ( .A(b[0]), .B(a[899]), .Z(n37373) );
  NAND U38589 ( .A(n37374), .B(n37373), .Z(n37415) );
  XNOR U38590 ( .A(n37414), .B(n37415), .Z(n37420) );
  XOR U38591 ( .A(n37421), .B(n37420), .Z(n37399) );
  NANDN U38592 ( .A(n37376), .B(n37375), .Z(n37380) );
  NANDN U38593 ( .A(n37378), .B(n37377), .Z(n37379) );
  AND U38594 ( .A(n37380), .B(n37379), .Z(n37398) );
  XNOR U38595 ( .A(n37399), .B(n37398), .Z(n37400) );
  NANDN U38596 ( .A(n37382), .B(n37381), .Z(n37386) );
  NAND U38597 ( .A(n37384), .B(n37383), .Z(n37385) );
  NAND U38598 ( .A(n37386), .B(n37385), .Z(n37401) );
  XNOR U38599 ( .A(n37400), .B(n37401), .Z(n37392) );
  XNOR U38600 ( .A(n37393), .B(n37392), .Z(n37394) );
  XNOR U38601 ( .A(n37395), .B(n37394), .Z(n37424) );
  XNOR U38602 ( .A(sreg[1916]), .B(n37424), .Z(n37426) );
  NANDN U38603 ( .A(sreg[1915]), .B(n37387), .Z(n37391) );
  NAND U38604 ( .A(n37389), .B(n37388), .Z(n37390) );
  NAND U38605 ( .A(n37391), .B(n37390), .Z(n37425) );
  XNOR U38606 ( .A(n37426), .B(n37425), .Z(c[1916]) );
  NANDN U38607 ( .A(n37393), .B(n37392), .Z(n37397) );
  NANDN U38608 ( .A(n37395), .B(n37394), .Z(n37396) );
  AND U38609 ( .A(n37397), .B(n37396), .Z(n37432) );
  NANDN U38610 ( .A(n37399), .B(n37398), .Z(n37403) );
  NANDN U38611 ( .A(n37401), .B(n37400), .Z(n37402) );
  AND U38612 ( .A(n37403), .B(n37402), .Z(n37430) );
  NAND U38613 ( .A(n42143), .B(n37404), .Z(n37406) );
  XNOR U38614 ( .A(a[895]), .B(n4199), .Z(n37441) );
  NAND U38615 ( .A(n42144), .B(n37441), .Z(n37405) );
  AND U38616 ( .A(n37406), .B(n37405), .Z(n37456) );
  XOR U38617 ( .A(a[899]), .B(n42012), .Z(n37444) );
  XNOR U38618 ( .A(n37456), .B(n37455), .Z(n37458) );
  AND U38619 ( .A(a[901]), .B(b[0]), .Z(n37408) );
  XNOR U38620 ( .A(n37408), .B(n4071), .Z(n37410) );
  NANDN U38621 ( .A(b[0]), .B(a[900]), .Z(n37409) );
  NAND U38622 ( .A(n37410), .B(n37409), .Z(n37452) );
  XOR U38623 ( .A(a[897]), .B(n42085), .Z(n37445) );
  AND U38624 ( .A(a[893]), .B(b[7]), .Z(n37449) );
  XNOR U38625 ( .A(n37450), .B(n37449), .Z(n37451) );
  XNOR U38626 ( .A(n37452), .B(n37451), .Z(n37457) );
  XOR U38627 ( .A(n37458), .B(n37457), .Z(n37436) );
  NANDN U38628 ( .A(n37413), .B(n37412), .Z(n37417) );
  NANDN U38629 ( .A(n37415), .B(n37414), .Z(n37416) );
  AND U38630 ( .A(n37417), .B(n37416), .Z(n37435) );
  XNOR U38631 ( .A(n37436), .B(n37435), .Z(n37437) );
  NANDN U38632 ( .A(n37419), .B(n37418), .Z(n37423) );
  NAND U38633 ( .A(n37421), .B(n37420), .Z(n37422) );
  NAND U38634 ( .A(n37423), .B(n37422), .Z(n37438) );
  XNOR U38635 ( .A(n37437), .B(n37438), .Z(n37429) );
  XNOR U38636 ( .A(n37430), .B(n37429), .Z(n37431) );
  XNOR U38637 ( .A(n37432), .B(n37431), .Z(n37461) );
  XNOR U38638 ( .A(sreg[1917]), .B(n37461), .Z(n37463) );
  NANDN U38639 ( .A(sreg[1916]), .B(n37424), .Z(n37428) );
  NAND U38640 ( .A(n37426), .B(n37425), .Z(n37427) );
  NAND U38641 ( .A(n37428), .B(n37427), .Z(n37462) );
  XNOR U38642 ( .A(n37463), .B(n37462), .Z(c[1917]) );
  NANDN U38643 ( .A(n37430), .B(n37429), .Z(n37434) );
  NANDN U38644 ( .A(n37432), .B(n37431), .Z(n37433) );
  AND U38645 ( .A(n37434), .B(n37433), .Z(n37469) );
  NANDN U38646 ( .A(n37436), .B(n37435), .Z(n37440) );
  NANDN U38647 ( .A(n37438), .B(n37437), .Z(n37439) );
  AND U38648 ( .A(n37440), .B(n37439), .Z(n37467) );
  NAND U38649 ( .A(n42143), .B(n37441), .Z(n37443) );
  XNOR U38650 ( .A(a[896]), .B(n4199), .Z(n37478) );
  NAND U38651 ( .A(n42144), .B(n37478), .Z(n37442) );
  AND U38652 ( .A(n37443), .B(n37442), .Z(n37493) );
  XOR U38653 ( .A(a[900]), .B(n42012), .Z(n37481) );
  XNOR U38654 ( .A(n37493), .B(n37492), .Z(n37495) );
  XOR U38655 ( .A(a[898]), .B(n42085), .Z(n37482) );
  AND U38656 ( .A(a[894]), .B(b[7]), .Z(n37486) );
  XNOR U38657 ( .A(n37487), .B(n37486), .Z(n37488) );
  AND U38658 ( .A(a[902]), .B(b[0]), .Z(n37446) );
  XNOR U38659 ( .A(n37446), .B(n4071), .Z(n37448) );
  NANDN U38660 ( .A(b[0]), .B(a[901]), .Z(n37447) );
  NAND U38661 ( .A(n37448), .B(n37447), .Z(n37489) );
  XNOR U38662 ( .A(n37488), .B(n37489), .Z(n37494) );
  XOR U38663 ( .A(n37495), .B(n37494), .Z(n37473) );
  NANDN U38664 ( .A(n37450), .B(n37449), .Z(n37454) );
  NANDN U38665 ( .A(n37452), .B(n37451), .Z(n37453) );
  AND U38666 ( .A(n37454), .B(n37453), .Z(n37472) );
  XNOR U38667 ( .A(n37473), .B(n37472), .Z(n37474) );
  NANDN U38668 ( .A(n37456), .B(n37455), .Z(n37460) );
  NAND U38669 ( .A(n37458), .B(n37457), .Z(n37459) );
  NAND U38670 ( .A(n37460), .B(n37459), .Z(n37475) );
  XNOR U38671 ( .A(n37474), .B(n37475), .Z(n37466) );
  XNOR U38672 ( .A(n37467), .B(n37466), .Z(n37468) );
  XNOR U38673 ( .A(n37469), .B(n37468), .Z(n37498) );
  XNOR U38674 ( .A(sreg[1918]), .B(n37498), .Z(n37500) );
  NANDN U38675 ( .A(sreg[1917]), .B(n37461), .Z(n37465) );
  NAND U38676 ( .A(n37463), .B(n37462), .Z(n37464) );
  NAND U38677 ( .A(n37465), .B(n37464), .Z(n37499) );
  XNOR U38678 ( .A(n37500), .B(n37499), .Z(c[1918]) );
  NANDN U38679 ( .A(n37467), .B(n37466), .Z(n37471) );
  NANDN U38680 ( .A(n37469), .B(n37468), .Z(n37470) );
  AND U38681 ( .A(n37471), .B(n37470), .Z(n37506) );
  NANDN U38682 ( .A(n37473), .B(n37472), .Z(n37477) );
  NANDN U38683 ( .A(n37475), .B(n37474), .Z(n37476) );
  AND U38684 ( .A(n37477), .B(n37476), .Z(n37504) );
  NAND U38685 ( .A(n42143), .B(n37478), .Z(n37480) );
  XNOR U38686 ( .A(a[897]), .B(n4200), .Z(n37515) );
  NAND U38687 ( .A(n42144), .B(n37515), .Z(n37479) );
  AND U38688 ( .A(n37480), .B(n37479), .Z(n37530) );
  XOR U38689 ( .A(a[901]), .B(n42012), .Z(n37518) );
  XNOR U38690 ( .A(n37530), .B(n37529), .Z(n37532) );
  XOR U38691 ( .A(a[899]), .B(n42085), .Z(n37519) );
  AND U38692 ( .A(a[895]), .B(b[7]), .Z(n37523) );
  XNOR U38693 ( .A(n37524), .B(n37523), .Z(n37525) );
  AND U38694 ( .A(a[903]), .B(b[0]), .Z(n37483) );
  XNOR U38695 ( .A(n37483), .B(n4071), .Z(n37485) );
  NANDN U38696 ( .A(b[0]), .B(a[902]), .Z(n37484) );
  NAND U38697 ( .A(n37485), .B(n37484), .Z(n37526) );
  XNOR U38698 ( .A(n37525), .B(n37526), .Z(n37531) );
  XOR U38699 ( .A(n37532), .B(n37531), .Z(n37510) );
  NANDN U38700 ( .A(n37487), .B(n37486), .Z(n37491) );
  NANDN U38701 ( .A(n37489), .B(n37488), .Z(n37490) );
  AND U38702 ( .A(n37491), .B(n37490), .Z(n37509) );
  XNOR U38703 ( .A(n37510), .B(n37509), .Z(n37511) );
  NANDN U38704 ( .A(n37493), .B(n37492), .Z(n37497) );
  NAND U38705 ( .A(n37495), .B(n37494), .Z(n37496) );
  NAND U38706 ( .A(n37497), .B(n37496), .Z(n37512) );
  XNOR U38707 ( .A(n37511), .B(n37512), .Z(n37503) );
  XNOR U38708 ( .A(n37504), .B(n37503), .Z(n37505) );
  XNOR U38709 ( .A(n37506), .B(n37505), .Z(n37535) );
  XNOR U38710 ( .A(sreg[1919]), .B(n37535), .Z(n37537) );
  NANDN U38711 ( .A(sreg[1918]), .B(n37498), .Z(n37502) );
  NAND U38712 ( .A(n37500), .B(n37499), .Z(n37501) );
  NAND U38713 ( .A(n37502), .B(n37501), .Z(n37536) );
  XNOR U38714 ( .A(n37537), .B(n37536), .Z(c[1919]) );
  NANDN U38715 ( .A(n37504), .B(n37503), .Z(n37508) );
  NANDN U38716 ( .A(n37506), .B(n37505), .Z(n37507) );
  AND U38717 ( .A(n37508), .B(n37507), .Z(n37543) );
  NANDN U38718 ( .A(n37510), .B(n37509), .Z(n37514) );
  NANDN U38719 ( .A(n37512), .B(n37511), .Z(n37513) );
  AND U38720 ( .A(n37514), .B(n37513), .Z(n37541) );
  NAND U38721 ( .A(n42143), .B(n37515), .Z(n37517) );
  XNOR U38722 ( .A(a[898]), .B(n4200), .Z(n37552) );
  NAND U38723 ( .A(n42144), .B(n37552), .Z(n37516) );
  AND U38724 ( .A(n37517), .B(n37516), .Z(n37567) );
  XOR U38725 ( .A(a[902]), .B(n42012), .Z(n37555) );
  XNOR U38726 ( .A(n37567), .B(n37566), .Z(n37569) );
  XOR U38727 ( .A(a[900]), .B(n42085), .Z(n37559) );
  AND U38728 ( .A(a[896]), .B(b[7]), .Z(n37560) );
  XNOR U38729 ( .A(n37561), .B(n37560), .Z(n37562) );
  AND U38730 ( .A(a[904]), .B(b[0]), .Z(n37520) );
  XNOR U38731 ( .A(n37520), .B(n4071), .Z(n37522) );
  NANDN U38732 ( .A(b[0]), .B(a[903]), .Z(n37521) );
  NAND U38733 ( .A(n37522), .B(n37521), .Z(n37563) );
  XNOR U38734 ( .A(n37562), .B(n37563), .Z(n37568) );
  XOR U38735 ( .A(n37569), .B(n37568), .Z(n37547) );
  NANDN U38736 ( .A(n37524), .B(n37523), .Z(n37528) );
  NANDN U38737 ( .A(n37526), .B(n37525), .Z(n37527) );
  AND U38738 ( .A(n37528), .B(n37527), .Z(n37546) );
  XNOR U38739 ( .A(n37547), .B(n37546), .Z(n37548) );
  NANDN U38740 ( .A(n37530), .B(n37529), .Z(n37534) );
  NAND U38741 ( .A(n37532), .B(n37531), .Z(n37533) );
  NAND U38742 ( .A(n37534), .B(n37533), .Z(n37549) );
  XNOR U38743 ( .A(n37548), .B(n37549), .Z(n37540) );
  XNOR U38744 ( .A(n37541), .B(n37540), .Z(n37542) );
  XNOR U38745 ( .A(n37543), .B(n37542), .Z(n37572) );
  XNOR U38746 ( .A(sreg[1920]), .B(n37572), .Z(n37574) );
  NANDN U38747 ( .A(sreg[1919]), .B(n37535), .Z(n37539) );
  NAND U38748 ( .A(n37537), .B(n37536), .Z(n37538) );
  NAND U38749 ( .A(n37539), .B(n37538), .Z(n37573) );
  XNOR U38750 ( .A(n37574), .B(n37573), .Z(c[1920]) );
  NANDN U38751 ( .A(n37541), .B(n37540), .Z(n37545) );
  NANDN U38752 ( .A(n37543), .B(n37542), .Z(n37544) );
  AND U38753 ( .A(n37545), .B(n37544), .Z(n37580) );
  NANDN U38754 ( .A(n37547), .B(n37546), .Z(n37551) );
  NANDN U38755 ( .A(n37549), .B(n37548), .Z(n37550) );
  AND U38756 ( .A(n37551), .B(n37550), .Z(n37578) );
  NAND U38757 ( .A(n42143), .B(n37552), .Z(n37554) );
  XNOR U38758 ( .A(a[899]), .B(n4200), .Z(n37589) );
  NAND U38759 ( .A(n42144), .B(n37589), .Z(n37553) );
  AND U38760 ( .A(n37554), .B(n37553), .Z(n37604) );
  XOR U38761 ( .A(a[903]), .B(n42012), .Z(n37592) );
  XNOR U38762 ( .A(n37604), .B(n37603), .Z(n37606) );
  AND U38763 ( .A(a[905]), .B(b[0]), .Z(n37556) );
  XNOR U38764 ( .A(n37556), .B(n4071), .Z(n37558) );
  NANDN U38765 ( .A(b[0]), .B(a[904]), .Z(n37557) );
  NAND U38766 ( .A(n37558), .B(n37557), .Z(n37600) );
  XOR U38767 ( .A(a[901]), .B(n42085), .Z(n37596) );
  AND U38768 ( .A(a[897]), .B(b[7]), .Z(n37597) );
  XNOR U38769 ( .A(n37598), .B(n37597), .Z(n37599) );
  XNOR U38770 ( .A(n37600), .B(n37599), .Z(n37605) );
  XOR U38771 ( .A(n37606), .B(n37605), .Z(n37584) );
  NANDN U38772 ( .A(n37561), .B(n37560), .Z(n37565) );
  NANDN U38773 ( .A(n37563), .B(n37562), .Z(n37564) );
  AND U38774 ( .A(n37565), .B(n37564), .Z(n37583) );
  XNOR U38775 ( .A(n37584), .B(n37583), .Z(n37585) );
  NANDN U38776 ( .A(n37567), .B(n37566), .Z(n37571) );
  NAND U38777 ( .A(n37569), .B(n37568), .Z(n37570) );
  NAND U38778 ( .A(n37571), .B(n37570), .Z(n37586) );
  XNOR U38779 ( .A(n37585), .B(n37586), .Z(n37577) );
  XNOR U38780 ( .A(n37578), .B(n37577), .Z(n37579) );
  XNOR U38781 ( .A(n37580), .B(n37579), .Z(n37609) );
  XNOR U38782 ( .A(sreg[1921]), .B(n37609), .Z(n37611) );
  NANDN U38783 ( .A(sreg[1920]), .B(n37572), .Z(n37576) );
  NAND U38784 ( .A(n37574), .B(n37573), .Z(n37575) );
  NAND U38785 ( .A(n37576), .B(n37575), .Z(n37610) );
  XNOR U38786 ( .A(n37611), .B(n37610), .Z(c[1921]) );
  NANDN U38787 ( .A(n37578), .B(n37577), .Z(n37582) );
  NANDN U38788 ( .A(n37580), .B(n37579), .Z(n37581) );
  AND U38789 ( .A(n37582), .B(n37581), .Z(n37617) );
  NANDN U38790 ( .A(n37584), .B(n37583), .Z(n37588) );
  NANDN U38791 ( .A(n37586), .B(n37585), .Z(n37587) );
  AND U38792 ( .A(n37588), .B(n37587), .Z(n37615) );
  NAND U38793 ( .A(n42143), .B(n37589), .Z(n37591) );
  XNOR U38794 ( .A(a[900]), .B(n4200), .Z(n37626) );
  NAND U38795 ( .A(n42144), .B(n37626), .Z(n37590) );
  AND U38796 ( .A(n37591), .B(n37590), .Z(n37641) );
  XOR U38797 ( .A(a[904]), .B(n42012), .Z(n37629) );
  XNOR U38798 ( .A(n37641), .B(n37640), .Z(n37643) );
  AND U38799 ( .A(a[906]), .B(b[0]), .Z(n37593) );
  XNOR U38800 ( .A(n37593), .B(n4071), .Z(n37595) );
  NANDN U38801 ( .A(b[0]), .B(a[905]), .Z(n37594) );
  NAND U38802 ( .A(n37595), .B(n37594), .Z(n37637) );
  XOR U38803 ( .A(a[902]), .B(n42085), .Z(n37630) );
  AND U38804 ( .A(a[898]), .B(b[7]), .Z(n37634) );
  XNOR U38805 ( .A(n37635), .B(n37634), .Z(n37636) );
  XNOR U38806 ( .A(n37637), .B(n37636), .Z(n37642) );
  XOR U38807 ( .A(n37643), .B(n37642), .Z(n37621) );
  NANDN U38808 ( .A(n37598), .B(n37597), .Z(n37602) );
  NANDN U38809 ( .A(n37600), .B(n37599), .Z(n37601) );
  AND U38810 ( .A(n37602), .B(n37601), .Z(n37620) );
  XNOR U38811 ( .A(n37621), .B(n37620), .Z(n37622) );
  NANDN U38812 ( .A(n37604), .B(n37603), .Z(n37608) );
  NAND U38813 ( .A(n37606), .B(n37605), .Z(n37607) );
  NAND U38814 ( .A(n37608), .B(n37607), .Z(n37623) );
  XNOR U38815 ( .A(n37622), .B(n37623), .Z(n37614) );
  XNOR U38816 ( .A(n37615), .B(n37614), .Z(n37616) );
  XNOR U38817 ( .A(n37617), .B(n37616), .Z(n37646) );
  XNOR U38818 ( .A(sreg[1922]), .B(n37646), .Z(n37648) );
  NANDN U38819 ( .A(sreg[1921]), .B(n37609), .Z(n37613) );
  NAND U38820 ( .A(n37611), .B(n37610), .Z(n37612) );
  NAND U38821 ( .A(n37613), .B(n37612), .Z(n37647) );
  XNOR U38822 ( .A(n37648), .B(n37647), .Z(c[1922]) );
  NANDN U38823 ( .A(n37615), .B(n37614), .Z(n37619) );
  NANDN U38824 ( .A(n37617), .B(n37616), .Z(n37618) );
  AND U38825 ( .A(n37619), .B(n37618), .Z(n37654) );
  NANDN U38826 ( .A(n37621), .B(n37620), .Z(n37625) );
  NANDN U38827 ( .A(n37623), .B(n37622), .Z(n37624) );
  AND U38828 ( .A(n37625), .B(n37624), .Z(n37652) );
  NAND U38829 ( .A(n42143), .B(n37626), .Z(n37628) );
  XNOR U38830 ( .A(a[901]), .B(n4200), .Z(n37663) );
  NAND U38831 ( .A(n42144), .B(n37663), .Z(n37627) );
  AND U38832 ( .A(n37628), .B(n37627), .Z(n37678) );
  XOR U38833 ( .A(a[905]), .B(n42012), .Z(n37666) );
  XNOR U38834 ( .A(n37678), .B(n37677), .Z(n37680) );
  XOR U38835 ( .A(a[903]), .B(n42085), .Z(n37670) );
  AND U38836 ( .A(a[899]), .B(b[7]), .Z(n37671) );
  XNOR U38837 ( .A(n37672), .B(n37671), .Z(n37673) );
  AND U38838 ( .A(a[907]), .B(b[0]), .Z(n37631) );
  XNOR U38839 ( .A(n37631), .B(n4071), .Z(n37633) );
  NANDN U38840 ( .A(b[0]), .B(a[906]), .Z(n37632) );
  NAND U38841 ( .A(n37633), .B(n37632), .Z(n37674) );
  XNOR U38842 ( .A(n37673), .B(n37674), .Z(n37679) );
  XOR U38843 ( .A(n37680), .B(n37679), .Z(n37658) );
  NANDN U38844 ( .A(n37635), .B(n37634), .Z(n37639) );
  NANDN U38845 ( .A(n37637), .B(n37636), .Z(n37638) );
  AND U38846 ( .A(n37639), .B(n37638), .Z(n37657) );
  XNOR U38847 ( .A(n37658), .B(n37657), .Z(n37659) );
  NANDN U38848 ( .A(n37641), .B(n37640), .Z(n37645) );
  NAND U38849 ( .A(n37643), .B(n37642), .Z(n37644) );
  NAND U38850 ( .A(n37645), .B(n37644), .Z(n37660) );
  XNOR U38851 ( .A(n37659), .B(n37660), .Z(n37651) );
  XNOR U38852 ( .A(n37652), .B(n37651), .Z(n37653) );
  XNOR U38853 ( .A(n37654), .B(n37653), .Z(n37683) );
  XNOR U38854 ( .A(sreg[1923]), .B(n37683), .Z(n37685) );
  NANDN U38855 ( .A(sreg[1922]), .B(n37646), .Z(n37650) );
  NAND U38856 ( .A(n37648), .B(n37647), .Z(n37649) );
  NAND U38857 ( .A(n37650), .B(n37649), .Z(n37684) );
  XNOR U38858 ( .A(n37685), .B(n37684), .Z(c[1923]) );
  NANDN U38859 ( .A(n37652), .B(n37651), .Z(n37656) );
  NANDN U38860 ( .A(n37654), .B(n37653), .Z(n37655) );
  AND U38861 ( .A(n37656), .B(n37655), .Z(n37691) );
  NANDN U38862 ( .A(n37658), .B(n37657), .Z(n37662) );
  NANDN U38863 ( .A(n37660), .B(n37659), .Z(n37661) );
  AND U38864 ( .A(n37662), .B(n37661), .Z(n37689) );
  NAND U38865 ( .A(n42143), .B(n37663), .Z(n37665) );
  XNOR U38866 ( .A(a[902]), .B(n4200), .Z(n37700) );
  NAND U38867 ( .A(n42144), .B(n37700), .Z(n37664) );
  AND U38868 ( .A(n37665), .B(n37664), .Z(n37715) );
  XOR U38869 ( .A(a[906]), .B(n42012), .Z(n37703) );
  XNOR U38870 ( .A(n37715), .B(n37714), .Z(n37717) );
  AND U38871 ( .A(a[908]), .B(b[0]), .Z(n37667) );
  XNOR U38872 ( .A(n37667), .B(n4071), .Z(n37669) );
  NANDN U38873 ( .A(b[0]), .B(a[907]), .Z(n37668) );
  NAND U38874 ( .A(n37669), .B(n37668), .Z(n37711) );
  XOR U38875 ( .A(a[904]), .B(n42085), .Z(n37707) );
  AND U38876 ( .A(a[900]), .B(b[7]), .Z(n37708) );
  XNOR U38877 ( .A(n37709), .B(n37708), .Z(n37710) );
  XNOR U38878 ( .A(n37711), .B(n37710), .Z(n37716) );
  XOR U38879 ( .A(n37717), .B(n37716), .Z(n37695) );
  NANDN U38880 ( .A(n37672), .B(n37671), .Z(n37676) );
  NANDN U38881 ( .A(n37674), .B(n37673), .Z(n37675) );
  AND U38882 ( .A(n37676), .B(n37675), .Z(n37694) );
  XNOR U38883 ( .A(n37695), .B(n37694), .Z(n37696) );
  NANDN U38884 ( .A(n37678), .B(n37677), .Z(n37682) );
  NAND U38885 ( .A(n37680), .B(n37679), .Z(n37681) );
  NAND U38886 ( .A(n37682), .B(n37681), .Z(n37697) );
  XNOR U38887 ( .A(n37696), .B(n37697), .Z(n37688) );
  XNOR U38888 ( .A(n37689), .B(n37688), .Z(n37690) );
  XNOR U38889 ( .A(n37691), .B(n37690), .Z(n37720) );
  XNOR U38890 ( .A(sreg[1924]), .B(n37720), .Z(n37722) );
  NANDN U38891 ( .A(sreg[1923]), .B(n37683), .Z(n37687) );
  NAND U38892 ( .A(n37685), .B(n37684), .Z(n37686) );
  NAND U38893 ( .A(n37687), .B(n37686), .Z(n37721) );
  XNOR U38894 ( .A(n37722), .B(n37721), .Z(c[1924]) );
  NANDN U38895 ( .A(n37689), .B(n37688), .Z(n37693) );
  NANDN U38896 ( .A(n37691), .B(n37690), .Z(n37692) );
  AND U38897 ( .A(n37693), .B(n37692), .Z(n37728) );
  NANDN U38898 ( .A(n37695), .B(n37694), .Z(n37699) );
  NANDN U38899 ( .A(n37697), .B(n37696), .Z(n37698) );
  AND U38900 ( .A(n37699), .B(n37698), .Z(n37726) );
  NAND U38901 ( .A(n42143), .B(n37700), .Z(n37702) );
  XNOR U38902 ( .A(a[903]), .B(n4200), .Z(n37737) );
  NAND U38903 ( .A(n42144), .B(n37737), .Z(n37701) );
  AND U38904 ( .A(n37702), .B(n37701), .Z(n37752) );
  XOR U38905 ( .A(a[907]), .B(n42012), .Z(n37740) );
  XNOR U38906 ( .A(n37752), .B(n37751), .Z(n37754) );
  AND U38907 ( .A(a[909]), .B(b[0]), .Z(n37704) );
  XNOR U38908 ( .A(n37704), .B(n4071), .Z(n37706) );
  NANDN U38909 ( .A(b[0]), .B(a[908]), .Z(n37705) );
  NAND U38910 ( .A(n37706), .B(n37705), .Z(n37748) );
  XOR U38911 ( .A(a[905]), .B(n42085), .Z(n37744) );
  AND U38912 ( .A(a[901]), .B(b[7]), .Z(n37745) );
  XNOR U38913 ( .A(n37746), .B(n37745), .Z(n37747) );
  XNOR U38914 ( .A(n37748), .B(n37747), .Z(n37753) );
  XOR U38915 ( .A(n37754), .B(n37753), .Z(n37732) );
  NANDN U38916 ( .A(n37709), .B(n37708), .Z(n37713) );
  NANDN U38917 ( .A(n37711), .B(n37710), .Z(n37712) );
  AND U38918 ( .A(n37713), .B(n37712), .Z(n37731) );
  XNOR U38919 ( .A(n37732), .B(n37731), .Z(n37733) );
  NANDN U38920 ( .A(n37715), .B(n37714), .Z(n37719) );
  NAND U38921 ( .A(n37717), .B(n37716), .Z(n37718) );
  NAND U38922 ( .A(n37719), .B(n37718), .Z(n37734) );
  XNOR U38923 ( .A(n37733), .B(n37734), .Z(n37725) );
  XNOR U38924 ( .A(n37726), .B(n37725), .Z(n37727) );
  XNOR U38925 ( .A(n37728), .B(n37727), .Z(n37757) );
  XNOR U38926 ( .A(sreg[1925]), .B(n37757), .Z(n37759) );
  NANDN U38927 ( .A(sreg[1924]), .B(n37720), .Z(n37724) );
  NAND U38928 ( .A(n37722), .B(n37721), .Z(n37723) );
  NAND U38929 ( .A(n37724), .B(n37723), .Z(n37758) );
  XNOR U38930 ( .A(n37759), .B(n37758), .Z(c[1925]) );
  NANDN U38931 ( .A(n37726), .B(n37725), .Z(n37730) );
  NANDN U38932 ( .A(n37728), .B(n37727), .Z(n37729) );
  AND U38933 ( .A(n37730), .B(n37729), .Z(n37765) );
  NANDN U38934 ( .A(n37732), .B(n37731), .Z(n37736) );
  NANDN U38935 ( .A(n37734), .B(n37733), .Z(n37735) );
  AND U38936 ( .A(n37736), .B(n37735), .Z(n37763) );
  NAND U38937 ( .A(n42143), .B(n37737), .Z(n37739) );
  XNOR U38938 ( .A(a[904]), .B(n4201), .Z(n37774) );
  NAND U38939 ( .A(n42144), .B(n37774), .Z(n37738) );
  AND U38940 ( .A(n37739), .B(n37738), .Z(n37789) );
  XOR U38941 ( .A(a[908]), .B(n42012), .Z(n37777) );
  XNOR U38942 ( .A(n37789), .B(n37788), .Z(n37791) );
  AND U38943 ( .A(a[910]), .B(b[0]), .Z(n37741) );
  XNOR U38944 ( .A(n37741), .B(n4071), .Z(n37743) );
  NANDN U38945 ( .A(b[0]), .B(a[909]), .Z(n37742) );
  NAND U38946 ( .A(n37743), .B(n37742), .Z(n37785) );
  XOR U38947 ( .A(a[906]), .B(n42085), .Z(n37778) );
  AND U38948 ( .A(a[902]), .B(b[7]), .Z(n37782) );
  XNOR U38949 ( .A(n37783), .B(n37782), .Z(n37784) );
  XNOR U38950 ( .A(n37785), .B(n37784), .Z(n37790) );
  XOR U38951 ( .A(n37791), .B(n37790), .Z(n37769) );
  NANDN U38952 ( .A(n37746), .B(n37745), .Z(n37750) );
  NANDN U38953 ( .A(n37748), .B(n37747), .Z(n37749) );
  AND U38954 ( .A(n37750), .B(n37749), .Z(n37768) );
  XNOR U38955 ( .A(n37769), .B(n37768), .Z(n37770) );
  NANDN U38956 ( .A(n37752), .B(n37751), .Z(n37756) );
  NAND U38957 ( .A(n37754), .B(n37753), .Z(n37755) );
  NAND U38958 ( .A(n37756), .B(n37755), .Z(n37771) );
  XNOR U38959 ( .A(n37770), .B(n37771), .Z(n37762) );
  XNOR U38960 ( .A(n37763), .B(n37762), .Z(n37764) );
  XNOR U38961 ( .A(n37765), .B(n37764), .Z(n37794) );
  XNOR U38962 ( .A(sreg[1926]), .B(n37794), .Z(n37796) );
  NANDN U38963 ( .A(sreg[1925]), .B(n37757), .Z(n37761) );
  NAND U38964 ( .A(n37759), .B(n37758), .Z(n37760) );
  NAND U38965 ( .A(n37761), .B(n37760), .Z(n37795) );
  XNOR U38966 ( .A(n37796), .B(n37795), .Z(c[1926]) );
  NANDN U38967 ( .A(n37763), .B(n37762), .Z(n37767) );
  NANDN U38968 ( .A(n37765), .B(n37764), .Z(n37766) );
  AND U38969 ( .A(n37767), .B(n37766), .Z(n37802) );
  NANDN U38970 ( .A(n37769), .B(n37768), .Z(n37773) );
  NANDN U38971 ( .A(n37771), .B(n37770), .Z(n37772) );
  AND U38972 ( .A(n37773), .B(n37772), .Z(n37800) );
  NAND U38973 ( .A(n42143), .B(n37774), .Z(n37776) );
  XNOR U38974 ( .A(a[905]), .B(n4201), .Z(n37811) );
  NAND U38975 ( .A(n42144), .B(n37811), .Z(n37775) );
  AND U38976 ( .A(n37776), .B(n37775), .Z(n37826) );
  XOR U38977 ( .A(a[909]), .B(n42012), .Z(n37814) );
  XNOR U38978 ( .A(n37826), .B(n37825), .Z(n37828) );
  XOR U38979 ( .A(a[907]), .B(n42085), .Z(n37818) );
  AND U38980 ( .A(a[903]), .B(b[7]), .Z(n37819) );
  XNOR U38981 ( .A(n37820), .B(n37819), .Z(n37821) );
  AND U38982 ( .A(a[911]), .B(b[0]), .Z(n37779) );
  XNOR U38983 ( .A(n37779), .B(n4071), .Z(n37781) );
  NANDN U38984 ( .A(b[0]), .B(a[910]), .Z(n37780) );
  NAND U38985 ( .A(n37781), .B(n37780), .Z(n37822) );
  XNOR U38986 ( .A(n37821), .B(n37822), .Z(n37827) );
  XOR U38987 ( .A(n37828), .B(n37827), .Z(n37806) );
  NANDN U38988 ( .A(n37783), .B(n37782), .Z(n37787) );
  NANDN U38989 ( .A(n37785), .B(n37784), .Z(n37786) );
  AND U38990 ( .A(n37787), .B(n37786), .Z(n37805) );
  XNOR U38991 ( .A(n37806), .B(n37805), .Z(n37807) );
  NANDN U38992 ( .A(n37789), .B(n37788), .Z(n37793) );
  NAND U38993 ( .A(n37791), .B(n37790), .Z(n37792) );
  NAND U38994 ( .A(n37793), .B(n37792), .Z(n37808) );
  XNOR U38995 ( .A(n37807), .B(n37808), .Z(n37799) );
  XNOR U38996 ( .A(n37800), .B(n37799), .Z(n37801) );
  XNOR U38997 ( .A(n37802), .B(n37801), .Z(n37831) );
  XNOR U38998 ( .A(sreg[1927]), .B(n37831), .Z(n37833) );
  NANDN U38999 ( .A(sreg[1926]), .B(n37794), .Z(n37798) );
  NAND U39000 ( .A(n37796), .B(n37795), .Z(n37797) );
  NAND U39001 ( .A(n37798), .B(n37797), .Z(n37832) );
  XNOR U39002 ( .A(n37833), .B(n37832), .Z(c[1927]) );
  NANDN U39003 ( .A(n37800), .B(n37799), .Z(n37804) );
  NANDN U39004 ( .A(n37802), .B(n37801), .Z(n37803) );
  AND U39005 ( .A(n37804), .B(n37803), .Z(n37839) );
  NANDN U39006 ( .A(n37806), .B(n37805), .Z(n37810) );
  NANDN U39007 ( .A(n37808), .B(n37807), .Z(n37809) );
  AND U39008 ( .A(n37810), .B(n37809), .Z(n37837) );
  NAND U39009 ( .A(n42143), .B(n37811), .Z(n37813) );
  XNOR U39010 ( .A(a[906]), .B(n4201), .Z(n37848) );
  NAND U39011 ( .A(n42144), .B(n37848), .Z(n37812) );
  AND U39012 ( .A(n37813), .B(n37812), .Z(n37863) );
  XOR U39013 ( .A(a[910]), .B(n42012), .Z(n37851) );
  XNOR U39014 ( .A(n37863), .B(n37862), .Z(n37865) );
  AND U39015 ( .A(a[912]), .B(b[0]), .Z(n37815) );
  XNOR U39016 ( .A(n37815), .B(n4071), .Z(n37817) );
  NANDN U39017 ( .A(b[0]), .B(a[911]), .Z(n37816) );
  NAND U39018 ( .A(n37817), .B(n37816), .Z(n37859) );
  XOR U39019 ( .A(a[908]), .B(n42085), .Z(n37855) );
  AND U39020 ( .A(a[904]), .B(b[7]), .Z(n37856) );
  XNOR U39021 ( .A(n37857), .B(n37856), .Z(n37858) );
  XNOR U39022 ( .A(n37859), .B(n37858), .Z(n37864) );
  XOR U39023 ( .A(n37865), .B(n37864), .Z(n37843) );
  NANDN U39024 ( .A(n37820), .B(n37819), .Z(n37824) );
  NANDN U39025 ( .A(n37822), .B(n37821), .Z(n37823) );
  AND U39026 ( .A(n37824), .B(n37823), .Z(n37842) );
  XNOR U39027 ( .A(n37843), .B(n37842), .Z(n37844) );
  NANDN U39028 ( .A(n37826), .B(n37825), .Z(n37830) );
  NAND U39029 ( .A(n37828), .B(n37827), .Z(n37829) );
  NAND U39030 ( .A(n37830), .B(n37829), .Z(n37845) );
  XNOR U39031 ( .A(n37844), .B(n37845), .Z(n37836) );
  XNOR U39032 ( .A(n37837), .B(n37836), .Z(n37838) );
  XNOR U39033 ( .A(n37839), .B(n37838), .Z(n37868) );
  XNOR U39034 ( .A(sreg[1928]), .B(n37868), .Z(n37870) );
  NANDN U39035 ( .A(sreg[1927]), .B(n37831), .Z(n37835) );
  NAND U39036 ( .A(n37833), .B(n37832), .Z(n37834) );
  NAND U39037 ( .A(n37835), .B(n37834), .Z(n37869) );
  XNOR U39038 ( .A(n37870), .B(n37869), .Z(c[1928]) );
  NANDN U39039 ( .A(n37837), .B(n37836), .Z(n37841) );
  NANDN U39040 ( .A(n37839), .B(n37838), .Z(n37840) );
  AND U39041 ( .A(n37841), .B(n37840), .Z(n37876) );
  NANDN U39042 ( .A(n37843), .B(n37842), .Z(n37847) );
  NANDN U39043 ( .A(n37845), .B(n37844), .Z(n37846) );
  AND U39044 ( .A(n37847), .B(n37846), .Z(n37874) );
  NAND U39045 ( .A(n42143), .B(n37848), .Z(n37850) );
  XNOR U39046 ( .A(a[907]), .B(n4201), .Z(n37885) );
  NAND U39047 ( .A(n42144), .B(n37885), .Z(n37849) );
  AND U39048 ( .A(n37850), .B(n37849), .Z(n37900) );
  XOR U39049 ( .A(a[911]), .B(n42012), .Z(n37888) );
  XNOR U39050 ( .A(n37900), .B(n37899), .Z(n37902) );
  AND U39051 ( .A(a[913]), .B(b[0]), .Z(n37852) );
  XNOR U39052 ( .A(n37852), .B(n4071), .Z(n37854) );
  NANDN U39053 ( .A(b[0]), .B(a[912]), .Z(n37853) );
  NAND U39054 ( .A(n37854), .B(n37853), .Z(n37896) );
  XOR U39055 ( .A(a[909]), .B(n42085), .Z(n37889) );
  AND U39056 ( .A(a[905]), .B(b[7]), .Z(n37893) );
  XNOR U39057 ( .A(n37894), .B(n37893), .Z(n37895) );
  XNOR U39058 ( .A(n37896), .B(n37895), .Z(n37901) );
  XOR U39059 ( .A(n37902), .B(n37901), .Z(n37880) );
  NANDN U39060 ( .A(n37857), .B(n37856), .Z(n37861) );
  NANDN U39061 ( .A(n37859), .B(n37858), .Z(n37860) );
  AND U39062 ( .A(n37861), .B(n37860), .Z(n37879) );
  XNOR U39063 ( .A(n37880), .B(n37879), .Z(n37881) );
  NANDN U39064 ( .A(n37863), .B(n37862), .Z(n37867) );
  NAND U39065 ( .A(n37865), .B(n37864), .Z(n37866) );
  NAND U39066 ( .A(n37867), .B(n37866), .Z(n37882) );
  XNOR U39067 ( .A(n37881), .B(n37882), .Z(n37873) );
  XNOR U39068 ( .A(n37874), .B(n37873), .Z(n37875) );
  XNOR U39069 ( .A(n37876), .B(n37875), .Z(n37905) );
  XNOR U39070 ( .A(sreg[1929]), .B(n37905), .Z(n37907) );
  NANDN U39071 ( .A(sreg[1928]), .B(n37868), .Z(n37872) );
  NAND U39072 ( .A(n37870), .B(n37869), .Z(n37871) );
  NAND U39073 ( .A(n37872), .B(n37871), .Z(n37906) );
  XNOR U39074 ( .A(n37907), .B(n37906), .Z(c[1929]) );
  NANDN U39075 ( .A(n37874), .B(n37873), .Z(n37878) );
  NANDN U39076 ( .A(n37876), .B(n37875), .Z(n37877) );
  AND U39077 ( .A(n37878), .B(n37877), .Z(n37913) );
  NANDN U39078 ( .A(n37880), .B(n37879), .Z(n37884) );
  NANDN U39079 ( .A(n37882), .B(n37881), .Z(n37883) );
  AND U39080 ( .A(n37884), .B(n37883), .Z(n37911) );
  NAND U39081 ( .A(n42143), .B(n37885), .Z(n37887) );
  XNOR U39082 ( .A(a[908]), .B(n4201), .Z(n37922) );
  NAND U39083 ( .A(n42144), .B(n37922), .Z(n37886) );
  AND U39084 ( .A(n37887), .B(n37886), .Z(n37937) );
  XOR U39085 ( .A(a[912]), .B(n42012), .Z(n37925) );
  XNOR U39086 ( .A(n37937), .B(n37936), .Z(n37939) );
  XOR U39087 ( .A(a[910]), .B(n42085), .Z(n37929) );
  AND U39088 ( .A(a[906]), .B(b[7]), .Z(n37930) );
  XNOR U39089 ( .A(n37931), .B(n37930), .Z(n37932) );
  AND U39090 ( .A(a[914]), .B(b[0]), .Z(n37890) );
  XNOR U39091 ( .A(n37890), .B(n4071), .Z(n37892) );
  NANDN U39092 ( .A(b[0]), .B(a[913]), .Z(n37891) );
  NAND U39093 ( .A(n37892), .B(n37891), .Z(n37933) );
  XNOR U39094 ( .A(n37932), .B(n37933), .Z(n37938) );
  XOR U39095 ( .A(n37939), .B(n37938), .Z(n37917) );
  NANDN U39096 ( .A(n37894), .B(n37893), .Z(n37898) );
  NANDN U39097 ( .A(n37896), .B(n37895), .Z(n37897) );
  AND U39098 ( .A(n37898), .B(n37897), .Z(n37916) );
  XNOR U39099 ( .A(n37917), .B(n37916), .Z(n37918) );
  NANDN U39100 ( .A(n37900), .B(n37899), .Z(n37904) );
  NAND U39101 ( .A(n37902), .B(n37901), .Z(n37903) );
  NAND U39102 ( .A(n37904), .B(n37903), .Z(n37919) );
  XNOR U39103 ( .A(n37918), .B(n37919), .Z(n37910) );
  XNOR U39104 ( .A(n37911), .B(n37910), .Z(n37912) );
  XNOR U39105 ( .A(n37913), .B(n37912), .Z(n37942) );
  XNOR U39106 ( .A(sreg[1930]), .B(n37942), .Z(n37944) );
  NANDN U39107 ( .A(sreg[1929]), .B(n37905), .Z(n37909) );
  NAND U39108 ( .A(n37907), .B(n37906), .Z(n37908) );
  NAND U39109 ( .A(n37909), .B(n37908), .Z(n37943) );
  XNOR U39110 ( .A(n37944), .B(n37943), .Z(c[1930]) );
  NANDN U39111 ( .A(n37911), .B(n37910), .Z(n37915) );
  NANDN U39112 ( .A(n37913), .B(n37912), .Z(n37914) );
  AND U39113 ( .A(n37915), .B(n37914), .Z(n37950) );
  NANDN U39114 ( .A(n37917), .B(n37916), .Z(n37921) );
  NANDN U39115 ( .A(n37919), .B(n37918), .Z(n37920) );
  AND U39116 ( .A(n37921), .B(n37920), .Z(n37948) );
  NAND U39117 ( .A(n42143), .B(n37922), .Z(n37924) );
  XNOR U39118 ( .A(a[909]), .B(n4201), .Z(n37959) );
  NAND U39119 ( .A(n42144), .B(n37959), .Z(n37923) );
  AND U39120 ( .A(n37924), .B(n37923), .Z(n37974) );
  XOR U39121 ( .A(a[913]), .B(n42012), .Z(n37962) );
  XNOR U39122 ( .A(n37974), .B(n37973), .Z(n37976) );
  AND U39123 ( .A(a[915]), .B(b[0]), .Z(n37926) );
  XNOR U39124 ( .A(n37926), .B(n4071), .Z(n37928) );
  NANDN U39125 ( .A(b[0]), .B(a[914]), .Z(n37927) );
  NAND U39126 ( .A(n37928), .B(n37927), .Z(n37970) );
  XOR U39127 ( .A(a[911]), .B(n42085), .Z(n37963) );
  AND U39128 ( .A(a[907]), .B(b[7]), .Z(n37967) );
  XNOR U39129 ( .A(n37968), .B(n37967), .Z(n37969) );
  XNOR U39130 ( .A(n37970), .B(n37969), .Z(n37975) );
  XOR U39131 ( .A(n37976), .B(n37975), .Z(n37954) );
  NANDN U39132 ( .A(n37931), .B(n37930), .Z(n37935) );
  NANDN U39133 ( .A(n37933), .B(n37932), .Z(n37934) );
  AND U39134 ( .A(n37935), .B(n37934), .Z(n37953) );
  XNOR U39135 ( .A(n37954), .B(n37953), .Z(n37955) );
  NANDN U39136 ( .A(n37937), .B(n37936), .Z(n37941) );
  NAND U39137 ( .A(n37939), .B(n37938), .Z(n37940) );
  NAND U39138 ( .A(n37941), .B(n37940), .Z(n37956) );
  XNOR U39139 ( .A(n37955), .B(n37956), .Z(n37947) );
  XNOR U39140 ( .A(n37948), .B(n37947), .Z(n37949) );
  XNOR U39141 ( .A(n37950), .B(n37949), .Z(n37979) );
  XNOR U39142 ( .A(sreg[1931]), .B(n37979), .Z(n37981) );
  NANDN U39143 ( .A(sreg[1930]), .B(n37942), .Z(n37946) );
  NAND U39144 ( .A(n37944), .B(n37943), .Z(n37945) );
  NAND U39145 ( .A(n37946), .B(n37945), .Z(n37980) );
  XNOR U39146 ( .A(n37981), .B(n37980), .Z(c[1931]) );
  NANDN U39147 ( .A(n37948), .B(n37947), .Z(n37952) );
  NANDN U39148 ( .A(n37950), .B(n37949), .Z(n37951) );
  AND U39149 ( .A(n37952), .B(n37951), .Z(n37987) );
  NANDN U39150 ( .A(n37954), .B(n37953), .Z(n37958) );
  NANDN U39151 ( .A(n37956), .B(n37955), .Z(n37957) );
  AND U39152 ( .A(n37958), .B(n37957), .Z(n37985) );
  NAND U39153 ( .A(n42143), .B(n37959), .Z(n37961) );
  XNOR U39154 ( .A(a[910]), .B(n4201), .Z(n37996) );
  NAND U39155 ( .A(n42144), .B(n37996), .Z(n37960) );
  AND U39156 ( .A(n37961), .B(n37960), .Z(n38011) );
  XOR U39157 ( .A(a[914]), .B(n42012), .Z(n37999) );
  XNOR U39158 ( .A(n38011), .B(n38010), .Z(n38013) );
  XOR U39159 ( .A(a[912]), .B(n42085), .Z(n38003) );
  AND U39160 ( .A(a[908]), .B(b[7]), .Z(n38004) );
  XNOR U39161 ( .A(n38005), .B(n38004), .Z(n38006) );
  AND U39162 ( .A(a[916]), .B(b[0]), .Z(n37964) );
  XNOR U39163 ( .A(n37964), .B(n4071), .Z(n37966) );
  NANDN U39164 ( .A(b[0]), .B(a[915]), .Z(n37965) );
  NAND U39165 ( .A(n37966), .B(n37965), .Z(n38007) );
  XNOR U39166 ( .A(n38006), .B(n38007), .Z(n38012) );
  XOR U39167 ( .A(n38013), .B(n38012), .Z(n37991) );
  NANDN U39168 ( .A(n37968), .B(n37967), .Z(n37972) );
  NANDN U39169 ( .A(n37970), .B(n37969), .Z(n37971) );
  AND U39170 ( .A(n37972), .B(n37971), .Z(n37990) );
  XNOR U39171 ( .A(n37991), .B(n37990), .Z(n37992) );
  NANDN U39172 ( .A(n37974), .B(n37973), .Z(n37978) );
  NAND U39173 ( .A(n37976), .B(n37975), .Z(n37977) );
  NAND U39174 ( .A(n37978), .B(n37977), .Z(n37993) );
  XNOR U39175 ( .A(n37992), .B(n37993), .Z(n37984) );
  XNOR U39176 ( .A(n37985), .B(n37984), .Z(n37986) );
  XNOR U39177 ( .A(n37987), .B(n37986), .Z(n38016) );
  XNOR U39178 ( .A(sreg[1932]), .B(n38016), .Z(n38018) );
  NANDN U39179 ( .A(sreg[1931]), .B(n37979), .Z(n37983) );
  NAND U39180 ( .A(n37981), .B(n37980), .Z(n37982) );
  NAND U39181 ( .A(n37983), .B(n37982), .Z(n38017) );
  XNOR U39182 ( .A(n38018), .B(n38017), .Z(c[1932]) );
  NANDN U39183 ( .A(n37985), .B(n37984), .Z(n37989) );
  NANDN U39184 ( .A(n37987), .B(n37986), .Z(n37988) );
  AND U39185 ( .A(n37989), .B(n37988), .Z(n38024) );
  NANDN U39186 ( .A(n37991), .B(n37990), .Z(n37995) );
  NANDN U39187 ( .A(n37993), .B(n37992), .Z(n37994) );
  AND U39188 ( .A(n37995), .B(n37994), .Z(n38022) );
  NAND U39189 ( .A(n42143), .B(n37996), .Z(n37998) );
  XNOR U39190 ( .A(a[911]), .B(n4202), .Z(n38033) );
  NAND U39191 ( .A(n42144), .B(n38033), .Z(n37997) );
  AND U39192 ( .A(n37998), .B(n37997), .Z(n38048) );
  XOR U39193 ( .A(a[915]), .B(n42012), .Z(n38036) );
  XNOR U39194 ( .A(n38048), .B(n38047), .Z(n38050) );
  AND U39195 ( .A(a[917]), .B(b[0]), .Z(n38000) );
  XNOR U39196 ( .A(n38000), .B(n4071), .Z(n38002) );
  NANDN U39197 ( .A(b[0]), .B(a[916]), .Z(n38001) );
  NAND U39198 ( .A(n38002), .B(n38001), .Z(n38044) );
  XOR U39199 ( .A(a[913]), .B(n42085), .Z(n38040) );
  AND U39200 ( .A(a[909]), .B(b[7]), .Z(n38041) );
  XNOR U39201 ( .A(n38042), .B(n38041), .Z(n38043) );
  XNOR U39202 ( .A(n38044), .B(n38043), .Z(n38049) );
  XOR U39203 ( .A(n38050), .B(n38049), .Z(n38028) );
  NANDN U39204 ( .A(n38005), .B(n38004), .Z(n38009) );
  NANDN U39205 ( .A(n38007), .B(n38006), .Z(n38008) );
  AND U39206 ( .A(n38009), .B(n38008), .Z(n38027) );
  XNOR U39207 ( .A(n38028), .B(n38027), .Z(n38029) );
  NANDN U39208 ( .A(n38011), .B(n38010), .Z(n38015) );
  NAND U39209 ( .A(n38013), .B(n38012), .Z(n38014) );
  NAND U39210 ( .A(n38015), .B(n38014), .Z(n38030) );
  XNOR U39211 ( .A(n38029), .B(n38030), .Z(n38021) );
  XNOR U39212 ( .A(n38022), .B(n38021), .Z(n38023) );
  XNOR U39213 ( .A(n38024), .B(n38023), .Z(n38053) );
  XNOR U39214 ( .A(sreg[1933]), .B(n38053), .Z(n38055) );
  NANDN U39215 ( .A(sreg[1932]), .B(n38016), .Z(n38020) );
  NAND U39216 ( .A(n38018), .B(n38017), .Z(n38019) );
  NAND U39217 ( .A(n38020), .B(n38019), .Z(n38054) );
  XNOR U39218 ( .A(n38055), .B(n38054), .Z(c[1933]) );
  NANDN U39219 ( .A(n38022), .B(n38021), .Z(n38026) );
  NANDN U39220 ( .A(n38024), .B(n38023), .Z(n38025) );
  AND U39221 ( .A(n38026), .B(n38025), .Z(n38061) );
  NANDN U39222 ( .A(n38028), .B(n38027), .Z(n38032) );
  NANDN U39223 ( .A(n38030), .B(n38029), .Z(n38031) );
  AND U39224 ( .A(n38032), .B(n38031), .Z(n38059) );
  NAND U39225 ( .A(n42143), .B(n38033), .Z(n38035) );
  XNOR U39226 ( .A(a[912]), .B(n4202), .Z(n38070) );
  NAND U39227 ( .A(n42144), .B(n38070), .Z(n38034) );
  AND U39228 ( .A(n38035), .B(n38034), .Z(n38085) );
  XOR U39229 ( .A(a[916]), .B(n42012), .Z(n38073) );
  XNOR U39230 ( .A(n38085), .B(n38084), .Z(n38087) );
  AND U39231 ( .A(a[918]), .B(b[0]), .Z(n38037) );
  XNOR U39232 ( .A(n38037), .B(n4071), .Z(n38039) );
  NANDN U39233 ( .A(b[0]), .B(a[917]), .Z(n38038) );
  NAND U39234 ( .A(n38039), .B(n38038), .Z(n38081) );
  XOR U39235 ( .A(a[914]), .B(n42085), .Z(n38077) );
  AND U39236 ( .A(a[910]), .B(b[7]), .Z(n38078) );
  XNOR U39237 ( .A(n38079), .B(n38078), .Z(n38080) );
  XNOR U39238 ( .A(n38081), .B(n38080), .Z(n38086) );
  XOR U39239 ( .A(n38087), .B(n38086), .Z(n38065) );
  NANDN U39240 ( .A(n38042), .B(n38041), .Z(n38046) );
  NANDN U39241 ( .A(n38044), .B(n38043), .Z(n38045) );
  AND U39242 ( .A(n38046), .B(n38045), .Z(n38064) );
  XNOR U39243 ( .A(n38065), .B(n38064), .Z(n38066) );
  NANDN U39244 ( .A(n38048), .B(n38047), .Z(n38052) );
  NAND U39245 ( .A(n38050), .B(n38049), .Z(n38051) );
  NAND U39246 ( .A(n38052), .B(n38051), .Z(n38067) );
  XNOR U39247 ( .A(n38066), .B(n38067), .Z(n38058) );
  XNOR U39248 ( .A(n38059), .B(n38058), .Z(n38060) );
  XNOR U39249 ( .A(n38061), .B(n38060), .Z(n38090) );
  XNOR U39250 ( .A(sreg[1934]), .B(n38090), .Z(n38092) );
  NANDN U39251 ( .A(sreg[1933]), .B(n38053), .Z(n38057) );
  NAND U39252 ( .A(n38055), .B(n38054), .Z(n38056) );
  NAND U39253 ( .A(n38057), .B(n38056), .Z(n38091) );
  XNOR U39254 ( .A(n38092), .B(n38091), .Z(c[1934]) );
  NANDN U39255 ( .A(n38059), .B(n38058), .Z(n38063) );
  NANDN U39256 ( .A(n38061), .B(n38060), .Z(n38062) );
  AND U39257 ( .A(n38063), .B(n38062), .Z(n38098) );
  NANDN U39258 ( .A(n38065), .B(n38064), .Z(n38069) );
  NANDN U39259 ( .A(n38067), .B(n38066), .Z(n38068) );
  AND U39260 ( .A(n38069), .B(n38068), .Z(n38096) );
  NAND U39261 ( .A(n42143), .B(n38070), .Z(n38072) );
  XNOR U39262 ( .A(a[913]), .B(n4202), .Z(n38107) );
  NAND U39263 ( .A(n42144), .B(n38107), .Z(n38071) );
  AND U39264 ( .A(n38072), .B(n38071), .Z(n38122) );
  XOR U39265 ( .A(a[917]), .B(n42012), .Z(n38110) );
  XNOR U39266 ( .A(n38122), .B(n38121), .Z(n38124) );
  AND U39267 ( .A(a[919]), .B(b[0]), .Z(n38074) );
  XNOR U39268 ( .A(n38074), .B(n4071), .Z(n38076) );
  NANDN U39269 ( .A(b[0]), .B(a[918]), .Z(n38075) );
  NAND U39270 ( .A(n38076), .B(n38075), .Z(n38118) );
  XOR U39271 ( .A(a[915]), .B(n42085), .Z(n38114) );
  AND U39272 ( .A(a[911]), .B(b[7]), .Z(n38115) );
  XNOR U39273 ( .A(n38116), .B(n38115), .Z(n38117) );
  XNOR U39274 ( .A(n38118), .B(n38117), .Z(n38123) );
  XOR U39275 ( .A(n38124), .B(n38123), .Z(n38102) );
  NANDN U39276 ( .A(n38079), .B(n38078), .Z(n38083) );
  NANDN U39277 ( .A(n38081), .B(n38080), .Z(n38082) );
  AND U39278 ( .A(n38083), .B(n38082), .Z(n38101) );
  XNOR U39279 ( .A(n38102), .B(n38101), .Z(n38103) );
  NANDN U39280 ( .A(n38085), .B(n38084), .Z(n38089) );
  NAND U39281 ( .A(n38087), .B(n38086), .Z(n38088) );
  NAND U39282 ( .A(n38089), .B(n38088), .Z(n38104) );
  XNOR U39283 ( .A(n38103), .B(n38104), .Z(n38095) );
  XNOR U39284 ( .A(n38096), .B(n38095), .Z(n38097) );
  XNOR U39285 ( .A(n38098), .B(n38097), .Z(n38127) );
  XNOR U39286 ( .A(sreg[1935]), .B(n38127), .Z(n38129) );
  NANDN U39287 ( .A(sreg[1934]), .B(n38090), .Z(n38094) );
  NAND U39288 ( .A(n38092), .B(n38091), .Z(n38093) );
  NAND U39289 ( .A(n38094), .B(n38093), .Z(n38128) );
  XNOR U39290 ( .A(n38129), .B(n38128), .Z(c[1935]) );
  NANDN U39291 ( .A(n38096), .B(n38095), .Z(n38100) );
  NANDN U39292 ( .A(n38098), .B(n38097), .Z(n38099) );
  AND U39293 ( .A(n38100), .B(n38099), .Z(n38135) );
  NANDN U39294 ( .A(n38102), .B(n38101), .Z(n38106) );
  NANDN U39295 ( .A(n38104), .B(n38103), .Z(n38105) );
  AND U39296 ( .A(n38106), .B(n38105), .Z(n38133) );
  NAND U39297 ( .A(n42143), .B(n38107), .Z(n38109) );
  XNOR U39298 ( .A(a[914]), .B(n4202), .Z(n38144) );
  NAND U39299 ( .A(n42144), .B(n38144), .Z(n38108) );
  AND U39300 ( .A(n38109), .B(n38108), .Z(n38159) );
  XOR U39301 ( .A(a[918]), .B(n42012), .Z(n38147) );
  XNOR U39302 ( .A(n38159), .B(n38158), .Z(n38161) );
  AND U39303 ( .A(a[920]), .B(b[0]), .Z(n38111) );
  XNOR U39304 ( .A(n38111), .B(n4071), .Z(n38113) );
  NANDN U39305 ( .A(b[0]), .B(a[919]), .Z(n38112) );
  NAND U39306 ( .A(n38113), .B(n38112), .Z(n38155) );
  XOR U39307 ( .A(a[916]), .B(n42085), .Z(n38151) );
  AND U39308 ( .A(a[912]), .B(b[7]), .Z(n38152) );
  XNOR U39309 ( .A(n38153), .B(n38152), .Z(n38154) );
  XNOR U39310 ( .A(n38155), .B(n38154), .Z(n38160) );
  XOR U39311 ( .A(n38161), .B(n38160), .Z(n38139) );
  NANDN U39312 ( .A(n38116), .B(n38115), .Z(n38120) );
  NANDN U39313 ( .A(n38118), .B(n38117), .Z(n38119) );
  AND U39314 ( .A(n38120), .B(n38119), .Z(n38138) );
  XNOR U39315 ( .A(n38139), .B(n38138), .Z(n38140) );
  NANDN U39316 ( .A(n38122), .B(n38121), .Z(n38126) );
  NAND U39317 ( .A(n38124), .B(n38123), .Z(n38125) );
  NAND U39318 ( .A(n38126), .B(n38125), .Z(n38141) );
  XNOR U39319 ( .A(n38140), .B(n38141), .Z(n38132) );
  XNOR U39320 ( .A(n38133), .B(n38132), .Z(n38134) );
  XNOR U39321 ( .A(n38135), .B(n38134), .Z(n38164) );
  XNOR U39322 ( .A(sreg[1936]), .B(n38164), .Z(n38166) );
  NANDN U39323 ( .A(sreg[1935]), .B(n38127), .Z(n38131) );
  NAND U39324 ( .A(n38129), .B(n38128), .Z(n38130) );
  NAND U39325 ( .A(n38131), .B(n38130), .Z(n38165) );
  XNOR U39326 ( .A(n38166), .B(n38165), .Z(c[1936]) );
  NANDN U39327 ( .A(n38133), .B(n38132), .Z(n38137) );
  NANDN U39328 ( .A(n38135), .B(n38134), .Z(n38136) );
  AND U39329 ( .A(n38137), .B(n38136), .Z(n38172) );
  NANDN U39330 ( .A(n38139), .B(n38138), .Z(n38143) );
  NANDN U39331 ( .A(n38141), .B(n38140), .Z(n38142) );
  AND U39332 ( .A(n38143), .B(n38142), .Z(n38170) );
  NAND U39333 ( .A(n42143), .B(n38144), .Z(n38146) );
  XNOR U39334 ( .A(a[915]), .B(n4202), .Z(n38181) );
  NAND U39335 ( .A(n42144), .B(n38181), .Z(n38145) );
  AND U39336 ( .A(n38146), .B(n38145), .Z(n38196) );
  XOR U39337 ( .A(a[919]), .B(n42012), .Z(n38184) );
  XNOR U39338 ( .A(n38196), .B(n38195), .Z(n38198) );
  AND U39339 ( .A(a[921]), .B(b[0]), .Z(n38148) );
  XNOR U39340 ( .A(n38148), .B(n4071), .Z(n38150) );
  NANDN U39341 ( .A(b[0]), .B(a[920]), .Z(n38149) );
  NAND U39342 ( .A(n38150), .B(n38149), .Z(n38192) );
  XOR U39343 ( .A(a[917]), .B(n42085), .Z(n38188) );
  AND U39344 ( .A(a[913]), .B(b[7]), .Z(n38189) );
  XNOR U39345 ( .A(n38190), .B(n38189), .Z(n38191) );
  XNOR U39346 ( .A(n38192), .B(n38191), .Z(n38197) );
  XOR U39347 ( .A(n38198), .B(n38197), .Z(n38176) );
  NANDN U39348 ( .A(n38153), .B(n38152), .Z(n38157) );
  NANDN U39349 ( .A(n38155), .B(n38154), .Z(n38156) );
  AND U39350 ( .A(n38157), .B(n38156), .Z(n38175) );
  XNOR U39351 ( .A(n38176), .B(n38175), .Z(n38177) );
  NANDN U39352 ( .A(n38159), .B(n38158), .Z(n38163) );
  NAND U39353 ( .A(n38161), .B(n38160), .Z(n38162) );
  NAND U39354 ( .A(n38163), .B(n38162), .Z(n38178) );
  XNOR U39355 ( .A(n38177), .B(n38178), .Z(n38169) );
  XNOR U39356 ( .A(n38170), .B(n38169), .Z(n38171) );
  XNOR U39357 ( .A(n38172), .B(n38171), .Z(n38201) );
  XNOR U39358 ( .A(sreg[1937]), .B(n38201), .Z(n38203) );
  NANDN U39359 ( .A(sreg[1936]), .B(n38164), .Z(n38168) );
  NAND U39360 ( .A(n38166), .B(n38165), .Z(n38167) );
  NAND U39361 ( .A(n38168), .B(n38167), .Z(n38202) );
  XNOR U39362 ( .A(n38203), .B(n38202), .Z(c[1937]) );
  NANDN U39363 ( .A(n38170), .B(n38169), .Z(n38174) );
  NANDN U39364 ( .A(n38172), .B(n38171), .Z(n38173) );
  AND U39365 ( .A(n38174), .B(n38173), .Z(n38209) );
  NANDN U39366 ( .A(n38176), .B(n38175), .Z(n38180) );
  NANDN U39367 ( .A(n38178), .B(n38177), .Z(n38179) );
  AND U39368 ( .A(n38180), .B(n38179), .Z(n38207) );
  NAND U39369 ( .A(n42143), .B(n38181), .Z(n38183) );
  XNOR U39370 ( .A(a[916]), .B(n4202), .Z(n38218) );
  NAND U39371 ( .A(n42144), .B(n38218), .Z(n38182) );
  AND U39372 ( .A(n38183), .B(n38182), .Z(n38233) );
  XOR U39373 ( .A(a[920]), .B(n42012), .Z(n38221) );
  XNOR U39374 ( .A(n38233), .B(n38232), .Z(n38235) );
  AND U39375 ( .A(a[922]), .B(b[0]), .Z(n38185) );
  XNOR U39376 ( .A(n38185), .B(n4071), .Z(n38187) );
  NANDN U39377 ( .A(b[0]), .B(a[921]), .Z(n38186) );
  NAND U39378 ( .A(n38187), .B(n38186), .Z(n38229) );
  XOR U39379 ( .A(a[918]), .B(n42085), .Z(n38225) );
  AND U39380 ( .A(a[914]), .B(b[7]), .Z(n38226) );
  XNOR U39381 ( .A(n38227), .B(n38226), .Z(n38228) );
  XNOR U39382 ( .A(n38229), .B(n38228), .Z(n38234) );
  XOR U39383 ( .A(n38235), .B(n38234), .Z(n38213) );
  NANDN U39384 ( .A(n38190), .B(n38189), .Z(n38194) );
  NANDN U39385 ( .A(n38192), .B(n38191), .Z(n38193) );
  AND U39386 ( .A(n38194), .B(n38193), .Z(n38212) );
  XNOR U39387 ( .A(n38213), .B(n38212), .Z(n38214) );
  NANDN U39388 ( .A(n38196), .B(n38195), .Z(n38200) );
  NAND U39389 ( .A(n38198), .B(n38197), .Z(n38199) );
  NAND U39390 ( .A(n38200), .B(n38199), .Z(n38215) );
  XNOR U39391 ( .A(n38214), .B(n38215), .Z(n38206) );
  XNOR U39392 ( .A(n38207), .B(n38206), .Z(n38208) );
  XNOR U39393 ( .A(n38209), .B(n38208), .Z(n38238) );
  XNOR U39394 ( .A(sreg[1938]), .B(n38238), .Z(n38240) );
  NANDN U39395 ( .A(sreg[1937]), .B(n38201), .Z(n38205) );
  NAND U39396 ( .A(n38203), .B(n38202), .Z(n38204) );
  NAND U39397 ( .A(n38205), .B(n38204), .Z(n38239) );
  XNOR U39398 ( .A(n38240), .B(n38239), .Z(c[1938]) );
  NANDN U39399 ( .A(n38207), .B(n38206), .Z(n38211) );
  NANDN U39400 ( .A(n38209), .B(n38208), .Z(n38210) );
  AND U39401 ( .A(n38211), .B(n38210), .Z(n38246) );
  NANDN U39402 ( .A(n38213), .B(n38212), .Z(n38217) );
  NANDN U39403 ( .A(n38215), .B(n38214), .Z(n38216) );
  AND U39404 ( .A(n38217), .B(n38216), .Z(n38244) );
  NAND U39405 ( .A(n42143), .B(n38218), .Z(n38220) );
  XNOR U39406 ( .A(a[917]), .B(n4202), .Z(n38255) );
  NAND U39407 ( .A(n42144), .B(n38255), .Z(n38219) );
  AND U39408 ( .A(n38220), .B(n38219), .Z(n38270) );
  XOR U39409 ( .A(a[921]), .B(n42012), .Z(n38258) );
  XNOR U39410 ( .A(n38270), .B(n38269), .Z(n38272) );
  AND U39411 ( .A(a[923]), .B(b[0]), .Z(n38222) );
  XNOR U39412 ( .A(n38222), .B(n4071), .Z(n38224) );
  NANDN U39413 ( .A(b[0]), .B(a[922]), .Z(n38223) );
  NAND U39414 ( .A(n38224), .B(n38223), .Z(n38266) );
  XOR U39415 ( .A(a[919]), .B(n42085), .Z(n38262) );
  AND U39416 ( .A(a[915]), .B(b[7]), .Z(n38263) );
  XNOR U39417 ( .A(n38264), .B(n38263), .Z(n38265) );
  XNOR U39418 ( .A(n38266), .B(n38265), .Z(n38271) );
  XOR U39419 ( .A(n38272), .B(n38271), .Z(n38250) );
  NANDN U39420 ( .A(n38227), .B(n38226), .Z(n38231) );
  NANDN U39421 ( .A(n38229), .B(n38228), .Z(n38230) );
  AND U39422 ( .A(n38231), .B(n38230), .Z(n38249) );
  XNOR U39423 ( .A(n38250), .B(n38249), .Z(n38251) );
  NANDN U39424 ( .A(n38233), .B(n38232), .Z(n38237) );
  NAND U39425 ( .A(n38235), .B(n38234), .Z(n38236) );
  NAND U39426 ( .A(n38237), .B(n38236), .Z(n38252) );
  XNOR U39427 ( .A(n38251), .B(n38252), .Z(n38243) );
  XNOR U39428 ( .A(n38244), .B(n38243), .Z(n38245) );
  XNOR U39429 ( .A(n38246), .B(n38245), .Z(n38275) );
  XNOR U39430 ( .A(sreg[1939]), .B(n38275), .Z(n38277) );
  NANDN U39431 ( .A(sreg[1938]), .B(n38238), .Z(n38242) );
  NAND U39432 ( .A(n38240), .B(n38239), .Z(n38241) );
  NAND U39433 ( .A(n38242), .B(n38241), .Z(n38276) );
  XNOR U39434 ( .A(n38277), .B(n38276), .Z(c[1939]) );
  NANDN U39435 ( .A(n38244), .B(n38243), .Z(n38248) );
  NANDN U39436 ( .A(n38246), .B(n38245), .Z(n38247) );
  AND U39437 ( .A(n38248), .B(n38247), .Z(n38283) );
  NANDN U39438 ( .A(n38250), .B(n38249), .Z(n38254) );
  NANDN U39439 ( .A(n38252), .B(n38251), .Z(n38253) );
  AND U39440 ( .A(n38254), .B(n38253), .Z(n38281) );
  NAND U39441 ( .A(n42143), .B(n38255), .Z(n38257) );
  XNOR U39442 ( .A(a[918]), .B(n4203), .Z(n38292) );
  NAND U39443 ( .A(n42144), .B(n38292), .Z(n38256) );
  AND U39444 ( .A(n38257), .B(n38256), .Z(n38307) );
  XOR U39445 ( .A(a[922]), .B(n42012), .Z(n38295) );
  XNOR U39446 ( .A(n38307), .B(n38306), .Z(n38309) );
  AND U39447 ( .A(a[924]), .B(b[0]), .Z(n38259) );
  XNOR U39448 ( .A(n38259), .B(n4071), .Z(n38261) );
  NANDN U39449 ( .A(b[0]), .B(a[923]), .Z(n38260) );
  NAND U39450 ( .A(n38261), .B(n38260), .Z(n38303) );
  XOR U39451 ( .A(a[920]), .B(n42085), .Z(n38296) );
  AND U39452 ( .A(a[916]), .B(b[7]), .Z(n38300) );
  XNOR U39453 ( .A(n38301), .B(n38300), .Z(n38302) );
  XNOR U39454 ( .A(n38303), .B(n38302), .Z(n38308) );
  XOR U39455 ( .A(n38309), .B(n38308), .Z(n38287) );
  NANDN U39456 ( .A(n38264), .B(n38263), .Z(n38268) );
  NANDN U39457 ( .A(n38266), .B(n38265), .Z(n38267) );
  AND U39458 ( .A(n38268), .B(n38267), .Z(n38286) );
  XNOR U39459 ( .A(n38287), .B(n38286), .Z(n38288) );
  NANDN U39460 ( .A(n38270), .B(n38269), .Z(n38274) );
  NAND U39461 ( .A(n38272), .B(n38271), .Z(n38273) );
  NAND U39462 ( .A(n38274), .B(n38273), .Z(n38289) );
  XNOR U39463 ( .A(n38288), .B(n38289), .Z(n38280) );
  XNOR U39464 ( .A(n38281), .B(n38280), .Z(n38282) );
  XNOR U39465 ( .A(n38283), .B(n38282), .Z(n38312) );
  XNOR U39466 ( .A(sreg[1940]), .B(n38312), .Z(n38314) );
  NANDN U39467 ( .A(sreg[1939]), .B(n38275), .Z(n38279) );
  NAND U39468 ( .A(n38277), .B(n38276), .Z(n38278) );
  NAND U39469 ( .A(n38279), .B(n38278), .Z(n38313) );
  XNOR U39470 ( .A(n38314), .B(n38313), .Z(c[1940]) );
  NANDN U39471 ( .A(n38281), .B(n38280), .Z(n38285) );
  NANDN U39472 ( .A(n38283), .B(n38282), .Z(n38284) );
  AND U39473 ( .A(n38285), .B(n38284), .Z(n38320) );
  NANDN U39474 ( .A(n38287), .B(n38286), .Z(n38291) );
  NANDN U39475 ( .A(n38289), .B(n38288), .Z(n38290) );
  AND U39476 ( .A(n38291), .B(n38290), .Z(n38318) );
  NAND U39477 ( .A(n42143), .B(n38292), .Z(n38294) );
  XNOR U39478 ( .A(a[919]), .B(n4203), .Z(n38329) );
  NAND U39479 ( .A(n42144), .B(n38329), .Z(n38293) );
  AND U39480 ( .A(n38294), .B(n38293), .Z(n38344) );
  XOR U39481 ( .A(a[923]), .B(n42012), .Z(n38332) );
  XNOR U39482 ( .A(n38344), .B(n38343), .Z(n38346) );
  XOR U39483 ( .A(a[921]), .B(n42085), .Z(n38333) );
  AND U39484 ( .A(a[917]), .B(b[7]), .Z(n38337) );
  XNOR U39485 ( .A(n38338), .B(n38337), .Z(n38339) );
  AND U39486 ( .A(a[925]), .B(b[0]), .Z(n38297) );
  XNOR U39487 ( .A(n38297), .B(n4071), .Z(n38299) );
  NANDN U39488 ( .A(b[0]), .B(a[924]), .Z(n38298) );
  NAND U39489 ( .A(n38299), .B(n38298), .Z(n38340) );
  XNOR U39490 ( .A(n38339), .B(n38340), .Z(n38345) );
  XOR U39491 ( .A(n38346), .B(n38345), .Z(n38324) );
  NANDN U39492 ( .A(n38301), .B(n38300), .Z(n38305) );
  NANDN U39493 ( .A(n38303), .B(n38302), .Z(n38304) );
  AND U39494 ( .A(n38305), .B(n38304), .Z(n38323) );
  XNOR U39495 ( .A(n38324), .B(n38323), .Z(n38325) );
  NANDN U39496 ( .A(n38307), .B(n38306), .Z(n38311) );
  NAND U39497 ( .A(n38309), .B(n38308), .Z(n38310) );
  NAND U39498 ( .A(n38311), .B(n38310), .Z(n38326) );
  XNOR U39499 ( .A(n38325), .B(n38326), .Z(n38317) );
  XNOR U39500 ( .A(n38318), .B(n38317), .Z(n38319) );
  XNOR U39501 ( .A(n38320), .B(n38319), .Z(n38349) );
  XNOR U39502 ( .A(sreg[1941]), .B(n38349), .Z(n38351) );
  NANDN U39503 ( .A(sreg[1940]), .B(n38312), .Z(n38316) );
  NAND U39504 ( .A(n38314), .B(n38313), .Z(n38315) );
  NAND U39505 ( .A(n38316), .B(n38315), .Z(n38350) );
  XNOR U39506 ( .A(n38351), .B(n38350), .Z(c[1941]) );
  NANDN U39507 ( .A(n38318), .B(n38317), .Z(n38322) );
  NANDN U39508 ( .A(n38320), .B(n38319), .Z(n38321) );
  AND U39509 ( .A(n38322), .B(n38321), .Z(n38357) );
  NANDN U39510 ( .A(n38324), .B(n38323), .Z(n38328) );
  NANDN U39511 ( .A(n38326), .B(n38325), .Z(n38327) );
  AND U39512 ( .A(n38328), .B(n38327), .Z(n38355) );
  NAND U39513 ( .A(n42143), .B(n38329), .Z(n38331) );
  XNOR U39514 ( .A(a[920]), .B(n4203), .Z(n38366) );
  NAND U39515 ( .A(n42144), .B(n38366), .Z(n38330) );
  AND U39516 ( .A(n38331), .B(n38330), .Z(n38381) );
  XOR U39517 ( .A(a[924]), .B(n42012), .Z(n38369) );
  XNOR U39518 ( .A(n38381), .B(n38380), .Z(n38383) );
  XOR U39519 ( .A(a[922]), .B(n42085), .Z(n38373) );
  AND U39520 ( .A(a[918]), .B(b[7]), .Z(n38374) );
  XNOR U39521 ( .A(n38375), .B(n38374), .Z(n38376) );
  AND U39522 ( .A(a[926]), .B(b[0]), .Z(n38334) );
  XNOR U39523 ( .A(n38334), .B(n4071), .Z(n38336) );
  NANDN U39524 ( .A(b[0]), .B(a[925]), .Z(n38335) );
  NAND U39525 ( .A(n38336), .B(n38335), .Z(n38377) );
  XNOR U39526 ( .A(n38376), .B(n38377), .Z(n38382) );
  XOR U39527 ( .A(n38383), .B(n38382), .Z(n38361) );
  NANDN U39528 ( .A(n38338), .B(n38337), .Z(n38342) );
  NANDN U39529 ( .A(n38340), .B(n38339), .Z(n38341) );
  AND U39530 ( .A(n38342), .B(n38341), .Z(n38360) );
  XNOR U39531 ( .A(n38361), .B(n38360), .Z(n38362) );
  NANDN U39532 ( .A(n38344), .B(n38343), .Z(n38348) );
  NAND U39533 ( .A(n38346), .B(n38345), .Z(n38347) );
  NAND U39534 ( .A(n38348), .B(n38347), .Z(n38363) );
  XNOR U39535 ( .A(n38362), .B(n38363), .Z(n38354) );
  XNOR U39536 ( .A(n38355), .B(n38354), .Z(n38356) );
  XNOR U39537 ( .A(n38357), .B(n38356), .Z(n38386) );
  XNOR U39538 ( .A(sreg[1942]), .B(n38386), .Z(n38388) );
  NANDN U39539 ( .A(sreg[1941]), .B(n38349), .Z(n38353) );
  NAND U39540 ( .A(n38351), .B(n38350), .Z(n38352) );
  NAND U39541 ( .A(n38353), .B(n38352), .Z(n38387) );
  XNOR U39542 ( .A(n38388), .B(n38387), .Z(c[1942]) );
  NANDN U39543 ( .A(n38355), .B(n38354), .Z(n38359) );
  NANDN U39544 ( .A(n38357), .B(n38356), .Z(n38358) );
  AND U39545 ( .A(n38359), .B(n38358), .Z(n38394) );
  NANDN U39546 ( .A(n38361), .B(n38360), .Z(n38365) );
  NANDN U39547 ( .A(n38363), .B(n38362), .Z(n38364) );
  AND U39548 ( .A(n38365), .B(n38364), .Z(n38392) );
  NAND U39549 ( .A(n42143), .B(n38366), .Z(n38368) );
  XNOR U39550 ( .A(a[921]), .B(n4203), .Z(n38403) );
  NAND U39551 ( .A(n42144), .B(n38403), .Z(n38367) );
  AND U39552 ( .A(n38368), .B(n38367), .Z(n38418) );
  XOR U39553 ( .A(a[925]), .B(n42012), .Z(n38406) );
  XNOR U39554 ( .A(n38418), .B(n38417), .Z(n38420) );
  AND U39555 ( .A(a[927]), .B(b[0]), .Z(n38370) );
  XNOR U39556 ( .A(n38370), .B(n4071), .Z(n38372) );
  NANDN U39557 ( .A(b[0]), .B(a[926]), .Z(n38371) );
  NAND U39558 ( .A(n38372), .B(n38371), .Z(n38414) );
  XOR U39559 ( .A(a[923]), .B(n42085), .Z(n38407) );
  AND U39560 ( .A(a[919]), .B(b[7]), .Z(n38411) );
  XNOR U39561 ( .A(n38412), .B(n38411), .Z(n38413) );
  XNOR U39562 ( .A(n38414), .B(n38413), .Z(n38419) );
  XOR U39563 ( .A(n38420), .B(n38419), .Z(n38398) );
  NANDN U39564 ( .A(n38375), .B(n38374), .Z(n38379) );
  NANDN U39565 ( .A(n38377), .B(n38376), .Z(n38378) );
  AND U39566 ( .A(n38379), .B(n38378), .Z(n38397) );
  XNOR U39567 ( .A(n38398), .B(n38397), .Z(n38399) );
  NANDN U39568 ( .A(n38381), .B(n38380), .Z(n38385) );
  NAND U39569 ( .A(n38383), .B(n38382), .Z(n38384) );
  NAND U39570 ( .A(n38385), .B(n38384), .Z(n38400) );
  XNOR U39571 ( .A(n38399), .B(n38400), .Z(n38391) );
  XNOR U39572 ( .A(n38392), .B(n38391), .Z(n38393) );
  XNOR U39573 ( .A(n38394), .B(n38393), .Z(n38423) );
  XNOR U39574 ( .A(sreg[1943]), .B(n38423), .Z(n38425) );
  NANDN U39575 ( .A(sreg[1942]), .B(n38386), .Z(n38390) );
  NAND U39576 ( .A(n38388), .B(n38387), .Z(n38389) );
  NAND U39577 ( .A(n38390), .B(n38389), .Z(n38424) );
  XNOR U39578 ( .A(n38425), .B(n38424), .Z(c[1943]) );
  NANDN U39579 ( .A(n38392), .B(n38391), .Z(n38396) );
  NANDN U39580 ( .A(n38394), .B(n38393), .Z(n38395) );
  AND U39581 ( .A(n38396), .B(n38395), .Z(n38431) );
  NANDN U39582 ( .A(n38398), .B(n38397), .Z(n38402) );
  NANDN U39583 ( .A(n38400), .B(n38399), .Z(n38401) );
  AND U39584 ( .A(n38402), .B(n38401), .Z(n38429) );
  NAND U39585 ( .A(n42143), .B(n38403), .Z(n38405) );
  XNOR U39586 ( .A(a[922]), .B(n4203), .Z(n38440) );
  NAND U39587 ( .A(n42144), .B(n38440), .Z(n38404) );
  AND U39588 ( .A(n38405), .B(n38404), .Z(n38455) );
  XOR U39589 ( .A(a[926]), .B(n42012), .Z(n38443) );
  XNOR U39590 ( .A(n38455), .B(n38454), .Z(n38457) );
  XOR U39591 ( .A(a[924]), .B(n42085), .Z(n38447) );
  AND U39592 ( .A(a[920]), .B(b[7]), .Z(n38448) );
  XNOR U39593 ( .A(n38449), .B(n38448), .Z(n38450) );
  AND U39594 ( .A(a[928]), .B(b[0]), .Z(n38408) );
  XNOR U39595 ( .A(n38408), .B(n4071), .Z(n38410) );
  NANDN U39596 ( .A(b[0]), .B(a[927]), .Z(n38409) );
  NAND U39597 ( .A(n38410), .B(n38409), .Z(n38451) );
  XNOR U39598 ( .A(n38450), .B(n38451), .Z(n38456) );
  XOR U39599 ( .A(n38457), .B(n38456), .Z(n38435) );
  NANDN U39600 ( .A(n38412), .B(n38411), .Z(n38416) );
  NANDN U39601 ( .A(n38414), .B(n38413), .Z(n38415) );
  AND U39602 ( .A(n38416), .B(n38415), .Z(n38434) );
  XNOR U39603 ( .A(n38435), .B(n38434), .Z(n38436) );
  NANDN U39604 ( .A(n38418), .B(n38417), .Z(n38422) );
  NAND U39605 ( .A(n38420), .B(n38419), .Z(n38421) );
  NAND U39606 ( .A(n38422), .B(n38421), .Z(n38437) );
  XNOR U39607 ( .A(n38436), .B(n38437), .Z(n38428) );
  XNOR U39608 ( .A(n38429), .B(n38428), .Z(n38430) );
  XNOR U39609 ( .A(n38431), .B(n38430), .Z(n38460) );
  XNOR U39610 ( .A(sreg[1944]), .B(n38460), .Z(n38462) );
  NANDN U39611 ( .A(sreg[1943]), .B(n38423), .Z(n38427) );
  NAND U39612 ( .A(n38425), .B(n38424), .Z(n38426) );
  NAND U39613 ( .A(n38427), .B(n38426), .Z(n38461) );
  XNOR U39614 ( .A(n38462), .B(n38461), .Z(c[1944]) );
  NANDN U39615 ( .A(n38429), .B(n38428), .Z(n38433) );
  NANDN U39616 ( .A(n38431), .B(n38430), .Z(n38432) );
  AND U39617 ( .A(n38433), .B(n38432), .Z(n38468) );
  NANDN U39618 ( .A(n38435), .B(n38434), .Z(n38439) );
  NANDN U39619 ( .A(n38437), .B(n38436), .Z(n38438) );
  AND U39620 ( .A(n38439), .B(n38438), .Z(n38466) );
  NAND U39621 ( .A(n42143), .B(n38440), .Z(n38442) );
  XNOR U39622 ( .A(a[923]), .B(n4203), .Z(n38477) );
  NAND U39623 ( .A(n42144), .B(n38477), .Z(n38441) );
  AND U39624 ( .A(n38442), .B(n38441), .Z(n38492) );
  XOR U39625 ( .A(a[927]), .B(n42012), .Z(n38480) );
  XNOR U39626 ( .A(n38492), .B(n38491), .Z(n38494) );
  AND U39627 ( .A(a[929]), .B(b[0]), .Z(n38444) );
  XNOR U39628 ( .A(n38444), .B(n4071), .Z(n38446) );
  NANDN U39629 ( .A(b[0]), .B(a[928]), .Z(n38445) );
  NAND U39630 ( .A(n38446), .B(n38445), .Z(n38488) );
  XOR U39631 ( .A(a[925]), .B(n42085), .Z(n38481) );
  AND U39632 ( .A(a[921]), .B(b[7]), .Z(n38485) );
  XNOR U39633 ( .A(n38486), .B(n38485), .Z(n38487) );
  XNOR U39634 ( .A(n38488), .B(n38487), .Z(n38493) );
  XOR U39635 ( .A(n38494), .B(n38493), .Z(n38472) );
  NANDN U39636 ( .A(n38449), .B(n38448), .Z(n38453) );
  NANDN U39637 ( .A(n38451), .B(n38450), .Z(n38452) );
  AND U39638 ( .A(n38453), .B(n38452), .Z(n38471) );
  XNOR U39639 ( .A(n38472), .B(n38471), .Z(n38473) );
  NANDN U39640 ( .A(n38455), .B(n38454), .Z(n38459) );
  NAND U39641 ( .A(n38457), .B(n38456), .Z(n38458) );
  NAND U39642 ( .A(n38459), .B(n38458), .Z(n38474) );
  XNOR U39643 ( .A(n38473), .B(n38474), .Z(n38465) );
  XNOR U39644 ( .A(n38466), .B(n38465), .Z(n38467) );
  XNOR U39645 ( .A(n38468), .B(n38467), .Z(n38497) );
  XNOR U39646 ( .A(sreg[1945]), .B(n38497), .Z(n38499) );
  NANDN U39647 ( .A(sreg[1944]), .B(n38460), .Z(n38464) );
  NAND U39648 ( .A(n38462), .B(n38461), .Z(n38463) );
  NAND U39649 ( .A(n38464), .B(n38463), .Z(n38498) );
  XNOR U39650 ( .A(n38499), .B(n38498), .Z(c[1945]) );
  NANDN U39651 ( .A(n38466), .B(n38465), .Z(n38470) );
  NANDN U39652 ( .A(n38468), .B(n38467), .Z(n38469) );
  AND U39653 ( .A(n38470), .B(n38469), .Z(n38505) );
  NANDN U39654 ( .A(n38472), .B(n38471), .Z(n38476) );
  NANDN U39655 ( .A(n38474), .B(n38473), .Z(n38475) );
  AND U39656 ( .A(n38476), .B(n38475), .Z(n38503) );
  NAND U39657 ( .A(n42143), .B(n38477), .Z(n38479) );
  XNOR U39658 ( .A(a[924]), .B(n4203), .Z(n38514) );
  NAND U39659 ( .A(n42144), .B(n38514), .Z(n38478) );
  AND U39660 ( .A(n38479), .B(n38478), .Z(n38529) );
  XOR U39661 ( .A(a[928]), .B(n42012), .Z(n38517) );
  XNOR U39662 ( .A(n38529), .B(n38528), .Z(n38531) );
  XOR U39663 ( .A(a[926]), .B(n42085), .Z(n38518) );
  AND U39664 ( .A(a[922]), .B(b[7]), .Z(n38522) );
  XNOR U39665 ( .A(n38523), .B(n38522), .Z(n38524) );
  AND U39666 ( .A(a[930]), .B(b[0]), .Z(n38482) );
  XNOR U39667 ( .A(n38482), .B(n4071), .Z(n38484) );
  NANDN U39668 ( .A(b[0]), .B(a[929]), .Z(n38483) );
  NAND U39669 ( .A(n38484), .B(n38483), .Z(n38525) );
  XNOR U39670 ( .A(n38524), .B(n38525), .Z(n38530) );
  XOR U39671 ( .A(n38531), .B(n38530), .Z(n38509) );
  NANDN U39672 ( .A(n38486), .B(n38485), .Z(n38490) );
  NANDN U39673 ( .A(n38488), .B(n38487), .Z(n38489) );
  AND U39674 ( .A(n38490), .B(n38489), .Z(n38508) );
  XNOR U39675 ( .A(n38509), .B(n38508), .Z(n38510) );
  NANDN U39676 ( .A(n38492), .B(n38491), .Z(n38496) );
  NAND U39677 ( .A(n38494), .B(n38493), .Z(n38495) );
  NAND U39678 ( .A(n38496), .B(n38495), .Z(n38511) );
  XNOR U39679 ( .A(n38510), .B(n38511), .Z(n38502) );
  XNOR U39680 ( .A(n38503), .B(n38502), .Z(n38504) );
  XNOR U39681 ( .A(n38505), .B(n38504), .Z(n38534) );
  XNOR U39682 ( .A(sreg[1946]), .B(n38534), .Z(n38536) );
  NANDN U39683 ( .A(sreg[1945]), .B(n38497), .Z(n38501) );
  NAND U39684 ( .A(n38499), .B(n38498), .Z(n38500) );
  NAND U39685 ( .A(n38501), .B(n38500), .Z(n38535) );
  XNOR U39686 ( .A(n38536), .B(n38535), .Z(c[1946]) );
  NANDN U39687 ( .A(n38503), .B(n38502), .Z(n38507) );
  NANDN U39688 ( .A(n38505), .B(n38504), .Z(n38506) );
  AND U39689 ( .A(n38507), .B(n38506), .Z(n38542) );
  NANDN U39690 ( .A(n38509), .B(n38508), .Z(n38513) );
  NANDN U39691 ( .A(n38511), .B(n38510), .Z(n38512) );
  AND U39692 ( .A(n38513), .B(n38512), .Z(n38540) );
  NAND U39693 ( .A(n42143), .B(n38514), .Z(n38516) );
  XNOR U39694 ( .A(a[925]), .B(n4204), .Z(n38551) );
  NAND U39695 ( .A(n42144), .B(n38551), .Z(n38515) );
  AND U39696 ( .A(n38516), .B(n38515), .Z(n38566) );
  XOR U39697 ( .A(a[929]), .B(n42012), .Z(n38554) );
  XNOR U39698 ( .A(n38566), .B(n38565), .Z(n38568) );
  XOR U39699 ( .A(a[927]), .B(n42085), .Z(n38558) );
  AND U39700 ( .A(a[923]), .B(b[7]), .Z(n38559) );
  XNOR U39701 ( .A(n38560), .B(n38559), .Z(n38561) );
  AND U39702 ( .A(a[931]), .B(b[0]), .Z(n38519) );
  XNOR U39703 ( .A(n38519), .B(n4071), .Z(n38521) );
  NANDN U39704 ( .A(b[0]), .B(a[930]), .Z(n38520) );
  NAND U39705 ( .A(n38521), .B(n38520), .Z(n38562) );
  XNOR U39706 ( .A(n38561), .B(n38562), .Z(n38567) );
  XOR U39707 ( .A(n38568), .B(n38567), .Z(n38546) );
  NANDN U39708 ( .A(n38523), .B(n38522), .Z(n38527) );
  NANDN U39709 ( .A(n38525), .B(n38524), .Z(n38526) );
  AND U39710 ( .A(n38527), .B(n38526), .Z(n38545) );
  XNOR U39711 ( .A(n38546), .B(n38545), .Z(n38547) );
  NANDN U39712 ( .A(n38529), .B(n38528), .Z(n38533) );
  NAND U39713 ( .A(n38531), .B(n38530), .Z(n38532) );
  NAND U39714 ( .A(n38533), .B(n38532), .Z(n38548) );
  XNOR U39715 ( .A(n38547), .B(n38548), .Z(n38539) );
  XNOR U39716 ( .A(n38540), .B(n38539), .Z(n38541) );
  XNOR U39717 ( .A(n38542), .B(n38541), .Z(n38571) );
  XNOR U39718 ( .A(sreg[1947]), .B(n38571), .Z(n38573) );
  NANDN U39719 ( .A(sreg[1946]), .B(n38534), .Z(n38538) );
  NAND U39720 ( .A(n38536), .B(n38535), .Z(n38537) );
  NAND U39721 ( .A(n38538), .B(n38537), .Z(n38572) );
  XNOR U39722 ( .A(n38573), .B(n38572), .Z(c[1947]) );
  NANDN U39723 ( .A(n38540), .B(n38539), .Z(n38544) );
  NANDN U39724 ( .A(n38542), .B(n38541), .Z(n38543) );
  AND U39725 ( .A(n38544), .B(n38543), .Z(n38579) );
  NANDN U39726 ( .A(n38546), .B(n38545), .Z(n38550) );
  NANDN U39727 ( .A(n38548), .B(n38547), .Z(n38549) );
  AND U39728 ( .A(n38550), .B(n38549), .Z(n38577) );
  NAND U39729 ( .A(n42143), .B(n38551), .Z(n38553) );
  XNOR U39730 ( .A(a[926]), .B(n4204), .Z(n38588) );
  NAND U39731 ( .A(n42144), .B(n38588), .Z(n38552) );
  AND U39732 ( .A(n38553), .B(n38552), .Z(n38603) );
  XOR U39733 ( .A(a[930]), .B(n42012), .Z(n38591) );
  XNOR U39734 ( .A(n38603), .B(n38602), .Z(n38605) );
  AND U39735 ( .A(a[932]), .B(b[0]), .Z(n38555) );
  XNOR U39736 ( .A(n38555), .B(n4071), .Z(n38557) );
  NANDN U39737 ( .A(b[0]), .B(a[931]), .Z(n38556) );
  NAND U39738 ( .A(n38557), .B(n38556), .Z(n38599) );
  XOR U39739 ( .A(a[928]), .B(n42085), .Z(n38595) );
  AND U39740 ( .A(a[924]), .B(b[7]), .Z(n38596) );
  XNOR U39741 ( .A(n38597), .B(n38596), .Z(n38598) );
  XNOR U39742 ( .A(n38599), .B(n38598), .Z(n38604) );
  XOR U39743 ( .A(n38605), .B(n38604), .Z(n38583) );
  NANDN U39744 ( .A(n38560), .B(n38559), .Z(n38564) );
  NANDN U39745 ( .A(n38562), .B(n38561), .Z(n38563) );
  AND U39746 ( .A(n38564), .B(n38563), .Z(n38582) );
  XNOR U39747 ( .A(n38583), .B(n38582), .Z(n38584) );
  NANDN U39748 ( .A(n38566), .B(n38565), .Z(n38570) );
  NAND U39749 ( .A(n38568), .B(n38567), .Z(n38569) );
  NAND U39750 ( .A(n38570), .B(n38569), .Z(n38585) );
  XNOR U39751 ( .A(n38584), .B(n38585), .Z(n38576) );
  XNOR U39752 ( .A(n38577), .B(n38576), .Z(n38578) );
  XNOR U39753 ( .A(n38579), .B(n38578), .Z(n38608) );
  XNOR U39754 ( .A(sreg[1948]), .B(n38608), .Z(n38610) );
  NANDN U39755 ( .A(sreg[1947]), .B(n38571), .Z(n38575) );
  NAND U39756 ( .A(n38573), .B(n38572), .Z(n38574) );
  NAND U39757 ( .A(n38575), .B(n38574), .Z(n38609) );
  XNOR U39758 ( .A(n38610), .B(n38609), .Z(c[1948]) );
  NANDN U39759 ( .A(n38577), .B(n38576), .Z(n38581) );
  NANDN U39760 ( .A(n38579), .B(n38578), .Z(n38580) );
  AND U39761 ( .A(n38581), .B(n38580), .Z(n38616) );
  NANDN U39762 ( .A(n38583), .B(n38582), .Z(n38587) );
  NANDN U39763 ( .A(n38585), .B(n38584), .Z(n38586) );
  AND U39764 ( .A(n38587), .B(n38586), .Z(n38614) );
  NAND U39765 ( .A(n42143), .B(n38588), .Z(n38590) );
  XNOR U39766 ( .A(a[927]), .B(n4204), .Z(n38625) );
  NAND U39767 ( .A(n42144), .B(n38625), .Z(n38589) );
  AND U39768 ( .A(n38590), .B(n38589), .Z(n38640) );
  XOR U39769 ( .A(a[931]), .B(n42012), .Z(n38628) );
  XNOR U39770 ( .A(n38640), .B(n38639), .Z(n38642) );
  AND U39771 ( .A(a[933]), .B(b[0]), .Z(n38592) );
  XNOR U39772 ( .A(n38592), .B(n4071), .Z(n38594) );
  NANDN U39773 ( .A(b[0]), .B(a[932]), .Z(n38593) );
  NAND U39774 ( .A(n38594), .B(n38593), .Z(n38636) );
  XOR U39775 ( .A(a[929]), .B(n42085), .Z(n38629) );
  AND U39776 ( .A(a[925]), .B(b[7]), .Z(n38633) );
  XNOR U39777 ( .A(n38634), .B(n38633), .Z(n38635) );
  XNOR U39778 ( .A(n38636), .B(n38635), .Z(n38641) );
  XOR U39779 ( .A(n38642), .B(n38641), .Z(n38620) );
  NANDN U39780 ( .A(n38597), .B(n38596), .Z(n38601) );
  NANDN U39781 ( .A(n38599), .B(n38598), .Z(n38600) );
  AND U39782 ( .A(n38601), .B(n38600), .Z(n38619) );
  XNOR U39783 ( .A(n38620), .B(n38619), .Z(n38621) );
  NANDN U39784 ( .A(n38603), .B(n38602), .Z(n38607) );
  NAND U39785 ( .A(n38605), .B(n38604), .Z(n38606) );
  NAND U39786 ( .A(n38607), .B(n38606), .Z(n38622) );
  XNOR U39787 ( .A(n38621), .B(n38622), .Z(n38613) );
  XNOR U39788 ( .A(n38614), .B(n38613), .Z(n38615) );
  XNOR U39789 ( .A(n38616), .B(n38615), .Z(n38645) );
  XNOR U39790 ( .A(sreg[1949]), .B(n38645), .Z(n38647) );
  NANDN U39791 ( .A(sreg[1948]), .B(n38608), .Z(n38612) );
  NAND U39792 ( .A(n38610), .B(n38609), .Z(n38611) );
  NAND U39793 ( .A(n38612), .B(n38611), .Z(n38646) );
  XNOR U39794 ( .A(n38647), .B(n38646), .Z(c[1949]) );
  NANDN U39795 ( .A(n38614), .B(n38613), .Z(n38618) );
  NANDN U39796 ( .A(n38616), .B(n38615), .Z(n38617) );
  AND U39797 ( .A(n38618), .B(n38617), .Z(n38653) );
  NANDN U39798 ( .A(n38620), .B(n38619), .Z(n38624) );
  NANDN U39799 ( .A(n38622), .B(n38621), .Z(n38623) );
  AND U39800 ( .A(n38624), .B(n38623), .Z(n38651) );
  NAND U39801 ( .A(n42143), .B(n38625), .Z(n38627) );
  XNOR U39802 ( .A(a[928]), .B(n4204), .Z(n38662) );
  NAND U39803 ( .A(n42144), .B(n38662), .Z(n38626) );
  AND U39804 ( .A(n38627), .B(n38626), .Z(n38677) );
  XOR U39805 ( .A(a[932]), .B(n42012), .Z(n38665) );
  XNOR U39806 ( .A(n38677), .B(n38676), .Z(n38679) );
  XOR U39807 ( .A(a[930]), .B(n42085), .Z(n38669) );
  AND U39808 ( .A(a[926]), .B(b[7]), .Z(n38670) );
  XNOR U39809 ( .A(n38671), .B(n38670), .Z(n38672) );
  AND U39810 ( .A(a[934]), .B(b[0]), .Z(n38630) );
  XNOR U39811 ( .A(n38630), .B(n4071), .Z(n38632) );
  NANDN U39812 ( .A(b[0]), .B(a[933]), .Z(n38631) );
  NAND U39813 ( .A(n38632), .B(n38631), .Z(n38673) );
  XNOR U39814 ( .A(n38672), .B(n38673), .Z(n38678) );
  XOR U39815 ( .A(n38679), .B(n38678), .Z(n38657) );
  NANDN U39816 ( .A(n38634), .B(n38633), .Z(n38638) );
  NANDN U39817 ( .A(n38636), .B(n38635), .Z(n38637) );
  AND U39818 ( .A(n38638), .B(n38637), .Z(n38656) );
  XNOR U39819 ( .A(n38657), .B(n38656), .Z(n38658) );
  NANDN U39820 ( .A(n38640), .B(n38639), .Z(n38644) );
  NAND U39821 ( .A(n38642), .B(n38641), .Z(n38643) );
  NAND U39822 ( .A(n38644), .B(n38643), .Z(n38659) );
  XNOR U39823 ( .A(n38658), .B(n38659), .Z(n38650) );
  XNOR U39824 ( .A(n38651), .B(n38650), .Z(n38652) );
  XNOR U39825 ( .A(n38653), .B(n38652), .Z(n38682) );
  XNOR U39826 ( .A(sreg[1950]), .B(n38682), .Z(n38684) );
  NANDN U39827 ( .A(sreg[1949]), .B(n38645), .Z(n38649) );
  NAND U39828 ( .A(n38647), .B(n38646), .Z(n38648) );
  NAND U39829 ( .A(n38649), .B(n38648), .Z(n38683) );
  XNOR U39830 ( .A(n38684), .B(n38683), .Z(c[1950]) );
  NANDN U39831 ( .A(n38651), .B(n38650), .Z(n38655) );
  NANDN U39832 ( .A(n38653), .B(n38652), .Z(n38654) );
  AND U39833 ( .A(n38655), .B(n38654), .Z(n38690) );
  NANDN U39834 ( .A(n38657), .B(n38656), .Z(n38661) );
  NANDN U39835 ( .A(n38659), .B(n38658), .Z(n38660) );
  AND U39836 ( .A(n38661), .B(n38660), .Z(n38688) );
  NAND U39837 ( .A(n42143), .B(n38662), .Z(n38664) );
  XNOR U39838 ( .A(a[929]), .B(n4204), .Z(n38699) );
  NAND U39839 ( .A(n42144), .B(n38699), .Z(n38663) );
  AND U39840 ( .A(n38664), .B(n38663), .Z(n38714) );
  XOR U39841 ( .A(a[933]), .B(n42012), .Z(n38702) );
  XNOR U39842 ( .A(n38714), .B(n38713), .Z(n38716) );
  AND U39843 ( .A(a[935]), .B(b[0]), .Z(n38666) );
  XNOR U39844 ( .A(n38666), .B(n4071), .Z(n38668) );
  NANDN U39845 ( .A(b[0]), .B(a[934]), .Z(n38667) );
  NAND U39846 ( .A(n38668), .B(n38667), .Z(n38710) );
  XOR U39847 ( .A(a[931]), .B(n42085), .Z(n38706) );
  AND U39848 ( .A(a[927]), .B(b[7]), .Z(n38707) );
  XNOR U39849 ( .A(n38708), .B(n38707), .Z(n38709) );
  XNOR U39850 ( .A(n38710), .B(n38709), .Z(n38715) );
  XOR U39851 ( .A(n38716), .B(n38715), .Z(n38694) );
  NANDN U39852 ( .A(n38671), .B(n38670), .Z(n38675) );
  NANDN U39853 ( .A(n38673), .B(n38672), .Z(n38674) );
  AND U39854 ( .A(n38675), .B(n38674), .Z(n38693) );
  XNOR U39855 ( .A(n38694), .B(n38693), .Z(n38695) );
  NANDN U39856 ( .A(n38677), .B(n38676), .Z(n38681) );
  NAND U39857 ( .A(n38679), .B(n38678), .Z(n38680) );
  NAND U39858 ( .A(n38681), .B(n38680), .Z(n38696) );
  XNOR U39859 ( .A(n38695), .B(n38696), .Z(n38687) );
  XNOR U39860 ( .A(n38688), .B(n38687), .Z(n38689) );
  XNOR U39861 ( .A(n38690), .B(n38689), .Z(n38719) );
  XNOR U39862 ( .A(sreg[1951]), .B(n38719), .Z(n38721) );
  NANDN U39863 ( .A(sreg[1950]), .B(n38682), .Z(n38686) );
  NAND U39864 ( .A(n38684), .B(n38683), .Z(n38685) );
  NAND U39865 ( .A(n38686), .B(n38685), .Z(n38720) );
  XNOR U39866 ( .A(n38721), .B(n38720), .Z(c[1951]) );
  NANDN U39867 ( .A(n38688), .B(n38687), .Z(n38692) );
  NANDN U39868 ( .A(n38690), .B(n38689), .Z(n38691) );
  AND U39869 ( .A(n38692), .B(n38691), .Z(n38727) );
  NANDN U39870 ( .A(n38694), .B(n38693), .Z(n38698) );
  NANDN U39871 ( .A(n38696), .B(n38695), .Z(n38697) );
  AND U39872 ( .A(n38698), .B(n38697), .Z(n38725) );
  NAND U39873 ( .A(n42143), .B(n38699), .Z(n38701) );
  XNOR U39874 ( .A(a[930]), .B(n4204), .Z(n38736) );
  NAND U39875 ( .A(n42144), .B(n38736), .Z(n38700) );
  AND U39876 ( .A(n38701), .B(n38700), .Z(n38751) );
  XOR U39877 ( .A(a[934]), .B(n42012), .Z(n38739) );
  XNOR U39878 ( .A(n38751), .B(n38750), .Z(n38753) );
  AND U39879 ( .A(a[936]), .B(b[0]), .Z(n38703) );
  XNOR U39880 ( .A(n38703), .B(n4071), .Z(n38705) );
  NANDN U39881 ( .A(b[0]), .B(a[935]), .Z(n38704) );
  NAND U39882 ( .A(n38705), .B(n38704), .Z(n38747) );
  XOR U39883 ( .A(a[932]), .B(n42085), .Z(n38743) );
  AND U39884 ( .A(a[928]), .B(b[7]), .Z(n38744) );
  XNOR U39885 ( .A(n38745), .B(n38744), .Z(n38746) );
  XNOR U39886 ( .A(n38747), .B(n38746), .Z(n38752) );
  XOR U39887 ( .A(n38753), .B(n38752), .Z(n38731) );
  NANDN U39888 ( .A(n38708), .B(n38707), .Z(n38712) );
  NANDN U39889 ( .A(n38710), .B(n38709), .Z(n38711) );
  AND U39890 ( .A(n38712), .B(n38711), .Z(n38730) );
  XNOR U39891 ( .A(n38731), .B(n38730), .Z(n38732) );
  NANDN U39892 ( .A(n38714), .B(n38713), .Z(n38718) );
  NAND U39893 ( .A(n38716), .B(n38715), .Z(n38717) );
  NAND U39894 ( .A(n38718), .B(n38717), .Z(n38733) );
  XNOR U39895 ( .A(n38732), .B(n38733), .Z(n38724) );
  XNOR U39896 ( .A(n38725), .B(n38724), .Z(n38726) );
  XNOR U39897 ( .A(n38727), .B(n38726), .Z(n38756) );
  XNOR U39898 ( .A(sreg[1952]), .B(n38756), .Z(n38758) );
  NANDN U39899 ( .A(sreg[1951]), .B(n38719), .Z(n38723) );
  NAND U39900 ( .A(n38721), .B(n38720), .Z(n38722) );
  NAND U39901 ( .A(n38723), .B(n38722), .Z(n38757) );
  XNOR U39902 ( .A(n38758), .B(n38757), .Z(c[1952]) );
  NANDN U39903 ( .A(n38725), .B(n38724), .Z(n38729) );
  NANDN U39904 ( .A(n38727), .B(n38726), .Z(n38728) );
  AND U39905 ( .A(n38729), .B(n38728), .Z(n38764) );
  NANDN U39906 ( .A(n38731), .B(n38730), .Z(n38735) );
  NANDN U39907 ( .A(n38733), .B(n38732), .Z(n38734) );
  AND U39908 ( .A(n38735), .B(n38734), .Z(n38762) );
  NAND U39909 ( .A(n42143), .B(n38736), .Z(n38738) );
  XNOR U39910 ( .A(a[931]), .B(n4204), .Z(n38773) );
  NAND U39911 ( .A(n42144), .B(n38773), .Z(n38737) );
  AND U39912 ( .A(n38738), .B(n38737), .Z(n38788) );
  XOR U39913 ( .A(a[935]), .B(n42012), .Z(n38776) );
  XNOR U39914 ( .A(n38788), .B(n38787), .Z(n38790) );
  AND U39915 ( .A(a[937]), .B(b[0]), .Z(n38740) );
  XNOR U39916 ( .A(n38740), .B(n4071), .Z(n38742) );
  NANDN U39917 ( .A(b[0]), .B(a[936]), .Z(n38741) );
  NAND U39918 ( .A(n38742), .B(n38741), .Z(n38784) );
  XOR U39919 ( .A(a[933]), .B(n42085), .Z(n38780) );
  AND U39920 ( .A(a[929]), .B(b[7]), .Z(n38781) );
  XNOR U39921 ( .A(n38782), .B(n38781), .Z(n38783) );
  XNOR U39922 ( .A(n38784), .B(n38783), .Z(n38789) );
  XOR U39923 ( .A(n38790), .B(n38789), .Z(n38768) );
  NANDN U39924 ( .A(n38745), .B(n38744), .Z(n38749) );
  NANDN U39925 ( .A(n38747), .B(n38746), .Z(n38748) );
  AND U39926 ( .A(n38749), .B(n38748), .Z(n38767) );
  XNOR U39927 ( .A(n38768), .B(n38767), .Z(n38769) );
  NANDN U39928 ( .A(n38751), .B(n38750), .Z(n38755) );
  NAND U39929 ( .A(n38753), .B(n38752), .Z(n38754) );
  NAND U39930 ( .A(n38755), .B(n38754), .Z(n38770) );
  XNOR U39931 ( .A(n38769), .B(n38770), .Z(n38761) );
  XNOR U39932 ( .A(n38762), .B(n38761), .Z(n38763) );
  XNOR U39933 ( .A(n38764), .B(n38763), .Z(n38793) );
  XNOR U39934 ( .A(sreg[1953]), .B(n38793), .Z(n38795) );
  NANDN U39935 ( .A(sreg[1952]), .B(n38756), .Z(n38760) );
  NAND U39936 ( .A(n38758), .B(n38757), .Z(n38759) );
  NAND U39937 ( .A(n38760), .B(n38759), .Z(n38794) );
  XNOR U39938 ( .A(n38795), .B(n38794), .Z(c[1953]) );
  NANDN U39939 ( .A(n38762), .B(n38761), .Z(n38766) );
  NANDN U39940 ( .A(n38764), .B(n38763), .Z(n38765) );
  AND U39941 ( .A(n38766), .B(n38765), .Z(n38801) );
  NANDN U39942 ( .A(n38768), .B(n38767), .Z(n38772) );
  NANDN U39943 ( .A(n38770), .B(n38769), .Z(n38771) );
  AND U39944 ( .A(n38772), .B(n38771), .Z(n38799) );
  NAND U39945 ( .A(n42143), .B(n38773), .Z(n38775) );
  XNOR U39946 ( .A(a[932]), .B(n4205), .Z(n38810) );
  NAND U39947 ( .A(n42144), .B(n38810), .Z(n38774) );
  AND U39948 ( .A(n38775), .B(n38774), .Z(n38825) );
  XOR U39949 ( .A(a[936]), .B(n42012), .Z(n38813) );
  XNOR U39950 ( .A(n38825), .B(n38824), .Z(n38827) );
  AND U39951 ( .A(a[938]), .B(b[0]), .Z(n38777) );
  XNOR U39952 ( .A(n38777), .B(n4071), .Z(n38779) );
  NANDN U39953 ( .A(b[0]), .B(a[937]), .Z(n38778) );
  NAND U39954 ( .A(n38779), .B(n38778), .Z(n38821) );
  XOR U39955 ( .A(a[934]), .B(n42085), .Z(n38817) );
  AND U39956 ( .A(a[930]), .B(b[7]), .Z(n38818) );
  XNOR U39957 ( .A(n38819), .B(n38818), .Z(n38820) );
  XNOR U39958 ( .A(n38821), .B(n38820), .Z(n38826) );
  XOR U39959 ( .A(n38827), .B(n38826), .Z(n38805) );
  NANDN U39960 ( .A(n38782), .B(n38781), .Z(n38786) );
  NANDN U39961 ( .A(n38784), .B(n38783), .Z(n38785) );
  AND U39962 ( .A(n38786), .B(n38785), .Z(n38804) );
  XNOR U39963 ( .A(n38805), .B(n38804), .Z(n38806) );
  NANDN U39964 ( .A(n38788), .B(n38787), .Z(n38792) );
  NAND U39965 ( .A(n38790), .B(n38789), .Z(n38791) );
  NAND U39966 ( .A(n38792), .B(n38791), .Z(n38807) );
  XNOR U39967 ( .A(n38806), .B(n38807), .Z(n38798) );
  XNOR U39968 ( .A(n38799), .B(n38798), .Z(n38800) );
  XNOR U39969 ( .A(n38801), .B(n38800), .Z(n38830) );
  XNOR U39970 ( .A(sreg[1954]), .B(n38830), .Z(n38832) );
  NANDN U39971 ( .A(sreg[1953]), .B(n38793), .Z(n38797) );
  NAND U39972 ( .A(n38795), .B(n38794), .Z(n38796) );
  NAND U39973 ( .A(n38797), .B(n38796), .Z(n38831) );
  XNOR U39974 ( .A(n38832), .B(n38831), .Z(c[1954]) );
  NANDN U39975 ( .A(n38799), .B(n38798), .Z(n38803) );
  NANDN U39976 ( .A(n38801), .B(n38800), .Z(n38802) );
  AND U39977 ( .A(n38803), .B(n38802), .Z(n38838) );
  NANDN U39978 ( .A(n38805), .B(n38804), .Z(n38809) );
  NANDN U39979 ( .A(n38807), .B(n38806), .Z(n38808) );
  AND U39980 ( .A(n38809), .B(n38808), .Z(n38836) );
  NAND U39981 ( .A(n42143), .B(n38810), .Z(n38812) );
  XNOR U39982 ( .A(a[933]), .B(n4205), .Z(n38847) );
  NAND U39983 ( .A(n42144), .B(n38847), .Z(n38811) );
  AND U39984 ( .A(n38812), .B(n38811), .Z(n38862) );
  XOR U39985 ( .A(a[937]), .B(n42012), .Z(n38850) );
  XNOR U39986 ( .A(n38862), .B(n38861), .Z(n38864) );
  AND U39987 ( .A(a[939]), .B(b[0]), .Z(n38814) );
  XNOR U39988 ( .A(n38814), .B(n4071), .Z(n38816) );
  NANDN U39989 ( .A(b[0]), .B(a[938]), .Z(n38815) );
  NAND U39990 ( .A(n38816), .B(n38815), .Z(n38858) );
  XOR U39991 ( .A(a[935]), .B(n42085), .Z(n38854) );
  AND U39992 ( .A(a[931]), .B(b[7]), .Z(n38855) );
  XNOR U39993 ( .A(n38856), .B(n38855), .Z(n38857) );
  XNOR U39994 ( .A(n38858), .B(n38857), .Z(n38863) );
  XOR U39995 ( .A(n38864), .B(n38863), .Z(n38842) );
  NANDN U39996 ( .A(n38819), .B(n38818), .Z(n38823) );
  NANDN U39997 ( .A(n38821), .B(n38820), .Z(n38822) );
  AND U39998 ( .A(n38823), .B(n38822), .Z(n38841) );
  XNOR U39999 ( .A(n38842), .B(n38841), .Z(n38843) );
  NANDN U40000 ( .A(n38825), .B(n38824), .Z(n38829) );
  NAND U40001 ( .A(n38827), .B(n38826), .Z(n38828) );
  NAND U40002 ( .A(n38829), .B(n38828), .Z(n38844) );
  XNOR U40003 ( .A(n38843), .B(n38844), .Z(n38835) );
  XNOR U40004 ( .A(n38836), .B(n38835), .Z(n38837) );
  XNOR U40005 ( .A(n38838), .B(n38837), .Z(n38867) );
  XNOR U40006 ( .A(sreg[1955]), .B(n38867), .Z(n38869) );
  NANDN U40007 ( .A(sreg[1954]), .B(n38830), .Z(n38834) );
  NAND U40008 ( .A(n38832), .B(n38831), .Z(n38833) );
  NAND U40009 ( .A(n38834), .B(n38833), .Z(n38868) );
  XNOR U40010 ( .A(n38869), .B(n38868), .Z(c[1955]) );
  NANDN U40011 ( .A(n38836), .B(n38835), .Z(n38840) );
  NANDN U40012 ( .A(n38838), .B(n38837), .Z(n38839) );
  AND U40013 ( .A(n38840), .B(n38839), .Z(n38875) );
  NANDN U40014 ( .A(n38842), .B(n38841), .Z(n38846) );
  NANDN U40015 ( .A(n38844), .B(n38843), .Z(n38845) );
  AND U40016 ( .A(n38846), .B(n38845), .Z(n38873) );
  NAND U40017 ( .A(n42143), .B(n38847), .Z(n38849) );
  XNOR U40018 ( .A(a[934]), .B(n4205), .Z(n38884) );
  NAND U40019 ( .A(n42144), .B(n38884), .Z(n38848) );
  AND U40020 ( .A(n38849), .B(n38848), .Z(n38899) );
  XOR U40021 ( .A(a[938]), .B(n42012), .Z(n38887) );
  XNOR U40022 ( .A(n38899), .B(n38898), .Z(n38901) );
  AND U40023 ( .A(a[940]), .B(b[0]), .Z(n38851) );
  XNOR U40024 ( .A(n38851), .B(n4071), .Z(n38853) );
  NANDN U40025 ( .A(b[0]), .B(a[939]), .Z(n38852) );
  NAND U40026 ( .A(n38853), .B(n38852), .Z(n38895) );
  XOR U40027 ( .A(a[936]), .B(n42085), .Z(n38891) );
  AND U40028 ( .A(a[932]), .B(b[7]), .Z(n38892) );
  XNOR U40029 ( .A(n38893), .B(n38892), .Z(n38894) );
  XNOR U40030 ( .A(n38895), .B(n38894), .Z(n38900) );
  XOR U40031 ( .A(n38901), .B(n38900), .Z(n38879) );
  NANDN U40032 ( .A(n38856), .B(n38855), .Z(n38860) );
  NANDN U40033 ( .A(n38858), .B(n38857), .Z(n38859) );
  AND U40034 ( .A(n38860), .B(n38859), .Z(n38878) );
  XNOR U40035 ( .A(n38879), .B(n38878), .Z(n38880) );
  NANDN U40036 ( .A(n38862), .B(n38861), .Z(n38866) );
  NAND U40037 ( .A(n38864), .B(n38863), .Z(n38865) );
  NAND U40038 ( .A(n38866), .B(n38865), .Z(n38881) );
  XNOR U40039 ( .A(n38880), .B(n38881), .Z(n38872) );
  XNOR U40040 ( .A(n38873), .B(n38872), .Z(n38874) );
  XNOR U40041 ( .A(n38875), .B(n38874), .Z(n38904) );
  XNOR U40042 ( .A(sreg[1956]), .B(n38904), .Z(n38906) );
  NANDN U40043 ( .A(sreg[1955]), .B(n38867), .Z(n38871) );
  NAND U40044 ( .A(n38869), .B(n38868), .Z(n38870) );
  NAND U40045 ( .A(n38871), .B(n38870), .Z(n38905) );
  XNOR U40046 ( .A(n38906), .B(n38905), .Z(c[1956]) );
  NANDN U40047 ( .A(n38873), .B(n38872), .Z(n38877) );
  NANDN U40048 ( .A(n38875), .B(n38874), .Z(n38876) );
  AND U40049 ( .A(n38877), .B(n38876), .Z(n38912) );
  NANDN U40050 ( .A(n38879), .B(n38878), .Z(n38883) );
  NANDN U40051 ( .A(n38881), .B(n38880), .Z(n38882) );
  AND U40052 ( .A(n38883), .B(n38882), .Z(n38910) );
  NAND U40053 ( .A(n42143), .B(n38884), .Z(n38886) );
  XNOR U40054 ( .A(a[935]), .B(n4205), .Z(n38921) );
  NAND U40055 ( .A(n42144), .B(n38921), .Z(n38885) );
  AND U40056 ( .A(n38886), .B(n38885), .Z(n38936) );
  XOR U40057 ( .A(a[939]), .B(n42012), .Z(n38924) );
  XNOR U40058 ( .A(n38936), .B(n38935), .Z(n38938) );
  AND U40059 ( .A(a[941]), .B(b[0]), .Z(n38888) );
  XNOR U40060 ( .A(n38888), .B(n4071), .Z(n38890) );
  NANDN U40061 ( .A(b[0]), .B(a[940]), .Z(n38889) );
  NAND U40062 ( .A(n38890), .B(n38889), .Z(n38932) );
  XOR U40063 ( .A(a[937]), .B(n42085), .Z(n38928) );
  AND U40064 ( .A(a[933]), .B(b[7]), .Z(n38929) );
  XNOR U40065 ( .A(n38930), .B(n38929), .Z(n38931) );
  XNOR U40066 ( .A(n38932), .B(n38931), .Z(n38937) );
  XOR U40067 ( .A(n38938), .B(n38937), .Z(n38916) );
  NANDN U40068 ( .A(n38893), .B(n38892), .Z(n38897) );
  NANDN U40069 ( .A(n38895), .B(n38894), .Z(n38896) );
  AND U40070 ( .A(n38897), .B(n38896), .Z(n38915) );
  XNOR U40071 ( .A(n38916), .B(n38915), .Z(n38917) );
  NANDN U40072 ( .A(n38899), .B(n38898), .Z(n38903) );
  NAND U40073 ( .A(n38901), .B(n38900), .Z(n38902) );
  NAND U40074 ( .A(n38903), .B(n38902), .Z(n38918) );
  XNOR U40075 ( .A(n38917), .B(n38918), .Z(n38909) );
  XNOR U40076 ( .A(n38910), .B(n38909), .Z(n38911) );
  XNOR U40077 ( .A(n38912), .B(n38911), .Z(n38941) );
  XNOR U40078 ( .A(sreg[1957]), .B(n38941), .Z(n38943) );
  NANDN U40079 ( .A(sreg[1956]), .B(n38904), .Z(n38908) );
  NAND U40080 ( .A(n38906), .B(n38905), .Z(n38907) );
  NAND U40081 ( .A(n38908), .B(n38907), .Z(n38942) );
  XNOR U40082 ( .A(n38943), .B(n38942), .Z(c[1957]) );
  NANDN U40083 ( .A(n38910), .B(n38909), .Z(n38914) );
  NANDN U40084 ( .A(n38912), .B(n38911), .Z(n38913) );
  AND U40085 ( .A(n38914), .B(n38913), .Z(n38949) );
  NANDN U40086 ( .A(n38916), .B(n38915), .Z(n38920) );
  NANDN U40087 ( .A(n38918), .B(n38917), .Z(n38919) );
  AND U40088 ( .A(n38920), .B(n38919), .Z(n38947) );
  NAND U40089 ( .A(n42143), .B(n38921), .Z(n38923) );
  XNOR U40090 ( .A(a[936]), .B(n4205), .Z(n38958) );
  NAND U40091 ( .A(n42144), .B(n38958), .Z(n38922) );
  AND U40092 ( .A(n38923), .B(n38922), .Z(n38973) );
  XOR U40093 ( .A(a[940]), .B(n42012), .Z(n38961) );
  XNOR U40094 ( .A(n38973), .B(n38972), .Z(n38975) );
  AND U40095 ( .A(a[942]), .B(b[0]), .Z(n38925) );
  XNOR U40096 ( .A(n38925), .B(n4071), .Z(n38927) );
  NANDN U40097 ( .A(b[0]), .B(a[941]), .Z(n38926) );
  NAND U40098 ( .A(n38927), .B(n38926), .Z(n38969) );
  XOR U40099 ( .A(a[938]), .B(n42085), .Z(n38962) );
  AND U40100 ( .A(a[934]), .B(b[7]), .Z(n38966) );
  XNOR U40101 ( .A(n38967), .B(n38966), .Z(n38968) );
  XNOR U40102 ( .A(n38969), .B(n38968), .Z(n38974) );
  XOR U40103 ( .A(n38975), .B(n38974), .Z(n38953) );
  NANDN U40104 ( .A(n38930), .B(n38929), .Z(n38934) );
  NANDN U40105 ( .A(n38932), .B(n38931), .Z(n38933) );
  AND U40106 ( .A(n38934), .B(n38933), .Z(n38952) );
  XNOR U40107 ( .A(n38953), .B(n38952), .Z(n38954) );
  NANDN U40108 ( .A(n38936), .B(n38935), .Z(n38940) );
  NAND U40109 ( .A(n38938), .B(n38937), .Z(n38939) );
  NAND U40110 ( .A(n38940), .B(n38939), .Z(n38955) );
  XNOR U40111 ( .A(n38954), .B(n38955), .Z(n38946) );
  XNOR U40112 ( .A(n38947), .B(n38946), .Z(n38948) );
  XNOR U40113 ( .A(n38949), .B(n38948), .Z(n38978) );
  XNOR U40114 ( .A(sreg[1958]), .B(n38978), .Z(n38980) );
  NANDN U40115 ( .A(sreg[1957]), .B(n38941), .Z(n38945) );
  NAND U40116 ( .A(n38943), .B(n38942), .Z(n38944) );
  NAND U40117 ( .A(n38945), .B(n38944), .Z(n38979) );
  XNOR U40118 ( .A(n38980), .B(n38979), .Z(c[1958]) );
  NANDN U40119 ( .A(n38947), .B(n38946), .Z(n38951) );
  NANDN U40120 ( .A(n38949), .B(n38948), .Z(n38950) );
  AND U40121 ( .A(n38951), .B(n38950), .Z(n38986) );
  NANDN U40122 ( .A(n38953), .B(n38952), .Z(n38957) );
  NANDN U40123 ( .A(n38955), .B(n38954), .Z(n38956) );
  AND U40124 ( .A(n38957), .B(n38956), .Z(n38984) );
  NAND U40125 ( .A(n42143), .B(n38958), .Z(n38960) );
  XNOR U40126 ( .A(a[937]), .B(n4205), .Z(n38995) );
  NAND U40127 ( .A(n42144), .B(n38995), .Z(n38959) );
  AND U40128 ( .A(n38960), .B(n38959), .Z(n39010) );
  XOR U40129 ( .A(a[941]), .B(n42012), .Z(n38998) );
  XNOR U40130 ( .A(n39010), .B(n39009), .Z(n39012) );
  XOR U40131 ( .A(a[939]), .B(n42085), .Z(n39002) );
  AND U40132 ( .A(a[935]), .B(b[7]), .Z(n39003) );
  XNOR U40133 ( .A(n39004), .B(n39003), .Z(n39005) );
  AND U40134 ( .A(a[943]), .B(b[0]), .Z(n38963) );
  XNOR U40135 ( .A(n38963), .B(n4071), .Z(n38965) );
  NANDN U40136 ( .A(b[0]), .B(a[942]), .Z(n38964) );
  NAND U40137 ( .A(n38965), .B(n38964), .Z(n39006) );
  XNOR U40138 ( .A(n39005), .B(n39006), .Z(n39011) );
  XOR U40139 ( .A(n39012), .B(n39011), .Z(n38990) );
  NANDN U40140 ( .A(n38967), .B(n38966), .Z(n38971) );
  NANDN U40141 ( .A(n38969), .B(n38968), .Z(n38970) );
  AND U40142 ( .A(n38971), .B(n38970), .Z(n38989) );
  XNOR U40143 ( .A(n38990), .B(n38989), .Z(n38991) );
  NANDN U40144 ( .A(n38973), .B(n38972), .Z(n38977) );
  NAND U40145 ( .A(n38975), .B(n38974), .Z(n38976) );
  NAND U40146 ( .A(n38977), .B(n38976), .Z(n38992) );
  XNOR U40147 ( .A(n38991), .B(n38992), .Z(n38983) );
  XNOR U40148 ( .A(n38984), .B(n38983), .Z(n38985) );
  XNOR U40149 ( .A(n38986), .B(n38985), .Z(n39015) );
  XNOR U40150 ( .A(sreg[1959]), .B(n39015), .Z(n39017) );
  NANDN U40151 ( .A(sreg[1958]), .B(n38978), .Z(n38982) );
  NAND U40152 ( .A(n38980), .B(n38979), .Z(n38981) );
  NAND U40153 ( .A(n38982), .B(n38981), .Z(n39016) );
  XNOR U40154 ( .A(n39017), .B(n39016), .Z(c[1959]) );
  NANDN U40155 ( .A(n38984), .B(n38983), .Z(n38988) );
  NANDN U40156 ( .A(n38986), .B(n38985), .Z(n38987) );
  AND U40157 ( .A(n38988), .B(n38987), .Z(n39023) );
  NANDN U40158 ( .A(n38990), .B(n38989), .Z(n38994) );
  NANDN U40159 ( .A(n38992), .B(n38991), .Z(n38993) );
  AND U40160 ( .A(n38994), .B(n38993), .Z(n39021) );
  NAND U40161 ( .A(n42143), .B(n38995), .Z(n38997) );
  XNOR U40162 ( .A(a[938]), .B(n4205), .Z(n39032) );
  NAND U40163 ( .A(n42144), .B(n39032), .Z(n38996) );
  AND U40164 ( .A(n38997), .B(n38996), .Z(n39047) );
  XOR U40165 ( .A(a[942]), .B(n42012), .Z(n39035) );
  XNOR U40166 ( .A(n39047), .B(n39046), .Z(n39049) );
  AND U40167 ( .A(a[944]), .B(b[0]), .Z(n38999) );
  XNOR U40168 ( .A(n38999), .B(n4071), .Z(n39001) );
  NANDN U40169 ( .A(b[0]), .B(a[943]), .Z(n39000) );
  NAND U40170 ( .A(n39001), .B(n39000), .Z(n39043) );
  XOR U40171 ( .A(a[940]), .B(n42085), .Z(n39039) );
  AND U40172 ( .A(a[936]), .B(b[7]), .Z(n39040) );
  XNOR U40173 ( .A(n39041), .B(n39040), .Z(n39042) );
  XNOR U40174 ( .A(n39043), .B(n39042), .Z(n39048) );
  XOR U40175 ( .A(n39049), .B(n39048), .Z(n39027) );
  NANDN U40176 ( .A(n39004), .B(n39003), .Z(n39008) );
  NANDN U40177 ( .A(n39006), .B(n39005), .Z(n39007) );
  AND U40178 ( .A(n39008), .B(n39007), .Z(n39026) );
  XNOR U40179 ( .A(n39027), .B(n39026), .Z(n39028) );
  NANDN U40180 ( .A(n39010), .B(n39009), .Z(n39014) );
  NAND U40181 ( .A(n39012), .B(n39011), .Z(n39013) );
  NAND U40182 ( .A(n39014), .B(n39013), .Z(n39029) );
  XNOR U40183 ( .A(n39028), .B(n39029), .Z(n39020) );
  XNOR U40184 ( .A(n39021), .B(n39020), .Z(n39022) );
  XNOR U40185 ( .A(n39023), .B(n39022), .Z(n39052) );
  XNOR U40186 ( .A(sreg[1960]), .B(n39052), .Z(n39054) );
  NANDN U40187 ( .A(sreg[1959]), .B(n39015), .Z(n39019) );
  NAND U40188 ( .A(n39017), .B(n39016), .Z(n39018) );
  NAND U40189 ( .A(n39019), .B(n39018), .Z(n39053) );
  XNOR U40190 ( .A(n39054), .B(n39053), .Z(c[1960]) );
  NANDN U40191 ( .A(n39021), .B(n39020), .Z(n39025) );
  NANDN U40192 ( .A(n39023), .B(n39022), .Z(n39024) );
  AND U40193 ( .A(n39025), .B(n39024), .Z(n39060) );
  NANDN U40194 ( .A(n39027), .B(n39026), .Z(n39031) );
  NANDN U40195 ( .A(n39029), .B(n39028), .Z(n39030) );
  AND U40196 ( .A(n39031), .B(n39030), .Z(n39058) );
  NAND U40197 ( .A(n42143), .B(n39032), .Z(n39034) );
  XNOR U40198 ( .A(a[939]), .B(n4206), .Z(n39069) );
  NAND U40199 ( .A(n42144), .B(n39069), .Z(n39033) );
  AND U40200 ( .A(n39034), .B(n39033), .Z(n39084) );
  XOR U40201 ( .A(a[943]), .B(n42012), .Z(n39072) );
  XNOR U40202 ( .A(n39084), .B(n39083), .Z(n39086) );
  AND U40203 ( .A(a[945]), .B(b[0]), .Z(n39036) );
  XNOR U40204 ( .A(n39036), .B(n4071), .Z(n39038) );
  NANDN U40205 ( .A(b[0]), .B(a[944]), .Z(n39037) );
  NAND U40206 ( .A(n39038), .B(n39037), .Z(n39080) );
  XOR U40207 ( .A(a[941]), .B(n42085), .Z(n39076) );
  AND U40208 ( .A(a[937]), .B(b[7]), .Z(n39077) );
  XNOR U40209 ( .A(n39078), .B(n39077), .Z(n39079) );
  XNOR U40210 ( .A(n39080), .B(n39079), .Z(n39085) );
  XOR U40211 ( .A(n39086), .B(n39085), .Z(n39064) );
  NANDN U40212 ( .A(n39041), .B(n39040), .Z(n39045) );
  NANDN U40213 ( .A(n39043), .B(n39042), .Z(n39044) );
  AND U40214 ( .A(n39045), .B(n39044), .Z(n39063) );
  XNOR U40215 ( .A(n39064), .B(n39063), .Z(n39065) );
  NANDN U40216 ( .A(n39047), .B(n39046), .Z(n39051) );
  NAND U40217 ( .A(n39049), .B(n39048), .Z(n39050) );
  NAND U40218 ( .A(n39051), .B(n39050), .Z(n39066) );
  XNOR U40219 ( .A(n39065), .B(n39066), .Z(n39057) );
  XNOR U40220 ( .A(n39058), .B(n39057), .Z(n39059) );
  XNOR U40221 ( .A(n39060), .B(n39059), .Z(n39089) );
  XNOR U40222 ( .A(sreg[1961]), .B(n39089), .Z(n39091) );
  NANDN U40223 ( .A(sreg[1960]), .B(n39052), .Z(n39056) );
  NAND U40224 ( .A(n39054), .B(n39053), .Z(n39055) );
  NAND U40225 ( .A(n39056), .B(n39055), .Z(n39090) );
  XNOR U40226 ( .A(n39091), .B(n39090), .Z(c[1961]) );
  NANDN U40227 ( .A(n39058), .B(n39057), .Z(n39062) );
  NANDN U40228 ( .A(n39060), .B(n39059), .Z(n39061) );
  AND U40229 ( .A(n39062), .B(n39061), .Z(n39097) );
  NANDN U40230 ( .A(n39064), .B(n39063), .Z(n39068) );
  NANDN U40231 ( .A(n39066), .B(n39065), .Z(n39067) );
  AND U40232 ( .A(n39068), .B(n39067), .Z(n39095) );
  NAND U40233 ( .A(n42143), .B(n39069), .Z(n39071) );
  XNOR U40234 ( .A(a[940]), .B(n4206), .Z(n39106) );
  NAND U40235 ( .A(n42144), .B(n39106), .Z(n39070) );
  AND U40236 ( .A(n39071), .B(n39070), .Z(n39121) );
  XOR U40237 ( .A(a[944]), .B(n42012), .Z(n39109) );
  XNOR U40238 ( .A(n39121), .B(n39120), .Z(n39123) );
  AND U40239 ( .A(a[946]), .B(b[0]), .Z(n39073) );
  XNOR U40240 ( .A(n39073), .B(n4071), .Z(n39075) );
  NANDN U40241 ( .A(b[0]), .B(a[945]), .Z(n39074) );
  NAND U40242 ( .A(n39075), .B(n39074), .Z(n39117) );
  XOR U40243 ( .A(a[942]), .B(n42085), .Z(n39110) );
  AND U40244 ( .A(a[938]), .B(b[7]), .Z(n39114) );
  XNOR U40245 ( .A(n39115), .B(n39114), .Z(n39116) );
  XNOR U40246 ( .A(n39117), .B(n39116), .Z(n39122) );
  XOR U40247 ( .A(n39123), .B(n39122), .Z(n39101) );
  NANDN U40248 ( .A(n39078), .B(n39077), .Z(n39082) );
  NANDN U40249 ( .A(n39080), .B(n39079), .Z(n39081) );
  AND U40250 ( .A(n39082), .B(n39081), .Z(n39100) );
  XNOR U40251 ( .A(n39101), .B(n39100), .Z(n39102) );
  NANDN U40252 ( .A(n39084), .B(n39083), .Z(n39088) );
  NAND U40253 ( .A(n39086), .B(n39085), .Z(n39087) );
  NAND U40254 ( .A(n39088), .B(n39087), .Z(n39103) );
  XNOR U40255 ( .A(n39102), .B(n39103), .Z(n39094) );
  XNOR U40256 ( .A(n39095), .B(n39094), .Z(n39096) );
  XNOR U40257 ( .A(n39097), .B(n39096), .Z(n39126) );
  XNOR U40258 ( .A(sreg[1962]), .B(n39126), .Z(n39128) );
  NANDN U40259 ( .A(sreg[1961]), .B(n39089), .Z(n39093) );
  NAND U40260 ( .A(n39091), .B(n39090), .Z(n39092) );
  NAND U40261 ( .A(n39093), .B(n39092), .Z(n39127) );
  XNOR U40262 ( .A(n39128), .B(n39127), .Z(c[1962]) );
  NANDN U40263 ( .A(n39095), .B(n39094), .Z(n39099) );
  NANDN U40264 ( .A(n39097), .B(n39096), .Z(n39098) );
  AND U40265 ( .A(n39099), .B(n39098), .Z(n39134) );
  NANDN U40266 ( .A(n39101), .B(n39100), .Z(n39105) );
  NANDN U40267 ( .A(n39103), .B(n39102), .Z(n39104) );
  AND U40268 ( .A(n39105), .B(n39104), .Z(n39132) );
  NAND U40269 ( .A(n42143), .B(n39106), .Z(n39108) );
  XNOR U40270 ( .A(a[941]), .B(n4206), .Z(n39143) );
  NAND U40271 ( .A(n42144), .B(n39143), .Z(n39107) );
  AND U40272 ( .A(n39108), .B(n39107), .Z(n39158) );
  XOR U40273 ( .A(a[945]), .B(n42012), .Z(n39146) );
  XNOR U40274 ( .A(n39158), .B(n39157), .Z(n39160) );
  XOR U40275 ( .A(a[943]), .B(n42085), .Z(n39147) );
  AND U40276 ( .A(a[939]), .B(b[7]), .Z(n39151) );
  XNOR U40277 ( .A(n39152), .B(n39151), .Z(n39153) );
  AND U40278 ( .A(a[947]), .B(b[0]), .Z(n39111) );
  XNOR U40279 ( .A(n39111), .B(n4071), .Z(n39113) );
  NANDN U40280 ( .A(b[0]), .B(a[946]), .Z(n39112) );
  NAND U40281 ( .A(n39113), .B(n39112), .Z(n39154) );
  XNOR U40282 ( .A(n39153), .B(n39154), .Z(n39159) );
  XOR U40283 ( .A(n39160), .B(n39159), .Z(n39138) );
  NANDN U40284 ( .A(n39115), .B(n39114), .Z(n39119) );
  NANDN U40285 ( .A(n39117), .B(n39116), .Z(n39118) );
  AND U40286 ( .A(n39119), .B(n39118), .Z(n39137) );
  XNOR U40287 ( .A(n39138), .B(n39137), .Z(n39139) );
  NANDN U40288 ( .A(n39121), .B(n39120), .Z(n39125) );
  NAND U40289 ( .A(n39123), .B(n39122), .Z(n39124) );
  NAND U40290 ( .A(n39125), .B(n39124), .Z(n39140) );
  XNOR U40291 ( .A(n39139), .B(n39140), .Z(n39131) );
  XNOR U40292 ( .A(n39132), .B(n39131), .Z(n39133) );
  XNOR U40293 ( .A(n39134), .B(n39133), .Z(n39163) );
  XNOR U40294 ( .A(sreg[1963]), .B(n39163), .Z(n39165) );
  NANDN U40295 ( .A(sreg[1962]), .B(n39126), .Z(n39130) );
  NAND U40296 ( .A(n39128), .B(n39127), .Z(n39129) );
  NAND U40297 ( .A(n39130), .B(n39129), .Z(n39164) );
  XNOR U40298 ( .A(n39165), .B(n39164), .Z(c[1963]) );
  NANDN U40299 ( .A(n39132), .B(n39131), .Z(n39136) );
  NANDN U40300 ( .A(n39134), .B(n39133), .Z(n39135) );
  AND U40301 ( .A(n39136), .B(n39135), .Z(n39171) );
  NANDN U40302 ( .A(n39138), .B(n39137), .Z(n39142) );
  NANDN U40303 ( .A(n39140), .B(n39139), .Z(n39141) );
  AND U40304 ( .A(n39142), .B(n39141), .Z(n39169) );
  NAND U40305 ( .A(n42143), .B(n39143), .Z(n39145) );
  XNOR U40306 ( .A(a[942]), .B(n4206), .Z(n39180) );
  NAND U40307 ( .A(n42144), .B(n39180), .Z(n39144) );
  AND U40308 ( .A(n39145), .B(n39144), .Z(n39195) );
  XOR U40309 ( .A(a[946]), .B(n42012), .Z(n39183) );
  XNOR U40310 ( .A(n39195), .B(n39194), .Z(n39197) );
  XOR U40311 ( .A(a[944]), .B(n42085), .Z(n39184) );
  AND U40312 ( .A(a[940]), .B(b[7]), .Z(n39188) );
  XNOR U40313 ( .A(n39189), .B(n39188), .Z(n39190) );
  AND U40314 ( .A(a[948]), .B(b[0]), .Z(n39148) );
  XNOR U40315 ( .A(n39148), .B(n4071), .Z(n39150) );
  NANDN U40316 ( .A(b[0]), .B(a[947]), .Z(n39149) );
  NAND U40317 ( .A(n39150), .B(n39149), .Z(n39191) );
  XNOR U40318 ( .A(n39190), .B(n39191), .Z(n39196) );
  XOR U40319 ( .A(n39197), .B(n39196), .Z(n39175) );
  NANDN U40320 ( .A(n39152), .B(n39151), .Z(n39156) );
  NANDN U40321 ( .A(n39154), .B(n39153), .Z(n39155) );
  AND U40322 ( .A(n39156), .B(n39155), .Z(n39174) );
  XNOR U40323 ( .A(n39175), .B(n39174), .Z(n39176) );
  NANDN U40324 ( .A(n39158), .B(n39157), .Z(n39162) );
  NAND U40325 ( .A(n39160), .B(n39159), .Z(n39161) );
  NAND U40326 ( .A(n39162), .B(n39161), .Z(n39177) );
  XNOR U40327 ( .A(n39176), .B(n39177), .Z(n39168) );
  XNOR U40328 ( .A(n39169), .B(n39168), .Z(n39170) );
  XNOR U40329 ( .A(n39171), .B(n39170), .Z(n39200) );
  XNOR U40330 ( .A(sreg[1964]), .B(n39200), .Z(n39202) );
  NANDN U40331 ( .A(sreg[1963]), .B(n39163), .Z(n39167) );
  NAND U40332 ( .A(n39165), .B(n39164), .Z(n39166) );
  NAND U40333 ( .A(n39167), .B(n39166), .Z(n39201) );
  XNOR U40334 ( .A(n39202), .B(n39201), .Z(c[1964]) );
  NANDN U40335 ( .A(n39169), .B(n39168), .Z(n39173) );
  NANDN U40336 ( .A(n39171), .B(n39170), .Z(n39172) );
  AND U40337 ( .A(n39173), .B(n39172), .Z(n39208) );
  NANDN U40338 ( .A(n39175), .B(n39174), .Z(n39179) );
  NANDN U40339 ( .A(n39177), .B(n39176), .Z(n39178) );
  AND U40340 ( .A(n39179), .B(n39178), .Z(n39206) );
  NAND U40341 ( .A(n42143), .B(n39180), .Z(n39182) );
  XNOR U40342 ( .A(a[943]), .B(n4206), .Z(n39217) );
  NAND U40343 ( .A(n42144), .B(n39217), .Z(n39181) );
  AND U40344 ( .A(n39182), .B(n39181), .Z(n39232) );
  XOR U40345 ( .A(a[947]), .B(n42012), .Z(n39220) );
  XNOR U40346 ( .A(n39232), .B(n39231), .Z(n39234) );
  XOR U40347 ( .A(a[945]), .B(n42085), .Z(n39224) );
  AND U40348 ( .A(a[941]), .B(b[7]), .Z(n39225) );
  XNOR U40349 ( .A(n39226), .B(n39225), .Z(n39227) );
  AND U40350 ( .A(a[949]), .B(b[0]), .Z(n39185) );
  XNOR U40351 ( .A(n39185), .B(n4071), .Z(n39187) );
  NANDN U40352 ( .A(b[0]), .B(a[948]), .Z(n39186) );
  NAND U40353 ( .A(n39187), .B(n39186), .Z(n39228) );
  XNOR U40354 ( .A(n39227), .B(n39228), .Z(n39233) );
  XOR U40355 ( .A(n39234), .B(n39233), .Z(n39212) );
  NANDN U40356 ( .A(n39189), .B(n39188), .Z(n39193) );
  NANDN U40357 ( .A(n39191), .B(n39190), .Z(n39192) );
  AND U40358 ( .A(n39193), .B(n39192), .Z(n39211) );
  XNOR U40359 ( .A(n39212), .B(n39211), .Z(n39213) );
  NANDN U40360 ( .A(n39195), .B(n39194), .Z(n39199) );
  NAND U40361 ( .A(n39197), .B(n39196), .Z(n39198) );
  NAND U40362 ( .A(n39199), .B(n39198), .Z(n39214) );
  XNOR U40363 ( .A(n39213), .B(n39214), .Z(n39205) );
  XNOR U40364 ( .A(n39206), .B(n39205), .Z(n39207) );
  XNOR U40365 ( .A(n39208), .B(n39207), .Z(n39237) );
  XNOR U40366 ( .A(sreg[1965]), .B(n39237), .Z(n39239) );
  NANDN U40367 ( .A(sreg[1964]), .B(n39200), .Z(n39204) );
  NAND U40368 ( .A(n39202), .B(n39201), .Z(n39203) );
  NAND U40369 ( .A(n39204), .B(n39203), .Z(n39238) );
  XNOR U40370 ( .A(n39239), .B(n39238), .Z(c[1965]) );
  NANDN U40371 ( .A(n39206), .B(n39205), .Z(n39210) );
  NANDN U40372 ( .A(n39208), .B(n39207), .Z(n39209) );
  AND U40373 ( .A(n39210), .B(n39209), .Z(n39245) );
  NANDN U40374 ( .A(n39212), .B(n39211), .Z(n39216) );
  NANDN U40375 ( .A(n39214), .B(n39213), .Z(n39215) );
  AND U40376 ( .A(n39216), .B(n39215), .Z(n39243) );
  NAND U40377 ( .A(n42143), .B(n39217), .Z(n39219) );
  XNOR U40378 ( .A(a[944]), .B(n4206), .Z(n39254) );
  NAND U40379 ( .A(n42144), .B(n39254), .Z(n39218) );
  AND U40380 ( .A(n39219), .B(n39218), .Z(n39269) );
  XOR U40381 ( .A(a[948]), .B(n42012), .Z(n39257) );
  XNOR U40382 ( .A(n39269), .B(n39268), .Z(n39271) );
  AND U40383 ( .A(a[950]), .B(b[0]), .Z(n39221) );
  XNOR U40384 ( .A(n39221), .B(n4071), .Z(n39223) );
  NANDN U40385 ( .A(b[0]), .B(a[949]), .Z(n39222) );
  NAND U40386 ( .A(n39223), .B(n39222), .Z(n39265) );
  XOR U40387 ( .A(a[946]), .B(n42085), .Z(n39258) );
  AND U40388 ( .A(a[942]), .B(b[7]), .Z(n39262) );
  XNOR U40389 ( .A(n39263), .B(n39262), .Z(n39264) );
  XNOR U40390 ( .A(n39265), .B(n39264), .Z(n39270) );
  XOR U40391 ( .A(n39271), .B(n39270), .Z(n39249) );
  NANDN U40392 ( .A(n39226), .B(n39225), .Z(n39230) );
  NANDN U40393 ( .A(n39228), .B(n39227), .Z(n39229) );
  AND U40394 ( .A(n39230), .B(n39229), .Z(n39248) );
  XNOR U40395 ( .A(n39249), .B(n39248), .Z(n39250) );
  NANDN U40396 ( .A(n39232), .B(n39231), .Z(n39236) );
  NAND U40397 ( .A(n39234), .B(n39233), .Z(n39235) );
  NAND U40398 ( .A(n39236), .B(n39235), .Z(n39251) );
  XNOR U40399 ( .A(n39250), .B(n39251), .Z(n39242) );
  XNOR U40400 ( .A(n39243), .B(n39242), .Z(n39244) );
  XNOR U40401 ( .A(n39245), .B(n39244), .Z(n39274) );
  XNOR U40402 ( .A(sreg[1966]), .B(n39274), .Z(n39276) );
  NANDN U40403 ( .A(sreg[1965]), .B(n39237), .Z(n39241) );
  NAND U40404 ( .A(n39239), .B(n39238), .Z(n39240) );
  NAND U40405 ( .A(n39241), .B(n39240), .Z(n39275) );
  XNOR U40406 ( .A(n39276), .B(n39275), .Z(c[1966]) );
  NANDN U40407 ( .A(n39243), .B(n39242), .Z(n39247) );
  NANDN U40408 ( .A(n39245), .B(n39244), .Z(n39246) );
  AND U40409 ( .A(n39247), .B(n39246), .Z(n39282) );
  NANDN U40410 ( .A(n39249), .B(n39248), .Z(n39253) );
  NANDN U40411 ( .A(n39251), .B(n39250), .Z(n39252) );
  AND U40412 ( .A(n39253), .B(n39252), .Z(n39280) );
  NAND U40413 ( .A(n42143), .B(n39254), .Z(n39256) );
  XNOR U40414 ( .A(a[945]), .B(n4206), .Z(n39291) );
  NAND U40415 ( .A(n42144), .B(n39291), .Z(n39255) );
  AND U40416 ( .A(n39256), .B(n39255), .Z(n39306) );
  XOR U40417 ( .A(a[949]), .B(n42012), .Z(n39294) );
  XNOR U40418 ( .A(n39306), .B(n39305), .Z(n39308) );
  XOR U40419 ( .A(a[947]), .B(n42085), .Z(n39298) );
  AND U40420 ( .A(a[943]), .B(b[7]), .Z(n39299) );
  XNOR U40421 ( .A(n39300), .B(n39299), .Z(n39301) );
  AND U40422 ( .A(a[951]), .B(b[0]), .Z(n39259) );
  XNOR U40423 ( .A(n39259), .B(n4071), .Z(n39261) );
  NANDN U40424 ( .A(b[0]), .B(a[950]), .Z(n39260) );
  NAND U40425 ( .A(n39261), .B(n39260), .Z(n39302) );
  XNOR U40426 ( .A(n39301), .B(n39302), .Z(n39307) );
  XOR U40427 ( .A(n39308), .B(n39307), .Z(n39286) );
  NANDN U40428 ( .A(n39263), .B(n39262), .Z(n39267) );
  NANDN U40429 ( .A(n39265), .B(n39264), .Z(n39266) );
  AND U40430 ( .A(n39267), .B(n39266), .Z(n39285) );
  XNOR U40431 ( .A(n39286), .B(n39285), .Z(n39287) );
  NANDN U40432 ( .A(n39269), .B(n39268), .Z(n39273) );
  NAND U40433 ( .A(n39271), .B(n39270), .Z(n39272) );
  NAND U40434 ( .A(n39273), .B(n39272), .Z(n39288) );
  XNOR U40435 ( .A(n39287), .B(n39288), .Z(n39279) );
  XNOR U40436 ( .A(n39280), .B(n39279), .Z(n39281) );
  XNOR U40437 ( .A(n39282), .B(n39281), .Z(n39311) );
  XNOR U40438 ( .A(sreg[1967]), .B(n39311), .Z(n39313) );
  NANDN U40439 ( .A(sreg[1966]), .B(n39274), .Z(n39278) );
  NAND U40440 ( .A(n39276), .B(n39275), .Z(n39277) );
  NAND U40441 ( .A(n39278), .B(n39277), .Z(n39312) );
  XNOR U40442 ( .A(n39313), .B(n39312), .Z(c[1967]) );
  NANDN U40443 ( .A(n39280), .B(n39279), .Z(n39284) );
  NANDN U40444 ( .A(n39282), .B(n39281), .Z(n39283) );
  AND U40445 ( .A(n39284), .B(n39283), .Z(n39319) );
  NANDN U40446 ( .A(n39286), .B(n39285), .Z(n39290) );
  NANDN U40447 ( .A(n39288), .B(n39287), .Z(n39289) );
  AND U40448 ( .A(n39290), .B(n39289), .Z(n39317) );
  NAND U40449 ( .A(n42143), .B(n39291), .Z(n39293) );
  XNOR U40450 ( .A(a[946]), .B(n4207), .Z(n39328) );
  NAND U40451 ( .A(n42144), .B(n39328), .Z(n39292) );
  AND U40452 ( .A(n39293), .B(n39292), .Z(n39343) );
  XOR U40453 ( .A(a[950]), .B(n42012), .Z(n39331) );
  XNOR U40454 ( .A(n39343), .B(n39342), .Z(n39345) );
  AND U40455 ( .A(a[952]), .B(b[0]), .Z(n39295) );
  XNOR U40456 ( .A(n39295), .B(n4071), .Z(n39297) );
  NANDN U40457 ( .A(b[0]), .B(a[951]), .Z(n39296) );
  NAND U40458 ( .A(n39297), .B(n39296), .Z(n39339) );
  XOR U40459 ( .A(a[948]), .B(n42085), .Z(n39332) );
  AND U40460 ( .A(a[944]), .B(b[7]), .Z(n39336) );
  XNOR U40461 ( .A(n39337), .B(n39336), .Z(n39338) );
  XNOR U40462 ( .A(n39339), .B(n39338), .Z(n39344) );
  XOR U40463 ( .A(n39345), .B(n39344), .Z(n39323) );
  NANDN U40464 ( .A(n39300), .B(n39299), .Z(n39304) );
  NANDN U40465 ( .A(n39302), .B(n39301), .Z(n39303) );
  AND U40466 ( .A(n39304), .B(n39303), .Z(n39322) );
  XNOR U40467 ( .A(n39323), .B(n39322), .Z(n39324) );
  NANDN U40468 ( .A(n39306), .B(n39305), .Z(n39310) );
  NAND U40469 ( .A(n39308), .B(n39307), .Z(n39309) );
  NAND U40470 ( .A(n39310), .B(n39309), .Z(n39325) );
  XNOR U40471 ( .A(n39324), .B(n39325), .Z(n39316) );
  XNOR U40472 ( .A(n39317), .B(n39316), .Z(n39318) );
  XNOR U40473 ( .A(n39319), .B(n39318), .Z(n39348) );
  XNOR U40474 ( .A(sreg[1968]), .B(n39348), .Z(n39350) );
  NANDN U40475 ( .A(sreg[1967]), .B(n39311), .Z(n39315) );
  NAND U40476 ( .A(n39313), .B(n39312), .Z(n39314) );
  NAND U40477 ( .A(n39315), .B(n39314), .Z(n39349) );
  XNOR U40478 ( .A(n39350), .B(n39349), .Z(c[1968]) );
  NANDN U40479 ( .A(n39317), .B(n39316), .Z(n39321) );
  NANDN U40480 ( .A(n39319), .B(n39318), .Z(n39320) );
  AND U40481 ( .A(n39321), .B(n39320), .Z(n39356) );
  NANDN U40482 ( .A(n39323), .B(n39322), .Z(n39327) );
  NANDN U40483 ( .A(n39325), .B(n39324), .Z(n39326) );
  AND U40484 ( .A(n39327), .B(n39326), .Z(n39354) );
  NAND U40485 ( .A(n42143), .B(n39328), .Z(n39330) );
  XNOR U40486 ( .A(a[947]), .B(n4207), .Z(n39365) );
  NAND U40487 ( .A(n42144), .B(n39365), .Z(n39329) );
  AND U40488 ( .A(n39330), .B(n39329), .Z(n39380) );
  XOR U40489 ( .A(a[951]), .B(n42012), .Z(n39368) );
  XNOR U40490 ( .A(n39380), .B(n39379), .Z(n39382) );
  XOR U40491 ( .A(a[949]), .B(n42085), .Z(n39372) );
  AND U40492 ( .A(a[945]), .B(b[7]), .Z(n39373) );
  XNOR U40493 ( .A(n39374), .B(n39373), .Z(n39375) );
  AND U40494 ( .A(a[953]), .B(b[0]), .Z(n39333) );
  XNOR U40495 ( .A(n39333), .B(n4071), .Z(n39335) );
  NANDN U40496 ( .A(b[0]), .B(a[952]), .Z(n39334) );
  NAND U40497 ( .A(n39335), .B(n39334), .Z(n39376) );
  XNOR U40498 ( .A(n39375), .B(n39376), .Z(n39381) );
  XOR U40499 ( .A(n39382), .B(n39381), .Z(n39360) );
  NANDN U40500 ( .A(n39337), .B(n39336), .Z(n39341) );
  NANDN U40501 ( .A(n39339), .B(n39338), .Z(n39340) );
  AND U40502 ( .A(n39341), .B(n39340), .Z(n39359) );
  XNOR U40503 ( .A(n39360), .B(n39359), .Z(n39361) );
  NANDN U40504 ( .A(n39343), .B(n39342), .Z(n39347) );
  NAND U40505 ( .A(n39345), .B(n39344), .Z(n39346) );
  NAND U40506 ( .A(n39347), .B(n39346), .Z(n39362) );
  XNOR U40507 ( .A(n39361), .B(n39362), .Z(n39353) );
  XNOR U40508 ( .A(n39354), .B(n39353), .Z(n39355) );
  XNOR U40509 ( .A(n39356), .B(n39355), .Z(n39385) );
  XNOR U40510 ( .A(sreg[1969]), .B(n39385), .Z(n39387) );
  NANDN U40511 ( .A(sreg[1968]), .B(n39348), .Z(n39352) );
  NAND U40512 ( .A(n39350), .B(n39349), .Z(n39351) );
  NAND U40513 ( .A(n39352), .B(n39351), .Z(n39386) );
  XNOR U40514 ( .A(n39387), .B(n39386), .Z(c[1969]) );
  NANDN U40515 ( .A(n39354), .B(n39353), .Z(n39358) );
  NANDN U40516 ( .A(n39356), .B(n39355), .Z(n39357) );
  AND U40517 ( .A(n39358), .B(n39357), .Z(n39393) );
  NANDN U40518 ( .A(n39360), .B(n39359), .Z(n39364) );
  NANDN U40519 ( .A(n39362), .B(n39361), .Z(n39363) );
  AND U40520 ( .A(n39364), .B(n39363), .Z(n39391) );
  NAND U40521 ( .A(n42143), .B(n39365), .Z(n39367) );
  XNOR U40522 ( .A(a[948]), .B(n4207), .Z(n39402) );
  NAND U40523 ( .A(n42144), .B(n39402), .Z(n39366) );
  AND U40524 ( .A(n39367), .B(n39366), .Z(n39417) );
  XOR U40525 ( .A(a[952]), .B(n42012), .Z(n39405) );
  XNOR U40526 ( .A(n39417), .B(n39416), .Z(n39419) );
  AND U40527 ( .A(a[954]), .B(b[0]), .Z(n39369) );
  XNOR U40528 ( .A(n39369), .B(n4071), .Z(n39371) );
  NANDN U40529 ( .A(b[0]), .B(a[953]), .Z(n39370) );
  NAND U40530 ( .A(n39371), .B(n39370), .Z(n39413) );
  XOR U40531 ( .A(a[950]), .B(n42085), .Z(n39409) );
  AND U40532 ( .A(a[946]), .B(b[7]), .Z(n39410) );
  XNOR U40533 ( .A(n39411), .B(n39410), .Z(n39412) );
  XNOR U40534 ( .A(n39413), .B(n39412), .Z(n39418) );
  XOR U40535 ( .A(n39419), .B(n39418), .Z(n39397) );
  NANDN U40536 ( .A(n39374), .B(n39373), .Z(n39378) );
  NANDN U40537 ( .A(n39376), .B(n39375), .Z(n39377) );
  AND U40538 ( .A(n39378), .B(n39377), .Z(n39396) );
  XNOR U40539 ( .A(n39397), .B(n39396), .Z(n39398) );
  NANDN U40540 ( .A(n39380), .B(n39379), .Z(n39384) );
  NAND U40541 ( .A(n39382), .B(n39381), .Z(n39383) );
  NAND U40542 ( .A(n39384), .B(n39383), .Z(n39399) );
  XNOR U40543 ( .A(n39398), .B(n39399), .Z(n39390) );
  XNOR U40544 ( .A(n39391), .B(n39390), .Z(n39392) );
  XNOR U40545 ( .A(n39393), .B(n39392), .Z(n39422) );
  XNOR U40546 ( .A(sreg[1970]), .B(n39422), .Z(n39424) );
  NANDN U40547 ( .A(sreg[1969]), .B(n39385), .Z(n39389) );
  NAND U40548 ( .A(n39387), .B(n39386), .Z(n39388) );
  NAND U40549 ( .A(n39389), .B(n39388), .Z(n39423) );
  XNOR U40550 ( .A(n39424), .B(n39423), .Z(c[1970]) );
  NANDN U40551 ( .A(n39391), .B(n39390), .Z(n39395) );
  NANDN U40552 ( .A(n39393), .B(n39392), .Z(n39394) );
  AND U40553 ( .A(n39395), .B(n39394), .Z(n39430) );
  NANDN U40554 ( .A(n39397), .B(n39396), .Z(n39401) );
  NANDN U40555 ( .A(n39399), .B(n39398), .Z(n39400) );
  AND U40556 ( .A(n39401), .B(n39400), .Z(n39428) );
  NAND U40557 ( .A(n42143), .B(n39402), .Z(n39404) );
  XNOR U40558 ( .A(a[949]), .B(n4207), .Z(n39439) );
  NAND U40559 ( .A(n42144), .B(n39439), .Z(n39403) );
  AND U40560 ( .A(n39404), .B(n39403), .Z(n39454) );
  XOR U40561 ( .A(a[953]), .B(n42012), .Z(n39442) );
  XNOR U40562 ( .A(n39454), .B(n39453), .Z(n39456) );
  AND U40563 ( .A(a[955]), .B(b[0]), .Z(n39406) );
  XNOR U40564 ( .A(n39406), .B(n4071), .Z(n39408) );
  NANDN U40565 ( .A(b[0]), .B(a[954]), .Z(n39407) );
  NAND U40566 ( .A(n39408), .B(n39407), .Z(n39450) );
  XOR U40567 ( .A(a[951]), .B(n42085), .Z(n39446) );
  AND U40568 ( .A(a[947]), .B(b[7]), .Z(n39447) );
  XNOR U40569 ( .A(n39448), .B(n39447), .Z(n39449) );
  XNOR U40570 ( .A(n39450), .B(n39449), .Z(n39455) );
  XOR U40571 ( .A(n39456), .B(n39455), .Z(n39434) );
  NANDN U40572 ( .A(n39411), .B(n39410), .Z(n39415) );
  NANDN U40573 ( .A(n39413), .B(n39412), .Z(n39414) );
  AND U40574 ( .A(n39415), .B(n39414), .Z(n39433) );
  XNOR U40575 ( .A(n39434), .B(n39433), .Z(n39435) );
  NANDN U40576 ( .A(n39417), .B(n39416), .Z(n39421) );
  NAND U40577 ( .A(n39419), .B(n39418), .Z(n39420) );
  NAND U40578 ( .A(n39421), .B(n39420), .Z(n39436) );
  XNOR U40579 ( .A(n39435), .B(n39436), .Z(n39427) );
  XNOR U40580 ( .A(n39428), .B(n39427), .Z(n39429) );
  XNOR U40581 ( .A(n39430), .B(n39429), .Z(n39459) );
  XNOR U40582 ( .A(sreg[1971]), .B(n39459), .Z(n39461) );
  NANDN U40583 ( .A(sreg[1970]), .B(n39422), .Z(n39426) );
  NAND U40584 ( .A(n39424), .B(n39423), .Z(n39425) );
  NAND U40585 ( .A(n39426), .B(n39425), .Z(n39460) );
  XNOR U40586 ( .A(n39461), .B(n39460), .Z(c[1971]) );
  NANDN U40587 ( .A(n39428), .B(n39427), .Z(n39432) );
  NANDN U40588 ( .A(n39430), .B(n39429), .Z(n39431) );
  AND U40589 ( .A(n39432), .B(n39431), .Z(n39467) );
  NANDN U40590 ( .A(n39434), .B(n39433), .Z(n39438) );
  NANDN U40591 ( .A(n39436), .B(n39435), .Z(n39437) );
  AND U40592 ( .A(n39438), .B(n39437), .Z(n39465) );
  NAND U40593 ( .A(n42143), .B(n39439), .Z(n39441) );
  XNOR U40594 ( .A(a[950]), .B(n4207), .Z(n39476) );
  NAND U40595 ( .A(n42144), .B(n39476), .Z(n39440) );
  AND U40596 ( .A(n39441), .B(n39440), .Z(n39491) );
  XOR U40597 ( .A(a[954]), .B(n42012), .Z(n39479) );
  XNOR U40598 ( .A(n39491), .B(n39490), .Z(n39493) );
  AND U40599 ( .A(a[956]), .B(b[0]), .Z(n39443) );
  XNOR U40600 ( .A(n39443), .B(n4071), .Z(n39445) );
  NANDN U40601 ( .A(b[0]), .B(a[955]), .Z(n39444) );
  NAND U40602 ( .A(n39445), .B(n39444), .Z(n39487) );
  XOR U40603 ( .A(a[952]), .B(n42085), .Z(n39483) );
  AND U40604 ( .A(a[948]), .B(b[7]), .Z(n39484) );
  XNOR U40605 ( .A(n39485), .B(n39484), .Z(n39486) );
  XNOR U40606 ( .A(n39487), .B(n39486), .Z(n39492) );
  XOR U40607 ( .A(n39493), .B(n39492), .Z(n39471) );
  NANDN U40608 ( .A(n39448), .B(n39447), .Z(n39452) );
  NANDN U40609 ( .A(n39450), .B(n39449), .Z(n39451) );
  AND U40610 ( .A(n39452), .B(n39451), .Z(n39470) );
  XNOR U40611 ( .A(n39471), .B(n39470), .Z(n39472) );
  NANDN U40612 ( .A(n39454), .B(n39453), .Z(n39458) );
  NAND U40613 ( .A(n39456), .B(n39455), .Z(n39457) );
  NAND U40614 ( .A(n39458), .B(n39457), .Z(n39473) );
  XNOR U40615 ( .A(n39472), .B(n39473), .Z(n39464) );
  XNOR U40616 ( .A(n39465), .B(n39464), .Z(n39466) );
  XNOR U40617 ( .A(n39467), .B(n39466), .Z(n39496) );
  XNOR U40618 ( .A(sreg[1972]), .B(n39496), .Z(n39498) );
  NANDN U40619 ( .A(sreg[1971]), .B(n39459), .Z(n39463) );
  NAND U40620 ( .A(n39461), .B(n39460), .Z(n39462) );
  NAND U40621 ( .A(n39463), .B(n39462), .Z(n39497) );
  XNOR U40622 ( .A(n39498), .B(n39497), .Z(c[1972]) );
  NANDN U40623 ( .A(n39465), .B(n39464), .Z(n39469) );
  NANDN U40624 ( .A(n39467), .B(n39466), .Z(n39468) );
  AND U40625 ( .A(n39469), .B(n39468), .Z(n39504) );
  NANDN U40626 ( .A(n39471), .B(n39470), .Z(n39475) );
  NANDN U40627 ( .A(n39473), .B(n39472), .Z(n39474) );
  AND U40628 ( .A(n39475), .B(n39474), .Z(n39502) );
  NAND U40629 ( .A(n42143), .B(n39476), .Z(n39478) );
  XNOR U40630 ( .A(a[951]), .B(n4207), .Z(n39513) );
  NAND U40631 ( .A(n42144), .B(n39513), .Z(n39477) );
  AND U40632 ( .A(n39478), .B(n39477), .Z(n39528) );
  XOR U40633 ( .A(a[955]), .B(n42012), .Z(n39516) );
  XNOR U40634 ( .A(n39528), .B(n39527), .Z(n39530) );
  AND U40635 ( .A(a[957]), .B(b[0]), .Z(n39480) );
  XNOR U40636 ( .A(n39480), .B(n4071), .Z(n39482) );
  NANDN U40637 ( .A(b[0]), .B(a[956]), .Z(n39481) );
  NAND U40638 ( .A(n39482), .B(n39481), .Z(n39524) );
  XOR U40639 ( .A(a[953]), .B(n42085), .Z(n39520) );
  AND U40640 ( .A(a[949]), .B(b[7]), .Z(n39521) );
  XNOR U40641 ( .A(n39522), .B(n39521), .Z(n39523) );
  XNOR U40642 ( .A(n39524), .B(n39523), .Z(n39529) );
  XOR U40643 ( .A(n39530), .B(n39529), .Z(n39508) );
  NANDN U40644 ( .A(n39485), .B(n39484), .Z(n39489) );
  NANDN U40645 ( .A(n39487), .B(n39486), .Z(n39488) );
  AND U40646 ( .A(n39489), .B(n39488), .Z(n39507) );
  XNOR U40647 ( .A(n39508), .B(n39507), .Z(n39509) );
  NANDN U40648 ( .A(n39491), .B(n39490), .Z(n39495) );
  NAND U40649 ( .A(n39493), .B(n39492), .Z(n39494) );
  NAND U40650 ( .A(n39495), .B(n39494), .Z(n39510) );
  XNOR U40651 ( .A(n39509), .B(n39510), .Z(n39501) );
  XNOR U40652 ( .A(n39502), .B(n39501), .Z(n39503) );
  XNOR U40653 ( .A(n39504), .B(n39503), .Z(n39533) );
  XNOR U40654 ( .A(sreg[1973]), .B(n39533), .Z(n39535) );
  NANDN U40655 ( .A(sreg[1972]), .B(n39496), .Z(n39500) );
  NAND U40656 ( .A(n39498), .B(n39497), .Z(n39499) );
  NAND U40657 ( .A(n39500), .B(n39499), .Z(n39534) );
  XNOR U40658 ( .A(n39535), .B(n39534), .Z(c[1973]) );
  NANDN U40659 ( .A(n39502), .B(n39501), .Z(n39506) );
  NANDN U40660 ( .A(n39504), .B(n39503), .Z(n39505) );
  AND U40661 ( .A(n39506), .B(n39505), .Z(n39541) );
  NANDN U40662 ( .A(n39508), .B(n39507), .Z(n39512) );
  NANDN U40663 ( .A(n39510), .B(n39509), .Z(n39511) );
  AND U40664 ( .A(n39512), .B(n39511), .Z(n39539) );
  NAND U40665 ( .A(n42143), .B(n39513), .Z(n39515) );
  XNOR U40666 ( .A(a[952]), .B(n4207), .Z(n39550) );
  NAND U40667 ( .A(n42144), .B(n39550), .Z(n39514) );
  AND U40668 ( .A(n39515), .B(n39514), .Z(n39565) );
  XOR U40669 ( .A(a[956]), .B(n42012), .Z(n39553) );
  XNOR U40670 ( .A(n39565), .B(n39564), .Z(n39567) );
  AND U40671 ( .A(a[958]), .B(b[0]), .Z(n39517) );
  XNOR U40672 ( .A(n39517), .B(n4071), .Z(n39519) );
  NANDN U40673 ( .A(b[0]), .B(a[957]), .Z(n39518) );
  NAND U40674 ( .A(n39519), .B(n39518), .Z(n39561) );
  XOR U40675 ( .A(a[954]), .B(n42085), .Z(n39557) );
  AND U40676 ( .A(a[950]), .B(b[7]), .Z(n39558) );
  XNOR U40677 ( .A(n39559), .B(n39558), .Z(n39560) );
  XNOR U40678 ( .A(n39561), .B(n39560), .Z(n39566) );
  XOR U40679 ( .A(n39567), .B(n39566), .Z(n39545) );
  NANDN U40680 ( .A(n39522), .B(n39521), .Z(n39526) );
  NANDN U40681 ( .A(n39524), .B(n39523), .Z(n39525) );
  AND U40682 ( .A(n39526), .B(n39525), .Z(n39544) );
  XNOR U40683 ( .A(n39545), .B(n39544), .Z(n39546) );
  NANDN U40684 ( .A(n39528), .B(n39527), .Z(n39532) );
  NAND U40685 ( .A(n39530), .B(n39529), .Z(n39531) );
  NAND U40686 ( .A(n39532), .B(n39531), .Z(n39547) );
  XNOR U40687 ( .A(n39546), .B(n39547), .Z(n39538) );
  XNOR U40688 ( .A(n39539), .B(n39538), .Z(n39540) );
  XNOR U40689 ( .A(n39541), .B(n39540), .Z(n39570) );
  XNOR U40690 ( .A(sreg[1974]), .B(n39570), .Z(n39572) );
  NANDN U40691 ( .A(sreg[1973]), .B(n39533), .Z(n39537) );
  NAND U40692 ( .A(n39535), .B(n39534), .Z(n39536) );
  NAND U40693 ( .A(n39537), .B(n39536), .Z(n39571) );
  XNOR U40694 ( .A(n39572), .B(n39571), .Z(c[1974]) );
  NANDN U40695 ( .A(n39539), .B(n39538), .Z(n39543) );
  NANDN U40696 ( .A(n39541), .B(n39540), .Z(n39542) );
  AND U40697 ( .A(n39543), .B(n39542), .Z(n39578) );
  NANDN U40698 ( .A(n39545), .B(n39544), .Z(n39549) );
  NANDN U40699 ( .A(n39547), .B(n39546), .Z(n39548) );
  AND U40700 ( .A(n39549), .B(n39548), .Z(n39576) );
  NAND U40701 ( .A(n42143), .B(n39550), .Z(n39552) );
  XNOR U40702 ( .A(a[953]), .B(n4208), .Z(n39587) );
  NAND U40703 ( .A(n42144), .B(n39587), .Z(n39551) );
  AND U40704 ( .A(n39552), .B(n39551), .Z(n39602) );
  XOR U40705 ( .A(a[957]), .B(n42012), .Z(n39590) );
  XNOR U40706 ( .A(n39602), .B(n39601), .Z(n39604) );
  AND U40707 ( .A(a[959]), .B(b[0]), .Z(n39554) );
  XNOR U40708 ( .A(n39554), .B(n4071), .Z(n39556) );
  NANDN U40709 ( .A(b[0]), .B(a[958]), .Z(n39555) );
  NAND U40710 ( .A(n39556), .B(n39555), .Z(n39598) );
  XOR U40711 ( .A(a[955]), .B(n42085), .Z(n39594) );
  AND U40712 ( .A(a[951]), .B(b[7]), .Z(n39595) );
  XNOR U40713 ( .A(n39596), .B(n39595), .Z(n39597) );
  XNOR U40714 ( .A(n39598), .B(n39597), .Z(n39603) );
  XOR U40715 ( .A(n39604), .B(n39603), .Z(n39582) );
  NANDN U40716 ( .A(n39559), .B(n39558), .Z(n39563) );
  NANDN U40717 ( .A(n39561), .B(n39560), .Z(n39562) );
  AND U40718 ( .A(n39563), .B(n39562), .Z(n39581) );
  XNOR U40719 ( .A(n39582), .B(n39581), .Z(n39583) );
  NANDN U40720 ( .A(n39565), .B(n39564), .Z(n39569) );
  NAND U40721 ( .A(n39567), .B(n39566), .Z(n39568) );
  NAND U40722 ( .A(n39569), .B(n39568), .Z(n39584) );
  XNOR U40723 ( .A(n39583), .B(n39584), .Z(n39575) );
  XNOR U40724 ( .A(n39576), .B(n39575), .Z(n39577) );
  XNOR U40725 ( .A(n39578), .B(n39577), .Z(n39607) );
  XNOR U40726 ( .A(sreg[1975]), .B(n39607), .Z(n39609) );
  NANDN U40727 ( .A(sreg[1974]), .B(n39570), .Z(n39574) );
  NAND U40728 ( .A(n39572), .B(n39571), .Z(n39573) );
  NAND U40729 ( .A(n39574), .B(n39573), .Z(n39608) );
  XNOR U40730 ( .A(n39609), .B(n39608), .Z(c[1975]) );
  NANDN U40731 ( .A(n39576), .B(n39575), .Z(n39580) );
  NANDN U40732 ( .A(n39578), .B(n39577), .Z(n39579) );
  AND U40733 ( .A(n39580), .B(n39579), .Z(n39615) );
  NANDN U40734 ( .A(n39582), .B(n39581), .Z(n39586) );
  NANDN U40735 ( .A(n39584), .B(n39583), .Z(n39585) );
  AND U40736 ( .A(n39586), .B(n39585), .Z(n39613) );
  NAND U40737 ( .A(n42143), .B(n39587), .Z(n39589) );
  XNOR U40738 ( .A(a[954]), .B(n4208), .Z(n39624) );
  NAND U40739 ( .A(n42144), .B(n39624), .Z(n39588) );
  AND U40740 ( .A(n39589), .B(n39588), .Z(n39639) );
  XOR U40741 ( .A(a[958]), .B(n42012), .Z(n39627) );
  XNOR U40742 ( .A(n39639), .B(n39638), .Z(n39641) );
  AND U40743 ( .A(a[960]), .B(b[0]), .Z(n39591) );
  XNOR U40744 ( .A(n39591), .B(n4071), .Z(n39593) );
  NANDN U40745 ( .A(b[0]), .B(a[959]), .Z(n39592) );
  NAND U40746 ( .A(n39593), .B(n39592), .Z(n39635) );
  XOR U40747 ( .A(a[956]), .B(n42085), .Z(n39631) );
  AND U40748 ( .A(a[952]), .B(b[7]), .Z(n39632) );
  XNOR U40749 ( .A(n39633), .B(n39632), .Z(n39634) );
  XNOR U40750 ( .A(n39635), .B(n39634), .Z(n39640) );
  XOR U40751 ( .A(n39641), .B(n39640), .Z(n39619) );
  NANDN U40752 ( .A(n39596), .B(n39595), .Z(n39600) );
  NANDN U40753 ( .A(n39598), .B(n39597), .Z(n39599) );
  AND U40754 ( .A(n39600), .B(n39599), .Z(n39618) );
  XNOR U40755 ( .A(n39619), .B(n39618), .Z(n39620) );
  NANDN U40756 ( .A(n39602), .B(n39601), .Z(n39606) );
  NAND U40757 ( .A(n39604), .B(n39603), .Z(n39605) );
  NAND U40758 ( .A(n39606), .B(n39605), .Z(n39621) );
  XNOR U40759 ( .A(n39620), .B(n39621), .Z(n39612) );
  XNOR U40760 ( .A(n39613), .B(n39612), .Z(n39614) );
  XNOR U40761 ( .A(n39615), .B(n39614), .Z(n39644) );
  XNOR U40762 ( .A(sreg[1976]), .B(n39644), .Z(n39646) );
  NANDN U40763 ( .A(sreg[1975]), .B(n39607), .Z(n39611) );
  NAND U40764 ( .A(n39609), .B(n39608), .Z(n39610) );
  NAND U40765 ( .A(n39611), .B(n39610), .Z(n39645) );
  XNOR U40766 ( .A(n39646), .B(n39645), .Z(c[1976]) );
  NANDN U40767 ( .A(n39613), .B(n39612), .Z(n39617) );
  NANDN U40768 ( .A(n39615), .B(n39614), .Z(n39616) );
  AND U40769 ( .A(n39617), .B(n39616), .Z(n39652) );
  NANDN U40770 ( .A(n39619), .B(n39618), .Z(n39623) );
  NANDN U40771 ( .A(n39621), .B(n39620), .Z(n39622) );
  AND U40772 ( .A(n39623), .B(n39622), .Z(n39650) );
  NAND U40773 ( .A(n42143), .B(n39624), .Z(n39626) );
  XNOR U40774 ( .A(a[955]), .B(n4208), .Z(n39661) );
  NAND U40775 ( .A(n42144), .B(n39661), .Z(n39625) );
  AND U40776 ( .A(n39626), .B(n39625), .Z(n39676) );
  XOR U40777 ( .A(a[959]), .B(n42012), .Z(n39664) );
  XNOR U40778 ( .A(n39676), .B(n39675), .Z(n39678) );
  AND U40779 ( .A(a[961]), .B(b[0]), .Z(n39628) );
  XNOR U40780 ( .A(n39628), .B(n4071), .Z(n39630) );
  NANDN U40781 ( .A(b[0]), .B(a[960]), .Z(n39629) );
  NAND U40782 ( .A(n39630), .B(n39629), .Z(n39672) );
  XOR U40783 ( .A(a[957]), .B(n42085), .Z(n39665) );
  AND U40784 ( .A(a[953]), .B(b[7]), .Z(n39669) );
  XNOR U40785 ( .A(n39670), .B(n39669), .Z(n39671) );
  XNOR U40786 ( .A(n39672), .B(n39671), .Z(n39677) );
  XOR U40787 ( .A(n39678), .B(n39677), .Z(n39656) );
  NANDN U40788 ( .A(n39633), .B(n39632), .Z(n39637) );
  NANDN U40789 ( .A(n39635), .B(n39634), .Z(n39636) );
  AND U40790 ( .A(n39637), .B(n39636), .Z(n39655) );
  XNOR U40791 ( .A(n39656), .B(n39655), .Z(n39657) );
  NANDN U40792 ( .A(n39639), .B(n39638), .Z(n39643) );
  NAND U40793 ( .A(n39641), .B(n39640), .Z(n39642) );
  NAND U40794 ( .A(n39643), .B(n39642), .Z(n39658) );
  XNOR U40795 ( .A(n39657), .B(n39658), .Z(n39649) );
  XNOR U40796 ( .A(n39650), .B(n39649), .Z(n39651) );
  XNOR U40797 ( .A(n39652), .B(n39651), .Z(n39681) );
  XNOR U40798 ( .A(sreg[1977]), .B(n39681), .Z(n39683) );
  NANDN U40799 ( .A(sreg[1976]), .B(n39644), .Z(n39648) );
  NAND U40800 ( .A(n39646), .B(n39645), .Z(n39647) );
  NAND U40801 ( .A(n39648), .B(n39647), .Z(n39682) );
  XNOR U40802 ( .A(n39683), .B(n39682), .Z(c[1977]) );
  NANDN U40803 ( .A(n39650), .B(n39649), .Z(n39654) );
  NANDN U40804 ( .A(n39652), .B(n39651), .Z(n39653) );
  AND U40805 ( .A(n39654), .B(n39653), .Z(n39689) );
  NANDN U40806 ( .A(n39656), .B(n39655), .Z(n39660) );
  NANDN U40807 ( .A(n39658), .B(n39657), .Z(n39659) );
  AND U40808 ( .A(n39660), .B(n39659), .Z(n39687) );
  NAND U40809 ( .A(n42143), .B(n39661), .Z(n39663) );
  XNOR U40810 ( .A(a[956]), .B(n4208), .Z(n39698) );
  NAND U40811 ( .A(n42144), .B(n39698), .Z(n39662) );
  AND U40812 ( .A(n39663), .B(n39662), .Z(n39713) );
  XOR U40813 ( .A(a[960]), .B(n42012), .Z(n39701) );
  XNOR U40814 ( .A(n39713), .B(n39712), .Z(n39715) );
  XOR U40815 ( .A(a[958]), .B(n42085), .Z(n39705) );
  AND U40816 ( .A(a[954]), .B(b[7]), .Z(n39706) );
  XNOR U40817 ( .A(n39707), .B(n39706), .Z(n39708) );
  AND U40818 ( .A(a[962]), .B(b[0]), .Z(n39666) );
  XNOR U40819 ( .A(n39666), .B(n4071), .Z(n39668) );
  NANDN U40820 ( .A(b[0]), .B(a[961]), .Z(n39667) );
  NAND U40821 ( .A(n39668), .B(n39667), .Z(n39709) );
  XNOR U40822 ( .A(n39708), .B(n39709), .Z(n39714) );
  XOR U40823 ( .A(n39715), .B(n39714), .Z(n39693) );
  NANDN U40824 ( .A(n39670), .B(n39669), .Z(n39674) );
  NANDN U40825 ( .A(n39672), .B(n39671), .Z(n39673) );
  AND U40826 ( .A(n39674), .B(n39673), .Z(n39692) );
  XNOR U40827 ( .A(n39693), .B(n39692), .Z(n39694) );
  NANDN U40828 ( .A(n39676), .B(n39675), .Z(n39680) );
  NAND U40829 ( .A(n39678), .B(n39677), .Z(n39679) );
  NAND U40830 ( .A(n39680), .B(n39679), .Z(n39695) );
  XNOR U40831 ( .A(n39694), .B(n39695), .Z(n39686) );
  XNOR U40832 ( .A(n39687), .B(n39686), .Z(n39688) );
  XNOR U40833 ( .A(n39689), .B(n39688), .Z(n39718) );
  XNOR U40834 ( .A(sreg[1978]), .B(n39718), .Z(n39720) );
  NANDN U40835 ( .A(sreg[1977]), .B(n39681), .Z(n39685) );
  NAND U40836 ( .A(n39683), .B(n39682), .Z(n39684) );
  NAND U40837 ( .A(n39685), .B(n39684), .Z(n39719) );
  XNOR U40838 ( .A(n39720), .B(n39719), .Z(c[1978]) );
  NANDN U40839 ( .A(n39687), .B(n39686), .Z(n39691) );
  NANDN U40840 ( .A(n39689), .B(n39688), .Z(n39690) );
  AND U40841 ( .A(n39691), .B(n39690), .Z(n39726) );
  NANDN U40842 ( .A(n39693), .B(n39692), .Z(n39697) );
  NANDN U40843 ( .A(n39695), .B(n39694), .Z(n39696) );
  AND U40844 ( .A(n39697), .B(n39696), .Z(n39724) );
  NAND U40845 ( .A(n42143), .B(n39698), .Z(n39700) );
  XNOR U40846 ( .A(a[957]), .B(n4208), .Z(n39735) );
  NAND U40847 ( .A(n42144), .B(n39735), .Z(n39699) );
  AND U40848 ( .A(n39700), .B(n39699), .Z(n39750) );
  XOR U40849 ( .A(a[961]), .B(n42012), .Z(n39738) );
  XNOR U40850 ( .A(n39750), .B(n39749), .Z(n39752) );
  AND U40851 ( .A(a[963]), .B(b[0]), .Z(n39702) );
  XNOR U40852 ( .A(n39702), .B(n4071), .Z(n39704) );
  NANDN U40853 ( .A(b[0]), .B(a[962]), .Z(n39703) );
  NAND U40854 ( .A(n39704), .B(n39703), .Z(n39746) );
  XOR U40855 ( .A(a[959]), .B(n42085), .Z(n39742) );
  AND U40856 ( .A(a[955]), .B(b[7]), .Z(n39743) );
  XNOR U40857 ( .A(n39744), .B(n39743), .Z(n39745) );
  XNOR U40858 ( .A(n39746), .B(n39745), .Z(n39751) );
  XOR U40859 ( .A(n39752), .B(n39751), .Z(n39730) );
  NANDN U40860 ( .A(n39707), .B(n39706), .Z(n39711) );
  NANDN U40861 ( .A(n39709), .B(n39708), .Z(n39710) );
  AND U40862 ( .A(n39711), .B(n39710), .Z(n39729) );
  XNOR U40863 ( .A(n39730), .B(n39729), .Z(n39731) );
  NANDN U40864 ( .A(n39713), .B(n39712), .Z(n39717) );
  NAND U40865 ( .A(n39715), .B(n39714), .Z(n39716) );
  NAND U40866 ( .A(n39717), .B(n39716), .Z(n39732) );
  XNOR U40867 ( .A(n39731), .B(n39732), .Z(n39723) );
  XNOR U40868 ( .A(n39724), .B(n39723), .Z(n39725) );
  XNOR U40869 ( .A(n39726), .B(n39725), .Z(n39755) );
  XNOR U40870 ( .A(sreg[1979]), .B(n39755), .Z(n39757) );
  NANDN U40871 ( .A(sreg[1978]), .B(n39718), .Z(n39722) );
  NAND U40872 ( .A(n39720), .B(n39719), .Z(n39721) );
  NAND U40873 ( .A(n39722), .B(n39721), .Z(n39756) );
  XNOR U40874 ( .A(n39757), .B(n39756), .Z(c[1979]) );
  NANDN U40875 ( .A(n39724), .B(n39723), .Z(n39728) );
  NANDN U40876 ( .A(n39726), .B(n39725), .Z(n39727) );
  AND U40877 ( .A(n39728), .B(n39727), .Z(n39763) );
  NANDN U40878 ( .A(n39730), .B(n39729), .Z(n39734) );
  NANDN U40879 ( .A(n39732), .B(n39731), .Z(n39733) );
  AND U40880 ( .A(n39734), .B(n39733), .Z(n39761) );
  NAND U40881 ( .A(n42143), .B(n39735), .Z(n39737) );
  XNOR U40882 ( .A(a[958]), .B(n4208), .Z(n39772) );
  NAND U40883 ( .A(n42144), .B(n39772), .Z(n39736) );
  AND U40884 ( .A(n39737), .B(n39736), .Z(n39787) );
  XOR U40885 ( .A(a[962]), .B(n42012), .Z(n39775) );
  XNOR U40886 ( .A(n39787), .B(n39786), .Z(n39789) );
  AND U40887 ( .A(a[964]), .B(b[0]), .Z(n39739) );
  XNOR U40888 ( .A(n39739), .B(n4071), .Z(n39741) );
  NANDN U40889 ( .A(b[0]), .B(a[963]), .Z(n39740) );
  NAND U40890 ( .A(n39741), .B(n39740), .Z(n39783) );
  XOR U40891 ( .A(a[960]), .B(n42085), .Z(n39779) );
  AND U40892 ( .A(a[956]), .B(b[7]), .Z(n39780) );
  XNOR U40893 ( .A(n39781), .B(n39780), .Z(n39782) );
  XNOR U40894 ( .A(n39783), .B(n39782), .Z(n39788) );
  XOR U40895 ( .A(n39789), .B(n39788), .Z(n39767) );
  NANDN U40896 ( .A(n39744), .B(n39743), .Z(n39748) );
  NANDN U40897 ( .A(n39746), .B(n39745), .Z(n39747) );
  AND U40898 ( .A(n39748), .B(n39747), .Z(n39766) );
  XNOR U40899 ( .A(n39767), .B(n39766), .Z(n39768) );
  NANDN U40900 ( .A(n39750), .B(n39749), .Z(n39754) );
  NAND U40901 ( .A(n39752), .B(n39751), .Z(n39753) );
  NAND U40902 ( .A(n39754), .B(n39753), .Z(n39769) );
  XNOR U40903 ( .A(n39768), .B(n39769), .Z(n39760) );
  XNOR U40904 ( .A(n39761), .B(n39760), .Z(n39762) );
  XNOR U40905 ( .A(n39763), .B(n39762), .Z(n39792) );
  XNOR U40906 ( .A(sreg[1980]), .B(n39792), .Z(n39794) );
  NANDN U40907 ( .A(sreg[1979]), .B(n39755), .Z(n39759) );
  NAND U40908 ( .A(n39757), .B(n39756), .Z(n39758) );
  NAND U40909 ( .A(n39759), .B(n39758), .Z(n39793) );
  XNOR U40910 ( .A(n39794), .B(n39793), .Z(c[1980]) );
  NANDN U40911 ( .A(n39761), .B(n39760), .Z(n39765) );
  NANDN U40912 ( .A(n39763), .B(n39762), .Z(n39764) );
  AND U40913 ( .A(n39765), .B(n39764), .Z(n39800) );
  NANDN U40914 ( .A(n39767), .B(n39766), .Z(n39771) );
  NANDN U40915 ( .A(n39769), .B(n39768), .Z(n39770) );
  AND U40916 ( .A(n39771), .B(n39770), .Z(n39798) );
  NAND U40917 ( .A(n42143), .B(n39772), .Z(n39774) );
  XNOR U40918 ( .A(a[959]), .B(n4208), .Z(n39809) );
  NAND U40919 ( .A(n42144), .B(n39809), .Z(n39773) );
  AND U40920 ( .A(n39774), .B(n39773), .Z(n39824) );
  XOR U40921 ( .A(a[963]), .B(n42012), .Z(n39812) );
  XNOR U40922 ( .A(n39824), .B(n39823), .Z(n39826) );
  AND U40923 ( .A(a[965]), .B(b[0]), .Z(n39776) );
  XNOR U40924 ( .A(n39776), .B(n4071), .Z(n39778) );
  NANDN U40925 ( .A(b[0]), .B(a[964]), .Z(n39777) );
  NAND U40926 ( .A(n39778), .B(n39777), .Z(n39820) );
  XOR U40927 ( .A(a[961]), .B(n42085), .Z(n39813) );
  AND U40928 ( .A(a[957]), .B(b[7]), .Z(n39817) );
  XNOR U40929 ( .A(n39818), .B(n39817), .Z(n39819) );
  XNOR U40930 ( .A(n39820), .B(n39819), .Z(n39825) );
  XOR U40931 ( .A(n39826), .B(n39825), .Z(n39804) );
  NANDN U40932 ( .A(n39781), .B(n39780), .Z(n39785) );
  NANDN U40933 ( .A(n39783), .B(n39782), .Z(n39784) );
  AND U40934 ( .A(n39785), .B(n39784), .Z(n39803) );
  XNOR U40935 ( .A(n39804), .B(n39803), .Z(n39805) );
  NANDN U40936 ( .A(n39787), .B(n39786), .Z(n39791) );
  NAND U40937 ( .A(n39789), .B(n39788), .Z(n39790) );
  NAND U40938 ( .A(n39791), .B(n39790), .Z(n39806) );
  XNOR U40939 ( .A(n39805), .B(n39806), .Z(n39797) );
  XNOR U40940 ( .A(n39798), .B(n39797), .Z(n39799) );
  XNOR U40941 ( .A(n39800), .B(n39799), .Z(n39829) );
  XNOR U40942 ( .A(sreg[1981]), .B(n39829), .Z(n39831) );
  NANDN U40943 ( .A(sreg[1980]), .B(n39792), .Z(n39796) );
  NAND U40944 ( .A(n39794), .B(n39793), .Z(n39795) );
  NAND U40945 ( .A(n39796), .B(n39795), .Z(n39830) );
  XNOR U40946 ( .A(n39831), .B(n39830), .Z(c[1981]) );
  NANDN U40947 ( .A(n39798), .B(n39797), .Z(n39802) );
  NANDN U40948 ( .A(n39800), .B(n39799), .Z(n39801) );
  AND U40949 ( .A(n39802), .B(n39801), .Z(n39837) );
  NANDN U40950 ( .A(n39804), .B(n39803), .Z(n39808) );
  NANDN U40951 ( .A(n39806), .B(n39805), .Z(n39807) );
  AND U40952 ( .A(n39808), .B(n39807), .Z(n39835) );
  NAND U40953 ( .A(n42143), .B(n39809), .Z(n39811) );
  XNOR U40954 ( .A(a[960]), .B(n4209), .Z(n39846) );
  NAND U40955 ( .A(n42144), .B(n39846), .Z(n39810) );
  AND U40956 ( .A(n39811), .B(n39810), .Z(n39861) );
  XOR U40957 ( .A(a[964]), .B(n42012), .Z(n39849) );
  XNOR U40958 ( .A(n39861), .B(n39860), .Z(n39863) );
  XOR U40959 ( .A(a[962]), .B(n42085), .Z(n39853) );
  AND U40960 ( .A(a[958]), .B(b[7]), .Z(n39854) );
  XNOR U40961 ( .A(n39855), .B(n39854), .Z(n39856) );
  AND U40962 ( .A(a[966]), .B(b[0]), .Z(n39814) );
  XNOR U40963 ( .A(n39814), .B(n4071), .Z(n39816) );
  NANDN U40964 ( .A(b[0]), .B(a[965]), .Z(n39815) );
  NAND U40965 ( .A(n39816), .B(n39815), .Z(n39857) );
  XNOR U40966 ( .A(n39856), .B(n39857), .Z(n39862) );
  XOR U40967 ( .A(n39863), .B(n39862), .Z(n39841) );
  NANDN U40968 ( .A(n39818), .B(n39817), .Z(n39822) );
  NANDN U40969 ( .A(n39820), .B(n39819), .Z(n39821) );
  AND U40970 ( .A(n39822), .B(n39821), .Z(n39840) );
  XNOR U40971 ( .A(n39841), .B(n39840), .Z(n39842) );
  NANDN U40972 ( .A(n39824), .B(n39823), .Z(n39828) );
  NAND U40973 ( .A(n39826), .B(n39825), .Z(n39827) );
  NAND U40974 ( .A(n39828), .B(n39827), .Z(n39843) );
  XNOR U40975 ( .A(n39842), .B(n39843), .Z(n39834) );
  XNOR U40976 ( .A(n39835), .B(n39834), .Z(n39836) );
  XNOR U40977 ( .A(n39837), .B(n39836), .Z(n39866) );
  XNOR U40978 ( .A(sreg[1982]), .B(n39866), .Z(n39868) );
  NANDN U40979 ( .A(sreg[1981]), .B(n39829), .Z(n39833) );
  NAND U40980 ( .A(n39831), .B(n39830), .Z(n39832) );
  NAND U40981 ( .A(n39833), .B(n39832), .Z(n39867) );
  XNOR U40982 ( .A(n39868), .B(n39867), .Z(c[1982]) );
  NANDN U40983 ( .A(n39835), .B(n39834), .Z(n39839) );
  NANDN U40984 ( .A(n39837), .B(n39836), .Z(n39838) );
  AND U40985 ( .A(n39839), .B(n39838), .Z(n39874) );
  NANDN U40986 ( .A(n39841), .B(n39840), .Z(n39845) );
  NANDN U40987 ( .A(n39843), .B(n39842), .Z(n39844) );
  AND U40988 ( .A(n39845), .B(n39844), .Z(n39872) );
  NAND U40989 ( .A(n42143), .B(n39846), .Z(n39848) );
  XNOR U40990 ( .A(a[961]), .B(n4209), .Z(n39883) );
  NAND U40991 ( .A(n42144), .B(n39883), .Z(n39847) );
  AND U40992 ( .A(n39848), .B(n39847), .Z(n39898) );
  XOR U40993 ( .A(a[965]), .B(n42012), .Z(n39886) );
  XNOR U40994 ( .A(n39898), .B(n39897), .Z(n39900) );
  AND U40995 ( .A(a[967]), .B(b[0]), .Z(n39850) );
  XNOR U40996 ( .A(n39850), .B(n4071), .Z(n39852) );
  NANDN U40997 ( .A(b[0]), .B(a[966]), .Z(n39851) );
  NAND U40998 ( .A(n39852), .B(n39851), .Z(n39894) );
  XOR U40999 ( .A(a[963]), .B(n42085), .Z(n39890) );
  AND U41000 ( .A(a[959]), .B(b[7]), .Z(n39891) );
  XNOR U41001 ( .A(n39892), .B(n39891), .Z(n39893) );
  XNOR U41002 ( .A(n39894), .B(n39893), .Z(n39899) );
  XOR U41003 ( .A(n39900), .B(n39899), .Z(n39878) );
  NANDN U41004 ( .A(n39855), .B(n39854), .Z(n39859) );
  NANDN U41005 ( .A(n39857), .B(n39856), .Z(n39858) );
  AND U41006 ( .A(n39859), .B(n39858), .Z(n39877) );
  XNOR U41007 ( .A(n39878), .B(n39877), .Z(n39879) );
  NANDN U41008 ( .A(n39861), .B(n39860), .Z(n39865) );
  NAND U41009 ( .A(n39863), .B(n39862), .Z(n39864) );
  NAND U41010 ( .A(n39865), .B(n39864), .Z(n39880) );
  XNOR U41011 ( .A(n39879), .B(n39880), .Z(n39871) );
  XNOR U41012 ( .A(n39872), .B(n39871), .Z(n39873) );
  XNOR U41013 ( .A(n39874), .B(n39873), .Z(n39903) );
  XNOR U41014 ( .A(sreg[1983]), .B(n39903), .Z(n39905) );
  NANDN U41015 ( .A(sreg[1982]), .B(n39866), .Z(n39870) );
  NAND U41016 ( .A(n39868), .B(n39867), .Z(n39869) );
  NAND U41017 ( .A(n39870), .B(n39869), .Z(n39904) );
  XNOR U41018 ( .A(n39905), .B(n39904), .Z(c[1983]) );
  NANDN U41019 ( .A(n39872), .B(n39871), .Z(n39876) );
  NANDN U41020 ( .A(n39874), .B(n39873), .Z(n39875) );
  AND U41021 ( .A(n39876), .B(n39875), .Z(n39911) );
  NANDN U41022 ( .A(n39878), .B(n39877), .Z(n39882) );
  NANDN U41023 ( .A(n39880), .B(n39879), .Z(n39881) );
  AND U41024 ( .A(n39882), .B(n39881), .Z(n39909) );
  NAND U41025 ( .A(n42143), .B(n39883), .Z(n39885) );
  XNOR U41026 ( .A(a[962]), .B(n4209), .Z(n39920) );
  NAND U41027 ( .A(n42144), .B(n39920), .Z(n39884) );
  AND U41028 ( .A(n39885), .B(n39884), .Z(n39935) );
  XOR U41029 ( .A(a[966]), .B(n42012), .Z(n39923) );
  XNOR U41030 ( .A(n39935), .B(n39934), .Z(n39937) );
  AND U41031 ( .A(a[968]), .B(b[0]), .Z(n39887) );
  XNOR U41032 ( .A(n39887), .B(n4071), .Z(n39889) );
  NANDN U41033 ( .A(b[0]), .B(a[967]), .Z(n39888) );
  NAND U41034 ( .A(n39889), .B(n39888), .Z(n39931) );
  XOR U41035 ( .A(a[964]), .B(n42085), .Z(n39924) );
  AND U41036 ( .A(a[960]), .B(b[7]), .Z(n39928) );
  XNOR U41037 ( .A(n39929), .B(n39928), .Z(n39930) );
  XNOR U41038 ( .A(n39931), .B(n39930), .Z(n39936) );
  XOR U41039 ( .A(n39937), .B(n39936), .Z(n39915) );
  NANDN U41040 ( .A(n39892), .B(n39891), .Z(n39896) );
  NANDN U41041 ( .A(n39894), .B(n39893), .Z(n39895) );
  AND U41042 ( .A(n39896), .B(n39895), .Z(n39914) );
  XNOR U41043 ( .A(n39915), .B(n39914), .Z(n39916) );
  NANDN U41044 ( .A(n39898), .B(n39897), .Z(n39902) );
  NAND U41045 ( .A(n39900), .B(n39899), .Z(n39901) );
  NAND U41046 ( .A(n39902), .B(n39901), .Z(n39917) );
  XNOR U41047 ( .A(n39916), .B(n39917), .Z(n39908) );
  XNOR U41048 ( .A(n39909), .B(n39908), .Z(n39910) );
  XNOR U41049 ( .A(n39911), .B(n39910), .Z(n39940) );
  XNOR U41050 ( .A(sreg[1984]), .B(n39940), .Z(n39942) );
  NANDN U41051 ( .A(sreg[1983]), .B(n39903), .Z(n39907) );
  NAND U41052 ( .A(n39905), .B(n39904), .Z(n39906) );
  NAND U41053 ( .A(n39907), .B(n39906), .Z(n39941) );
  XNOR U41054 ( .A(n39942), .B(n39941), .Z(c[1984]) );
  NANDN U41055 ( .A(n39909), .B(n39908), .Z(n39913) );
  NANDN U41056 ( .A(n39911), .B(n39910), .Z(n39912) );
  AND U41057 ( .A(n39913), .B(n39912), .Z(n39948) );
  NANDN U41058 ( .A(n39915), .B(n39914), .Z(n39919) );
  NANDN U41059 ( .A(n39917), .B(n39916), .Z(n39918) );
  AND U41060 ( .A(n39919), .B(n39918), .Z(n39946) );
  NAND U41061 ( .A(n42143), .B(n39920), .Z(n39922) );
  XNOR U41062 ( .A(a[963]), .B(n4209), .Z(n39957) );
  NAND U41063 ( .A(n42144), .B(n39957), .Z(n39921) );
  AND U41064 ( .A(n39922), .B(n39921), .Z(n39972) );
  XOR U41065 ( .A(a[967]), .B(n42012), .Z(n39960) );
  XNOR U41066 ( .A(n39972), .B(n39971), .Z(n39974) );
  XOR U41067 ( .A(a[965]), .B(n42085), .Z(n39964) );
  AND U41068 ( .A(a[961]), .B(b[7]), .Z(n39965) );
  XNOR U41069 ( .A(n39966), .B(n39965), .Z(n39967) );
  AND U41070 ( .A(a[969]), .B(b[0]), .Z(n39925) );
  XNOR U41071 ( .A(n39925), .B(n4071), .Z(n39927) );
  NANDN U41072 ( .A(b[0]), .B(a[968]), .Z(n39926) );
  NAND U41073 ( .A(n39927), .B(n39926), .Z(n39968) );
  XNOR U41074 ( .A(n39967), .B(n39968), .Z(n39973) );
  XOR U41075 ( .A(n39974), .B(n39973), .Z(n39952) );
  NANDN U41076 ( .A(n39929), .B(n39928), .Z(n39933) );
  NANDN U41077 ( .A(n39931), .B(n39930), .Z(n39932) );
  AND U41078 ( .A(n39933), .B(n39932), .Z(n39951) );
  XNOR U41079 ( .A(n39952), .B(n39951), .Z(n39953) );
  NANDN U41080 ( .A(n39935), .B(n39934), .Z(n39939) );
  NAND U41081 ( .A(n39937), .B(n39936), .Z(n39938) );
  NAND U41082 ( .A(n39939), .B(n39938), .Z(n39954) );
  XNOR U41083 ( .A(n39953), .B(n39954), .Z(n39945) );
  XNOR U41084 ( .A(n39946), .B(n39945), .Z(n39947) );
  XNOR U41085 ( .A(n39948), .B(n39947), .Z(n39977) );
  XNOR U41086 ( .A(sreg[1985]), .B(n39977), .Z(n39979) );
  NANDN U41087 ( .A(sreg[1984]), .B(n39940), .Z(n39944) );
  NAND U41088 ( .A(n39942), .B(n39941), .Z(n39943) );
  NAND U41089 ( .A(n39944), .B(n39943), .Z(n39978) );
  XNOR U41090 ( .A(n39979), .B(n39978), .Z(c[1985]) );
  NANDN U41091 ( .A(n39946), .B(n39945), .Z(n39950) );
  NANDN U41092 ( .A(n39948), .B(n39947), .Z(n39949) );
  AND U41093 ( .A(n39950), .B(n39949), .Z(n39985) );
  NANDN U41094 ( .A(n39952), .B(n39951), .Z(n39956) );
  NANDN U41095 ( .A(n39954), .B(n39953), .Z(n39955) );
  AND U41096 ( .A(n39956), .B(n39955), .Z(n39983) );
  NAND U41097 ( .A(n42143), .B(n39957), .Z(n39959) );
  XNOR U41098 ( .A(a[964]), .B(n4209), .Z(n39994) );
  NAND U41099 ( .A(n42144), .B(n39994), .Z(n39958) );
  AND U41100 ( .A(n39959), .B(n39958), .Z(n40009) );
  XOR U41101 ( .A(a[968]), .B(n42012), .Z(n39997) );
  XNOR U41102 ( .A(n40009), .B(n40008), .Z(n40011) );
  AND U41103 ( .A(a[970]), .B(b[0]), .Z(n39961) );
  XNOR U41104 ( .A(n39961), .B(n4071), .Z(n39963) );
  NANDN U41105 ( .A(b[0]), .B(a[969]), .Z(n39962) );
  NAND U41106 ( .A(n39963), .B(n39962), .Z(n40005) );
  XOR U41107 ( .A(a[966]), .B(n42085), .Z(n39998) );
  AND U41108 ( .A(a[962]), .B(b[7]), .Z(n40002) );
  XNOR U41109 ( .A(n40003), .B(n40002), .Z(n40004) );
  XNOR U41110 ( .A(n40005), .B(n40004), .Z(n40010) );
  XOR U41111 ( .A(n40011), .B(n40010), .Z(n39989) );
  NANDN U41112 ( .A(n39966), .B(n39965), .Z(n39970) );
  NANDN U41113 ( .A(n39968), .B(n39967), .Z(n39969) );
  AND U41114 ( .A(n39970), .B(n39969), .Z(n39988) );
  XNOR U41115 ( .A(n39989), .B(n39988), .Z(n39990) );
  NANDN U41116 ( .A(n39972), .B(n39971), .Z(n39976) );
  NAND U41117 ( .A(n39974), .B(n39973), .Z(n39975) );
  NAND U41118 ( .A(n39976), .B(n39975), .Z(n39991) );
  XNOR U41119 ( .A(n39990), .B(n39991), .Z(n39982) );
  XNOR U41120 ( .A(n39983), .B(n39982), .Z(n39984) );
  XNOR U41121 ( .A(n39985), .B(n39984), .Z(n40014) );
  XNOR U41122 ( .A(sreg[1986]), .B(n40014), .Z(n40016) );
  NANDN U41123 ( .A(sreg[1985]), .B(n39977), .Z(n39981) );
  NAND U41124 ( .A(n39979), .B(n39978), .Z(n39980) );
  NAND U41125 ( .A(n39981), .B(n39980), .Z(n40015) );
  XNOR U41126 ( .A(n40016), .B(n40015), .Z(c[1986]) );
  NANDN U41127 ( .A(n39983), .B(n39982), .Z(n39987) );
  NANDN U41128 ( .A(n39985), .B(n39984), .Z(n39986) );
  AND U41129 ( .A(n39987), .B(n39986), .Z(n40022) );
  NANDN U41130 ( .A(n39989), .B(n39988), .Z(n39993) );
  NANDN U41131 ( .A(n39991), .B(n39990), .Z(n39992) );
  AND U41132 ( .A(n39993), .B(n39992), .Z(n40020) );
  NAND U41133 ( .A(n42143), .B(n39994), .Z(n39996) );
  XNOR U41134 ( .A(a[965]), .B(n4209), .Z(n40031) );
  NAND U41135 ( .A(n42144), .B(n40031), .Z(n39995) );
  AND U41136 ( .A(n39996), .B(n39995), .Z(n40046) );
  XOR U41137 ( .A(a[969]), .B(n42012), .Z(n40034) );
  XNOR U41138 ( .A(n40046), .B(n40045), .Z(n40048) );
  XOR U41139 ( .A(a[967]), .B(n42085), .Z(n40035) );
  AND U41140 ( .A(a[963]), .B(b[7]), .Z(n40039) );
  XNOR U41141 ( .A(n40040), .B(n40039), .Z(n40041) );
  AND U41142 ( .A(a[971]), .B(b[0]), .Z(n39999) );
  XNOR U41143 ( .A(n39999), .B(n4071), .Z(n40001) );
  NANDN U41144 ( .A(b[0]), .B(a[970]), .Z(n40000) );
  NAND U41145 ( .A(n40001), .B(n40000), .Z(n40042) );
  XNOR U41146 ( .A(n40041), .B(n40042), .Z(n40047) );
  XOR U41147 ( .A(n40048), .B(n40047), .Z(n40026) );
  NANDN U41148 ( .A(n40003), .B(n40002), .Z(n40007) );
  NANDN U41149 ( .A(n40005), .B(n40004), .Z(n40006) );
  AND U41150 ( .A(n40007), .B(n40006), .Z(n40025) );
  XNOR U41151 ( .A(n40026), .B(n40025), .Z(n40027) );
  NANDN U41152 ( .A(n40009), .B(n40008), .Z(n40013) );
  NAND U41153 ( .A(n40011), .B(n40010), .Z(n40012) );
  NAND U41154 ( .A(n40013), .B(n40012), .Z(n40028) );
  XNOR U41155 ( .A(n40027), .B(n40028), .Z(n40019) );
  XNOR U41156 ( .A(n40020), .B(n40019), .Z(n40021) );
  XNOR U41157 ( .A(n40022), .B(n40021), .Z(n40051) );
  XNOR U41158 ( .A(sreg[1987]), .B(n40051), .Z(n40053) );
  NANDN U41159 ( .A(sreg[1986]), .B(n40014), .Z(n40018) );
  NAND U41160 ( .A(n40016), .B(n40015), .Z(n40017) );
  NAND U41161 ( .A(n40018), .B(n40017), .Z(n40052) );
  XNOR U41162 ( .A(n40053), .B(n40052), .Z(c[1987]) );
  NANDN U41163 ( .A(n40020), .B(n40019), .Z(n40024) );
  NANDN U41164 ( .A(n40022), .B(n40021), .Z(n40023) );
  AND U41165 ( .A(n40024), .B(n40023), .Z(n40059) );
  NANDN U41166 ( .A(n40026), .B(n40025), .Z(n40030) );
  NANDN U41167 ( .A(n40028), .B(n40027), .Z(n40029) );
  AND U41168 ( .A(n40030), .B(n40029), .Z(n40057) );
  NAND U41169 ( .A(n42143), .B(n40031), .Z(n40033) );
  XNOR U41170 ( .A(a[966]), .B(n4209), .Z(n40068) );
  NAND U41171 ( .A(n42144), .B(n40068), .Z(n40032) );
  AND U41172 ( .A(n40033), .B(n40032), .Z(n40083) );
  XOR U41173 ( .A(a[970]), .B(n42012), .Z(n40071) );
  XNOR U41174 ( .A(n40083), .B(n40082), .Z(n40085) );
  XOR U41175 ( .A(a[968]), .B(n42085), .Z(n40072) );
  AND U41176 ( .A(a[964]), .B(b[7]), .Z(n40076) );
  XNOR U41177 ( .A(n40077), .B(n40076), .Z(n40078) );
  AND U41178 ( .A(a[972]), .B(b[0]), .Z(n40036) );
  XNOR U41179 ( .A(n40036), .B(n4071), .Z(n40038) );
  NANDN U41180 ( .A(b[0]), .B(a[971]), .Z(n40037) );
  NAND U41181 ( .A(n40038), .B(n40037), .Z(n40079) );
  XNOR U41182 ( .A(n40078), .B(n40079), .Z(n40084) );
  XOR U41183 ( .A(n40085), .B(n40084), .Z(n40063) );
  NANDN U41184 ( .A(n40040), .B(n40039), .Z(n40044) );
  NANDN U41185 ( .A(n40042), .B(n40041), .Z(n40043) );
  AND U41186 ( .A(n40044), .B(n40043), .Z(n40062) );
  XNOR U41187 ( .A(n40063), .B(n40062), .Z(n40064) );
  NANDN U41188 ( .A(n40046), .B(n40045), .Z(n40050) );
  NAND U41189 ( .A(n40048), .B(n40047), .Z(n40049) );
  NAND U41190 ( .A(n40050), .B(n40049), .Z(n40065) );
  XNOR U41191 ( .A(n40064), .B(n40065), .Z(n40056) );
  XNOR U41192 ( .A(n40057), .B(n40056), .Z(n40058) );
  XNOR U41193 ( .A(n40059), .B(n40058), .Z(n40088) );
  XNOR U41194 ( .A(sreg[1988]), .B(n40088), .Z(n40090) );
  NANDN U41195 ( .A(sreg[1987]), .B(n40051), .Z(n40055) );
  NAND U41196 ( .A(n40053), .B(n40052), .Z(n40054) );
  NAND U41197 ( .A(n40055), .B(n40054), .Z(n40089) );
  XNOR U41198 ( .A(n40090), .B(n40089), .Z(c[1988]) );
  NANDN U41199 ( .A(n40057), .B(n40056), .Z(n40061) );
  NANDN U41200 ( .A(n40059), .B(n40058), .Z(n40060) );
  AND U41201 ( .A(n40061), .B(n40060), .Z(n40096) );
  NANDN U41202 ( .A(n40063), .B(n40062), .Z(n40067) );
  NANDN U41203 ( .A(n40065), .B(n40064), .Z(n40066) );
  AND U41204 ( .A(n40067), .B(n40066), .Z(n40094) );
  NAND U41205 ( .A(n42143), .B(n40068), .Z(n40070) );
  XNOR U41206 ( .A(a[967]), .B(n4210), .Z(n40105) );
  NAND U41207 ( .A(n42144), .B(n40105), .Z(n40069) );
  AND U41208 ( .A(n40070), .B(n40069), .Z(n40120) );
  XOR U41209 ( .A(a[971]), .B(n42012), .Z(n40108) );
  XNOR U41210 ( .A(n40120), .B(n40119), .Z(n40122) );
  XOR U41211 ( .A(a[969]), .B(n42085), .Z(n40112) );
  AND U41212 ( .A(a[965]), .B(b[7]), .Z(n40113) );
  XNOR U41213 ( .A(n40114), .B(n40113), .Z(n40115) );
  AND U41214 ( .A(a[973]), .B(b[0]), .Z(n40073) );
  XNOR U41215 ( .A(n40073), .B(n4071), .Z(n40075) );
  NANDN U41216 ( .A(b[0]), .B(a[972]), .Z(n40074) );
  NAND U41217 ( .A(n40075), .B(n40074), .Z(n40116) );
  XNOR U41218 ( .A(n40115), .B(n40116), .Z(n40121) );
  XOR U41219 ( .A(n40122), .B(n40121), .Z(n40100) );
  NANDN U41220 ( .A(n40077), .B(n40076), .Z(n40081) );
  NANDN U41221 ( .A(n40079), .B(n40078), .Z(n40080) );
  AND U41222 ( .A(n40081), .B(n40080), .Z(n40099) );
  XNOR U41223 ( .A(n40100), .B(n40099), .Z(n40101) );
  NANDN U41224 ( .A(n40083), .B(n40082), .Z(n40087) );
  NAND U41225 ( .A(n40085), .B(n40084), .Z(n40086) );
  NAND U41226 ( .A(n40087), .B(n40086), .Z(n40102) );
  XNOR U41227 ( .A(n40101), .B(n40102), .Z(n40093) );
  XNOR U41228 ( .A(n40094), .B(n40093), .Z(n40095) );
  XNOR U41229 ( .A(n40096), .B(n40095), .Z(n40125) );
  XNOR U41230 ( .A(sreg[1989]), .B(n40125), .Z(n40127) );
  NANDN U41231 ( .A(sreg[1988]), .B(n40088), .Z(n40092) );
  NAND U41232 ( .A(n40090), .B(n40089), .Z(n40091) );
  NAND U41233 ( .A(n40092), .B(n40091), .Z(n40126) );
  XNOR U41234 ( .A(n40127), .B(n40126), .Z(c[1989]) );
  NANDN U41235 ( .A(n40094), .B(n40093), .Z(n40098) );
  NANDN U41236 ( .A(n40096), .B(n40095), .Z(n40097) );
  AND U41237 ( .A(n40098), .B(n40097), .Z(n40133) );
  NANDN U41238 ( .A(n40100), .B(n40099), .Z(n40104) );
  NANDN U41239 ( .A(n40102), .B(n40101), .Z(n40103) );
  AND U41240 ( .A(n40104), .B(n40103), .Z(n40131) );
  NAND U41241 ( .A(n42143), .B(n40105), .Z(n40107) );
  XNOR U41242 ( .A(a[968]), .B(n4210), .Z(n40142) );
  NAND U41243 ( .A(n42144), .B(n40142), .Z(n40106) );
  AND U41244 ( .A(n40107), .B(n40106), .Z(n40157) );
  XOR U41245 ( .A(a[972]), .B(n42012), .Z(n40145) );
  XNOR U41246 ( .A(n40157), .B(n40156), .Z(n40159) );
  AND U41247 ( .A(a[974]), .B(b[0]), .Z(n40109) );
  XNOR U41248 ( .A(n40109), .B(n4071), .Z(n40111) );
  NANDN U41249 ( .A(b[0]), .B(a[973]), .Z(n40110) );
  NAND U41250 ( .A(n40111), .B(n40110), .Z(n40153) );
  XOR U41251 ( .A(a[970]), .B(n42085), .Z(n40149) );
  AND U41252 ( .A(a[966]), .B(b[7]), .Z(n40150) );
  XNOR U41253 ( .A(n40151), .B(n40150), .Z(n40152) );
  XNOR U41254 ( .A(n40153), .B(n40152), .Z(n40158) );
  XOR U41255 ( .A(n40159), .B(n40158), .Z(n40137) );
  NANDN U41256 ( .A(n40114), .B(n40113), .Z(n40118) );
  NANDN U41257 ( .A(n40116), .B(n40115), .Z(n40117) );
  AND U41258 ( .A(n40118), .B(n40117), .Z(n40136) );
  XNOR U41259 ( .A(n40137), .B(n40136), .Z(n40138) );
  NANDN U41260 ( .A(n40120), .B(n40119), .Z(n40124) );
  NAND U41261 ( .A(n40122), .B(n40121), .Z(n40123) );
  NAND U41262 ( .A(n40124), .B(n40123), .Z(n40139) );
  XNOR U41263 ( .A(n40138), .B(n40139), .Z(n40130) );
  XNOR U41264 ( .A(n40131), .B(n40130), .Z(n40132) );
  XNOR U41265 ( .A(n40133), .B(n40132), .Z(n40162) );
  XNOR U41266 ( .A(sreg[1990]), .B(n40162), .Z(n40164) );
  NANDN U41267 ( .A(sreg[1989]), .B(n40125), .Z(n40129) );
  NAND U41268 ( .A(n40127), .B(n40126), .Z(n40128) );
  NAND U41269 ( .A(n40129), .B(n40128), .Z(n40163) );
  XNOR U41270 ( .A(n40164), .B(n40163), .Z(c[1990]) );
  NANDN U41271 ( .A(n40131), .B(n40130), .Z(n40135) );
  NANDN U41272 ( .A(n40133), .B(n40132), .Z(n40134) );
  AND U41273 ( .A(n40135), .B(n40134), .Z(n40170) );
  NANDN U41274 ( .A(n40137), .B(n40136), .Z(n40141) );
  NANDN U41275 ( .A(n40139), .B(n40138), .Z(n40140) );
  AND U41276 ( .A(n40141), .B(n40140), .Z(n40168) );
  NAND U41277 ( .A(n42143), .B(n40142), .Z(n40144) );
  XNOR U41278 ( .A(a[969]), .B(n4210), .Z(n40179) );
  NAND U41279 ( .A(n42144), .B(n40179), .Z(n40143) );
  AND U41280 ( .A(n40144), .B(n40143), .Z(n40194) );
  XOR U41281 ( .A(a[973]), .B(n42012), .Z(n40182) );
  XNOR U41282 ( .A(n40194), .B(n40193), .Z(n40196) );
  AND U41283 ( .A(a[975]), .B(b[0]), .Z(n40146) );
  XNOR U41284 ( .A(n40146), .B(n4071), .Z(n40148) );
  NANDN U41285 ( .A(b[0]), .B(a[974]), .Z(n40147) );
  NAND U41286 ( .A(n40148), .B(n40147), .Z(n40190) );
  XOR U41287 ( .A(a[971]), .B(n42085), .Z(n40186) );
  AND U41288 ( .A(a[967]), .B(b[7]), .Z(n40187) );
  XNOR U41289 ( .A(n40188), .B(n40187), .Z(n40189) );
  XNOR U41290 ( .A(n40190), .B(n40189), .Z(n40195) );
  XOR U41291 ( .A(n40196), .B(n40195), .Z(n40174) );
  NANDN U41292 ( .A(n40151), .B(n40150), .Z(n40155) );
  NANDN U41293 ( .A(n40153), .B(n40152), .Z(n40154) );
  AND U41294 ( .A(n40155), .B(n40154), .Z(n40173) );
  XNOR U41295 ( .A(n40174), .B(n40173), .Z(n40175) );
  NANDN U41296 ( .A(n40157), .B(n40156), .Z(n40161) );
  NAND U41297 ( .A(n40159), .B(n40158), .Z(n40160) );
  NAND U41298 ( .A(n40161), .B(n40160), .Z(n40176) );
  XNOR U41299 ( .A(n40175), .B(n40176), .Z(n40167) );
  XNOR U41300 ( .A(n40168), .B(n40167), .Z(n40169) );
  XNOR U41301 ( .A(n40170), .B(n40169), .Z(n40199) );
  XNOR U41302 ( .A(sreg[1991]), .B(n40199), .Z(n40201) );
  NANDN U41303 ( .A(sreg[1990]), .B(n40162), .Z(n40166) );
  NAND U41304 ( .A(n40164), .B(n40163), .Z(n40165) );
  NAND U41305 ( .A(n40166), .B(n40165), .Z(n40200) );
  XNOR U41306 ( .A(n40201), .B(n40200), .Z(c[1991]) );
  NANDN U41307 ( .A(n40168), .B(n40167), .Z(n40172) );
  NANDN U41308 ( .A(n40170), .B(n40169), .Z(n40171) );
  AND U41309 ( .A(n40172), .B(n40171), .Z(n40207) );
  NANDN U41310 ( .A(n40174), .B(n40173), .Z(n40178) );
  NANDN U41311 ( .A(n40176), .B(n40175), .Z(n40177) );
  AND U41312 ( .A(n40178), .B(n40177), .Z(n40205) );
  NAND U41313 ( .A(n42143), .B(n40179), .Z(n40181) );
  XNOR U41314 ( .A(a[970]), .B(n4210), .Z(n40216) );
  NAND U41315 ( .A(n42144), .B(n40216), .Z(n40180) );
  AND U41316 ( .A(n40181), .B(n40180), .Z(n40231) );
  XOR U41317 ( .A(a[974]), .B(n42012), .Z(n40219) );
  XNOR U41318 ( .A(n40231), .B(n40230), .Z(n40233) );
  AND U41319 ( .A(a[976]), .B(b[0]), .Z(n40183) );
  XNOR U41320 ( .A(n40183), .B(n4071), .Z(n40185) );
  NANDN U41321 ( .A(b[0]), .B(a[975]), .Z(n40184) );
  NAND U41322 ( .A(n40185), .B(n40184), .Z(n40227) );
  XOR U41323 ( .A(a[972]), .B(n42085), .Z(n40223) );
  AND U41324 ( .A(a[968]), .B(b[7]), .Z(n40224) );
  XNOR U41325 ( .A(n40225), .B(n40224), .Z(n40226) );
  XNOR U41326 ( .A(n40227), .B(n40226), .Z(n40232) );
  XOR U41327 ( .A(n40233), .B(n40232), .Z(n40211) );
  NANDN U41328 ( .A(n40188), .B(n40187), .Z(n40192) );
  NANDN U41329 ( .A(n40190), .B(n40189), .Z(n40191) );
  AND U41330 ( .A(n40192), .B(n40191), .Z(n40210) );
  XNOR U41331 ( .A(n40211), .B(n40210), .Z(n40212) );
  NANDN U41332 ( .A(n40194), .B(n40193), .Z(n40198) );
  NAND U41333 ( .A(n40196), .B(n40195), .Z(n40197) );
  NAND U41334 ( .A(n40198), .B(n40197), .Z(n40213) );
  XNOR U41335 ( .A(n40212), .B(n40213), .Z(n40204) );
  XNOR U41336 ( .A(n40205), .B(n40204), .Z(n40206) );
  XNOR U41337 ( .A(n40207), .B(n40206), .Z(n40236) );
  XNOR U41338 ( .A(sreg[1992]), .B(n40236), .Z(n40238) );
  NANDN U41339 ( .A(sreg[1991]), .B(n40199), .Z(n40203) );
  NAND U41340 ( .A(n40201), .B(n40200), .Z(n40202) );
  NAND U41341 ( .A(n40203), .B(n40202), .Z(n40237) );
  XNOR U41342 ( .A(n40238), .B(n40237), .Z(c[1992]) );
  NANDN U41343 ( .A(n40205), .B(n40204), .Z(n40209) );
  NANDN U41344 ( .A(n40207), .B(n40206), .Z(n40208) );
  AND U41345 ( .A(n40209), .B(n40208), .Z(n40244) );
  NANDN U41346 ( .A(n40211), .B(n40210), .Z(n40215) );
  NANDN U41347 ( .A(n40213), .B(n40212), .Z(n40214) );
  AND U41348 ( .A(n40215), .B(n40214), .Z(n40242) );
  NAND U41349 ( .A(n42143), .B(n40216), .Z(n40218) );
  XNOR U41350 ( .A(a[971]), .B(n4210), .Z(n40253) );
  NAND U41351 ( .A(n42144), .B(n40253), .Z(n40217) );
  AND U41352 ( .A(n40218), .B(n40217), .Z(n40268) );
  XOR U41353 ( .A(a[975]), .B(n42012), .Z(n40256) );
  XNOR U41354 ( .A(n40268), .B(n40267), .Z(n40270) );
  AND U41355 ( .A(a[977]), .B(b[0]), .Z(n40220) );
  XNOR U41356 ( .A(n40220), .B(n4071), .Z(n40222) );
  NANDN U41357 ( .A(b[0]), .B(a[976]), .Z(n40221) );
  NAND U41358 ( .A(n40222), .B(n40221), .Z(n40264) );
  XOR U41359 ( .A(a[973]), .B(n42085), .Z(n40260) );
  AND U41360 ( .A(a[969]), .B(b[7]), .Z(n40261) );
  XNOR U41361 ( .A(n40262), .B(n40261), .Z(n40263) );
  XNOR U41362 ( .A(n40264), .B(n40263), .Z(n40269) );
  XOR U41363 ( .A(n40270), .B(n40269), .Z(n40248) );
  NANDN U41364 ( .A(n40225), .B(n40224), .Z(n40229) );
  NANDN U41365 ( .A(n40227), .B(n40226), .Z(n40228) );
  AND U41366 ( .A(n40229), .B(n40228), .Z(n40247) );
  XNOR U41367 ( .A(n40248), .B(n40247), .Z(n40249) );
  NANDN U41368 ( .A(n40231), .B(n40230), .Z(n40235) );
  NAND U41369 ( .A(n40233), .B(n40232), .Z(n40234) );
  NAND U41370 ( .A(n40235), .B(n40234), .Z(n40250) );
  XNOR U41371 ( .A(n40249), .B(n40250), .Z(n40241) );
  XNOR U41372 ( .A(n40242), .B(n40241), .Z(n40243) );
  XNOR U41373 ( .A(n40244), .B(n40243), .Z(n40273) );
  XNOR U41374 ( .A(sreg[1993]), .B(n40273), .Z(n40275) );
  NANDN U41375 ( .A(sreg[1992]), .B(n40236), .Z(n40240) );
  NAND U41376 ( .A(n40238), .B(n40237), .Z(n40239) );
  NAND U41377 ( .A(n40240), .B(n40239), .Z(n40274) );
  XNOR U41378 ( .A(n40275), .B(n40274), .Z(c[1993]) );
  NANDN U41379 ( .A(n40242), .B(n40241), .Z(n40246) );
  NANDN U41380 ( .A(n40244), .B(n40243), .Z(n40245) );
  AND U41381 ( .A(n40246), .B(n40245), .Z(n40281) );
  NANDN U41382 ( .A(n40248), .B(n40247), .Z(n40252) );
  NANDN U41383 ( .A(n40250), .B(n40249), .Z(n40251) );
  AND U41384 ( .A(n40252), .B(n40251), .Z(n40279) );
  NAND U41385 ( .A(n42143), .B(n40253), .Z(n40255) );
  XNOR U41386 ( .A(a[972]), .B(n4210), .Z(n40290) );
  NAND U41387 ( .A(n42144), .B(n40290), .Z(n40254) );
  AND U41388 ( .A(n40255), .B(n40254), .Z(n40305) );
  XOR U41389 ( .A(a[976]), .B(n42012), .Z(n40293) );
  XNOR U41390 ( .A(n40305), .B(n40304), .Z(n40307) );
  AND U41391 ( .A(a[978]), .B(b[0]), .Z(n40257) );
  XNOR U41392 ( .A(n40257), .B(n4071), .Z(n40259) );
  NANDN U41393 ( .A(b[0]), .B(a[977]), .Z(n40258) );
  NAND U41394 ( .A(n40259), .B(n40258), .Z(n40301) );
  XOR U41395 ( .A(a[974]), .B(n42085), .Z(n40294) );
  AND U41396 ( .A(a[970]), .B(b[7]), .Z(n40298) );
  XNOR U41397 ( .A(n40299), .B(n40298), .Z(n40300) );
  XNOR U41398 ( .A(n40301), .B(n40300), .Z(n40306) );
  XOR U41399 ( .A(n40307), .B(n40306), .Z(n40285) );
  NANDN U41400 ( .A(n40262), .B(n40261), .Z(n40266) );
  NANDN U41401 ( .A(n40264), .B(n40263), .Z(n40265) );
  AND U41402 ( .A(n40266), .B(n40265), .Z(n40284) );
  XNOR U41403 ( .A(n40285), .B(n40284), .Z(n40286) );
  NANDN U41404 ( .A(n40268), .B(n40267), .Z(n40272) );
  NAND U41405 ( .A(n40270), .B(n40269), .Z(n40271) );
  NAND U41406 ( .A(n40272), .B(n40271), .Z(n40287) );
  XNOR U41407 ( .A(n40286), .B(n40287), .Z(n40278) );
  XNOR U41408 ( .A(n40279), .B(n40278), .Z(n40280) );
  XNOR U41409 ( .A(n40281), .B(n40280), .Z(n40310) );
  XNOR U41410 ( .A(sreg[1994]), .B(n40310), .Z(n40312) );
  NANDN U41411 ( .A(sreg[1993]), .B(n40273), .Z(n40277) );
  NAND U41412 ( .A(n40275), .B(n40274), .Z(n40276) );
  NAND U41413 ( .A(n40277), .B(n40276), .Z(n40311) );
  XNOR U41414 ( .A(n40312), .B(n40311), .Z(c[1994]) );
  NANDN U41415 ( .A(n40279), .B(n40278), .Z(n40283) );
  NANDN U41416 ( .A(n40281), .B(n40280), .Z(n40282) );
  AND U41417 ( .A(n40283), .B(n40282), .Z(n40318) );
  NANDN U41418 ( .A(n40285), .B(n40284), .Z(n40289) );
  NANDN U41419 ( .A(n40287), .B(n40286), .Z(n40288) );
  AND U41420 ( .A(n40289), .B(n40288), .Z(n40316) );
  NAND U41421 ( .A(n42143), .B(n40290), .Z(n40292) );
  XNOR U41422 ( .A(a[973]), .B(n4210), .Z(n40327) );
  NAND U41423 ( .A(n42144), .B(n40327), .Z(n40291) );
  AND U41424 ( .A(n40292), .B(n40291), .Z(n40342) );
  XOR U41425 ( .A(a[977]), .B(n42012), .Z(n40330) );
  XNOR U41426 ( .A(n40342), .B(n40341), .Z(n40344) );
  XOR U41427 ( .A(a[975]), .B(n42085), .Z(n40334) );
  AND U41428 ( .A(a[971]), .B(b[7]), .Z(n40335) );
  XNOR U41429 ( .A(n40336), .B(n40335), .Z(n40337) );
  AND U41430 ( .A(a[979]), .B(b[0]), .Z(n40295) );
  XNOR U41431 ( .A(n40295), .B(n4071), .Z(n40297) );
  NANDN U41432 ( .A(b[0]), .B(a[978]), .Z(n40296) );
  NAND U41433 ( .A(n40297), .B(n40296), .Z(n40338) );
  XNOR U41434 ( .A(n40337), .B(n40338), .Z(n40343) );
  XOR U41435 ( .A(n40344), .B(n40343), .Z(n40322) );
  NANDN U41436 ( .A(n40299), .B(n40298), .Z(n40303) );
  NANDN U41437 ( .A(n40301), .B(n40300), .Z(n40302) );
  AND U41438 ( .A(n40303), .B(n40302), .Z(n40321) );
  XNOR U41439 ( .A(n40322), .B(n40321), .Z(n40323) );
  NANDN U41440 ( .A(n40305), .B(n40304), .Z(n40309) );
  NAND U41441 ( .A(n40307), .B(n40306), .Z(n40308) );
  NAND U41442 ( .A(n40309), .B(n40308), .Z(n40324) );
  XNOR U41443 ( .A(n40323), .B(n40324), .Z(n40315) );
  XNOR U41444 ( .A(n40316), .B(n40315), .Z(n40317) );
  XNOR U41445 ( .A(n40318), .B(n40317), .Z(n40347) );
  XNOR U41446 ( .A(sreg[1995]), .B(n40347), .Z(n40349) );
  NANDN U41447 ( .A(sreg[1994]), .B(n40310), .Z(n40314) );
  NAND U41448 ( .A(n40312), .B(n40311), .Z(n40313) );
  NAND U41449 ( .A(n40314), .B(n40313), .Z(n40348) );
  XNOR U41450 ( .A(n40349), .B(n40348), .Z(c[1995]) );
  NANDN U41451 ( .A(n40316), .B(n40315), .Z(n40320) );
  NANDN U41452 ( .A(n40318), .B(n40317), .Z(n40319) );
  AND U41453 ( .A(n40320), .B(n40319), .Z(n40355) );
  NANDN U41454 ( .A(n40322), .B(n40321), .Z(n40326) );
  NANDN U41455 ( .A(n40324), .B(n40323), .Z(n40325) );
  AND U41456 ( .A(n40326), .B(n40325), .Z(n40353) );
  NAND U41457 ( .A(n42143), .B(n40327), .Z(n40329) );
  XNOR U41458 ( .A(a[974]), .B(n4211), .Z(n40364) );
  NAND U41459 ( .A(n42144), .B(n40364), .Z(n40328) );
  AND U41460 ( .A(n40329), .B(n40328), .Z(n40379) );
  XOR U41461 ( .A(a[978]), .B(n42012), .Z(n40367) );
  XNOR U41462 ( .A(n40379), .B(n40378), .Z(n40381) );
  AND U41463 ( .A(a[980]), .B(b[0]), .Z(n40331) );
  XNOR U41464 ( .A(n40331), .B(n4071), .Z(n40333) );
  NANDN U41465 ( .A(b[0]), .B(a[979]), .Z(n40332) );
  NAND U41466 ( .A(n40333), .B(n40332), .Z(n40375) );
  XOR U41467 ( .A(a[976]), .B(n42085), .Z(n40368) );
  AND U41468 ( .A(a[972]), .B(b[7]), .Z(n40372) );
  XNOR U41469 ( .A(n40373), .B(n40372), .Z(n40374) );
  XNOR U41470 ( .A(n40375), .B(n40374), .Z(n40380) );
  XOR U41471 ( .A(n40381), .B(n40380), .Z(n40359) );
  NANDN U41472 ( .A(n40336), .B(n40335), .Z(n40340) );
  NANDN U41473 ( .A(n40338), .B(n40337), .Z(n40339) );
  AND U41474 ( .A(n40340), .B(n40339), .Z(n40358) );
  XNOR U41475 ( .A(n40359), .B(n40358), .Z(n40360) );
  NANDN U41476 ( .A(n40342), .B(n40341), .Z(n40346) );
  NAND U41477 ( .A(n40344), .B(n40343), .Z(n40345) );
  NAND U41478 ( .A(n40346), .B(n40345), .Z(n40361) );
  XNOR U41479 ( .A(n40360), .B(n40361), .Z(n40352) );
  XNOR U41480 ( .A(n40353), .B(n40352), .Z(n40354) );
  XNOR U41481 ( .A(n40355), .B(n40354), .Z(n40384) );
  XNOR U41482 ( .A(sreg[1996]), .B(n40384), .Z(n40386) );
  NANDN U41483 ( .A(sreg[1995]), .B(n40347), .Z(n40351) );
  NAND U41484 ( .A(n40349), .B(n40348), .Z(n40350) );
  NAND U41485 ( .A(n40351), .B(n40350), .Z(n40385) );
  XNOR U41486 ( .A(n40386), .B(n40385), .Z(c[1996]) );
  NANDN U41487 ( .A(n40353), .B(n40352), .Z(n40357) );
  NANDN U41488 ( .A(n40355), .B(n40354), .Z(n40356) );
  AND U41489 ( .A(n40357), .B(n40356), .Z(n40392) );
  NANDN U41490 ( .A(n40359), .B(n40358), .Z(n40363) );
  NANDN U41491 ( .A(n40361), .B(n40360), .Z(n40362) );
  AND U41492 ( .A(n40363), .B(n40362), .Z(n40390) );
  NAND U41493 ( .A(n42143), .B(n40364), .Z(n40366) );
  XNOR U41494 ( .A(a[975]), .B(n4211), .Z(n40401) );
  NAND U41495 ( .A(n42144), .B(n40401), .Z(n40365) );
  AND U41496 ( .A(n40366), .B(n40365), .Z(n40416) );
  XOR U41497 ( .A(a[979]), .B(n42012), .Z(n40404) );
  XNOR U41498 ( .A(n40416), .B(n40415), .Z(n40418) );
  XOR U41499 ( .A(a[977]), .B(n42085), .Z(n40408) );
  AND U41500 ( .A(a[973]), .B(b[7]), .Z(n40409) );
  XNOR U41501 ( .A(n40410), .B(n40409), .Z(n40411) );
  AND U41502 ( .A(a[981]), .B(b[0]), .Z(n40369) );
  XNOR U41503 ( .A(n40369), .B(n4071), .Z(n40371) );
  NANDN U41504 ( .A(b[0]), .B(a[980]), .Z(n40370) );
  NAND U41505 ( .A(n40371), .B(n40370), .Z(n40412) );
  XNOR U41506 ( .A(n40411), .B(n40412), .Z(n40417) );
  XOR U41507 ( .A(n40418), .B(n40417), .Z(n40396) );
  NANDN U41508 ( .A(n40373), .B(n40372), .Z(n40377) );
  NANDN U41509 ( .A(n40375), .B(n40374), .Z(n40376) );
  AND U41510 ( .A(n40377), .B(n40376), .Z(n40395) );
  XNOR U41511 ( .A(n40396), .B(n40395), .Z(n40397) );
  NANDN U41512 ( .A(n40379), .B(n40378), .Z(n40383) );
  NAND U41513 ( .A(n40381), .B(n40380), .Z(n40382) );
  NAND U41514 ( .A(n40383), .B(n40382), .Z(n40398) );
  XNOR U41515 ( .A(n40397), .B(n40398), .Z(n40389) );
  XNOR U41516 ( .A(n40390), .B(n40389), .Z(n40391) );
  XNOR U41517 ( .A(n40392), .B(n40391), .Z(n40421) );
  XNOR U41518 ( .A(sreg[1997]), .B(n40421), .Z(n40423) );
  NANDN U41519 ( .A(sreg[1996]), .B(n40384), .Z(n40388) );
  NAND U41520 ( .A(n40386), .B(n40385), .Z(n40387) );
  NAND U41521 ( .A(n40388), .B(n40387), .Z(n40422) );
  XNOR U41522 ( .A(n40423), .B(n40422), .Z(c[1997]) );
  NANDN U41523 ( .A(n40390), .B(n40389), .Z(n40394) );
  NANDN U41524 ( .A(n40392), .B(n40391), .Z(n40393) );
  AND U41525 ( .A(n40394), .B(n40393), .Z(n40429) );
  NANDN U41526 ( .A(n40396), .B(n40395), .Z(n40400) );
  NANDN U41527 ( .A(n40398), .B(n40397), .Z(n40399) );
  AND U41528 ( .A(n40400), .B(n40399), .Z(n40427) );
  NAND U41529 ( .A(n42143), .B(n40401), .Z(n40403) );
  XNOR U41530 ( .A(a[976]), .B(n4211), .Z(n40438) );
  NAND U41531 ( .A(n42144), .B(n40438), .Z(n40402) );
  AND U41532 ( .A(n40403), .B(n40402), .Z(n40453) );
  XOR U41533 ( .A(a[980]), .B(n42012), .Z(n40441) );
  XNOR U41534 ( .A(n40453), .B(n40452), .Z(n40455) );
  AND U41535 ( .A(a[982]), .B(b[0]), .Z(n40405) );
  XNOR U41536 ( .A(n40405), .B(n4071), .Z(n40407) );
  NANDN U41537 ( .A(b[0]), .B(a[981]), .Z(n40406) );
  NAND U41538 ( .A(n40407), .B(n40406), .Z(n40449) );
  XOR U41539 ( .A(a[978]), .B(n42085), .Z(n40445) );
  AND U41540 ( .A(a[974]), .B(b[7]), .Z(n40446) );
  XNOR U41541 ( .A(n40447), .B(n40446), .Z(n40448) );
  XNOR U41542 ( .A(n40449), .B(n40448), .Z(n40454) );
  XOR U41543 ( .A(n40455), .B(n40454), .Z(n40433) );
  NANDN U41544 ( .A(n40410), .B(n40409), .Z(n40414) );
  NANDN U41545 ( .A(n40412), .B(n40411), .Z(n40413) );
  AND U41546 ( .A(n40414), .B(n40413), .Z(n40432) );
  XNOR U41547 ( .A(n40433), .B(n40432), .Z(n40434) );
  NANDN U41548 ( .A(n40416), .B(n40415), .Z(n40420) );
  NAND U41549 ( .A(n40418), .B(n40417), .Z(n40419) );
  NAND U41550 ( .A(n40420), .B(n40419), .Z(n40435) );
  XNOR U41551 ( .A(n40434), .B(n40435), .Z(n40426) );
  XNOR U41552 ( .A(n40427), .B(n40426), .Z(n40428) );
  XNOR U41553 ( .A(n40429), .B(n40428), .Z(n40458) );
  XNOR U41554 ( .A(sreg[1998]), .B(n40458), .Z(n40460) );
  NANDN U41555 ( .A(sreg[1997]), .B(n40421), .Z(n40425) );
  NAND U41556 ( .A(n40423), .B(n40422), .Z(n40424) );
  NAND U41557 ( .A(n40425), .B(n40424), .Z(n40459) );
  XNOR U41558 ( .A(n40460), .B(n40459), .Z(c[1998]) );
  NANDN U41559 ( .A(n40427), .B(n40426), .Z(n40431) );
  NANDN U41560 ( .A(n40429), .B(n40428), .Z(n40430) );
  AND U41561 ( .A(n40431), .B(n40430), .Z(n40466) );
  NANDN U41562 ( .A(n40433), .B(n40432), .Z(n40437) );
  NANDN U41563 ( .A(n40435), .B(n40434), .Z(n40436) );
  AND U41564 ( .A(n40437), .B(n40436), .Z(n40464) );
  NAND U41565 ( .A(n42143), .B(n40438), .Z(n40440) );
  XNOR U41566 ( .A(a[977]), .B(n4211), .Z(n40475) );
  NAND U41567 ( .A(n42144), .B(n40475), .Z(n40439) );
  AND U41568 ( .A(n40440), .B(n40439), .Z(n40490) );
  XOR U41569 ( .A(a[981]), .B(n42012), .Z(n40478) );
  XNOR U41570 ( .A(n40490), .B(n40489), .Z(n40492) );
  AND U41571 ( .A(a[983]), .B(b[0]), .Z(n40442) );
  XNOR U41572 ( .A(n40442), .B(n4071), .Z(n40444) );
  NANDN U41573 ( .A(b[0]), .B(a[982]), .Z(n40443) );
  NAND U41574 ( .A(n40444), .B(n40443), .Z(n40486) );
  XOR U41575 ( .A(a[979]), .B(n42085), .Z(n40482) );
  AND U41576 ( .A(a[975]), .B(b[7]), .Z(n40483) );
  XNOR U41577 ( .A(n40484), .B(n40483), .Z(n40485) );
  XNOR U41578 ( .A(n40486), .B(n40485), .Z(n40491) );
  XOR U41579 ( .A(n40492), .B(n40491), .Z(n40470) );
  NANDN U41580 ( .A(n40447), .B(n40446), .Z(n40451) );
  NANDN U41581 ( .A(n40449), .B(n40448), .Z(n40450) );
  AND U41582 ( .A(n40451), .B(n40450), .Z(n40469) );
  XNOR U41583 ( .A(n40470), .B(n40469), .Z(n40471) );
  NANDN U41584 ( .A(n40453), .B(n40452), .Z(n40457) );
  NAND U41585 ( .A(n40455), .B(n40454), .Z(n40456) );
  NAND U41586 ( .A(n40457), .B(n40456), .Z(n40472) );
  XNOR U41587 ( .A(n40471), .B(n40472), .Z(n40463) );
  XNOR U41588 ( .A(n40464), .B(n40463), .Z(n40465) );
  XNOR U41589 ( .A(n40466), .B(n40465), .Z(n40495) );
  XNOR U41590 ( .A(sreg[1999]), .B(n40495), .Z(n40497) );
  NANDN U41591 ( .A(sreg[1998]), .B(n40458), .Z(n40462) );
  NAND U41592 ( .A(n40460), .B(n40459), .Z(n40461) );
  NAND U41593 ( .A(n40462), .B(n40461), .Z(n40496) );
  XNOR U41594 ( .A(n40497), .B(n40496), .Z(c[1999]) );
  NANDN U41595 ( .A(n40464), .B(n40463), .Z(n40468) );
  NANDN U41596 ( .A(n40466), .B(n40465), .Z(n40467) );
  AND U41597 ( .A(n40468), .B(n40467), .Z(n40503) );
  NANDN U41598 ( .A(n40470), .B(n40469), .Z(n40474) );
  NANDN U41599 ( .A(n40472), .B(n40471), .Z(n40473) );
  AND U41600 ( .A(n40474), .B(n40473), .Z(n40501) );
  NAND U41601 ( .A(n42143), .B(n40475), .Z(n40477) );
  XNOR U41602 ( .A(a[978]), .B(n4211), .Z(n40512) );
  NAND U41603 ( .A(n42144), .B(n40512), .Z(n40476) );
  AND U41604 ( .A(n40477), .B(n40476), .Z(n40527) );
  XOR U41605 ( .A(a[982]), .B(n42012), .Z(n40515) );
  XNOR U41606 ( .A(n40527), .B(n40526), .Z(n40529) );
  AND U41607 ( .A(a[984]), .B(b[0]), .Z(n40479) );
  XNOR U41608 ( .A(n40479), .B(n4071), .Z(n40481) );
  NANDN U41609 ( .A(b[0]), .B(a[983]), .Z(n40480) );
  NAND U41610 ( .A(n40481), .B(n40480), .Z(n40523) );
  XOR U41611 ( .A(a[980]), .B(n42085), .Z(n40519) );
  AND U41612 ( .A(a[976]), .B(b[7]), .Z(n40520) );
  XNOR U41613 ( .A(n40521), .B(n40520), .Z(n40522) );
  XNOR U41614 ( .A(n40523), .B(n40522), .Z(n40528) );
  XOR U41615 ( .A(n40529), .B(n40528), .Z(n40507) );
  NANDN U41616 ( .A(n40484), .B(n40483), .Z(n40488) );
  NANDN U41617 ( .A(n40486), .B(n40485), .Z(n40487) );
  AND U41618 ( .A(n40488), .B(n40487), .Z(n40506) );
  XNOR U41619 ( .A(n40507), .B(n40506), .Z(n40508) );
  NANDN U41620 ( .A(n40490), .B(n40489), .Z(n40494) );
  NAND U41621 ( .A(n40492), .B(n40491), .Z(n40493) );
  NAND U41622 ( .A(n40494), .B(n40493), .Z(n40509) );
  XNOR U41623 ( .A(n40508), .B(n40509), .Z(n40500) );
  XNOR U41624 ( .A(n40501), .B(n40500), .Z(n40502) );
  XNOR U41625 ( .A(n40503), .B(n40502), .Z(n40532) );
  XNOR U41626 ( .A(sreg[2000]), .B(n40532), .Z(n40534) );
  NANDN U41627 ( .A(sreg[1999]), .B(n40495), .Z(n40499) );
  NAND U41628 ( .A(n40497), .B(n40496), .Z(n40498) );
  NAND U41629 ( .A(n40499), .B(n40498), .Z(n40533) );
  XNOR U41630 ( .A(n40534), .B(n40533), .Z(c[2000]) );
  NANDN U41631 ( .A(n40501), .B(n40500), .Z(n40505) );
  NANDN U41632 ( .A(n40503), .B(n40502), .Z(n40504) );
  AND U41633 ( .A(n40505), .B(n40504), .Z(n40540) );
  NANDN U41634 ( .A(n40507), .B(n40506), .Z(n40511) );
  NANDN U41635 ( .A(n40509), .B(n40508), .Z(n40510) );
  AND U41636 ( .A(n40511), .B(n40510), .Z(n40538) );
  NAND U41637 ( .A(n42143), .B(n40512), .Z(n40514) );
  XNOR U41638 ( .A(a[979]), .B(n4211), .Z(n40549) );
  NAND U41639 ( .A(n42144), .B(n40549), .Z(n40513) );
  AND U41640 ( .A(n40514), .B(n40513), .Z(n40564) );
  XOR U41641 ( .A(a[983]), .B(n42012), .Z(n40552) );
  XNOR U41642 ( .A(n40564), .B(n40563), .Z(n40566) );
  AND U41643 ( .A(a[985]), .B(b[0]), .Z(n40516) );
  XNOR U41644 ( .A(n40516), .B(n4071), .Z(n40518) );
  NANDN U41645 ( .A(b[0]), .B(a[984]), .Z(n40517) );
  NAND U41646 ( .A(n40518), .B(n40517), .Z(n40560) );
  XOR U41647 ( .A(a[981]), .B(n42085), .Z(n40556) );
  AND U41648 ( .A(a[977]), .B(b[7]), .Z(n40557) );
  XNOR U41649 ( .A(n40558), .B(n40557), .Z(n40559) );
  XNOR U41650 ( .A(n40560), .B(n40559), .Z(n40565) );
  XOR U41651 ( .A(n40566), .B(n40565), .Z(n40544) );
  NANDN U41652 ( .A(n40521), .B(n40520), .Z(n40525) );
  NANDN U41653 ( .A(n40523), .B(n40522), .Z(n40524) );
  AND U41654 ( .A(n40525), .B(n40524), .Z(n40543) );
  XNOR U41655 ( .A(n40544), .B(n40543), .Z(n40545) );
  NANDN U41656 ( .A(n40527), .B(n40526), .Z(n40531) );
  NAND U41657 ( .A(n40529), .B(n40528), .Z(n40530) );
  NAND U41658 ( .A(n40531), .B(n40530), .Z(n40546) );
  XNOR U41659 ( .A(n40545), .B(n40546), .Z(n40537) );
  XNOR U41660 ( .A(n40538), .B(n40537), .Z(n40539) );
  XNOR U41661 ( .A(n40540), .B(n40539), .Z(n40569) );
  XNOR U41662 ( .A(sreg[2001]), .B(n40569), .Z(n40571) );
  NANDN U41663 ( .A(sreg[2000]), .B(n40532), .Z(n40536) );
  NAND U41664 ( .A(n40534), .B(n40533), .Z(n40535) );
  NAND U41665 ( .A(n40536), .B(n40535), .Z(n40570) );
  XNOR U41666 ( .A(n40571), .B(n40570), .Z(c[2001]) );
  NANDN U41667 ( .A(n40538), .B(n40537), .Z(n40542) );
  NANDN U41668 ( .A(n40540), .B(n40539), .Z(n40541) );
  AND U41669 ( .A(n40542), .B(n40541), .Z(n40577) );
  NANDN U41670 ( .A(n40544), .B(n40543), .Z(n40548) );
  NANDN U41671 ( .A(n40546), .B(n40545), .Z(n40547) );
  AND U41672 ( .A(n40548), .B(n40547), .Z(n40575) );
  NAND U41673 ( .A(n42143), .B(n40549), .Z(n40551) );
  XNOR U41674 ( .A(a[980]), .B(n4211), .Z(n40586) );
  NAND U41675 ( .A(n42144), .B(n40586), .Z(n40550) );
  AND U41676 ( .A(n40551), .B(n40550), .Z(n40601) );
  XOR U41677 ( .A(a[984]), .B(n42012), .Z(n40589) );
  XNOR U41678 ( .A(n40601), .B(n40600), .Z(n40603) );
  AND U41679 ( .A(a[986]), .B(b[0]), .Z(n40553) );
  XNOR U41680 ( .A(n40553), .B(n4071), .Z(n40555) );
  NANDN U41681 ( .A(b[0]), .B(a[985]), .Z(n40554) );
  NAND U41682 ( .A(n40555), .B(n40554), .Z(n40597) );
  XOR U41683 ( .A(a[982]), .B(n42085), .Z(n40593) );
  AND U41684 ( .A(a[978]), .B(b[7]), .Z(n40594) );
  XNOR U41685 ( .A(n40595), .B(n40594), .Z(n40596) );
  XNOR U41686 ( .A(n40597), .B(n40596), .Z(n40602) );
  XOR U41687 ( .A(n40603), .B(n40602), .Z(n40581) );
  NANDN U41688 ( .A(n40558), .B(n40557), .Z(n40562) );
  NANDN U41689 ( .A(n40560), .B(n40559), .Z(n40561) );
  AND U41690 ( .A(n40562), .B(n40561), .Z(n40580) );
  XNOR U41691 ( .A(n40581), .B(n40580), .Z(n40582) );
  NANDN U41692 ( .A(n40564), .B(n40563), .Z(n40568) );
  NAND U41693 ( .A(n40566), .B(n40565), .Z(n40567) );
  NAND U41694 ( .A(n40568), .B(n40567), .Z(n40583) );
  XNOR U41695 ( .A(n40582), .B(n40583), .Z(n40574) );
  XNOR U41696 ( .A(n40575), .B(n40574), .Z(n40576) );
  XNOR U41697 ( .A(n40577), .B(n40576), .Z(n40606) );
  XNOR U41698 ( .A(sreg[2002]), .B(n40606), .Z(n40608) );
  NANDN U41699 ( .A(sreg[2001]), .B(n40569), .Z(n40573) );
  NAND U41700 ( .A(n40571), .B(n40570), .Z(n40572) );
  NAND U41701 ( .A(n40573), .B(n40572), .Z(n40607) );
  XNOR U41702 ( .A(n40608), .B(n40607), .Z(c[2002]) );
  NANDN U41703 ( .A(n40575), .B(n40574), .Z(n40579) );
  NANDN U41704 ( .A(n40577), .B(n40576), .Z(n40578) );
  AND U41705 ( .A(n40579), .B(n40578), .Z(n40614) );
  NANDN U41706 ( .A(n40581), .B(n40580), .Z(n40585) );
  NANDN U41707 ( .A(n40583), .B(n40582), .Z(n40584) );
  AND U41708 ( .A(n40585), .B(n40584), .Z(n40612) );
  NAND U41709 ( .A(n42143), .B(n40586), .Z(n40588) );
  XNOR U41710 ( .A(a[981]), .B(n4212), .Z(n40623) );
  NAND U41711 ( .A(n42144), .B(n40623), .Z(n40587) );
  AND U41712 ( .A(n40588), .B(n40587), .Z(n40638) );
  XOR U41713 ( .A(a[985]), .B(n42012), .Z(n40626) );
  XNOR U41714 ( .A(n40638), .B(n40637), .Z(n40640) );
  AND U41715 ( .A(a[987]), .B(b[0]), .Z(n40590) );
  XNOR U41716 ( .A(n40590), .B(n4071), .Z(n40592) );
  NANDN U41717 ( .A(b[0]), .B(a[986]), .Z(n40591) );
  NAND U41718 ( .A(n40592), .B(n40591), .Z(n40634) );
  XOR U41719 ( .A(a[983]), .B(n42085), .Z(n40630) );
  AND U41720 ( .A(a[979]), .B(b[7]), .Z(n40631) );
  XNOR U41721 ( .A(n40632), .B(n40631), .Z(n40633) );
  XNOR U41722 ( .A(n40634), .B(n40633), .Z(n40639) );
  XOR U41723 ( .A(n40640), .B(n40639), .Z(n40618) );
  NANDN U41724 ( .A(n40595), .B(n40594), .Z(n40599) );
  NANDN U41725 ( .A(n40597), .B(n40596), .Z(n40598) );
  AND U41726 ( .A(n40599), .B(n40598), .Z(n40617) );
  XNOR U41727 ( .A(n40618), .B(n40617), .Z(n40619) );
  NANDN U41728 ( .A(n40601), .B(n40600), .Z(n40605) );
  NAND U41729 ( .A(n40603), .B(n40602), .Z(n40604) );
  NAND U41730 ( .A(n40605), .B(n40604), .Z(n40620) );
  XNOR U41731 ( .A(n40619), .B(n40620), .Z(n40611) );
  XNOR U41732 ( .A(n40612), .B(n40611), .Z(n40613) );
  XNOR U41733 ( .A(n40614), .B(n40613), .Z(n40643) );
  XNOR U41734 ( .A(sreg[2003]), .B(n40643), .Z(n40645) );
  NANDN U41735 ( .A(sreg[2002]), .B(n40606), .Z(n40610) );
  NAND U41736 ( .A(n40608), .B(n40607), .Z(n40609) );
  NAND U41737 ( .A(n40610), .B(n40609), .Z(n40644) );
  XNOR U41738 ( .A(n40645), .B(n40644), .Z(c[2003]) );
  NANDN U41739 ( .A(n40612), .B(n40611), .Z(n40616) );
  NANDN U41740 ( .A(n40614), .B(n40613), .Z(n40615) );
  AND U41741 ( .A(n40616), .B(n40615), .Z(n40651) );
  NANDN U41742 ( .A(n40618), .B(n40617), .Z(n40622) );
  NANDN U41743 ( .A(n40620), .B(n40619), .Z(n40621) );
  AND U41744 ( .A(n40622), .B(n40621), .Z(n40649) );
  NAND U41745 ( .A(n42143), .B(n40623), .Z(n40625) );
  XNOR U41746 ( .A(a[982]), .B(n4212), .Z(n40660) );
  NAND U41747 ( .A(n42144), .B(n40660), .Z(n40624) );
  AND U41748 ( .A(n40625), .B(n40624), .Z(n40675) );
  XOR U41749 ( .A(a[986]), .B(n42012), .Z(n40663) );
  XNOR U41750 ( .A(n40675), .B(n40674), .Z(n40677) );
  AND U41751 ( .A(a[988]), .B(b[0]), .Z(n40627) );
  XNOR U41752 ( .A(n40627), .B(n4071), .Z(n40629) );
  NANDN U41753 ( .A(b[0]), .B(a[987]), .Z(n40628) );
  NAND U41754 ( .A(n40629), .B(n40628), .Z(n40671) );
  XOR U41755 ( .A(a[984]), .B(n42085), .Z(n40664) );
  AND U41756 ( .A(a[980]), .B(b[7]), .Z(n40668) );
  XNOR U41757 ( .A(n40669), .B(n40668), .Z(n40670) );
  XNOR U41758 ( .A(n40671), .B(n40670), .Z(n40676) );
  XOR U41759 ( .A(n40677), .B(n40676), .Z(n40655) );
  NANDN U41760 ( .A(n40632), .B(n40631), .Z(n40636) );
  NANDN U41761 ( .A(n40634), .B(n40633), .Z(n40635) );
  AND U41762 ( .A(n40636), .B(n40635), .Z(n40654) );
  XNOR U41763 ( .A(n40655), .B(n40654), .Z(n40656) );
  NANDN U41764 ( .A(n40638), .B(n40637), .Z(n40642) );
  NAND U41765 ( .A(n40640), .B(n40639), .Z(n40641) );
  NAND U41766 ( .A(n40642), .B(n40641), .Z(n40657) );
  XNOR U41767 ( .A(n40656), .B(n40657), .Z(n40648) );
  XNOR U41768 ( .A(n40649), .B(n40648), .Z(n40650) );
  XNOR U41769 ( .A(n40651), .B(n40650), .Z(n40680) );
  XNOR U41770 ( .A(sreg[2004]), .B(n40680), .Z(n40682) );
  NANDN U41771 ( .A(sreg[2003]), .B(n40643), .Z(n40647) );
  NAND U41772 ( .A(n40645), .B(n40644), .Z(n40646) );
  NAND U41773 ( .A(n40647), .B(n40646), .Z(n40681) );
  XNOR U41774 ( .A(n40682), .B(n40681), .Z(c[2004]) );
  NANDN U41775 ( .A(n40649), .B(n40648), .Z(n40653) );
  NANDN U41776 ( .A(n40651), .B(n40650), .Z(n40652) );
  AND U41777 ( .A(n40653), .B(n40652), .Z(n40688) );
  NANDN U41778 ( .A(n40655), .B(n40654), .Z(n40659) );
  NANDN U41779 ( .A(n40657), .B(n40656), .Z(n40658) );
  AND U41780 ( .A(n40659), .B(n40658), .Z(n40686) );
  NAND U41781 ( .A(n42143), .B(n40660), .Z(n40662) );
  XNOR U41782 ( .A(a[983]), .B(n4212), .Z(n40697) );
  NAND U41783 ( .A(n42144), .B(n40697), .Z(n40661) );
  AND U41784 ( .A(n40662), .B(n40661), .Z(n40712) );
  XOR U41785 ( .A(a[987]), .B(n42012), .Z(n40700) );
  XNOR U41786 ( .A(n40712), .B(n40711), .Z(n40714) );
  XOR U41787 ( .A(a[985]), .B(n42085), .Z(n40704) );
  AND U41788 ( .A(a[981]), .B(b[7]), .Z(n40705) );
  XNOR U41789 ( .A(n40706), .B(n40705), .Z(n40707) );
  AND U41790 ( .A(a[989]), .B(b[0]), .Z(n40665) );
  XNOR U41791 ( .A(n40665), .B(n4071), .Z(n40667) );
  NANDN U41792 ( .A(b[0]), .B(a[988]), .Z(n40666) );
  NAND U41793 ( .A(n40667), .B(n40666), .Z(n40708) );
  XNOR U41794 ( .A(n40707), .B(n40708), .Z(n40713) );
  XOR U41795 ( .A(n40714), .B(n40713), .Z(n40692) );
  NANDN U41796 ( .A(n40669), .B(n40668), .Z(n40673) );
  NANDN U41797 ( .A(n40671), .B(n40670), .Z(n40672) );
  AND U41798 ( .A(n40673), .B(n40672), .Z(n40691) );
  XNOR U41799 ( .A(n40692), .B(n40691), .Z(n40693) );
  NANDN U41800 ( .A(n40675), .B(n40674), .Z(n40679) );
  NAND U41801 ( .A(n40677), .B(n40676), .Z(n40678) );
  NAND U41802 ( .A(n40679), .B(n40678), .Z(n40694) );
  XNOR U41803 ( .A(n40693), .B(n40694), .Z(n40685) );
  XNOR U41804 ( .A(n40686), .B(n40685), .Z(n40687) );
  XNOR U41805 ( .A(n40688), .B(n40687), .Z(n40717) );
  XNOR U41806 ( .A(sreg[2005]), .B(n40717), .Z(n40719) );
  NANDN U41807 ( .A(sreg[2004]), .B(n40680), .Z(n40684) );
  NAND U41808 ( .A(n40682), .B(n40681), .Z(n40683) );
  NAND U41809 ( .A(n40684), .B(n40683), .Z(n40718) );
  XNOR U41810 ( .A(n40719), .B(n40718), .Z(c[2005]) );
  NANDN U41811 ( .A(n40686), .B(n40685), .Z(n40690) );
  NANDN U41812 ( .A(n40688), .B(n40687), .Z(n40689) );
  AND U41813 ( .A(n40690), .B(n40689), .Z(n40725) );
  NANDN U41814 ( .A(n40692), .B(n40691), .Z(n40696) );
  NANDN U41815 ( .A(n40694), .B(n40693), .Z(n40695) );
  AND U41816 ( .A(n40696), .B(n40695), .Z(n40723) );
  NAND U41817 ( .A(n42143), .B(n40697), .Z(n40699) );
  XNOR U41818 ( .A(a[984]), .B(n4212), .Z(n40734) );
  NAND U41819 ( .A(n42144), .B(n40734), .Z(n40698) );
  AND U41820 ( .A(n40699), .B(n40698), .Z(n40749) );
  XOR U41821 ( .A(a[988]), .B(n42012), .Z(n40737) );
  XNOR U41822 ( .A(n40749), .B(n40748), .Z(n40751) );
  AND U41823 ( .A(a[990]), .B(b[0]), .Z(n40701) );
  XNOR U41824 ( .A(n40701), .B(n4071), .Z(n40703) );
  NANDN U41825 ( .A(b[0]), .B(a[989]), .Z(n40702) );
  NAND U41826 ( .A(n40703), .B(n40702), .Z(n40745) );
  XOR U41827 ( .A(a[986]), .B(n42085), .Z(n40738) );
  AND U41828 ( .A(a[982]), .B(b[7]), .Z(n40742) );
  XNOR U41829 ( .A(n40743), .B(n40742), .Z(n40744) );
  XNOR U41830 ( .A(n40745), .B(n40744), .Z(n40750) );
  XOR U41831 ( .A(n40751), .B(n40750), .Z(n40729) );
  NANDN U41832 ( .A(n40706), .B(n40705), .Z(n40710) );
  NANDN U41833 ( .A(n40708), .B(n40707), .Z(n40709) );
  AND U41834 ( .A(n40710), .B(n40709), .Z(n40728) );
  XNOR U41835 ( .A(n40729), .B(n40728), .Z(n40730) );
  NANDN U41836 ( .A(n40712), .B(n40711), .Z(n40716) );
  NAND U41837 ( .A(n40714), .B(n40713), .Z(n40715) );
  NAND U41838 ( .A(n40716), .B(n40715), .Z(n40731) );
  XNOR U41839 ( .A(n40730), .B(n40731), .Z(n40722) );
  XNOR U41840 ( .A(n40723), .B(n40722), .Z(n40724) );
  XNOR U41841 ( .A(n40725), .B(n40724), .Z(n40754) );
  XNOR U41842 ( .A(sreg[2006]), .B(n40754), .Z(n40756) );
  NANDN U41843 ( .A(sreg[2005]), .B(n40717), .Z(n40721) );
  NAND U41844 ( .A(n40719), .B(n40718), .Z(n40720) );
  NAND U41845 ( .A(n40721), .B(n40720), .Z(n40755) );
  XNOR U41846 ( .A(n40756), .B(n40755), .Z(c[2006]) );
  NANDN U41847 ( .A(n40723), .B(n40722), .Z(n40727) );
  NANDN U41848 ( .A(n40725), .B(n40724), .Z(n40726) );
  AND U41849 ( .A(n40727), .B(n40726), .Z(n40762) );
  NANDN U41850 ( .A(n40729), .B(n40728), .Z(n40733) );
  NANDN U41851 ( .A(n40731), .B(n40730), .Z(n40732) );
  AND U41852 ( .A(n40733), .B(n40732), .Z(n40760) );
  NAND U41853 ( .A(n42143), .B(n40734), .Z(n40736) );
  XNOR U41854 ( .A(a[985]), .B(n4212), .Z(n40771) );
  NAND U41855 ( .A(n42144), .B(n40771), .Z(n40735) );
  AND U41856 ( .A(n40736), .B(n40735), .Z(n40786) );
  XOR U41857 ( .A(a[989]), .B(n42012), .Z(n40774) );
  XNOR U41858 ( .A(n40786), .B(n40785), .Z(n40788) );
  XOR U41859 ( .A(a[987]), .B(n42085), .Z(n40775) );
  AND U41860 ( .A(a[983]), .B(b[7]), .Z(n40779) );
  XNOR U41861 ( .A(n40780), .B(n40779), .Z(n40781) );
  AND U41862 ( .A(a[991]), .B(b[0]), .Z(n40739) );
  XNOR U41863 ( .A(n40739), .B(n4071), .Z(n40741) );
  NANDN U41864 ( .A(b[0]), .B(a[990]), .Z(n40740) );
  NAND U41865 ( .A(n40741), .B(n40740), .Z(n40782) );
  XNOR U41866 ( .A(n40781), .B(n40782), .Z(n40787) );
  XOR U41867 ( .A(n40788), .B(n40787), .Z(n40766) );
  NANDN U41868 ( .A(n40743), .B(n40742), .Z(n40747) );
  NANDN U41869 ( .A(n40745), .B(n40744), .Z(n40746) );
  AND U41870 ( .A(n40747), .B(n40746), .Z(n40765) );
  XNOR U41871 ( .A(n40766), .B(n40765), .Z(n40767) );
  NANDN U41872 ( .A(n40749), .B(n40748), .Z(n40753) );
  NAND U41873 ( .A(n40751), .B(n40750), .Z(n40752) );
  NAND U41874 ( .A(n40753), .B(n40752), .Z(n40768) );
  XNOR U41875 ( .A(n40767), .B(n40768), .Z(n40759) );
  XNOR U41876 ( .A(n40760), .B(n40759), .Z(n40761) );
  XNOR U41877 ( .A(n40762), .B(n40761), .Z(n40791) );
  XNOR U41878 ( .A(sreg[2007]), .B(n40791), .Z(n40793) );
  NANDN U41879 ( .A(sreg[2006]), .B(n40754), .Z(n40758) );
  NAND U41880 ( .A(n40756), .B(n40755), .Z(n40757) );
  NAND U41881 ( .A(n40758), .B(n40757), .Z(n40792) );
  XNOR U41882 ( .A(n40793), .B(n40792), .Z(c[2007]) );
  NANDN U41883 ( .A(n40760), .B(n40759), .Z(n40764) );
  NANDN U41884 ( .A(n40762), .B(n40761), .Z(n40763) );
  AND U41885 ( .A(n40764), .B(n40763), .Z(n40799) );
  NANDN U41886 ( .A(n40766), .B(n40765), .Z(n40770) );
  NANDN U41887 ( .A(n40768), .B(n40767), .Z(n40769) );
  AND U41888 ( .A(n40770), .B(n40769), .Z(n40797) );
  NAND U41889 ( .A(n42143), .B(n40771), .Z(n40773) );
  XNOR U41890 ( .A(a[986]), .B(n4212), .Z(n40808) );
  NAND U41891 ( .A(n42144), .B(n40808), .Z(n40772) );
  AND U41892 ( .A(n40773), .B(n40772), .Z(n40823) );
  XOR U41893 ( .A(a[990]), .B(n42012), .Z(n40811) );
  XNOR U41894 ( .A(n40823), .B(n40822), .Z(n40825) );
  XOR U41895 ( .A(a[988]), .B(n42085), .Z(n40815) );
  AND U41896 ( .A(a[984]), .B(b[7]), .Z(n40816) );
  XNOR U41897 ( .A(n40817), .B(n40816), .Z(n40818) );
  AND U41898 ( .A(a[992]), .B(b[0]), .Z(n40776) );
  XNOR U41899 ( .A(n40776), .B(n4071), .Z(n40778) );
  NANDN U41900 ( .A(b[0]), .B(a[991]), .Z(n40777) );
  NAND U41901 ( .A(n40778), .B(n40777), .Z(n40819) );
  XNOR U41902 ( .A(n40818), .B(n40819), .Z(n40824) );
  XOR U41903 ( .A(n40825), .B(n40824), .Z(n40803) );
  NANDN U41904 ( .A(n40780), .B(n40779), .Z(n40784) );
  NANDN U41905 ( .A(n40782), .B(n40781), .Z(n40783) );
  AND U41906 ( .A(n40784), .B(n40783), .Z(n40802) );
  XNOR U41907 ( .A(n40803), .B(n40802), .Z(n40804) );
  NANDN U41908 ( .A(n40786), .B(n40785), .Z(n40790) );
  NAND U41909 ( .A(n40788), .B(n40787), .Z(n40789) );
  NAND U41910 ( .A(n40790), .B(n40789), .Z(n40805) );
  XNOR U41911 ( .A(n40804), .B(n40805), .Z(n40796) );
  XNOR U41912 ( .A(n40797), .B(n40796), .Z(n40798) );
  XNOR U41913 ( .A(n40799), .B(n40798), .Z(n40828) );
  XNOR U41914 ( .A(sreg[2008]), .B(n40828), .Z(n40830) );
  NANDN U41915 ( .A(sreg[2007]), .B(n40791), .Z(n40795) );
  NAND U41916 ( .A(n40793), .B(n40792), .Z(n40794) );
  NAND U41917 ( .A(n40795), .B(n40794), .Z(n40829) );
  XNOR U41918 ( .A(n40830), .B(n40829), .Z(c[2008]) );
  NANDN U41919 ( .A(n40797), .B(n40796), .Z(n40801) );
  NANDN U41920 ( .A(n40799), .B(n40798), .Z(n40800) );
  AND U41921 ( .A(n40801), .B(n40800), .Z(n40836) );
  NANDN U41922 ( .A(n40803), .B(n40802), .Z(n40807) );
  NANDN U41923 ( .A(n40805), .B(n40804), .Z(n40806) );
  AND U41924 ( .A(n40807), .B(n40806), .Z(n40834) );
  NAND U41925 ( .A(n42143), .B(n40808), .Z(n40810) );
  XNOR U41926 ( .A(a[987]), .B(n4212), .Z(n40845) );
  NAND U41927 ( .A(n42144), .B(n40845), .Z(n40809) );
  AND U41928 ( .A(n40810), .B(n40809), .Z(n40860) );
  XOR U41929 ( .A(a[991]), .B(n42012), .Z(n40848) );
  XNOR U41930 ( .A(n40860), .B(n40859), .Z(n40862) );
  AND U41931 ( .A(a[993]), .B(b[0]), .Z(n40812) );
  XNOR U41932 ( .A(n40812), .B(n4071), .Z(n40814) );
  NANDN U41933 ( .A(b[0]), .B(a[992]), .Z(n40813) );
  NAND U41934 ( .A(n40814), .B(n40813), .Z(n40856) );
  XOR U41935 ( .A(a[989]), .B(n42085), .Z(n40849) );
  AND U41936 ( .A(a[985]), .B(b[7]), .Z(n40853) );
  XNOR U41937 ( .A(n40854), .B(n40853), .Z(n40855) );
  XNOR U41938 ( .A(n40856), .B(n40855), .Z(n40861) );
  XOR U41939 ( .A(n40862), .B(n40861), .Z(n40840) );
  NANDN U41940 ( .A(n40817), .B(n40816), .Z(n40821) );
  NANDN U41941 ( .A(n40819), .B(n40818), .Z(n40820) );
  AND U41942 ( .A(n40821), .B(n40820), .Z(n40839) );
  XNOR U41943 ( .A(n40840), .B(n40839), .Z(n40841) );
  NANDN U41944 ( .A(n40823), .B(n40822), .Z(n40827) );
  NAND U41945 ( .A(n40825), .B(n40824), .Z(n40826) );
  NAND U41946 ( .A(n40827), .B(n40826), .Z(n40842) );
  XNOR U41947 ( .A(n40841), .B(n40842), .Z(n40833) );
  XNOR U41948 ( .A(n40834), .B(n40833), .Z(n40835) );
  XNOR U41949 ( .A(n40836), .B(n40835), .Z(n40865) );
  XNOR U41950 ( .A(sreg[2009]), .B(n40865), .Z(n40867) );
  NANDN U41951 ( .A(sreg[2008]), .B(n40828), .Z(n40832) );
  NAND U41952 ( .A(n40830), .B(n40829), .Z(n40831) );
  NAND U41953 ( .A(n40832), .B(n40831), .Z(n40866) );
  XNOR U41954 ( .A(n40867), .B(n40866), .Z(c[2009]) );
  NANDN U41955 ( .A(n40834), .B(n40833), .Z(n40838) );
  NANDN U41956 ( .A(n40836), .B(n40835), .Z(n40837) );
  AND U41957 ( .A(n40838), .B(n40837), .Z(n40873) );
  NANDN U41958 ( .A(n40840), .B(n40839), .Z(n40844) );
  NANDN U41959 ( .A(n40842), .B(n40841), .Z(n40843) );
  AND U41960 ( .A(n40844), .B(n40843), .Z(n40871) );
  NAND U41961 ( .A(n42143), .B(n40845), .Z(n40847) );
  XNOR U41962 ( .A(a[988]), .B(n4213), .Z(n40882) );
  NAND U41963 ( .A(n42144), .B(n40882), .Z(n40846) );
  AND U41964 ( .A(n40847), .B(n40846), .Z(n40897) );
  XOR U41965 ( .A(a[992]), .B(n42012), .Z(n40885) );
  XNOR U41966 ( .A(n40897), .B(n40896), .Z(n40899) );
  XOR U41967 ( .A(a[990]), .B(n42085), .Z(n40886) );
  AND U41968 ( .A(a[986]), .B(b[7]), .Z(n40890) );
  XNOR U41969 ( .A(n40891), .B(n40890), .Z(n40892) );
  AND U41970 ( .A(a[994]), .B(b[0]), .Z(n40850) );
  XNOR U41971 ( .A(n40850), .B(n4071), .Z(n40852) );
  NANDN U41972 ( .A(b[0]), .B(a[993]), .Z(n40851) );
  NAND U41973 ( .A(n40852), .B(n40851), .Z(n40893) );
  XNOR U41974 ( .A(n40892), .B(n40893), .Z(n40898) );
  XOR U41975 ( .A(n40899), .B(n40898), .Z(n40877) );
  NANDN U41976 ( .A(n40854), .B(n40853), .Z(n40858) );
  NANDN U41977 ( .A(n40856), .B(n40855), .Z(n40857) );
  AND U41978 ( .A(n40858), .B(n40857), .Z(n40876) );
  XNOR U41979 ( .A(n40877), .B(n40876), .Z(n40878) );
  NANDN U41980 ( .A(n40860), .B(n40859), .Z(n40864) );
  NAND U41981 ( .A(n40862), .B(n40861), .Z(n40863) );
  NAND U41982 ( .A(n40864), .B(n40863), .Z(n40879) );
  XNOR U41983 ( .A(n40878), .B(n40879), .Z(n40870) );
  XNOR U41984 ( .A(n40871), .B(n40870), .Z(n40872) );
  XNOR U41985 ( .A(n40873), .B(n40872), .Z(n40902) );
  XNOR U41986 ( .A(sreg[2010]), .B(n40902), .Z(n40904) );
  NANDN U41987 ( .A(sreg[2009]), .B(n40865), .Z(n40869) );
  NAND U41988 ( .A(n40867), .B(n40866), .Z(n40868) );
  NAND U41989 ( .A(n40869), .B(n40868), .Z(n40903) );
  XNOR U41990 ( .A(n40904), .B(n40903), .Z(c[2010]) );
  NANDN U41991 ( .A(n40871), .B(n40870), .Z(n40875) );
  NANDN U41992 ( .A(n40873), .B(n40872), .Z(n40874) );
  AND U41993 ( .A(n40875), .B(n40874), .Z(n40910) );
  NANDN U41994 ( .A(n40877), .B(n40876), .Z(n40881) );
  NANDN U41995 ( .A(n40879), .B(n40878), .Z(n40880) );
  AND U41996 ( .A(n40881), .B(n40880), .Z(n40908) );
  NAND U41997 ( .A(n42143), .B(n40882), .Z(n40884) );
  XNOR U41998 ( .A(a[989]), .B(n4213), .Z(n40919) );
  NAND U41999 ( .A(n42144), .B(n40919), .Z(n40883) );
  AND U42000 ( .A(n40884), .B(n40883), .Z(n40934) );
  XOR U42001 ( .A(a[993]), .B(n42012), .Z(n40922) );
  XNOR U42002 ( .A(n40934), .B(n40933), .Z(n40936) );
  XOR U42003 ( .A(a[991]), .B(n42085), .Z(n40926) );
  AND U42004 ( .A(a[987]), .B(b[7]), .Z(n40927) );
  XNOR U42005 ( .A(n40928), .B(n40927), .Z(n40929) );
  AND U42006 ( .A(a[995]), .B(b[0]), .Z(n40887) );
  XNOR U42007 ( .A(n40887), .B(n4071), .Z(n40889) );
  NANDN U42008 ( .A(b[0]), .B(a[994]), .Z(n40888) );
  NAND U42009 ( .A(n40889), .B(n40888), .Z(n40930) );
  XNOR U42010 ( .A(n40929), .B(n40930), .Z(n40935) );
  XOR U42011 ( .A(n40936), .B(n40935), .Z(n40914) );
  NANDN U42012 ( .A(n40891), .B(n40890), .Z(n40895) );
  NANDN U42013 ( .A(n40893), .B(n40892), .Z(n40894) );
  AND U42014 ( .A(n40895), .B(n40894), .Z(n40913) );
  XNOR U42015 ( .A(n40914), .B(n40913), .Z(n40915) );
  NANDN U42016 ( .A(n40897), .B(n40896), .Z(n40901) );
  NAND U42017 ( .A(n40899), .B(n40898), .Z(n40900) );
  NAND U42018 ( .A(n40901), .B(n40900), .Z(n40916) );
  XNOR U42019 ( .A(n40915), .B(n40916), .Z(n40907) );
  XNOR U42020 ( .A(n40908), .B(n40907), .Z(n40909) );
  XNOR U42021 ( .A(n40910), .B(n40909), .Z(n40939) );
  XNOR U42022 ( .A(sreg[2011]), .B(n40939), .Z(n40941) );
  NANDN U42023 ( .A(sreg[2010]), .B(n40902), .Z(n40906) );
  NAND U42024 ( .A(n40904), .B(n40903), .Z(n40905) );
  NAND U42025 ( .A(n40906), .B(n40905), .Z(n40940) );
  XNOR U42026 ( .A(n40941), .B(n40940), .Z(c[2011]) );
  NANDN U42027 ( .A(n40908), .B(n40907), .Z(n40912) );
  NANDN U42028 ( .A(n40910), .B(n40909), .Z(n40911) );
  AND U42029 ( .A(n40912), .B(n40911), .Z(n40947) );
  NANDN U42030 ( .A(n40914), .B(n40913), .Z(n40918) );
  NANDN U42031 ( .A(n40916), .B(n40915), .Z(n40917) );
  AND U42032 ( .A(n40918), .B(n40917), .Z(n40945) );
  NAND U42033 ( .A(n42143), .B(n40919), .Z(n40921) );
  XNOR U42034 ( .A(a[990]), .B(n4213), .Z(n40956) );
  NAND U42035 ( .A(n42144), .B(n40956), .Z(n40920) );
  AND U42036 ( .A(n40921), .B(n40920), .Z(n40971) );
  XOR U42037 ( .A(a[994]), .B(n42012), .Z(n40959) );
  XNOR U42038 ( .A(n40971), .B(n40970), .Z(n40973) );
  AND U42039 ( .A(a[996]), .B(b[0]), .Z(n40923) );
  XNOR U42040 ( .A(n40923), .B(n4071), .Z(n40925) );
  NANDN U42041 ( .A(b[0]), .B(a[995]), .Z(n40924) );
  NAND U42042 ( .A(n40925), .B(n40924), .Z(n40967) );
  XOR U42043 ( .A(a[992]), .B(n42085), .Z(n40960) );
  AND U42044 ( .A(a[988]), .B(b[7]), .Z(n40964) );
  XNOR U42045 ( .A(n40965), .B(n40964), .Z(n40966) );
  XNOR U42046 ( .A(n40967), .B(n40966), .Z(n40972) );
  XOR U42047 ( .A(n40973), .B(n40972), .Z(n40951) );
  NANDN U42048 ( .A(n40928), .B(n40927), .Z(n40932) );
  NANDN U42049 ( .A(n40930), .B(n40929), .Z(n40931) );
  AND U42050 ( .A(n40932), .B(n40931), .Z(n40950) );
  XNOR U42051 ( .A(n40951), .B(n40950), .Z(n40952) );
  NANDN U42052 ( .A(n40934), .B(n40933), .Z(n40938) );
  NAND U42053 ( .A(n40936), .B(n40935), .Z(n40937) );
  NAND U42054 ( .A(n40938), .B(n40937), .Z(n40953) );
  XNOR U42055 ( .A(n40952), .B(n40953), .Z(n40944) );
  XNOR U42056 ( .A(n40945), .B(n40944), .Z(n40946) );
  XNOR U42057 ( .A(n40947), .B(n40946), .Z(n40976) );
  XNOR U42058 ( .A(sreg[2012]), .B(n40976), .Z(n40978) );
  NANDN U42059 ( .A(sreg[2011]), .B(n40939), .Z(n40943) );
  NAND U42060 ( .A(n40941), .B(n40940), .Z(n40942) );
  NAND U42061 ( .A(n40943), .B(n40942), .Z(n40977) );
  XNOR U42062 ( .A(n40978), .B(n40977), .Z(c[2012]) );
  NANDN U42063 ( .A(n40945), .B(n40944), .Z(n40949) );
  NANDN U42064 ( .A(n40947), .B(n40946), .Z(n40948) );
  AND U42065 ( .A(n40949), .B(n40948), .Z(n40984) );
  NANDN U42066 ( .A(n40951), .B(n40950), .Z(n40955) );
  NANDN U42067 ( .A(n40953), .B(n40952), .Z(n40954) );
  AND U42068 ( .A(n40955), .B(n40954), .Z(n40982) );
  NAND U42069 ( .A(n42143), .B(n40956), .Z(n40958) );
  XNOR U42070 ( .A(a[991]), .B(n4213), .Z(n40993) );
  NAND U42071 ( .A(n42144), .B(n40993), .Z(n40957) );
  AND U42072 ( .A(n40958), .B(n40957), .Z(n41008) );
  XOR U42073 ( .A(a[995]), .B(n42012), .Z(n40996) );
  XNOR U42074 ( .A(n41008), .B(n41007), .Z(n41010) );
  XOR U42075 ( .A(a[993]), .B(n42085), .Z(n41000) );
  AND U42076 ( .A(a[989]), .B(b[7]), .Z(n41001) );
  XNOR U42077 ( .A(n41002), .B(n41001), .Z(n41003) );
  AND U42078 ( .A(a[997]), .B(b[0]), .Z(n40961) );
  XNOR U42079 ( .A(n40961), .B(n4071), .Z(n40963) );
  NANDN U42080 ( .A(b[0]), .B(a[996]), .Z(n40962) );
  NAND U42081 ( .A(n40963), .B(n40962), .Z(n41004) );
  XNOR U42082 ( .A(n41003), .B(n41004), .Z(n41009) );
  XOR U42083 ( .A(n41010), .B(n41009), .Z(n40988) );
  NANDN U42084 ( .A(n40965), .B(n40964), .Z(n40969) );
  NANDN U42085 ( .A(n40967), .B(n40966), .Z(n40968) );
  AND U42086 ( .A(n40969), .B(n40968), .Z(n40987) );
  XNOR U42087 ( .A(n40988), .B(n40987), .Z(n40989) );
  NANDN U42088 ( .A(n40971), .B(n40970), .Z(n40975) );
  NAND U42089 ( .A(n40973), .B(n40972), .Z(n40974) );
  NAND U42090 ( .A(n40975), .B(n40974), .Z(n40990) );
  XNOR U42091 ( .A(n40989), .B(n40990), .Z(n40981) );
  XNOR U42092 ( .A(n40982), .B(n40981), .Z(n40983) );
  XNOR U42093 ( .A(n40984), .B(n40983), .Z(n41013) );
  XNOR U42094 ( .A(sreg[2013]), .B(n41013), .Z(n41015) );
  NANDN U42095 ( .A(sreg[2012]), .B(n40976), .Z(n40980) );
  NAND U42096 ( .A(n40978), .B(n40977), .Z(n40979) );
  NAND U42097 ( .A(n40980), .B(n40979), .Z(n41014) );
  XNOR U42098 ( .A(n41015), .B(n41014), .Z(c[2013]) );
  NANDN U42099 ( .A(n40982), .B(n40981), .Z(n40986) );
  NANDN U42100 ( .A(n40984), .B(n40983), .Z(n40985) );
  AND U42101 ( .A(n40986), .B(n40985), .Z(n41021) );
  NANDN U42102 ( .A(n40988), .B(n40987), .Z(n40992) );
  NANDN U42103 ( .A(n40990), .B(n40989), .Z(n40991) );
  AND U42104 ( .A(n40992), .B(n40991), .Z(n41019) );
  NAND U42105 ( .A(n42143), .B(n40993), .Z(n40995) );
  XNOR U42106 ( .A(a[992]), .B(n4213), .Z(n41030) );
  NAND U42107 ( .A(n42144), .B(n41030), .Z(n40994) );
  AND U42108 ( .A(n40995), .B(n40994), .Z(n41045) );
  XOR U42109 ( .A(a[996]), .B(n42012), .Z(n41033) );
  XNOR U42110 ( .A(n41045), .B(n41044), .Z(n41047) );
  AND U42111 ( .A(a[998]), .B(b[0]), .Z(n40997) );
  XNOR U42112 ( .A(n40997), .B(n4071), .Z(n40999) );
  NANDN U42113 ( .A(b[0]), .B(a[997]), .Z(n40998) );
  NAND U42114 ( .A(n40999), .B(n40998), .Z(n41041) );
  XOR U42115 ( .A(a[994]), .B(n42085), .Z(n41034) );
  AND U42116 ( .A(a[990]), .B(b[7]), .Z(n41038) );
  XNOR U42117 ( .A(n41039), .B(n41038), .Z(n41040) );
  XNOR U42118 ( .A(n41041), .B(n41040), .Z(n41046) );
  XOR U42119 ( .A(n41047), .B(n41046), .Z(n41025) );
  NANDN U42120 ( .A(n41002), .B(n41001), .Z(n41006) );
  NANDN U42121 ( .A(n41004), .B(n41003), .Z(n41005) );
  AND U42122 ( .A(n41006), .B(n41005), .Z(n41024) );
  XNOR U42123 ( .A(n41025), .B(n41024), .Z(n41026) );
  NANDN U42124 ( .A(n41008), .B(n41007), .Z(n41012) );
  NAND U42125 ( .A(n41010), .B(n41009), .Z(n41011) );
  NAND U42126 ( .A(n41012), .B(n41011), .Z(n41027) );
  XNOR U42127 ( .A(n41026), .B(n41027), .Z(n41018) );
  XNOR U42128 ( .A(n41019), .B(n41018), .Z(n41020) );
  XNOR U42129 ( .A(n41021), .B(n41020), .Z(n41050) );
  XNOR U42130 ( .A(sreg[2014]), .B(n41050), .Z(n41052) );
  NANDN U42131 ( .A(sreg[2013]), .B(n41013), .Z(n41017) );
  NAND U42132 ( .A(n41015), .B(n41014), .Z(n41016) );
  NAND U42133 ( .A(n41017), .B(n41016), .Z(n41051) );
  XNOR U42134 ( .A(n41052), .B(n41051), .Z(c[2014]) );
  NANDN U42135 ( .A(n41019), .B(n41018), .Z(n41023) );
  NANDN U42136 ( .A(n41021), .B(n41020), .Z(n41022) );
  AND U42137 ( .A(n41023), .B(n41022), .Z(n41058) );
  NANDN U42138 ( .A(n41025), .B(n41024), .Z(n41029) );
  NANDN U42139 ( .A(n41027), .B(n41026), .Z(n41028) );
  AND U42140 ( .A(n41029), .B(n41028), .Z(n41056) );
  NAND U42141 ( .A(n42143), .B(n41030), .Z(n41032) );
  XNOR U42142 ( .A(a[993]), .B(n4213), .Z(n41067) );
  NAND U42143 ( .A(n42144), .B(n41067), .Z(n41031) );
  AND U42144 ( .A(n41032), .B(n41031), .Z(n41082) );
  XOR U42145 ( .A(a[997]), .B(n42012), .Z(n41070) );
  XNOR U42146 ( .A(n41082), .B(n41081), .Z(n41084) );
  XOR U42147 ( .A(a[995]), .B(n42085), .Z(n41071) );
  AND U42148 ( .A(a[991]), .B(b[7]), .Z(n41075) );
  XNOR U42149 ( .A(n41076), .B(n41075), .Z(n41077) );
  AND U42150 ( .A(a[999]), .B(b[0]), .Z(n41035) );
  XNOR U42151 ( .A(n41035), .B(n4071), .Z(n41037) );
  NANDN U42152 ( .A(b[0]), .B(a[998]), .Z(n41036) );
  NAND U42153 ( .A(n41037), .B(n41036), .Z(n41078) );
  XNOR U42154 ( .A(n41077), .B(n41078), .Z(n41083) );
  XOR U42155 ( .A(n41084), .B(n41083), .Z(n41062) );
  NANDN U42156 ( .A(n41039), .B(n41038), .Z(n41043) );
  NANDN U42157 ( .A(n41041), .B(n41040), .Z(n41042) );
  AND U42158 ( .A(n41043), .B(n41042), .Z(n41061) );
  XNOR U42159 ( .A(n41062), .B(n41061), .Z(n41063) );
  NANDN U42160 ( .A(n41045), .B(n41044), .Z(n41049) );
  NAND U42161 ( .A(n41047), .B(n41046), .Z(n41048) );
  NAND U42162 ( .A(n41049), .B(n41048), .Z(n41064) );
  XNOR U42163 ( .A(n41063), .B(n41064), .Z(n41055) );
  XNOR U42164 ( .A(n41056), .B(n41055), .Z(n41057) );
  XNOR U42165 ( .A(n41058), .B(n41057), .Z(n41087) );
  XNOR U42166 ( .A(sreg[2015]), .B(n41087), .Z(n41089) );
  NANDN U42167 ( .A(sreg[2014]), .B(n41050), .Z(n41054) );
  NAND U42168 ( .A(n41052), .B(n41051), .Z(n41053) );
  NAND U42169 ( .A(n41054), .B(n41053), .Z(n41088) );
  XNOR U42170 ( .A(n41089), .B(n41088), .Z(c[2015]) );
  NANDN U42171 ( .A(n41056), .B(n41055), .Z(n41060) );
  NANDN U42172 ( .A(n41058), .B(n41057), .Z(n41059) );
  AND U42173 ( .A(n41060), .B(n41059), .Z(n41095) );
  NANDN U42174 ( .A(n41062), .B(n41061), .Z(n41066) );
  NANDN U42175 ( .A(n41064), .B(n41063), .Z(n41065) );
  AND U42176 ( .A(n41066), .B(n41065), .Z(n41093) );
  NAND U42177 ( .A(n42143), .B(n41067), .Z(n41069) );
  XNOR U42178 ( .A(a[994]), .B(n4213), .Z(n41104) );
  NAND U42179 ( .A(n42144), .B(n41104), .Z(n41068) );
  AND U42180 ( .A(n41069), .B(n41068), .Z(n41119) );
  XOR U42181 ( .A(a[998]), .B(n42012), .Z(n41107) );
  XNOR U42182 ( .A(n41119), .B(n41118), .Z(n41121) );
  XOR U42183 ( .A(a[996]), .B(n42085), .Z(n41108) );
  AND U42184 ( .A(a[992]), .B(b[7]), .Z(n41112) );
  XNOR U42185 ( .A(n41113), .B(n41112), .Z(n41114) );
  AND U42186 ( .A(a[1000]), .B(b[0]), .Z(n41072) );
  XNOR U42187 ( .A(n41072), .B(n4071), .Z(n41074) );
  NANDN U42188 ( .A(b[0]), .B(a[999]), .Z(n41073) );
  NAND U42189 ( .A(n41074), .B(n41073), .Z(n41115) );
  XNOR U42190 ( .A(n41114), .B(n41115), .Z(n41120) );
  XOR U42191 ( .A(n41121), .B(n41120), .Z(n41099) );
  NANDN U42192 ( .A(n41076), .B(n41075), .Z(n41080) );
  NANDN U42193 ( .A(n41078), .B(n41077), .Z(n41079) );
  AND U42194 ( .A(n41080), .B(n41079), .Z(n41098) );
  XNOR U42195 ( .A(n41099), .B(n41098), .Z(n41100) );
  NANDN U42196 ( .A(n41082), .B(n41081), .Z(n41086) );
  NAND U42197 ( .A(n41084), .B(n41083), .Z(n41085) );
  NAND U42198 ( .A(n41086), .B(n41085), .Z(n41101) );
  XNOR U42199 ( .A(n41100), .B(n41101), .Z(n41092) );
  XNOR U42200 ( .A(n41093), .B(n41092), .Z(n41094) );
  XNOR U42201 ( .A(n41095), .B(n41094), .Z(n41124) );
  XNOR U42202 ( .A(sreg[2016]), .B(n41124), .Z(n41126) );
  NANDN U42203 ( .A(sreg[2015]), .B(n41087), .Z(n41091) );
  NAND U42204 ( .A(n41089), .B(n41088), .Z(n41090) );
  NAND U42205 ( .A(n41091), .B(n41090), .Z(n41125) );
  XNOR U42206 ( .A(n41126), .B(n41125), .Z(c[2016]) );
  NANDN U42207 ( .A(n41093), .B(n41092), .Z(n41097) );
  NANDN U42208 ( .A(n41095), .B(n41094), .Z(n41096) );
  AND U42209 ( .A(n41097), .B(n41096), .Z(n41132) );
  NANDN U42210 ( .A(n41099), .B(n41098), .Z(n41103) );
  NANDN U42211 ( .A(n41101), .B(n41100), .Z(n41102) );
  AND U42212 ( .A(n41103), .B(n41102), .Z(n41130) );
  NAND U42213 ( .A(n42143), .B(n41104), .Z(n41106) );
  XNOR U42214 ( .A(a[995]), .B(n4214), .Z(n41141) );
  NAND U42215 ( .A(n42144), .B(n41141), .Z(n41105) );
  AND U42216 ( .A(n41106), .B(n41105), .Z(n41156) );
  XOR U42217 ( .A(a[999]), .B(n42012), .Z(n41144) );
  XNOR U42218 ( .A(n41156), .B(n41155), .Z(n41158) );
  XOR U42219 ( .A(a[997]), .B(n42085), .Z(n41148) );
  AND U42220 ( .A(a[993]), .B(b[7]), .Z(n41149) );
  XNOR U42221 ( .A(n41150), .B(n41149), .Z(n41151) );
  AND U42222 ( .A(a[1001]), .B(b[0]), .Z(n41109) );
  XNOR U42223 ( .A(n41109), .B(n4071), .Z(n41111) );
  NANDN U42224 ( .A(b[0]), .B(a[1000]), .Z(n41110) );
  NAND U42225 ( .A(n41111), .B(n41110), .Z(n41152) );
  XNOR U42226 ( .A(n41151), .B(n41152), .Z(n41157) );
  XOR U42227 ( .A(n41158), .B(n41157), .Z(n41136) );
  NANDN U42228 ( .A(n41113), .B(n41112), .Z(n41117) );
  NANDN U42229 ( .A(n41115), .B(n41114), .Z(n41116) );
  AND U42230 ( .A(n41117), .B(n41116), .Z(n41135) );
  XNOR U42231 ( .A(n41136), .B(n41135), .Z(n41137) );
  NANDN U42232 ( .A(n41119), .B(n41118), .Z(n41123) );
  NAND U42233 ( .A(n41121), .B(n41120), .Z(n41122) );
  NAND U42234 ( .A(n41123), .B(n41122), .Z(n41138) );
  XNOR U42235 ( .A(n41137), .B(n41138), .Z(n41129) );
  XNOR U42236 ( .A(n41130), .B(n41129), .Z(n41131) );
  XNOR U42237 ( .A(n41132), .B(n41131), .Z(n41161) );
  XNOR U42238 ( .A(sreg[2017]), .B(n41161), .Z(n41163) );
  NANDN U42239 ( .A(sreg[2016]), .B(n41124), .Z(n41128) );
  NAND U42240 ( .A(n41126), .B(n41125), .Z(n41127) );
  NAND U42241 ( .A(n41128), .B(n41127), .Z(n41162) );
  XNOR U42242 ( .A(n41163), .B(n41162), .Z(c[2017]) );
  NANDN U42243 ( .A(n41130), .B(n41129), .Z(n41134) );
  NANDN U42244 ( .A(n41132), .B(n41131), .Z(n41133) );
  AND U42245 ( .A(n41134), .B(n41133), .Z(n41169) );
  NANDN U42246 ( .A(n41136), .B(n41135), .Z(n41140) );
  NANDN U42247 ( .A(n41138), .B(n41137), .Z(n41139) );
  AND U42248 ( .A(n41140), .B(n41139), .Z(n41167) );
  NAND U42249 ( .A(n42143), .B(n41141), .Z(n41143) );
  XNOR U42250 ( .A(a[996]), .B(n4214), .Z(n41178) );
  NAND U42251 ( .A(n42144), .B(n41178), .Z(n41142) );
  AND U42252 ( .A(n41143), .B(n41142), .Z(n41193) );
  XOR U42253 ( .A(a[1000]), .B(n42012), .Z(n41181) );
  XNOR U42254 ( .A(n41193), .B(n41192), .Z(n41195) );
  AND U42255 ( .A(a[1002]), .B(b[0]), .Z(n41145) );
  XNOR U42256 ( .A(n41145), .B(n4071), .Z(n41147) );
  NANDN U42257 ( .A(b[0]), .B(a[1001]), .Z(n41146) );
  NAND U42258 ( .A(n41147), .B(n41146), .Z(n41189) );
  XOR U42259 ( .A(a[998]), .B(n42085), .Z(n41185) );
  AND U42260 ( .A(a[994]), .B(b[7]), .Z(n41186) );
  XNOR U42261 ( .A(n41187), .B(n41186), .Z(n41188) );
  XNOR U42262 ( .A(n41189), .B(n41188), .Z(n41194) );
  XOR U42263 ( .A(n41195), .B(n41194), .Z(n41173) );
  NANDN U42264 ( .A(n41150), .B(n41149), .Z(n41154) );
  NANDN U42265 ( .A(n41152), .B(n41151), .Z(n41153) );
  AND U42266 ( .A(n41154), .B(n41153), .Z(n41172) );
  XNOR U42267 ( .A(n41173), .B(n41172), .Z(n41174) );
  NANDN U42268 ( .A(n41156), .B(n41155), .Z(n41160) );
  NAND U42269 ( .A(n41158), .B(n41157), .Z(n41159) );
  NAND U42270 ( .A(n41160), .B(n41159), .Z(n41175) );
  XNOR U42271 ( .A(n41174), .B(n41175), .Z(n41166) );
  XNOR U42272 ( .A(n41167), .B(n41166), .Z(n41168) );
  XNOR U42273 ( .A(n41169), .B(n41168), .Z(n41198) );
  XNOR U42274 ( .A(sreg[2018]), .B(n41198), .Z(n41200) );
  NANDN U42275 ( .A(sreg[2017]), .B(n41161), .Z(n41165) );
  NAND U42276 ( .A(n41163), .B(n41162), .Z(n41164) );
  NAND U42277 ( .A(n41165), .B(n41164), .Z(n41199) );
  XNOR U42278 ( .A(n41200), .B(n41199), .Z(c[2018]) );
  NANDN U42279 ( .A(n41167), .B(n41166), .Z(n41171) );
  NANDN U42280 ( .A(n41169), .B(n41168), .Z(n41170) );
  AND U42281 ( .A(n41171), .B(n41170), .Z(n41206) );
  NANDN U42282 ( .A(n41173), .B(n41172), .Z(n41177) );
  NANDN U42283 ( .A(n41175), .B(n41174), .Z(n41176) );
  AND U42284 ( .A(n41177), .B(n41176), .Z(n41204) );
  NAND U42285 ( .A(n42143), .B(n41178), .Z(n41180) );
  XNOR U42286 ( .A(a[997]), .B(n4214), .Z(n41215) );
  NAND U42287 ( .A(n42144), .B(n41215), .Z(n41179) );
  AND U42288 ( .A(n41180), .B(n41179), .Z(n41230) );
  XOR U42289 ( .A(a[1001]), .B(n42012), .Z(n41218) );
  XNOR U42290 ( .A(n41230), .B(n41229), .Z(n41232) );
  AND U42291 ( .A(a[1003]), .B(b[0]), .Z(n41182) );
  XNOR U42292 ( .A(n41182), .B(n4071), .Z(n41184) );
  NANDN U42293 ( .A(b[0]), .B(a[1002]), .Z(n41183) );
  NAND U42294 ( .A(n41184), .B(n41183), .Z(n41226) );
  XOR U42295 ( .A(a[999]), .B(n42085), .Z(n41219) );
  AND U42296 ( .A(a[995]), .B(b[7]), .Z(n41223) );
  XNOR U42297 ( .A(n41224), .B(n41223), .Z(n41225) );
  XNOR U42298 ( .A(n41226), .B(n41225), .Z(n41231) );
  XOR U42299 ( .A(n41232), .B(n41231), .Z(n41210) );
  NANDN U42300 ( .A(n41187), .B(n41186), .Z(n41191) );
  NANDN U42301 ( .A(n41189), .B(n41188), .Z(n41190) );
  AND U42302 ( .A(n41191), .B(n41190), .Z(n41209) );
  XNOR U42303 ( .A(n41210), .B(n41209), .Z(n41211) );
  NANDN U42304 ( .A(n41193), .B(n41192), .Z(n41197) );
  NAND U42305 ( .A(n41195), .B(n41194), .Z(n41196) );
  NAND U42306 ( .A(n41197), .B(n41196), .Z(n41212) );
  XNOR U42307 ( .A(n41211), .B(n41212), .Z(n41203) );
  XNOR U42308 ( .A(n41204), .B(n41203), .Z(n41205) );
  XNOR U42309 ( .A(n41206), .B(n41205), .Z(n41235) );
  XNOR U42310 ( .A(sreg[2019]), .B(n41235), .Z(n41237) );
  NANDN U42311 ( .A(sreg[2018]), .B(n41198), .Z(n41202) );
  NAND U42312 ( .A(n41200), .B(n41199), .Z(n41201) );
  NAND U42313 ( .A(n41202), .B(n41201), .Z(n41236) );
  XNOR U42314 ( .A(n41237), .B(n41236), .Z(c[2019]) );
  NANDN U42315 ( .A(n41204), .B(n41203), .Z(n41208) );
  NANDN U42316 ( .A(n41206), .B(n41205), .Z(n41207) );
  AND U42317 ( .A(n41208), .B(n41207), .Z(n41243) );
  NANDN U42318 ( .A(n41210), .B(n41209), .Z(n41214) );
  NANDN U42319 ( .A(n41212), .B(n41211), .Z(n41213) );
  AND U42320 ( .A(n41214), .B(n41213), .Z(n41241) );
  NAND U42321 ( .A(n42143), .B(n41215), .Z(n41217) );
  XNOR U42322 ( .A(a[998]), .B(n4214), .Z(n41252) );
  NAND U42323 ( .A(n42144), .B(n41252), .Z(n41216) );
  AND U42324 ( .A(n41217), .B(n41216), .Z(n41267) );
  XOR U42325 ( .A(a[1002]), .B(n42012), .Z(n41255) );
  XNOR U42326 ( .A(n41267), .B(n41266), .Z(n41269) );
  XOR U42327 ( .A(a[1000]), .B(n42085), .Z(n41259) );
  AND U42328 ( .A(a[996]), .B(b[7]), .Z(n41260) );
  XNOR U42329 ( .A(n41261), .B(n41260), .Z(n41262) );
  AND U42330 ( .A(a[1004]), .B(b[0]), .Z(n41220) );
  XNOR U42331 ( .A(n41220), .B(n4071), .Z(n41222) );
  NANDN U42332 ( .A(b[0]), .B(a[1003]), .Z(n41221) );
  NAND U42333 ( .A(n41222), .B(n41221), .Z(n41263) );
  XNOR U42334 ( .A(n41262), .B(n41263), .Z(n41268) );
  XOR U42335 ( .A(n41269), .B(n41268), .Z(n41247) );
  NANDN U42336 ( .A(n41224), .B(n41223), .Z(n41228) );
  NANDN U42337 ( .A(n41226), .B(n41225), .Z(n41227) );
  AND U42338 ( .A(n41228), .B(n41227), .Z(n41246) );
  XNOR U42339 ( .A(n41247), .B(n41246), .Z(n41248) );
  NANDN U42340 ( .A(n41230), .B(n41229), .Z(n41234) );
  NAND U42341 ( .A(n41232), .B(n41231), .Z(n41233) );
  NAND U42342 ( .A(n41234), .B(n41233), .Z(n41249) );
  XNOR U42343 ( .A(n41248), .B(n41249), .Z(n41240) );
  XNOR U42344 ( .A(n41241), .B(n41240), .Z(n41242) );
  XNOR U42345 ( .A(n41243), .B(n41242), .Z(n41272) );
  XNOR U42346 ( .A(sreg[2020]), .B(n41272), .Z(n41274) );
  NANDN U42347 ( .A(sreg[2019]), .B(n41235), .Z(n41239) );
  NAND U42348 ( .A(n41237), .B(n41236), .Z(n41238) );
  NAND U42349 ( .A(n41239), .B(n41238), .Z(n41273) );
  XNOR U42350 ( .A(n41274), .B(n41273), .Z(c[2020]) );
  NANDN U42351 ( .A(n41241), .B(n41240), .Z(n41245) );
  NANDN U42352 ( .A(n41243), .B(n41242), .Z(n41244) );
  AND U42353 ( .A(n41245), .B(n41244), .Z(n41280) );
  NANDN U42354 ( .A(n41247), .B(n41246), .Z(n41251) );
  NANDN U42355 ( .A(n41249), .B(n41248), .Z(n41250) );
  AND U42356 ( .A(n41251), .B(n41250), .Z(n41278) );
  NAND U42357 ( .A(n42143), .B(n41252), .Z(n41254) );
  XNOR U42358 ( .A(a[999]), .B(n4214), .Z(n41289) );
  NAND U42359 ( .A(n42144), .B(n41289), .Z(n41253) );
  AND U42360 ( .A(n41254), .B(n41253), .Z(n41304) );
  XOR U42361 ( .A(a[1003]), .B(n42012), .Z(n41292) );
  XNOR U42362 ( .A(n41304), .B(n41303), .Z(n41306) );
  AND U42363 ( .A(a[1005]), .B(b[0]), .Z(n41256) );
  XNOR U42364 ( .A(n41256), .B(n4071), .Z(n41258) );
  NANDN U42365 ( .A(b[0]), .B(a[1004]), .Z(n41257) );
  NAND U42366 ( .A(n41258), .B(n41257), .Z(n41300) );
  XOR U42367 ( .A(a[1001]), .B(n42085), .Z(n41293) );
  AND U42368 ( .A(a[997]), .B(b[7]), .Z(n41297) );
  XNOR U42369 ( .A(n41298), .B(n41297), .Z(n41299) );
  XNOR U42370 ( .A(n41300), .B(n41299), .Z(n41305) );
  XOR U42371 ( .A(n41306), .B(n41305), .Z(n41284) );
  NANDN U42372 ( .A(n41261), .B(n41260), .Z(n41265) );
  NANDN U42373 ( .A(n41263), .B(n41262), .Z(n41264) );
  AND U42374 ( .A(n41265), .B(n41264), .Z(n41283) );
  XNOR U42375 ( .A(n41284), .B(n41283), .Z(n41285) );
  NANDN U42376 ( .A(n41267), .B(n41266), .Z(n41271) );
  NAND U42377 ( .A(n41269), .B(n41268), .Z(n41270) );
  NAND U42378 ( .A(n41271), .B(n41270), .Z(n41286) );
  XNOR U42379 ( .A(n41285), .B(n41286), .Z(n41277) );
  XNOR U42380 ( .A(n41278), .B(n41277), .Z(n41279) );
  XNOR U42381 ( .A(n41280), .B(n41279), .Z(n41309) );
  XNOR U42382 ( .A(sreg[2021]), .B(n41309), .Z(n41311) );
  NANDN U42383 ( .A(sreg[2020]), .B(n41272), .Z(n41276) );
  NAND U42384 ( .A(n41274), .B(n41273), .Z(n41275) );
  NAND U42385 ( .A(n41276), .B(n41275), .Z(n41310) );
  XNOR U42386 ( .A(n41311), .B(n41310), .Z(c[2021]) );
  NANDN U42387 ( .A(n41278), .B(n41277), .Z(n41282) );
  NANDN U42388 ( .A(n41280), .B(n41279), .Z(n41281) );
  AND U42389 ( .A(n41282), .B(n41281), .Z(n41317) );
  NANDN U42390 ( .A(n41284), .B(n41283), .Z(n41288) );
  NANDN U42391 ( .A(n41286), .B(n41285), .Z(n41287) );
  AND U42392 ( .A(n41288), .B(n41287), .Z(n41315) );
  NAND U42393 ( .A(n42143), .B(n41289), .Z(n41291) );
  XNOR U42394 ( .A(a[1000]), .B(n4214), .Z(n41326) );
  NAND U42395 ( .A(n42144), .B(n41326), .Z(n41290) );
  AND U42396 ( .A(n41291), .B(n41290), .Z(n41341) );
  XOR U42397 ( .A(a[1004]), .B(n42012), .Z(n41329) );
  XNOR U42398 ( .A(n41341), .B(n41340), .Z(n41343) );
  XOR U42399 ( .A(a[1002]), .B(n42085), .Z(n41333) );
  AND U42400 ( .A(a[998]), .B(b[7]), .Z(n41334) );
  XNOR U42401 ( .A(n41335), .B(n41334), .Z(n41336) );
  AND U42402 ( .A(a[1006]), .B(b[0]), .Z(n41294) );
  XNOR U42403 ( .A(n41294), .B(n4071), .Z(n41296) );
  NANDN U42404 ( .A(b[0]), .B(a[1005]), .Z(n41295) );
  NAND U42405 ( .A(n41296), .B(n41295), .Z(n41337) );
  XNOR U42406 ( .A(n41336), .B(n41337), .Z(n41342) );
  XOR U42407 ( .A(n41343), .B(n41342), .Z(n41321) );
  NANDN U42408 ( .A(n41298), .B(n41297), .Z(n41302) );
  NANDN U42409 ( .A(n41300), .B(n41299), .Z(n41301) );
  AND U42410 ( .A(n41302), .B(n41301), .Z(n41320) );
  XNOR U42411 ( .A(n41321), .B(n41320), .Z(n41322) );
  NANDN U42412 ( .A(n41304), .B(n41303), .Z(n41308) );
  NAND U42413 ( .A(n41306), .B(n41305), .Z(n41307) );
  NAND U42414 ( .A(n41308), .B(n41307), .Z(n41323) );
  XNOR U42415 ( .A(n41322), .B(n41323), .Z(n41314) );
  XNOR U42416 ( .A(n41315), .B(n41314), .Z(n41316) );
  XNOR U42417 ( .A(n41317), .B(n41316), .Z(n41346) );
  XNOR U42418 ( .A(sreg[2022]), .B(n41346), .Z(n41348) );
  NANDN U42419 ( .A(sreg[2021]), .B(n41309), .Z(n41313) );
  NAND U42420 ( .A(n41311), .B(n41310), .Z(n41312) );
  NAND U42421 ( .A(n41313), .B(n41312), .Z(n41347) );
  XNOR U42422 ( .A(n41348), .B(n41347), .Z(c[2022]) );
  NANDN U42423 ( .A(n41315), .B(n41314), .Z(n41319) );
  NANDN U42424 ( .A(n41317), .B(n41316), .Z(n41318) );
  AND U42425 ( .A(n41319), .B(n41318), .Z(n41354) );
  NANDN U42426 ( .A(n41321), .B(n41320), .Z(n41325) );
  NANDN U42427 ( .A(n41323), .B(n41322), .Z(n41324) );
  AND U42428 ( .A(n41325), .B(n41324), .Z(n41352) );
  NAND U42429 ( .A(n42143), .B(n41326), .Z(n41328) );
  XNOR U42430 ( .A(a[1001]), .B(n4214), .Z(n41363) );
  NAND U42431 ( .A(n42144), .B(n41363), .Z(n41327) );
  AND U42432 ( .A(n41328), .B(n41327), .Z(n41378) );
  XOR U42433 ( .A(a[1005]), .B(n42012), .Z(n41366) );
  XNOR U42434 ( .A(n41378), .B(n41377), .Z(n41380) );
  AND U42435 ( .A(a[1007]), .B(b[0]), .Z(n41330) );
  XNOR U42436 ( .A(n41330), .B(n4071), .Z(n41332) );
  NANDN U42437 ( .A(b[0]), .B(a[1006]), .Z(n41331) );
  NAND U42438 ( .A(n41332), .B(n41331), .Z(n41374) );
  XOR U42439 ( .A(a[1003]), .B(n42085), .Z(n41367) );
  AND U42440 ( .A(a[999]), .B(b[7]), .Z(n41371) );
  XNOR U42441 ( .A(n41372), .B(n41371), .Z(n41373) );
  XNOR U42442 ( .A(n41374), .B(n41373), .Z(n41379) );
  XOR U42443 ( .A(n41380), .B(n41379), .Z(n41358) );
  NANDN U42444 ( .A(n41335), .B(n41334), .Z(n41339) );
  NANDN U42445 ( .A(n41337), .B(n41336), .Z(n41338) );
  AND U42446 ( .A(n41339), .B(n41338), .Z(n41357) );
  XNOR U42447 ( .A(n41358), .B(n41357), .Z(n41359) );
  NANDN U42448 ( .A(n41341), .B(n41340), .Z(n41345) );
  NAND U42449 ( .A(n41343), .B(n41342), .Z(n41344) );
  NAND U42450 ( .A(n41345), .B(n41344), .Z(n41360) );
  XNOR U42451 ( .A(n41359), .B(n41360), .Z(n41351) );
  XNOR U42452 ( .A(n41352), .B(n41351), .Z(n41353) );
  XNOR U42453 ( .A(n41354), .B(n41353), .Z(n41383) );
  XNOR U42454 ( .A(sreg[2023]), .B(n41383), .Z(n41385) );
  NANDN U42455 ( .A(sreg[2022]), .B(n41346), .Z(n41350) );
  NAND U42456 ( .A(n41348), .B(n41347), .Z(n41349) );
  NAND U42457 ( .A(n41350), .B(n41349), .Z(n41384) );
  XNOR U42458 ( .A(n41385), .B(n41384), .Z(c[2023]) );
  NANDN U42459 ( .A(n41352), .B(n41351), .Z(n41356) );
  NANDN U42460 ( .A(n41354), .B(n41353), .Z(n41355) );
  AND U42461 ( .A(n41356), .B(n41355), .Z(n41391) );
  NANDN U42462 ( .A(n41358), .B(n41357), .Z(n41362) );
  NANDN U42463 ( .A(n41360), .B(n41359), .Z(n41361) );
  AND U42464 ( .A(n41362), .B(n41361), .Z(n41389) );
  NAND U42465 ( .A(n42143), .B(n41363), .Z(n41365) );
  XNOR U42466 ( .A(a[1002]), .B(n4215), .Z(n41400) );
  NAND U42467 ( .A(n42144), .B(n41400), .Z(n41364) );
  AND U42468 ( .A(n41365), .B(n41364), .Z(n41415) );
  XOR U42469 ( .A(a[1006]), .B(n42012), .Z(n41403) );
  XNOR U42470 ( .A(n41415), .B(n41414), .Z(n41417) );
  XOR U42471 ( .A(a[1004]), .B(n42085), .Z(n41407) );
  AND U42472 ( .A(a[1000]), .B(b[7]), .Z(n41408) );
  XNOR U42473 ( .A(n41409), .B(n41408), .Z(n41410) );
  AND U42474 ( .A(a[1008]), .B(b[0]), .Z(n41368) );
  XNOR U42475 ( .A(n41368), .B(n4071), .Z(n41370) );
  NANDN U42476 ( .A(b[0]), .B(a[1007]), .Z(n41369) );
  NAND U42477 ( .A(n41370), .B(n41369), .Z(n41411) );
  XNOR U42478 ( .A(n41410), .B(n41411), .Z(n41416) );
  XOR U42479 ( .A(n41417), .B(n41416), .Z(n41395) );
  NANDN U42480 ( .A(n41372), .B(n41371), .Z(n41376) );
  NANDN U42481 ( .A(n41374), .B(n41373), .Z(n41375) );
  AND U42482 ( .A(n41376), .B(n41375), .Z(n41394) );
  XNOR U42483 ( .A(n41395), .B(n41394), .Z(n41396) );
  NANDN U42484 ( .A(n41378), .B(n41377), .Z(n41382) );
  NAND U42485 ( .A(n41380), .B(n41379), .Z(n41381) );
  NAND U42486 ( .A(n41382), .B(n41381), .Z(n41397) );
  XNOR U42487 ( .A(n41396), .B(n41397), .Z(n41388) );
  XNOR U42488 ( .A(n41389), .B(n41388), .Z(n41390) );
  XNOR U42489 ( .A(n41391), .B(n41390), .Z(n41420) );
  XNOR U42490 ( .A(sreg[2024]), .B(n41420), .Z(n41422) );
  NANDN U42491 ( .A(sreg[2023]), .B(n41383), .Z(n41387) );
  NAND U42492 ( .A(n41385), .B(n41384), .Z(n41386) );
  NAND U42493 ( .A(n41387), .B(n41386), .Z(n41421) );
  XNOR U42494 ( .A(n41422), .B(n41421), .Z(c[2024]) );
  NANDN U42495 ( .A(n41389), .B(n41388), .Z(n41393) );
  NANDN U42496 ( .A(n41391), .B(n41390), .Z(n41392) );
  AND U42497 ( .A(n41393), .B(n41392), .Z(n41428) );
  NANDN U42498 ( .A(n41395), .B(n41394), .Z(n41399) );
  NANDN U42499 ( .A(n41397), .B(n41396), .Z(n41398) );
  AND U42500 ( .A(n41399), .B(n41398), .Z(n41426) );
  NAND U42501 ( .A(n42143), .B(n41400), .Z(n41402) );
  XNOR U42502 ( .A(a[1003]), .B(n4215), .Z(n41437) );
  NAND U42503 ( .A(n42144), .B(n41437), .Z(n41401) );
  AND U42504 ( .A(n41402), .B(n41401), .Z(n41452) );
  XOR U42505 ( .A(a[1007]), .B(n42012), .Z(n41440) );
  XNOR U42506 ( .A(n41452), .B(n41451), .Z(n41454) );
  AND U42507 ( .A(a[1009]), .B(b[0]), .Z(n41404) );
  XNOR U42508 ( .A(n41404), .B(n4071), .Z(n41406) );
  NANDN U42509 ( .A(b[0]), .B(a[1008]), .Z(n41405) );
  NAND U42510 ( .A(n41406), .B(n41405), .Z(n41448) );
  XOR U42511 ( .A(a[1005]), .B(n42085), .Z(n41444) );
  AND U42512 ( .A(a[1001]), .B(b[7]), .Z(n41445) );
  XNOR U42513 ( .A(n41446), .B(n41445), .Z(n41447) );
  XNOR U42514 ( .A(n41448), .B(n41447), .Z(n41453) );
  XOR U42515 ( .A(n41454), .B(n41453), .Z(n41432) );
  NANDN U42516 ( .A(n41409), .B(n41408), .Z(n41413) );
  NANDN U42517 ( .A(n41411), .B(n41410), .Z(n41412) );
  AND U42518 ( .A(n41413), .B(n41412), .Z(n41431) );
  XNOR U42519 ( .A(n41432), .B(n41431), .Z(n41433) );
  NANDN U42520 ( .A(n41415), .B(n41414), .Z(n41419) );
  NAND U42521 ( .A(n41417), .B(n41416), .Z(n41418) );
  NAND U42522 ( .A(n41419), .B(n41418), .Z(n41434) );
  XNOR U42523 ( .A(n41433), .B(n41434), .Z(n41425) );
  XNOR U42524 ( .A(n41426), .B(n41425), .Z(n41427) );
  XNOR U42525 ( .A(n41428), .B(n41427), .Z(n41457) );
  XNOR U42526 ( .A(sreg[2025]), .B(n41457), .Z(n41459) );
  NANDN U42527 ( .A(sreg[2024]), .B(n41420), .Z(n41424) );
  NAND U42528 ( .A(n41422), .B(n41421), .Z(n41423) );
  NAND U42529 ( .A(n41424), .B(n41423), .Z(n41458) );
  XNOR U42530 ( .A(n41459), .B(n41458), .Z(c[2025]) );
  NANDN U42531 ( .A(n41426), .B(n41425), .Z(n41430) );
  NANDN U42532 ( .A(n41428), .B(n41427), .Z(n41429) );
  AND U42533 ( .A(n41430), .B(n41429), .Z(n41465) );
  NANDN U42534 ( .A(n41432), .B(n41431), .Z(n41436) );
  NANDN U42535 ( .A(n41434), .B(n41433), .Z(n41435) );
  AND U42536 ( .A(n41436), .B(n41435), .Z(n41463) );
  NAND U42537 ( .A(n42143), .B(n41437), .Z(n41439) );
  XNOR U42538 ( .A(a[1004]), .B(n4215), .Z(n41474) );
  NAND U42539 ( .A(n42144), .B(n41474), .Z(n41438) );
  AND U42540 ( .A(n41439), .B(n41438), .Z(n41489) );
  XOR U42541 ( .A(a[1008]), .B(n42012), .Z(n41477) );
  XNOR U42542 ( .A(n41489), .B(n41488), .Z(n41491) );
  AND U42543 ( .A(a[1010]), .B(b[0]), .Z(n41441) );
  XNOR U42544 ( .A(n41441), .B(n4071), .Z(n41443) );
  NANDN U42545 ( .A(b[0]), .B(a[1009]), .Z(n41442) );
  NAND U42546 ( .A(n41443), .B(n41442), .Z(n41485) );
  XOR U42547 ( .A(a[1006]), .B(n42085), .Z(n41481) );
  AND U42548 ( .A(a[1002]), .B(b[7]), .Z(n41482) );
  XNOR U42549 ( .A(n41483), .B(n41482), .Z(n41484) );
  XNOR U42550 ( .A(n41485), .B(n41484), .Z(n41490) );
  XOR U42551 ( .A(n41491), .B(n41490), .Z(n41469) );
  NANDN U42552 ( .A(n41446), .B(n41445), .Z(n41450) );
  NANDN U42553 ( .A(n41448), .B(n41447), .Z(n41449) );
  AND U42554 ( .A(n41450), .B(n41449), .Z(n41468) );
  XNOR U42555 ( .A(n41469), .B(n41468), .Z(n41470) );
  NANDN U42556 ( .A(n41452), .B(n41451), .Z(n41456) );
  NAND U42557 ( .A(n41454), .B(n41453), .Z(n41455) );
  NAND U42558 ( .A(n41456), .B(n41455), .Z(n41471) );
  XNOR U42559 ( .A(n41470), .B(n41471), .Z(n41462) );
  XNOR U42560 ( .A(n41463), .B(n41462), .Z(n41464) );
  XNOR U42561 ( .A(n41465), .B(n41464), .Z(n41494) );
  XNOR U42562 ( .A(sreg[2026]), .B(n41494), .Z(n41496) );
  NANDN U42563 ( .A(sreg[2025]), .B(n41457), .Z(n41461) );
  NAND U42564 ( .A(n41459), .B(n41458), .Z(n41460) );
  NAND U42565 ( .A(n41461), .B(n41460), .Z(n41495) );
  XNOR U42566 ( .A(n41496), .B(n41495), .Z(c[2026]) );
  NANDN U42567 ( .A(n41463), .B(n41462), .Z(n41467) );
  NANDN U42568 ( .A(n41465), .B(n41464), .Z(n41466) );
  AND U42569 ( .A(n41467), .B(n41466), .Z(n41502) );
  NANDN U42570 ( .A(n41469), .B(n41468), .Z(n41473) );
  NANDN U42571 ( .A(n41471), .B(n41470), .Z(n41472) );
  AND U42572 ( .A(n41473), .B(n41472), .Z(n41500) );
  NAND U42573 ( .A(n42143), .B(n41474), .Z(n41476) );
  XNOR U42574 ( .A(a[1005]), .B(n4215), .Z(n41511) );
  NAND U42575 ( .A(n42144), .B(n41511), .Z(n41475) );
  AND U42576 ( .A(n41476), .B(n41475), .Z(n41526) );
  XOR U42577 ( .A(a[1009]), .B(n42012), .Z(n41514) );
  XNOR U42578 ( .A(n41526), .B(n41525), .Z(n41528) );
  AND U42579 ( .A(a[1011]), .B(b[0]), .Z(n41478) );
  XNOR U42580 ( .A(n41478), .B(n4071), .Z(n41480) );
  NANDN U42581 ( .A(b[0]), .B(a[1010]), .Z(n41479) );
  NAND U42582 ( .A(n41480), .B(n41479), .Z(n41522) );
  XOR U42583 ( .A(a[1007]), .B(n42085), .Z(n41518) );
  AND U42584 ( .A(a[1003]), .B(b[7]), .Z(n41519) );
  XNOR U42585 ( .A(n41520), .B(n41519), .Z(n41521) );
  XNOR U42586 ( .A(n41522), .B(n41521), .Z(n41527) );
  XOR U42587 ( .A(n41528), .B(n41527), .Z(n41506) );
  NANDN U42588 ( .A(n41483), .B(n41482), .Z(n41487) );
  NANDN U42589 ( .A(n41485), .B(n41484), .Z(n41486) );
  AND U42590 ( .A(n41487), .B(n41486), .Z(n41505) );
  XNOR U42591 ( .A(n41506), .B(n41505), .Z(n41507) );
  NANDN U42592 ( .A(n41489), .B(n41488), .Z(n41493) );
  NAND U42593 ( .A(n41491), .B(n41490), .Z(n41492) );
  NAND U42594 ( .A(n41493), .B(n41492), .Z(n41508) );
  XNOR U42595 ( .A(n41507), .B(n41508), .Z(n41499) );
  XNOR U42596 ( .A(n41500), .B(n41499), .Z(n41501) );
  XNOR U42597 ( .A(n41502), .B(n41501), .Z(n41531) );
  XNOR U42598 ( .A(sreg[2027]), .B(n41531), .Z(n41533) );
  NANDN U42599 ( .A(sreg[2026]), .B(n41494), .Z(n41498) );
  NAND U42600 ( .A(n41496), .B(n41495), .Z(n41497) );
  NAND U42601 ( .A(n41498), .B(n41497), .Z(n41532) );
  XNOR U42602 ( .A(n41533), .B(n41532), .Z(c[2027]) );
  NANDN U42603 ( .A(n41500), .B(n41499), .Z(n41504) );
  NANDN U42604 ( .A(n41502), .B(n41501), .Z(n41503) );
  AND U42605 ( .A(n41504), .B(n41503), .Z(n41539) );
  NANDN U42606 ( .A(n41506), .B(n41505), .Z(n41510) );
  NANDN U42607 ( .A(n41508), .B(n41507), .Z(n41509) );
  AND U42608 ( .A(n41510), .B(n41509), .Z(n41537) );
  NAND U42609 ( .A(n42143), .B(n41511), .Z(n41513) );
  XNOR U42610 ( .A(a[1006]), .B(n4215), .Z(n41548) );
  NAND U42611 ( .A(n42144), .B(n41548), .Z(n41512) );
  AND U42612 ( .A(n41513), .B(n41512), .Z(n41563) );
  XOR U42613 ( .A(a[1010]), .B(n42012), .Z(n41551) );
  XNOR U42614 ( .A(n41563), .B(n41562), .Z(n41565) );
  AND U42615 ( .A(a[1012]), .B(b[0]), .Z(n41515) );
  XNOR U42616 ( .A(n41515), .B(n4071), .Z(n41517) );
  NANDN U42617 ( .A(b[0]), .B(a[1011]), .Z(n41516) );
  NAND U42618 ( .A(n41517), .B(n41516), .Z(n41559) );
  XOR U42619 ( .A(a[1008]), .B(n42085), .Z(n41555) );
  AND U42620 ( .A(a[1004]), .B(b[7]), .Z(n41556) );
  XNOR U42621 ( .A(n41557), .B(n41556), .Z(n41558) );
  XNOR U42622 ( .A(n41559), .B(n41558), .Z(n41564) );
  XOR U42623 ( .A(n41565), .B(n41564), .Z(n41543) );
  NANDN U42624 ( .A(n41520), .B(n41519), .Z(n41524) );
  NANDN U42625 ( .A(n41522), .B(n41521), .Z(n41523) );
  AND U42626 ( .A(n41524), .B(n41523), .Z(n41542) );
  XNOR U42627 ( .A(n41543), .B(n41542), .Z(n41544) );
  NANDN U42628 ( .A(n41526), .B(n41525), .Z(n41530) );
  NAND U42629 ( .A(n41528), .B(n41527), .Z(n41529) );
  NAND U42630 ( .A(n41530), .B(n41529), .Z(n41545) );
  XNOR U42631 ( .A(n41544), .B(n41545), .Z(n41536) );
  XNOR U42632 ( .A(n41537), .B(n41536), .Z(n41538) );
  XNOR U42633 ( .A(n41539), .B(n41538), .Z(n41568) );
  XNOR U42634 ( .A(sreg[2028]), .B(n41568), .Z(n41570) );
  NANDN U42635 ( .A(sreg[2027]), .B(n41531), .Z(n41535) );
  NAND U42636 ( .A(n41533), .B(n41532), .Z(n41534) );
  NAND U42637 ( .A(n41535), .B(n41534), .Z(n41569) );
  XNOR U42638 ( .A(n41570), .B(n41569), .Z(c[2028]) );
  NANDN U42639 ( .A(n41537), .B(n41536), .Z(n41541) );
  NANDN U42640 ( .A(n41539), .B(n41538), .Z(n41540) );
  AND U42641 ( .A(n41541), .B(n41540), .Z(n41576) );
  NANDN U42642 ( .A(n41543), .B(n41542), .Z(n41547) );
  NANDN U42643 ( .A(n41545), .B(n41544), .Z(n41546) );
  AND U42644 ( .A(n41547), .B(n41546), .Z(n41574) );
  NAND U42645 ( .A(n42143), .B(n41548), .Z(n41550) );
  XNOR U42646 ( .A(a[1007]), .B(n4215), .Z(n41585) );
  NAND U42647 ( .A(n42144), .B(n41585), .Z(n41549) );
  AND U42648 ( .A(n41550), .B(n41549), .Z(n41600) );
  XOR U42649 ( .A(a[1011]), .B(n42012), .Z(n41588) );
  XNOR U42650 ( .A(n41600), .B(n41599), .Z(n41602) );
  AND U42651 ( .A(a[1013]), .B(b[0]), .Z(n41552) );
  XNOR U42652 ( .A(n41552), .B(n4071), .Z(n41554) );
  NANDN U42653 ( .A(b[0]), .B(a[1012]), .Z(n41553) );
  NAND U42654 ( .A(n41554), .B(n41553), .Z(n41596) );
  XOR U42655 ( .A(a[1009]), .B(n42085), .Z(n41592) );
  AND U42656 ( .A(a[1005]), .B(b[7]), .Z(n41593) );
  XNOR U42657 ( .A(n41594), .B(n41593), .Z(n41595) );
  XNOR U42658 ( .A(n41596), .B(n41595), .Z(n41601) );
  XOR U42659 ( .A(n41602), .B(n41601), .Z(n41580) );
  NANDN U42660 ( .A(n41557), .B(n41556), .Z(n41561) );
  NANDN U42661 ( .A(n41559), .B(n41558), .Z(n41560) );
  AND U42662 ( .A(n41561), .B(n41560), .Z(n41579) );
  XNOR U42663 ( .A(n41580), .B(n41579), .Z(n41581) );
  NANDN U42664 ( .A(n41563), .B(n41562), .Z(n41567) );
  NAND U42665 ( .A(n41565), .B(n41564), .Z(n41566) );
  NAND U42666 ( .A(n41567), .B(n41566), .Z(n41582) );
  XNOR U42667 ( .A(n41581), .B(n41582), .Z(n41573) );
  XNOR U42668 ( .A(n41574), .B(n41573), .Z(n41575) );
  XNOR U42669 ( .A(n41576), .B(n41575), .Z(n41605) );
  XNOR U42670 ( .A(sreg[2029]), .B(n41605), .Z(n41607) );
  NANDN U42671 ( .A(sreg[2028]), .B(n41568), .Z(n41572) );
  NAND U42672 ( .A(n41570), .B(n41569), .Z(n41571) );
  NAND U42673 ( .A(n41572), .B(n41571), .Z(n41606) );
  XNOR U42674 ( .A(n41607), .B(n41606), .Z(c[2029]) );
  NANDN U42675 ( .A(n41574), .B(n41573), .Z(n41578) );
  NANDN U42676 ( .A(n41576), .B(n41575), .Z(n41577) );
  AND U42677 ( .A(n41578), .B(n41577), .Z(n41613) );
  NANDN U42678 ( .A(n41580), .B(n41579), .Z(n41584) );
  NANDN U42679 ( .A(n41582), .B(n41581), .Z(n41583) );
  AND U42680 ( .A(n41584), .B(n41583), .Z(n41611) );
  NAND U42681 ( .A(n42143), .B(n41585), .Z(n41587) );
  XNOR U42682 ( .A(a[1008]), .B(n4215), .Z(n41622) );
  NAND U42683 ( .A(n42144), .B(n41622), .Z(n41586) );
  AND U42684 ( .A(n41587), .B(n41586), .Z(n41637) );
  XOR U42685 ( .A(a[1012]), .B(n42012), .Z(n41625) );
  XNOR U42686 ( .A(n41637), .B(n41636), .Z(n41639) );
  AND U42687 ( .A(a[1014]), .B(b[0]), .Z(n41589) );
  XNOR U42688 ( .A(n41589), .B(n4071), .Z(n41591) );
  NANDN U42689 ( .A(b[0]), .B(a[1013]), .Z(n41590) );
  NAND U42690 ( .A(n41591), .B(n41590), .Z(n41633) );
  XOR U42691 ( .A(a[1010]), .B(n42085), .Z(n41626) );
  AND U42692 ( .A(a[1006]), .B(b[7]), .Z(n41630) );
  XNOR U42693 ( .A(n41631), .B(n41630), .Z(n41632) );
  XNOR U42694 ( .A(n41633), .B(n41632), .Z(n41638) );
  XOR U42695 ( .A(n41639), .B(n41638), .Z(n41617) );
  NANDN U42696 ( .A(n41594), .B(n41593), .Z(n41598) );
  NANDN U42697 ( .A(n41596), .B(n41595), .Z(n41597) );
  AND U42698 ( .A(n41598), .B(n41597), .Z(n41616) );
  XNOR U42699 ( .A(n41617), .B(n41616), .Z(n41618) );
  NANDN U42700 ( .A(n41600), .B(n41599), .Z(n41604) );
  NAND U42701 ( .A(n41602), .B(n41601), .Z(n41603) );
  NAND U42702 ( .A(n41604), .B(n41603), .Z(n41619) );
  XNOR U42703 ( .A(n41618), .B(n41619), .Z(n41610) );
  XNOR U42704 ( .A(n41611), .B(n41610), .Z(n41612) );
  XNOR U42705 ( .A(n41613), .B(n41612), .Z(n41642) );
  XNOR U42706 ( .A(sreg[2030]), .B(n41642), .Z(n41644) );
  NANDN U42707 ( .A(sreg[2029]), .B(n41605), .Z(n41609) );
  NAND U42708 ( .A(n41607), .B(n41606), .Z(n41608) );
  NAND U42709 ( .A(n41609), .B(n41608), .Z(n41643) );
  XNOR U42710 ( .A(n41644), .B(n41643), .Z(c[2030]) );
  NANDN U42711 ( .A(n41611), .B(n41610), .Z(n41615) );
  NANDN U42712 ( .A(n41613), .B(n41612), .Z(n41614) );
  AND U42713 ( .A(n41615), .B(n41614), .Z(n41650) );
  NANDN U42714 ( .A(n41617), .B(n41616), .Z(n41621) );
  NANDN U42715 ( .A(n41619), .B(n41618), .Z(n41620) );
  AND U42716 ( .A(n41621), .B(n41620), .Z(n41648) );
  NAND U42717 ( .A(n42143), .B(n41622), .Z(n41624) );
  XNOR U42718 ( .A(a[1009]), .B(n4216), .Z(n41659) );
  NAND U42719 ( .A(n42144), .B(n41659), .Z(n41623) );
  AND U42720 ( .A(n41624), .B(n41623), .Z(n41674) );
  XOR U42721 ( .A(a[1013]), .B(n42012), .Z(n41662) );
  XNOR U42722 ( .A(n41674), .B(n41673), .Z(n41676) );
  XOR U42723 ( .A(a[1011]), .B(n42085), .Z(n41666) );
  AND U42724 ( .A(a[1007]), .B(b[7]), .Z(n41667) );
  XNOR U42725 ( .A(n41668), .B(n41667), .Z(n41669) );
  AND U42726 ( .A(a[1015]), .B(b[0]), .Z(n41627) );
  XNOR U42727 ( .A(n41627), .B(n4071), .Z(n41629) );
  NANDN U42728 ( .A(b[0]), .B(a[1014]), .Z(n41628) );
  NAND U42729 ( .A(n41629), .B(n41628), .Z(n41670) );
  XNOR U42730 ( .A(n41669), .B(n41670), .Z(n41675) );
  XOR U42731 ( .A(n41676), .B(n41675), .Z(n41654) );
  NANDN U42732 ( .A(n41631), .B(n41630), .Z(n41635) );
  NANDN U42733 ( .A(n41633), .B(n41632), .Z(n41634) );
  AND U42734 ( .A(n41635), .B(n41634), .Z(n41653) );
  XNOR U42735 ( .A(n41654), .B(n41653), .Z(n41655) );
  NANDN U42736 ( .A(n41637), .B(n41636), .Z(n41641) );
  NAND U42737 ( .A(n41639), .B(n41638), .Z(n41640) );
  NAND U42738 ( .A(n41641), .B(n41640), .Z(n41656) );
  XNOR U42739 ( .A(n41655), .B(n41656), .Z(n41647) );
  XNOR U42740 ( .A(n41648), .B(n41647), .Z(n41649) );
  XNOR U42741 ( .A(n41650), .B(n41649), .Z(n41679) );
  XNOR U42742 ( .A(sreg[2031]), .B(n41679), .Z(n41681) );
  NANDN U42743 ( .A(sreg[2030]), .B(n41642), .Z(n41646) );
  NAND U42744 ( .A(n41644), .B(n41643), .Z(n41645) );
  NAND U42745 ( .A(n41646), .B(n41645), .Z(n41680) );
  XNOR U42746 ( .A(n41681), .B(n41680), .Z(c[2031]) );
  NANDN U42747 ( .A(n41648), .B(n41647), .Z(n41652) );
  NANDN U42748 ( .A(n41650), .B(n41649), .Z(n41651) );
  AND U42749 ( .A(n41652), .B(n41651), .Z(n41687) );
  NANDN U42750 ( .A(n41654), .B(n41653), .Z(n41658) );
  NANDN U42751 ( .A(n41656), .B(n41655), .Z(n41657) );
  AND U42752 ( .A(n41658), .B(n41657), .Z(n41685) );
  NAND U42753 ( .A(n42143), .B(n41659), .Z(n41661) );
  XNOR U42754 ( .A(a[1010]), .B(n4216), .Z(n41696) );
  NAND U42755 ( .A(n42144), .B(n41696), .Z(n41660) );
  AND U42756 ( .A(n41661), .B(n41660), .Z(n41711) );
  XOR U42757 ( .A(a[1014]), .B(n42012), .Z(n41699) );
  XNOR U42758 ( .A(n41711), .B(n41710), .Z(n41713) );
  AND U42759 ( .A(a[1016]), .B(b[0]), .Z(n41663) );
  XNOR U42760 ( .A(n41663), .B(n4071), .Z(n41665) );
  NANDN U42761 ( .A(b[0]), .B(a[1015]), .Z(n41664) );
  NAND U42762 ( .A(n41665), .B(n41664), .Z(n41707) );
  XOR U42763 ( .A(a[1012]), .B(n42085), .Z(n41700) );
  AND U42764 ( .A(a[1008]), .B(b[7]), .Z(n41704) );
  XNOR U42765 ( .A(n41705), .B(n41704), .Z(n41706) );
  XNOR U42766 ( .A(n41707), .B(n41706), .Z(n41712) );
  XOR U42767 ( .A(n41713), .B(n41712), .Z(n41691) );
  NANDN U42768 ( .A(n41668), .B(n41667), .Z(n41672) );
  NANDN U42769 ( .A(n41670), .B(n41669), .Z(n41671) );
  AND U42770 ( .A(n41672), .B(n41671), .Z(n41690) );
  XNOR U42771 ( .A(n41691), .B(n41690), .Z(n41692) );
  NANDN U42772 ( .A(n41674), .B(n41673), .Z(n41678) );
  NAND U42773 ( .A(n41676), .B(n41675), .Z(n41677) );
  NAND U42774 ( .A(n41678), .B(n41677), .Z(n41693) );
  XNOR U42775 ( .A(n41692), .B(n41693), .Z(n41684) );
  XNOR U42776 ( .A(n41685), .B(n41684), .Z(n41686) );
  XNOR U42777 ( .A(n41687), .B(n41686), .Z(n41716) );
  XNOR U42778 ( .A(sreg[2032]), .B(n41716), .Z(n41718) );
  NANDN U42779 ( .A(sreg[2031]), .B(n41679), .Z(n41683) );
  NAND U42780 ( .A(n41681), .B(n41680), .Z(n41682) );
  NAND U42781 ( .A(n41683), .B(n41682), .Z(n41717) );
  XNOR U42782 ( .A(n41718), .B(n41717), .Z(c[2032]) );
  NANDN U42783 ( .A(n41685), .B(n41684), .Z(n41689) );
  NANDN U42784 ( .A(n41687), .B(n41686), .Z(n41688) );
  AND U42785 ( .A(n41689), .B(n41688), .Z(n41724) );
  NANDN U42786 ( .A(n41691), .B(n41690), .Z(n41695) );
  NANDN U42787 ( .A(n41693), .B(n41692), .Z(n41694) );
  AND U42788 ( .A(n41695), .B(n41694), .Z(n41722) );
  NAND U42789 ( .A(n42143), .B(n41696), .Z(n41698) );
  XNOR U42790 ( .A(a[1011]), .B(n4216), .Z(n41733) );
  NAND U42791 ( .A(n42144), .B(n41733), .Z(n41697) );
  AND U42792 ( .A(n41698), .B(n41697), .Z(n41748) );
  XOR U42793 ( .A(a[1015]), .B(n42012), .Z(n41736) );
  XNOR U42794 ( .A(n41748), .B(n41747), .Z(n41750) );
  XOR U42795 ( .A(a[1013]), .B(n42085), .Z(n41737) );
  AND U42796 ( .A(a[1009]), .B(b[7]), .Z(n41741) );
  XNOR U42797 ( .A(n41742), .B(n41741), .Z(n41743) );
  AND U42798 ( .A(a[1017]), .B(b[0]), .Z(n41701) );
  XNOR U42799 ( .A(n41701), .B(n4071), .Z(n41703) );
  NANDN U42800 ( .A(b[0]), .B(a[1016]), .Z(n41702) );
  NAND U42801 ( .A(n41703), .B(n41702), .Z(n41744) );
  XNOR U42802 ( .A(n41743), .B(n41744), .Z(n41749) );
  XOR U42803 ( .A(n41750), .B(n41749), .Z(n41728) );
  NANDN U42804 ( .A(n41705), .B(n41704), .Z(n41709) );
  NANDN U42805 ( .A(n41707), .B(n41706), .Z(n41708) );
  AND U42806 ( .A(n41709), .B(n41708), .Z(n41727) );
  XNOR U42807 ( .A(n41728), .B(n41727), .Z(n41729) );
  NANDN U42808 ( .A(n41711), .B(n41710), .Z(n41715) );
  NAND U42809 ( .A(n41713), .B(n41712), .Z(n41714) );
  NAND U42810 ( .A(n41715), .B(n41714), .Z(n41730) );
  XNOR U42811 ( .A(n41729), .B(n41730), .Z(n41721) );
  XNOR U42812 ( .A(n41722), .B(n41721), .Z(n41723) );
  XNOR U42813 ( .A(n41724), .B(n41723), .Z(n41753) );
  XNOR U42814 ( .A(sreg[2033]), .B(n41753), .Z(n41755) );
  NANDN U42815 ( .A(sreg[2032]), .B(n41716), .Z(n41720) );
  NAND U42816 ( .A(n41718), .B(n41717), .Z(n41719) );
  NAND U42817 ( .A(n41720), .B(n41719), .Z(n41754) );
  XNOR U42818 ( .A(n41755), .B(n41754), .Z(c[2033]) );
  NANDN U42819 ( .A(n41722), .B(n41721), .Z(n41726) );
  NANDN U42820 ( .A(n41724), .B(n41723), .Z(n41725) );
  AND U42821 ( .A(n41726), .B(n41725), .Z(n41761) );
  NANDN U42822 ( .A(n41728), .B(n41727), .Z(n41732) );
  NANDN U42823 ( .A(n41730), .B(n41729), .Z(n41731) );
  AND U42824 ( .A(n41732), .B(n41731), .Z(n41759) );
  NAND U42825 ( .A(n42143), .B(n41733), .Z(n41735) );
  XNOR U42826 ( .A(a[1012]), .B(n4216), .Z(n41770) );
  NAND U42827 ( .A(n42144), .B(n41770), .Z(n41734) );
  AND U42828 ( .A(n41735), .B(n41734), .Z(n41785) );
  XOR U42829 ( .A(a[1016]), .B(n42012), .Z(n41773) );
  XNOR U42830 ( .A(n41785), .B(n41784), .Z(n41787) );
  XOR U42831 ( .A(a[1014]), .B(n42085), .Z(n41777) );
  AND U42832 ( .A(a[1010]), .B(b[7]), .Z(n41778) );
  XNOR U42833 ( .A(n41779), .B(n41778), .Z(n41780) );
  AND U42834 ( .A(a[1018]), .B(b[0]), .Z(n41738) );
  XNOR U42835 ( .A(n41738), .B(n4071), .Z(n41740) );
  NANDN U42836 ( .A(b[0]), .B(a[1017]), .Z(n41739) );
  NAND U42837 ( .A(n41740), .B(n41739), .Z(n41781) );
  XNOR U42838 ( .A(n41780), .B(n41781), .Z(n41786) );
  XOR U42839 ( .A(n41787), .B(n41786), .Z(n41765) );
  NANDN U42840 ( .A(n41742), .B(n41741), .Z(n41746) );
  NANDN U42841 ( .A(n41744), .B(n41743), .Z(n41745) );
  AND U42842 ( .A(n41746), .B(n41745), .Z(n41764) );
  XNOR U42843 ( .A(n41765), .B(n41764), .Z(n41766) );
  NANDN U42844 ( .A(n41748), .B(n41747), .Z(n41752) );
  NAND U42845 ( .A(n41750), .B(n41749), .Z(n41751) );
  NAND U42846 ( .A(n41752), .B(n41751), .Z(n41767) );
  XNOR U42847 ( .A(n41766), .B(n41767), .Z(n41758) );
  XNOR U42848 ( .A(n41759), .B(n41758), .Z(n41760) );
  XNOR U42849 ( .A(n41761), .B(n41760), .Z(n41790) );
  XNOR U42850 ( .A(sreg[2034]), .B(n41790), .Z(n41792) );
  NANDN U42851 ( .A(sreg[2033]), .B(n41753), .Z(n41757) );
  NAND U42852 ( .A(n41755), .B(n41754), .Z(n41756) );
  NAND U42853 ( .A(n41757), .B(n41756), .Z(n41791) );
  XNOR U42854 ( .A(n41792), .B(n41791), .Z(c[2034]) );
  NANDN U42855 ( .A(n41759), .B(n41758), .Z(n41763) );
  NANDN U42856 ( .A(n41761), .B(n41760), .Z(n41762) );
  AND U42857 ( .A(n41763), .B(n41762), .Z(n41798) );
  NANDN U42858 ( .A(n41765), .B(n41764), .Z(n41769) );
  NANDN U42859 ( .A(n41767), .B(n41766), .Z(n41768) );
  AND U42860 ( .A(n41769), .B(n41768), .Z(n41796) );
  NAND U42861 ( .A(n42143), .B(n41770), .Z(n41772) );
  XNOR U42862 ( .A(a[1013]), .B(n4216), .Z(n41807) );
  NAND U42863 ( .A(n42144), .B(n41807), .Z(n41771) );
  AND U42864 ( .A(n41772), .B(n41771), .Z(n41822) );
  XOR U42865 ( .A(a[1017]), .B(n42012), .Z(n41810) );
  XNOR U42866 ( .A(n41822), .B(n41821), .Z(n41824) );
  AND U42867 ( .A(a[1019]), .B(b[0]), .Z(n41774) );
  XNOR U42868 ( .A(n41774), .B(n4071), .Z(n41776) );
  NANDN U42869 ( .A(b[0]), .B(a[1018]), .Z(n41775) );
  NAND U42870 ( .A(n41776), .B(n41775), .Z(n41818) );
  XOR U42871 ( .A(a[1015]), .B(n42085), .Z(n41811) );
  AND U42872 ( .A(a[1011]), .B(b[7]), .Z(n41815) );
  XNOR U42873 ( .A(n41816), .B(n41815), .Z(n41817) );
  XNOR U42874 ( .A(n41818), .B(n41817), .Z(n41823) );
  XOR U42875 ( .A(n41824), .B(n41823), .Z(n41802) );
  NANDN U42876 ( .A(n41779), .B(n41778), .Z(n41783) );
  NANDN U42877 ( .A(n41781), .B(n41780), .Z(n41782) );
  AND U42878 ( .A(n41783), .B(n41782), .Z(n41801) );
  XNOR U42879 ( .A(n41802), .B(n41801), .Z(n41803) );
  NANDN U42880 ( .A(n41785), .B(n41784), .Z(n41789) );
  NAND U42881 ( .A(n41787), .B(n41786), .Z(n41788) );
  NAND U42882 ( .A(n41789), .B(n41788), .Z(n41804) );
  XNOR U42883 ( .A(n41803), .B(n41804), .Z(n41795) );
  XNOR U42884 ( .A(n41796), .B(n41795), .Z(n41797) );
  XNOR U42885 ( .A(n41798), .B(n41797), .Z(n41827) );
  XNOR U42886 ( .A(sreg[2035]), .B(n41827), .Z(n41829) );
  NANDN U42887 ( .A(sreg[2034]), .B(n41790), .Z(n41794) );
  NAND U42888 ( .A(n41792), .B(n41791), .Z(n41793) );
  NAND U42889 ( .A(n41794), .B(n41793), .Z(n41828) );
  XNOR U42890 ( .A(n41829), .B(n41828), .Z(c[2035]) );
  NANDN U42891 ( .A(n41796), .B(n41795), .Z(n41800) );
  NANDN U42892 ( .A(n41798), .B(n41797), .Z(n41799) );
  AND U42893 ( .A(n41800), .B(n41799), .Z(n41835) );
  NANDN U42894 ( .A(n41802), .B(n41801), .Z(n41806) );
  NANDN U42895 ( .A(n41804), .B(n41803), .Z(n41805) );
  AND U42896 ( .A(n41806), .B(n41805), .Z(n41833) );
  NAND U42897 ( .A(n42143), .B(n41807), .Z(n41809) );
  XNOR U42898 ( .A(a[1014]), .B(n4216), .Z(n41844) );
  NAND U42899 ( .A(n42144), .B(n41844), .Z(n41808) );
  AND U42900 ( .A(n41809), .B(n41808), .Z(n41859) );
  XOR U42901 ( .A(a[1018]), .B(n42012), .Z(n41847) );
  XNOR U42902 ( .A(n41859), .B(n41858), .Z(n41861) );
  XOR U42903 ( .A(a[1016]), .B(n42085), .Z(n41848) );
  AND U42904 ( .A(a[1012]), .B(b[7]), .Z(n41852) );
  XNOR U42905 ( .A(n41853), .B(n41852), .Z(n41854) );
  AND U42906 ( .A(a[1020]), .B(b[0]), .Z(n41812) );
  XNOR U42907 ( .A(n41812), .B(n4071), .Z(n41814) );
  NANDN U42908 ( .A(b[0]), .B(a[1019]), .Z(n41813) );
  NAND U42909 ( .A(n41814), .B(n41813), .Z(n41855) );
  XNOR U42910 ( .A(n41854), .B(n41855), .Z(n41860) );
  XOR U42911 ( .A(n41861), .B(n41860), .Z(n41839) );
  NANDN U42912 ( .A(n41816), .B(n41815), .Z(n41820) );
  NANDN U42913 ( .A(n41818), .B(n41817), .Z(n41819) );
  AND U42914 ( .A(n41820), .B(n41819), .Z(n41838) );
  XNOR U42915 ( .A(n41839), .B(n41838), .Z(n41840) );
  NANDN U42916 ( .A(n41822), .B(n41821), .Z(n41826) );
  NAND U42917 ( .A(n41824), .B(n41823), .Z(n41825) );
  NAND U42918 ( .A(n41826), .B(n41825), .Z(n41841) );
  XNOR U42919 ( .A(n41840), .B(n41841), .Z(n41832) );
  XNOR U42920 ( .A(n41833), .B(n41832), .Z(n41834) );
  XNOR U42921 ( .A(n41835), .B(n41834), .Z(n41864) );
  XNOR U42922 ( .A(sreg[2036]), .B(n41864), .Z(n41866) );
  NANDN U42923 ( .A(sreg[2035]), .B(n41827), .Z(n41831) );
  NAND U42924 ( .A(n41829), .B(n41828), .Z(n41830) );
  NAND U42925 ( .A(n41831), .B(n41830), .Z(n41865) );
  XNOR U42926 ( .A(n41866), .B(n41865), .Z(c[2036]) );
  NANDN U42927 ( .A(n41833), .B(n41832), .Z(n41837) );
  NANDN U42928 ( .A(n41835), .B(n41834), .Z(n41836) );
  AND U42929 ( .A(n41837), .B(n41836), .Z(n41872) );
  NANDN U42930 ( .A(n41839), .B(n41838), .Z(n41843) );
  NANDN U42931 ( .A(n41841), .B(n41840), .Z(n41842) );
  AND U42932 ( .A(n41843), .B(n41842), .Z(n41870) );
  NAND U42933 ( .A(n42143), .B(n41844), .Z(n41846) );
  XNOR U42934 ( .A(a[1015]), .B(n4216), .Z(n41881) );
  NAND U42935 ( .A(n42144), .B(n41881), .Z(n41845) );
  AND U42936 ( .A(n41846), .B(n41845), .Z(n41900) );
  XNOR U42937 ( .A(a[1019]), .B(n42012), .Z(n41884) );
  XNOR U42938 ( .A(n41900), .B(n41899), .Z(n41902) );
  XNOR U42939 ( .A(a[1017]), .B(n42085), .Z(n41890) );
  AND U42940 ( .A(a[1013]), .B(b[7]), .Z(n41893) );
  XNOR U42941 ( .A(n41894), .B(n41893), .Z(n41895) );
  AND U42942 ( .A(a[1021]), .B(b[0]), .Z(n41849) );
  XNOR U42943 ( .A(n41849), .B(n4071), .Z(n41851) );
  NANDN U42944 ( .A(b[0]), .B(a[1020]), .Z(n41850) );
  NAND U42945 ( .A(n41851), .B(n41850), .Z(n41896) );
  XNOR U42946 ( .A(n41895), .B(n41896), .Z(n41901) );
  XOR U42947 ( .A(n41902), .B(n41901), .Z(n41876) );
  NANDN U42948 ( .A(n41853), .B(n41852), .Z(n41857) );
  NANDN U42949 ( .A(n41855), .B(n41854), .Z(n41856) );
  AND U42950 ( .A(n41857), .B(n41856), .Z(n41875) );
  XNOR U42951 ( .A(n41876), .B(n41875), .Z(n41877) );
  NANDN U42952 ( .A(n41859), .B(n41858), .Z(n41863) );
  NAND U42953 ( .A(n41861), .B(n41860), .Z(n41862) );
  NAND U42954 ( .A(n41863), .B(n41862), .Z(n41878) );
  XNOR U42955 ( .A(n41877), .B(n41878), .Z(n41869) );
  XNOR U42956 ( .A(n41870), .B(n41869), .Z(n41871) );
  XNOR U42957 ( .A(n41872), .B(n41871), .Z(n41905) );
  XNOR U42958 ( .A(sreg[2037]), .B(n41905), .Z(n41907) );
  NANDN U42959 ( .A(sreg[2036]), .B(n41864), .Z(n41868) );
  NAND U42960 ( .A(n41866), .B(n41865), .Z(n41867) );
  NAND U42961 ( .A(n41868), .B(n41867), .Z(n41906) );
  XNOR U42962 ( .A(n41907), .B(n41906), .Z(c[2037]) );
  NANDN U42963 ( .A(n41870), .B(n41869), .Z(n41874) );
  NANDN U42964 ( .A(n41872), .B(n41871), .Z(n41873) );
  AND U42965 ( .A(n41874), .B(n41873), .Z(n41913) );
  NANDN U42966 ( .A(n41876), .B(n41875), .Z(n41880) );
  NANDN U42967 ( .A(n41878), .B(n41877), .Z(n41879) );
  AND U42968 ( .A(n41880), .B(n41879), .Z(n41911) );
  NAND U42969 ( .A(n42143), .B(n41881), .Z(n41883) );
  XNOR U42970 ( .A(a[1016]), .B(n4217), .Z(n41934) );
  NAND U42971 ( .A(n42144), .B(n41934), .Z(n41882) );
  NAND U42972 ( .A(n41883), .B(n41882), .Z(n41923) );
  XNOR U42973 ( .A(a[1020]), .B(n42012), .Z(n41937) );
  NANDN U42974 ( .A(n4064), .B(n41937), .Z(n41886) );
  NAND U42975 ( .A(n42047), .B(n41884), .Z(n41885) );
  NAND U42976 ( .A(n41886), .B(n41885), .Z(n41922) );
  AND U42977 ( .A(a[1022]), .B(b[0]), .Z(n41887) );
  XNOR U42978 ( .A(n41887), .B(n4071), .Z(n41889) );
  NANDN U42979 ( .A(b[0]), .B(a[1021]), .Z(n41888) );
  NAND U42980 ( .A(n41889), .B(n41888), .Z(n41931) );
  XNOR U42981 ( .A(a[1018]), .B(n42085), .Z(n41943) );
  NANDN U42982 ( .A(n4065), .B(n41943), .Z(n41892) );
  NAND U42983 ( .A(n41890), .B(n42115), .Z(n41891) );
  NAND U42984 ( .A(n41892), .B(n41891), .Z(n41929) );
  AND U42985 ( .A(a[1014]), .B(b[7]), .Z(n41928) );
  XNOR U42986 ( .A(n41931), .B(n41930), .Z(n41924) );
  XNOR U42987 ( .A(n41925), .B(n41924), .Z(n41917) );
  NANDN U42988 ( .A(n41894), .B(n41893), .Z(n41898) );
  NANDN U42989 ( .A(n41896), .B(n41895), .Z(n41897) );
  AND U42990 ( .A(n41898), .B(n41897), .Z(n41916) );
  NANDN U42991 ( .A(n41900), .B(n41899), .Z(n41904) );
  NAND U42992 ( .A(n41902), .B(n41901), .Z(n41903) );
  AND U42993 ( .A(n41904), .B(n41903), .Z(n41919) );
  XNOR U42994 ( .A(n41911), .B(n41910), .Z(n41912) );
  XNOR U42995 ( .A(n41913), .B(n41912), .Z(n41946) );
  XNOR U42996 ( .A(sreg[2038]), .B(n41946), .Z(n41948) );
  NANDN U42997 ( .A(sreg[2037]), .B(n41905), .Z(n41909) );
  NAND U42998 ( .A(n41907), .B(n41906), .Z(n41908) );
  NAND U42999 ( .A(n41909), .B(n41908), .Z(n41947) );
  XNOR U43000 ( .A(n41948), .B(n41947), .Z(c[2038]) );
  NANDN U43001 ( .A(n41911), .B(n41910), .Z(n41915) );
  NANDN U43002 ( .A(n41913), .B(n41912), .Z(n41914) );
  NAND U43003 ( .A(n41915), .B(n41914), .Z(n41959) );
  NAND U43004 ( .A(n41917), .B(n41916), .Z(n41921) );
  NAND U43005 ( .A(n41919), .B(n41918), .Z(n41920) );
  NAND U43006 ( .A(n41921), .B(n41920), .Z(n41957) );
  NAND U43007 ( .A(n41923), .B(n41922), .Z(n41927) );
  NAND U43008 ( .A(n41925), .B(n41924), .Z(n41926) );
  AND U43009 ( .A(n41927), .B(n41926), .Z(n41988) );
  NAND U43010 ( .A(n41929), .B(n41928), .Z(n41933) );
  NANDN U43011 ( .A(n41931), .B(n41930), .Z(n41932) );
  NAND U43012 ( .A(n41933), .B(n41932), .Z(n41986) );
  NAND U43013 ( .A(n42143), .B(n41934), .Z(n41936) );
  XNOR U43014 ( .A(a[1017]), .B(n4217), .Z(n41974) );
  NAND U43015 ( .A(n42144), .B(n41974), .Z(n41935) );
  NAND U43016 ( .A(n41936), .B(n41935), .Z(n41965) );
  XNOR U43017 ( .A(a[1021]), .B(n42012), .Z(n41977) );
  NANDN U43018 ( .A(n4064), .B(n41977), .Z(n41939) );
  NAND U43019 ( .A(n42047), .B(n41937), .Z(n41938) );
  NAND U43020 ( .A(n41939), .B(n41938), .Z(n41963) );
  AND U43021 ( .A(a[1023]), .B(b[0]), .Z(n41940) );
  XNOR U43022 ( .A(n41940), .B(n4071), .Z(n41942) );
  NANDN U43023 ( .A(b[0]), .B(a[1022]), .Z(n41941) );
  NAND U43024 ( .A(n41942), .B(n41941), .Z(n41971) );
  XNOR U43025 ( .A(a[1019]), .B(n42085), .Z(n41980) );
  NANDN U43026 ( .A(n4065), .B(n41980), .Z(n41945) );
  NAND U43027 ( .A(n41943), .B(n42115), .Z(n41944) );
  NAND U43028 ( .A(n41945), .B(n41944), .Z(n41969) );
  AND U43029 ( .A(a[1015]), .B(b[7]), .Z(n41968) );
  XNOR U43030 ( .A(n41971), .B(n41970), .Z(n41962) );
  XOR U43031 ( .A(n41988), .B(n41987), .Z(n41956) );
  XNOR U43032 ( .A(sreg[2039]), .B(n41951), .Z(n41953) );
  NANDN U43033 ( .A(sreg[2038]), .B(n41946), .Z(n41950) );
  NAND U43034 ( .A(n41948), .B(n41947), .Z(n41949) );
  NAND U43035 ( .A(n41950), .B(n41949), .Z(n41952) );
  XNOR U43036 ( .A(n41953), .B(n41952), .Z(c[2039]) );
  NANDN U43037 ( .A(sreg[2039]), .B(n41951), .Z(n41955) );
  NAND U43038 ( .A(n41953), .B(n41952), .Z(n41954) );
  AND U43039 ( .A(n41955), .B(n41954), .Z(n41992) );
  NAND U43040 ( .A(n41957), .B(n41956), .Z(n41961) );
  NAND U43041 ( .A(n41959), .B(n41958), .Z(n41960) );
  AND U43042 ( .A(n41961), .B(n41960), .Z(n41996) );
  NAND U43043 ( .A(n41963), .B(n41962), .Z(n41967) );
  NAND U43044 ( .A(n41965), .B(n41964), .Z(n41966) );
  NAND U43045 ( .A(n41967), .B(n41966), .Z(n42024) );
  NAND U43046 ( .A(n41969), .B(n41968), .Z(n41973) );
  NANDN U43047 ( .A(n41971), .B(n41970), .Z(n41972) );
  NAND U43048 ( .A(n41973), .B(n41972), .Z(n42022) );
  NAND U43049 ( .A(n42143), .B(n41974), .Z(n41976) );
  XNOR U43050 ( .A(a[1018]), .B(n4217), .Z(n42005) );
  NAND U43051 ( .A(n42144), .B(n42005), .Z(n41975) );
  NAND U43052 ( .A(n41976), .B(n41975), .Z(n42002) );
  XNOR U43053 ( .A(b[3]), .B(a[1022]), .Z(n42011) );
  OR U43054 ( .A(n42011), .B(n4064), .Z(n41979) );
  NAND U43055 ( .A(n42047), .B(n41977), .Z(n41978) );
  NAND U43056 ( .A(n41979), .B(n41978), .Z(n42000) );
  XNOR U43057 ( .A(a[1020]), .B(n42085), .Z(n42008) );
  NANDN U43058 ( .A(n4065), .B(n42008), .Z(n41982) );
  NAND U43059 ( .A(n41980), .B(n42115), .Z(n41981) );
  NAND U43060 ( .A(n41982), .B(n41981), .Z(n42018) );
  NAND U43061 ( .A(b[1]), .B(b[0]), .Z(n41984) );
  NANDN U43062 ( .A(a[1023]), .B(b[1]), .Z(n41983) );
  NAND U43063 ( .A(n41984), .B(n41983), .Z(n42016) );
  AND U43064 ( .A(a[1016]), .B(b[7]), .Z(n42015) );
  NAND U43065 ( .A(n41986), .B(n41985), .Z(n41990) );
  NANDN U43066 ( .A(n41988), .B(n41987), .Z(n41989) );
  AND U43067 ( .A(n41990), .B(n41989), .Z(n41994) );
  XOR U43068 ( .A(n41993), .B(n41994), .Z(n41995) );
  XOR U43069 ( .A(n41996), .B(n41995), .Z(n41991) );
  XOR U43070 ( .A(n41992), .B(n41991), .Z(c[2040]) );
  AND U43071 ( .A(n41992), .B(n41991), .Z(n42028) );
  NAND U43072 ( .A(n41994), .B(n41993), .Z(n41998) );
  NANDN U43073 ( .A(n41996), .B(n41995), .Z(n41997) );
  AND U43074 ( .A(n41998), .B(n41997), .Z(n42032) );
  NAND U43075 ( .A(n42000), .B(n41999), .Z(n42004) );
  NAND U43076 ( .A(n42002), .B(n42001), .Z(n42003) );
  NAND U43077 ( .A(n42004), .B(n42003), .Z(n42038) );
  NAND U43078 ( .A(n42143), .B(n42005), .Z(n42007) );
  XNOR U43079 ( .A(a[1019]), .B(n4217), .Z(n42050) );
  NAND U43080 ( .A(n42144), .B(n42050), .Z(n42006) );
  NAND U43081 ( .A(n42007), .B(n42006), .Z(n42058) );
  AND U43082 ( .A(a[1017]), .B(b[7]), .Z(n42122) );
  XNOR U43083 ( .A(a[1021]), .B(n42085), .Z(n42053) );
  NANDN U43084 ( .A(n4065), .B(n42053), .Z(n42010) );
  NAND U43085 ( .A(n42008), .B(n42115), .Z(n42009) );
  NAND U43086 ( .A(n42010), .B(n42009), .Z(n42056) );
  XNOR U43087 ( .A(n42122), .B(n42056), .Z(n42057) );
  OR U43088 ( .A(n42011), .B(n4066), .Z(n42014) );
  XNOR U43089 ( .A(a[1023]), .B(n42012), .Z(n42046) );
  NANDN U43090 ( .A(n4064), .B(n42046), .Z(n42013) );
  AND U43091 ( .A(n42014), .B(n42013), .Z(n42041) );
  XOR U43092 ( .A(b[1]), .B(n42041), .Z(n42043) );
  XNOR U43093 ( .A(n42042), .B(n42043), .Z(n42036) );
  NAND U43094 ( .A(n42016), .B(n42015), .Z(n42020) );
  NAND U43095 ( .A(n42018), .B(n42017), .Z(n42019) );
  NAND U43096 ( .A(n42020), .B(n42019), .Z(n42035) );
  XOR U43097 ( .A(n42036), .B(n42035), .Z(n42037) );
  NAND U43098 ( .A(n42022), .B(n42021), .Z(n42026) );
  NAND U43099 ( .A(n42024), .B(n42023), .Z(n42025) );
  AND U43100 ( .A(n42026), .B(n42025), .Z(n42030) );
  XOR U43101 ( .A(n42029), .B(n42030), .Z(n42031) );
  XOR U43102 ( .A(n42032), .B(n42031), .Z(n42027) );
  XOR U43103 ( .A(n42028), .B(n42027), .Z(c[2041]) );
  AND U43104 ( .A(n42028), .B(n42027), .Z(n42062) );
  NAND U43105 ( .A(n42030), .B(n42029), .Z(n42034) );
  NANDN U43106 ( .A(n42032), .B(n42031), .Z(n42033) );
  AND U43107 ( .A(n42034), .B(n42033), .Z(n42066) );
  NAND U43108 ( .A(n42036), .B(n42035), .Z(n42040) );
  NAND U43109 ( .A(n42038), .B(n42037), .Z(n42039) );
  AND U43110 ( .A(n42040), .B(n42039), .Z(n42064) );
  NAND U43111 ( .A(b[1]), .B(n42041), .Z(n42045) );
  NAND U43112 ( .A(n42043), .B(n42042), .Z(n42044) );
  NAND U43113 ( .A(n42045), .B(n42044), .Z(n42072) );
  NAND U43114 ( .A(n42047), .B(n42046), .Z(n42049) );
  NAND U43115 ( .A(n4067), .B(b[3]), .Z(n42048) );
  NAND U43116 ( .A(n42049), .B(n42048), .Z(n42089) );
  AND U43117 ( .A(a[1018]), .B(b[7]), .Z(n42088) );
  XNOR U43118 ( .A(n42122), .B(n42090), .Z(n42077) );
  NAND U43119 ( .A(n42143), .B(n42050), .Z(n42052) );
  XNOR U43120 ( .A(a[1020]), .B(n4217), .Z(n42081) );
  NAND U43121 ( .A(n42144), .B(n42081), .Z(n42051) );
  NAND U43122 ( .A(n42052), .B(n42051), .Z(n42075) );
  XNOR U43123 ( .A(a[1022]), .B(n42085), .Z(n42084) );
  NANDN U43124 ( .A(n4065), .B(n42084), .Z(n42055) );
  NAND U43125 ( .A(n42053), .B(n42115), .Z(n42054) );
  AND U43126 ( .A(n42055), .B(n42054), .Z(n42076) );
  XOR U43127 ( .A(n42075), .B(n42076), .Z(n42078) );
  XOR U43128 ( .A(n42077), .B(n42078), .Z(n42069) );
  IV U43129 ( .A(n42122), .Z(n42091) );
  NAND U43130 ( .A(n42091), .B(n42056), .Z(n42060) );
  NAND U43131 ( .A(n42058), .B(n42057), .Z(n42059) );
  AND U43132 ( .A(n42060), .B(n42059), .Z(n42070) );
  XOR U43133 ( .A(n42069), .B(n42070), .Z(n42071) );
  XOR U43134 ( .A(n42064), .B(n42063), .Z(n42065) );
  XOR U43135 ( .A(n42066), .B(n42065), .Z(n42061) );
  XOR U43136 ( .A(n42062), .B(n42061), .Z(c[2042]) );
  AND U43137 ( .A(n42062), .B(n42061), .Z(n42095) );
  NAND U43138 ( .A(n42064), .B(n42063), .Z(n42068) );
  NANDN U43139 ( .A(n42066), .B(n42065), .Z(n42067) );
  AND U43140 ( .A(n42068), .B(n42067), .Z(n42099) );
  NAND U43141 ( .A(n42070), .B(n42069), .Z(n42074) );
  NAND U43142 ( .A(n42072), .B(n42071), .Z(n42073) );
  NAND U43143 ( .A(n42074), .B(n42073), .Z(n42097) );
  NANDN U43144 ( .A(n42076), .B(n42075), .Z(n42080) );
  NANDN U43145 ( .A(n42078), .B(n42077), .Z(n42079) );
  AND U43146 ( .A(n42080), .B(n42079), .Z(n42105) );
  NAND U43147 ( .A(n42143), .B(n42081), .Z(n42083) );
  XNOR U43148 ( .A(a[1021]), .B(n4217), .Z(n42118) );
  NAND U43149 ( .A(n42144), .B(n42118), .Z(n42082) );
  NAND U43150 ( .A(n42083), .B(n42082), .Z(n42109) );
  NAND U43151 ( .A(n42084), .B(n42115), .Z(n42087) );
  XNOR U43152 ( .A(a[1023]), .B(n42085), .Z(n42114) );
  NANDN U43153 ( .A(n4065), .B(n42114), .Z(n42086) );
  NAND U43154 ( .A(n42087), .B(n42086), .Z(n42108) );
  AND U43155 ( .A(a[1019]), .B(b[7]), .Z(n42121) );
  XNOR U43156 ( .A(n42091), .B(n42121), .Z(n42123) );
  XNOR U43157 ( .A(n42124), .B(n42123), .Z(n42110) );
  XNOR U43158 ( .A(n42111), .B(n42110), .Z(n42103) );
  NAND U43159 ( .A(n42089), .B(n42088), .Z(n42093) );
  NAND U43160 ( .A(n42091), .B(n42090), .Z(n42092) );
  AND U43161 ( .A(n42093), .B(n42092), .Z(n42102) );
  XOR U43162 ( .A(n42105), .B(n42104), .Z(n42096) );
  XOR U43163 ( .A(n42099), .B(n42098), .Z(n42094) );
  XOR U43164 ( .A(n42095), .B(n42094), .Z(c[2043]) );
  AND U43165 ( .A(n42095), .B(n42094), .Z(n42128) );
  NAND U43166 ( .A(n42097), .B(n42096), .Z(n42101) );
  NANDN U43167 ( .A(n42099), .B(n42098), .Z(n42100) );
  AND U43168 ( .A(n42101), .B(n42100), .Z(n42132) );
  NAND U43169 ( .A(n42103), .B(n42102), .Z(n42107) );
  NAND U43170 ( .A(n42105), .B(n42104), .Z(n42106) );
  NAND U43171 ( .A(n42107), .B(n42106), .Z(n42130) );
  NAND U43172 ( .A(n42109), .B(n42108), .Z(n42113) );
  NAND U43173 ( .A(n42111), .B(n42110), .Z(n42112) );
  AND U43174 ( .A(n42113), .B(n42112), .Z(n42138) );
  AND U43175 ( .A(a[1020]), .B(b[7]), .Z(n42156) );
  NAND U43176 ( .A(n42115), .B(n42114), .Z(n42117) );
  NAND U43177 ( .A(n4068), .B(b[5]), .Z(n42116) );
  NAND U43178 ( .A(n42117), .B(n42116), .Z(n42147) );
  XNOR U43179 ( .A(n42156), .B(n42147), .Z(n42149) );
  NAND U43180 ( .A(n42143), .B(n42118), .Z(n42120) );
  XNOR U43181 ( .A(a[1022]), .B(n4217), .Z(n42142) );
  NAND U43182 ( .A(n42144), .B(n42142), .Z(n42119) );
  NAND U43183 ( .A(n42120), .B(n42119), .Z(n42148) );
  XNOR U43184 ( .A(n42149), .B(n42148), .Z(n42136) );
  NAND U43185 ( .A(n42122), .B(n42121), .Z(n42126) );
  NANDN U43186 ( .A(n42124), .B(n42123), .Z(n42125) );
  AND U43187 ( .A(n42126), .B(n42125), .Z(n42135) );
  XOR U43188 ( .A(n42138), .B(n42137), .Z(n42129) );
  XOR U43189 ( .A(n42132), .B(n42131), .Z(n42127) );
  XOR U43190 ( .A(n42128), .B(n42127), .Z(c[2044]) );
  AND U43191 ( .A(n42128), .B(n42127), .Z(n42153) );
  NAND U43192 ( .A(n42130), .B(n42129), .Z(n42134) );
  NANDN U43193 ( .A(n42132), .B(n42131), .Z(n42133) );
  AND U43194 ( .A(n42134), .B(n42133), .Z(n42166) );
  NAND U43195 ( .A(n42136), .B(n42135), .Z(n42140) );
  NAND U43196 ( .A(n42138), .B(n42137), .Z(n42139) );
  NAND U43197 ( .A(n42140), .B(n42139), .Z(n42164) );
  AND U43198 ( .A(a[1021]), .B(b[7]), .Z(n42155) );
  XOR U43199 ( .A(n42141), .B(n42155), .Z(n42157) );
  XNOR U43200 ( .A(n42156), .B(n42157), .Z(n42169) );
  NAND U43201 ( .A(n42143), .B(n42142), .Z(n42146) );
  NAND U43202 ( .A(n42144), .B(n42160), .Z(n42145) );
  NAND U43203 ( .A(n42146), .B(n42145), .Z(n42170) );
  NANDN U43204 ( .A(n42156), .B(n42147), .Z(n42151) );
  NAND U43205 ( .A(n42149), .B(n42148), .Z(n42150) );
  NAND U43206 ( .A(n42151), .B(n42150), .Z(n42171) );
  XNOR U43207 ( .A(n42172), .B(n42171), .Z(n42163) );
  XOR U43208 ( .A(n42166), .B(n42165), .Z(n42152) );
  XOR U43209 ( .A(n42153), .B(n42152), .Z(c[2045]) );
  AND U43210 ( .A(n42153), .B(n42152), .Z(n42176) );
  AND U43211 ( .A(n42155), .B(n42154), .Z(n42159) );
  NANDN U43212 ( .A(n42157), .B(n42156), .Z(n42158) );
  NANDN U43213 ( .A(n42159), .B(n42158), .Z(n42191) );
  AND U43214 ( .A(a[1022]), .B(b[7]), .Z(n42189) );
  NANDN U43215 ( .A(n4069), .B(n42160), .Z(n42162) );
  NANDN U43216 ( .A(n4070), .B(b[7]), .Z(n42161) );
  AND U43217 ( .A(n42162), .B(n42161), .Z(n42188) );
  XOR U43218 ( .A(n42189), .B(n42188), .Z(n42190) );
  NAND U43219 ( .A(n42164), .B(n42163), .Z(n42168) );
  NANDN U43220 ( .A(n42166), .B(n42165), .Z(n42167) );
  NAND U43221 ( .A(n42168), .B(n42167), .Z(n42177) );
  NAND U43222 ( .A(n42170), .B(n42169), .Z(n42174) );
  NAND U43223 ( .A(n42172), .B(n42171), .Z(n42173) );
  AND U43224 ( .A(n42174), .B(n42173), .Z(n42178) );
  XNOR U43225 ( .A(n42179), .B(n42180), .Z(n42175) );
  XOR U43226 ( .A(n42176), .B(n42175), .Z(c[2046]) );
  NAND U43227 ( .A(n42176), .B(n42175), .Z(n42184) );
  AND U43228 ( .A(n42178), .B(n42177), .Z(n42182) );
  AND U43229 ( .A(n42180), .B(n42179), .Z(n42181) );
  OR U43230 ( .A(n42182), .B(n42181), .Z(n42183) );
  AND U43231 ( .A(n42184), .B(n42183), .Z(n42197) );
  XNOR U43232 ( .A(a[1022]), .B(a[1023]), .Z(n42185) );
  XNOR U43233 ( .A(n42186), .B(n42185), .Z(n42187) );
  ANDN U43234 ( .B(b[7]), .A(n42187), .Z(n42195) );
  NOR U43235 ( .A(n42189), .B(n42188), .Z(n42193) );
  AND U43236 ( .A(n42191), .B(n42190), .Z(n42192) );
  OR U43237 ( .A(n42193), .B(n42192), .Z(n42194) );
  XNOR U43238 ( .A(n42195), .B(n42194), .Z(n42196) );
  XNOR U43239 ( .A(n42197), .B(n42196), .Z(c[2047]) );
endmodule

