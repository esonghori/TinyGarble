
module modexp_2N_NN_N1024_CC2097152 ( clk, rst, m, e, n, c );
  input [1023:0] m;
  input [1023:0] e;
  input [1023:0] n;
  output [1023:0] c;
  input clk, rst;
  wire   first_one, mul_pow, n6, n8, \modmult_1/xin[1023] ,
         \modmult_1/xin[1022] , \modmult_1/xin[1021] , \modmult_1/xin[1020] ,
         \modmult_1/xin[1019] , \modmult_1/xin[1018] , \modmult_1/xin[1017] ,
         \modmult_1/xin[1016] , \modmult_1/xin[1015] , \modmult_1/xin[1014] ,
         \modmult_1/xin[1013] , \modmult_1/xin[1012] , \modmult_1/xin[1011] ,
         \modmult_1/xin[1010] , \modmult_1/xin[1009] , \modmult_1/xin[1008] ,
         \modmult_1/xin[1007] , \modmult_1/xin[1006] , \modmult_1/xin[1005] ,
         \modmult_1/xin[1004] , \modmult_1/xin[1003] , \modmult_1/xin[1002] ,
         \modmult_1/xin[1001] , \modmult_1/xin[1000] , \modmult_1/xin[999] ,
         \modmult_1/xin[998] , \modmult_1/xin[997] , \modmult_1/xin[996] ,
         \modmult_1/xin[995] , \modmult_1/xin[994] , \modmult_1/xin[993] ,
         \modmult_1/xin[992] , \modmult_1/xin[991] , \modmult_1/xin[990] ,
         \modmult_1/xin[989] , \modmult_1/xin[988] , \modmult_1/xin[987] ,
         \modmult_1/xin[986] , \modmult_1/xin[985] , \modmult_1/xin[984] ,
         \modmult_1/xin[983] , \modmult_1/xin[982] , \modmult_1/xin[981] ,
         \modmult_1/xin[980] , \modmult_1/xin[979] , \modmult_1/xin[978] ,
         \modmult_1/xin[977] , \modmult_1/xin[976] , \modmult_1/xin[975] ,
         \modmult_1/xin[974] , \modmult_1/xin[973] , \modmult_1/xin[972] ,
         \modmult_1/xin[971] , \modmult_1/xin[970] , \modmult_1/xin[969] ,
         \modmult_1/xin[968] , \modmult_1/xin[967] , \modmult_1/xin[966] ,
         \modmult_1/xin[965] , \modmult_1/xin[964] , \modmult_1/xin[963] ,
         \modmult_1/xin[962] , \modmult_1/xin[961] , \modmult_1/xin[960] ,
         \modmult_1/xin[959] , \modmult_1/xin[958] , \modmult_1/xin[957] ,
         \modmult_1/xin[956] , \modmult_1/xin[955] , \modmult_1/xin[954] ,
         \modmult_1/xin[953] , \modmult_1/xin[952] , \modmult_1/xin[951] ,
         \modmult_1/xin[950] , \modmult_1/xin[949] , \modmult_1/xin[948] ,
         \modmult_1/xin[947] , \modmult_1/xin[946] , \modmult_1/xin[945] ,
         \modmult_1/xin[944] , \modmult_1/xin[943] , \modmult_1/xin[942] ,
         \modmult_1/xin[941] , \modmult_1/xin[940] , \modmult_1/xin[939] ,
         \modmult_1/xin[938] , \modmult_1/xin[937] , \modmult_1/xin[936] ,
         \modmult_1/xin[935] , \modmult_1/xin[934] , \modmult_1/xin[933] ,
         \modmult_1/xin[932] , \modmult_1/xin[931] , \modmult_1/xin[930] ,
         \modmult_1/xin[929] , \modmult_1/xin[928] , \modmult_1/xin[927] ,
         \modmult_1/xin[926] , \modmult_1/xin[925] , \modmult_1/xin[924] ,
         \modmult_1/xin[923] , \modmult_1/xin[922] , \modmult_1/xin[921] ,
         \modmult_1/xin[920] , \modmult_1/xin[919] , \modmult_1/xin[918] ,
         \modmult_1/xin[917] , \modmult_1/xin[916] , \modmult_1/xin[915] ,
         \modmult_1/xin[914] , \modmult_1/xin[913] , \modmult_1/xin[912] ,
         \modmult_1/xin[911] , \modmult_1/xin[910] , \modmult_1/xin[909] ,
         \modmult_1/xin[908] , \modmult_1/xin[907] , \modmult_1/xin[906] ,
         \modmult_1/xin[905] , \modmult_1/xin[904] , \modmult_1/xin[903] ,
         \modmult_1/xin[902] , \modmult_1/xin[901] , \modmult_1/xin[900] ,
         \modmult_1/xin[899] , \modmult_1/xin[898] , \modmult_1/xin[897] ,
         \modmult_1/xin[896] , \modmult_1/xin[895] , \modmult_1/xin[894] ,
         \modmult_1/xin[893] , \modmult_1/xin[892] , \modmult_1/xin[891] ,
         \modmult_1/xin[890] , \modmult_1/xin[889] , \modmult_1/xin[888] ,
         \modmult_1/xin[887] , \modmult_1/xin[886] , \modmult_1/xin[885] ,
         \modmult_1/xin[884] , \modmult_1/xin[883] , \modmult_1/xin[882] ,
         \modmult_1/xin[881] , \modmult_1/xin[880] , \modmult_1/xin[879] ,
         \modmult_1/xin[878] , \modmult_1/xin[877] , \modmult_1/xin[876] ,
         \modmult_1/xin[875] , \modmult_1/xin[874] , \modmult_1/xin[873] ,
         \modmult_1/xin[872] , \modmult_1/xin[871] , \modmult_1/xin[870] ,
         \modmult_1/xin[869] , \modmult_1/xin[868] , \modmult_1/xin[867] ,
         \modmult_1/xin[866] , \modmult_1/xin[865] , \modmult_1/xin[864] ,
         \modmult_1/xin[863] , \modmult_1/xin[862] , \modmult_1/xin[861] ,
         \modmult_1/xin[860] , \modmult_1/xin[859] , \modmult_1/xin[858] ,
         \modmult_1/xin[857] , \modmult_1/xin[856] , \modmult_1/xin[855] ,
         \modmult_1/xin[854] , \modmult_1/xin[853] , \modmult_1/xin[852] ,
         \modmult_1/xin[851] , \modmult_1/xin[850] , \modmult_1/xin[849] ,
         \modmult_1/xin[848] , \modmult_1/xin[847] , \modmult_1/xin[846] ,
         \modmult_1/xin[845] , \modmult_1/xin[844] , \modmult_1/xin[843] ,
         \modmult_1/xin[842] , \modmult_1/xin[841] , \modmult_1/xin[840] ,
         \modmult_1/xin[839] , \modmult_1/xin[838] , \modmult_1/xin[837] ,
         \modmult_1/xin[836] , \modmult_1/xin[835] , \modmult_1/xin[834] ,
         \modmult_1/xin[833] , \modmult_1/xin[832] , \modmult_1/xin[831] ,
         \modmult_1/xin[830] , \modmult_1/xin[829] , \modmult_1/xin[828] ,
         \modmult_1/xin[827] , \modmult_1/xin[826] , \modmult_1/xin[825] ,
         \modmult_1/xin[824] , \modmult_1/xin[823] , \modmult_1/xin[822] ,
         \modmult_1/xin[821] , \modmult_1/xin[820] , \modmult_1/xin[819] ,
         \modmult_1/xin[818] , \modmult_1/xin[817] , \modmult_1/xin[816] ,
         \modmult_1/xin[815] , \modmult_1/xin[814] , \modmult_1/xin[813] ,
         \modmult_1/xin[812] , \modmult_1/xin[811] , \modmult_1/xin[810] ,
         \modmult_1/xin[809] , \modmult_1/xin[808] , \modmult_1/xin[807] ,
         \modmult_1/xin[806] , \modmult_1/xin[805] , \modmult_1/xin[804] ,
         \modmult_1/xin[803] , \modmult_1/xin[802] , \modmult_1/xin[801] ,
         \modmult_1/xin[800] , \modmult_1/xin[799] , \modmult_1/xin[798] ,
         \modmult_1/xin[797] , \modmult_1/xin[796] , \modmult_1/xin[795] ,
         \modmult_1/xin[794] , \modmult_1/xin[793] , \modmult_1/xin[792] ,
         \modmult_1/xin[791] , \modmult_1/xin[790] , \modmult_1/xin[789] ,
         \modmult_1/xin[788] , \modmult_1/xin[787] , \modmult_1/xin[786] ,
         \modmult_1/xin[785] , \modmult_1/xin[784] , \modmult_1/xin[783] ,
         \modmult_1/xin[782] , \modmult_1/xin[781] , \modmult_1/xin[780] ,
         \modmult_1/xin[779] , \modmult_1/xin[778] , \modmult_1/xin[777] ,
         \modmult_1/xin[776] , \modmult_1/xin[775] , \modmult_1/xin[774] ,
         \modmult_1/xin[773] , \modmult_1/xin[772] , \modmult_1/xin[771] ,
         \modmult_1/xin[770] , \modmult_1/xin[769] , \modmult_1/xin[768] ,
         \modmult_1/xin[767] , \modmult_1/xin[766] , \modmult_1/xin[765] ,
         \modmult_1/xin[764] , \modmult_1/xin[763] , \modmult_1/xin[762] ,
         \modmult_1/xin[761] , \modmult_1/xin[760] , \modmult_1/xin[759] ,
         \modmult_1/xin[758] , \modmult_1/xin[757] , \modmult_1/xin[756] ,
         \modmult_1/xin[755] , \modmult_1/xin[754] , \modmult_1/xin[753] ,
         \modmult_1/xin[752] , \modmult_1/xin[751] , \modmult_1/xin[750] ,
         \modmult_1/xin[749] , \modmult_1/xin[748] , \modmult_1/xin[747] ,
         \modmult_1/xin[746] , \modmult_1/xin[745] , \modmult_1/xin[744] ,
         \modmult_1/xin[743] , \modmult_1/xin[742] , \modmult_1/xin[741] ,
         \modmult_1/xin[740] , \modmult_1/xin[739] , \modmult_1/xin[738] ,
         \modmult_1/xin[737] , \modmult_1/xin[736] , \modmult_1/xin[735] ,
         \modmult_1/xin[734] , \modmult_1/xin[733] , \modmult_1/xin[732] ,
         \modmult_1/xin[731] , \modmult_1/xin[730] , \modmult_1/xin[729] ,
         \modmult_1/xin[728] , \modmult_1/xin[727] , \modmult_1/xin[726] ,
         \modmult_1/xin[725] , \modmult_1/xin[724] , \modmult_1/xin[723] ,
         \modmult_1/xin[722] , \modmult_1/xin[721] , \modmult_1/xin[720] ,
         \modmult_1/xin[719] , \modmult_1/xin[718] , \modmult_1/xin[717] ,
         \modmult_1/xin[716] , \modmult_1/xin[715] , \modmult_1/xin[714] ,
         \modmult_1/xin[713] , \modmult_1/xin[712] , \modmult_1/xin[711] ,
         \modmult_1/xin[710] , \modmult_1/xin[709] , \modmult_1/xin[708] ,
         \modmult_1/xin[707] , \modmult_1/xin[706] , \modmult_1/xin[705] ,
         \modmult_1/xin[704] , \modmult_1/xin[703] , \modmult_1/xin[702] ,
         \modmult_1/xin[701] , \modmult_1/xin[700] , \modmult_1/xin[699] ,
         \modmult_1/xin[698] , \modmult_1/xin[697] , \modmult_1/xin[696] ,
         \modmult_1/xin[695] , \modmult_1/xin[694] , \modmult_1/xin[693] ,
         \modmult_1/xin[692] , \modmult_1/xin[691] , \modmult_1/xin[690] ,
         \modmult_1/xin[689] , \modmult_1/xin[688] , \modmult_1/xin[687] ,
         \modmult_1/xin[686] , \modmult_1/xin[685] , \modmult_1/xin[684] ,
         \modmult_1/xin[683] , \modmult_1/xin[682] , \modmult_1/xin[681] ,
         \modmult_1/xin[680] , \modmult_1/xin[679] , \modmult_1/xin[678] ,
         \modmult_1/xin[677] , \modmult_1/xin[676] , \modmult_1/xin[675] ,
         \modmult_1/xin[674] , \modmult_1/xin[673] , \modmult_1/xin[672] ,
         \modmult_1/xin[671] , \modmult_1/xin[670] , \modmult_1/xin[669] ,
         \modmult_1/xin[668] , \modmult_1/xin[667] , \modmult_1/xin[666] ,
         \modmult_1/xin[665] , \modmult_1/xin[664] , \modmult_1/xin[663] ,
         \modmult_1/xin[662] , \modmult_1/xin[661] , \modmult_1/xin[660] ,
         \modmult_1/xin[659] , \modmult_1/xin[658] , \modmult_1/xin[657] ,
         \modmult_1/xin[656] , \modmult_1/xin[655] , \modmult_1/xin[654] ,
         \modmult_1/xin[653] , \modmult_1/xin[652] , \modmult_1/xin[651] ,
         \modmult_1/xin[650] , \modmult_1/xin[649] , \modmult_1/xin[648] ,
         \modmult_1/xin[647] , \modmult_1/xin[646] , \modmult_1/xin[645] ,
         \modmult_1/xin[644] , \modmult_1/xin[643] , \modmult_1/xin[642] ,
         \modmult_1/xin[641] , \modmult_1/xin[640] , \modmult_1/xin[639] ,
         \modmult_1/xin[638] , \modmult_1/xin[637] , \modmult_1/xin[636] ,
         \modmult_1/xin[635] , \modmult_1/xin[634] , \modmult_1/xin[633] ,
         \modmult_1/xin[632] , \modmult_1/xin[631] , \modmult_1/xin[630] ,
         \modmult_1/xin[629] , \modmult_1/xin[628] , \modmult_1/xin[627] ,
         \modmult_1/xin[626] , \modmult_1/xin[625] , \modmult_1/xin[624] ,
         \modmult_1/xin[623] , \modmult_1/xin[622] , \modmult_1/xin[621] ,
         \modmult_1/xin[620] , \modmult_1/xin[619] , \modmult_1/xin[618] ,
         \modmult_1/xin[617] , \modmult_1/xin[616] , \modmult_1/xin[615] ,
         \modmult_1/xin[614] , \modmult_1/xin[613] , \modmult_1/xin[612] ,
         \modmult_1/xin[611] , \modmult_1/xin[610] , \modmult_1/xin[609] ,
         \modmult_1/xin[608] , \modmult_1/xin[607] , \modmult_1/xin[606] ,
         \modmult_1/xin[605] , \modmult_1/xin[604] , \modmult_1/xin[603] ,
         \modmult_1/xin[602] , \modmult_1/xin[601] , \modmult_1/xin[600] ,
         \modmult_1/xin[599] , \modmult_1/xin[598] , \modmult_1/xin[597] ,
         \modmult_1/xin[596] , \modmult_1/xin[595] , \modmult_1/xin[594] ,
         \modmult_1/xin[593] , \modmult_1/xin[592] , \modmult_1/xin[591] ,
         \modmult_1/xin[590] , \modmult_1/xin[589] , \modmult_1/xin[588] ,
         \modmult_1/xin[587] , \modmult_1/xin[586] , \modmult_1/xin[585] ,
         \modmult_1/xin[584] , \modmult_1/xin[583] , \modmult_1/xin[582] ,
         \modmult_1/xin[581] , \modmult_1/xin[580] , \modmult_1/xin[579] ,
         \modmult_1/xin[578] , \modmult_1/xin[577] , \modmult_1/xin[576] ,
         \modmult_1/xin[575] , \modmult_1/xin[574] , \modmult_1/xin[573] ,
         \modmult_1/xin[572] , \modmult_1/xin[571] , \modmult_1/xin[570] ,
         \modmult_1/xin[569] , \modmult_1/xin[568] , \modmult_1/xin[567] ,
         \modmult_1/xin[566] , \modmult_1/xin[565] , \modmult_1/xin[564] ,
         \modmult_1/xin[563] , \modmult_1/xin[562] , \modmult_1/xin[561] ,
         \modmult_1/xin[560] , \modmult_1/xin[559] , \modmult_1/xin[558] ,
         \modmult_1/xin[557] , \modmult_1/xin[556] , \modmult_1/xin[555] ,
         \modmult_1/xin[554] , \modmult_1/xin[553] , \modmult_1/xin[552] ,
         \modmult_1/xin[551] , \modmult_1/xin[550] , \modmult_1/xin[549] ,
         \modmult_1/xin[548] , \modmult_1/xin[547] , \modmult_1/xin[546] ,
         \modmult_1/xin[545] , \modmult_1/xin[544] , \modmult_1/xin[543] ,
         \modmult_1/xin[542] , \modmult_1/xin[541] , \modmult_1/xin[540] ,
         \modmult_1/xin[539] , \modmult_1/xin[538] , \modmult_1/xin[537] ,
         \modmult_1/xin[536] , \modmult_1/xin[535] , \modmult_1/xin[534] ,
         \modmult_1/xin[533] , \modmult_1/xin[532] , \modmult_1/xin[531] ,
         \modmult_1/xin[530] , \modmult_1/xin[529] , \modmult_1/xin[528] ,
         \modmult_1/xin[527] , \modmult_1/xin[526] , \modmult_1/xin[525] ,
         \modmult_1/xin[524] , \modmult_1/xin[523] , \modmult_1/xin[522] ,
         \modmult_1/xin[521] , \modmult_1/xin[520] , \modmult_1/xin[519] ,
         \modmult_1/xin[518] , \modmult_1/xin[517] , \modmult_1/xin[516] ,
         \modmult_1/xin[515] , \modmult_1/xin[514] , \modmult_1/xin[513] ,
         \modmult_1/xin[512] , \modmult_1/xin[511] , \modmult_1/xin[510] ,
         \modmult_1/xin[509] , \modmult_1/xin[508] , \modmult_1/xin[507] ,
         \modmult_1/xin[506] , \modmult_1/xin[505] , \modmult_1/xin[504] ,
         \modmult_1/xin[503] , \modmult_1/xin[502] , \modmult_1/xin[501] ,
         \modmult_1/xin[500] , \modmult_1/xin[499] , \modmult_1/xin[498] ,
         \modmult_1/xin[497] , \modmult_1/xin[496] , \modmult_1/xin[495] ,
         \modmult_1/xin[494] , \modmult_1/xin[493] , \modmult_1/xin[492] ,
         \modmult_1/xin[491] , \modmult_1/xin[490] , \modmult_1/xin[489] ,
         \modmult_1/xin[488] , \modmult_1/xin[487] , \modmult_1/xin[486] ,
         \modmult_1/xin[485] , \modmult_1/xin[484] , \modmult_1/xin[483] ,
         \modmult_1/xin[482] , \modmult_1/xin[481] , \modmult_1/xin[480] ,
         \modmult_1/xin[479] , \modmult_1/xin[478] , \modmult_1/xin[477] ,
         \modmult_1/xin[476] , \modmult_1/xin[475] , \modmult_1/xin[474] ,
         \modmult_1/xin[473] , \modmult_1/xin[472] , \modmult_1/xin[471] ,
         \modmult_1/xin[470] , \modmult_1/xin[469] , \modmult_1/xin[468] ,
         \modmult_1/xin[467] , \modmult_1/xin[466] , \modmult_1/xin[465] ,
         \modmult_1/xin[464] , \modmult_1/xin[463] , \modmult_1/xin[462] ,
         \modmult_1/xin[461] , \modmult_1/xin[460] , \modmult_1/xin[459] ,
         \modmult_1/xin[458] , \modmult_1/xin[457] , \modmult_1/xin[456] ,
         \modmult_1/xin[455] , \modmult_1/xin[454] , \modmult_1/xin[453] ,
         \modmult_1/xin[452] , \modmult_1/xin[451] , \modmult_1/xin[450] ,
         \modmult_1/xin[449] , \modmult_1/xin[448] , \modmult_1/xin[447] ,
         \modmult_1/xin[446] , \modmult_1/xin[445] , \modmult_1/xin[444] ,
         \modmult_1/xin[443] , \modmult_1/xin[442] , \modmult_1/xin[441] ,
         \modmult_1/xin[440] , \modmult_1/xin[439] , \modmult_1/xin[438] ,
         \modmult_1/xin[437] , \modmult_1/xin[436] , \modmult_1/xin[435] ,
         \modmult_1/xin[434] , \modmult_1/xin[433] , \modmult_1/xin[432] ,
         \modmult_1/xin[431] , \modmult_1/xin[430] , \modmult_1/xin[429] ,
         \modmult_1/xin[428] , \modmult_1/xin[427] , \modmult_1/xin[426] ,
         \modmult_1/xin[425] , \modmult_1/xin[424] , \modmult_1/xin[423] ,
         \modmult_1/xin[422] , \modmult_1/xin[421] , \modmult_1/xin[420] ,
         \modmult_1/xin[419] , \modmult_1/xin[418] , \modmult_1/xin[417] ,
         \modmult_1/xin[416] , \modmult_1/xin[415] , \modmult_1/xin[414] ,
         \modmult_1/xin[413] , \modmult_1/xin[412] , \modmult_1/xin[411] ,
         \modmult_1/xin[410] , \modmult_1/xin[409] , \modmult_1/xin[408] ,
         \modmult_1/xin[407] , \modmult_1/xin[406] , \modmult_1/xin[405] ,
         \modmult_1/xin[404] , \modmult_1/xin[403] , \modmult_1/xin[402] ,
         \modmult_1/xin[401] , \modmult_1/xin[400] , \modmult_1/xin[399] ,
         \modmult_1/xin[398] , \modmult_1/xin[397] , \modmult_1/xin[396] ,
         \modmult_1/xin[395] , \modmult_1/xin[394] , \modmult_1/xin[393] ,
         \modmult_1/xin[392] , \modmult_1/xin[391] , \modmult_1/xin[390] ,
         \modmult_1/xin[389] , \modmult_1/xin[388] , \modmult_1/xin[387] ,
         \modmult_1/xin[386] , \modmult_1/xin[385] , \modmult_1/xin[384] ,
         \modmult_1/xin[383] , \modmult_1/xin[382] , \modmult_1/xin[381] ,
         \modmult_1/xin[380] , \modmult_1/xin[379] , \modmult_1/xin[378] ,
         \modmult_1/xin[377] , \modmult_1/xin[376] , \modmult_1/xin[375] ,
         \modmult_1/xin[374] , \modmult_1/xin[373] , \modmult_1/xin[372] ,
         \modmult_1/xin[371] , \modmult_1/xin[370] , \modmult_1/xin[369] ,
         \modmult_1/xin[368] , \modmult_1/xin[367] , \modmult_1/xin[366] ,
         \modmult_1/xin[365] , \modmult_1/xin[364] , \modmult_1/xin[363] ,
         \modmult_1/xin[362] , \modmult_1/xin[361] , \modmult_1/xin[360] ,
         \modmult_1/xin[359] , \modmult_1/xin[358] , \modmult_1/xin[357] ,
         \modmult_1/xin[356] , \modmult_1/xin[355] , \modmult_1/xin[354] ,
         \modmult_1/xin[353] , \modmult_1/xin[352] , \modmult_1/xin[351] ,
         \modmult_1/xin[350] , \modmult_1/xin[349] , \modmult_1/xin[348] ,
         \modmult_1/xin[347] , \modmult_1/xin[346] , \modmult_1/xin[345] ,
         \modmult_1/xin[344] , \modmult_1/xin[343] , \modmult_1/xin[342] ,
         \modmult_1/xin[341] , \modmult_1/xin[340] , \modmult_1/xin[339] ,
         \modmult_1/xin[338] , \modmult_1/xin[337] , \modmult_1/xin[336] ,
         \modmult_1/xin[335] , \modmult_1/xin[334] , \modmult_1/xin[333] ,
         \modmult_1/xin[332] , \modmult_1/xin[331] , \modmult_1/xin[330] ,
         \modmult_1/xin[329] , \modmult_1/xin[328] , \modmult_1/xin[327] ,
         \modmult_1/xin[326] , \modmult_1/xin[325] , \modmult_1/xin[324] ,
         \modmult_1/xin[323] , \modmult_1/xin[322] , \modmult_1/xin[321] ,
         \modmult_1/xin[320] , \modmult_1/xin[319] , \modmult_1/xin[318] ,
         \modmult_1/xin[317] , \modmult_1/xin[316] , \modmult_1/xin[315] ,
         \modmult_1/xin[314] , \modmult_1/xin[313] , \modmult_1/xin[312] ,
         \modmult_1/xin[311] , \modmult_1/xin[310] , \modmult_1/xin[309] ,
         \modmult_1/xin[308] , \modmult_1/xin[307] , \modmult_1/xin[306] ,
         \modmult_1/xin[305] , \modmult_1/xin[304] , \modmult_1/xin[303] ,
         \modmult_1/xin[302] , \modmult_1/xin[301] , \modmult_1/xin[300] ,
         \modmult_1/xin[299] , \modmult_1/xin[298] , \modmult_1/xin[297] ,
         \modmult_1/xin[296] , \modmult_1/xin[295] , \modmult_1/xin[294] ,
         \modmult_1/xin[293] , \modmult_1/xin[292] , \modmult_1/xin[291] ,
         \modmult_1/xin[290] , \modmult_1/xin[289] , \modmult_1/xin[288] ,
         \modmult_1/xin[287] , \modmult_1/xin[286] , \modmult_1/xin[285] ,
         \modmult_1/xin[284] , \modmult_1/xin[283] , \modmult_1/xin[282] ,
         \modmult_1/xin[281] , \modmult_1/xin[280] , \modmult_1/xin[279] ,
         \modmult_1/xin[278] , \modmult_1/xin[277] , \modmult_1/xin[276] ,
         \modmult_1/xin[275] , \modmult_1/xin[274] , \modmult_1/xin[273] ,
         \modmult_1/xin[272] , \modmult_1/xin[271] , \modmult_1/xin[270] ,
         \modmult_1/xin[269] , \modmult_1/xin[268] , \modmult_1/xin[267] ,
         \modmult_1/xin[266] , \modmult_1/xin[265] , \modmult_1/xin[264] ,
         \modmult_1/xin[263] , \modmult_1/xin[262] , \modmult_1/xin[261] ,
         \modmult_1/xin[260] , \modmult_1/xin[259] , \modmult_1/xin[258] ,
         \modmult_1/xin[257] , \modmult_1/xin[256] , \modmult_1/xin[255] ,
         \modmult_1/xin[254] , \modmult_1/xin[253] , \modmult_1/xin[252] ,
         \modmult_1/xin[251] , \modmult_1/xin[250] , \modmult_1/xin[249] ,
         \modmult_1/xin[248] , \modmult_1/xin[247] , \modmult_1/xin[246] ,
         \modmult_1/xin[245] , \modmult_1/xin[244] , \modmult_1/xin[243] ,
         \modmult_1/xin[242] , \modmult_1/xin[241] , \modmult_1/xin[240] ,
         \modmult_1/xin[239] , \modmult_1/xin[238] , \modmult_1/xin[237] ,
         \modmult_1/xin[236] , \modmult_1/xin[235] , \modmult_1/xin[234] ,
         \modmult_1/xin[233] , \modmult_1/xin[232] , \modmult_1/xin[231] ,
         \modmult_1/xin[230] , \modmult_1/xin[229] , \modmult_1/xin[228] ,
         \modmult_1/xin[227] , \modmult_1/xin[226] , \modmult_1/xin[225] ,
         \modmult_1/xin[224] , \modmult_1/xin[223] , \modmult_1/xin[222] ,
         \modmult_1/xin[221] , \modmult_1/xin[220] , \modmult_1/xin[219] ,
         \modmult_1/xin[218] , \modmult_1/xin[217] , \modmult_1/xin[216] ,
         \modmult_1/xin[215] , \modmult_1/xin[214] , \modmult_1/xin[213] ,
         \modmult_1/xin[212] , \modmult_1/xin[211] , \modmult_1/xin[210] ,
         \modmult_1/xin[209] , \modmult_1/xin[208] , \modmult_1/xin[207] ,
         \modmult_1/xin[206] , \modmult_1/xin[205] , \modmult_1/xin[204] ,
         \modmult_1/xin[203] , \modmult_1/xin[202] , \modmult_1/xin[201] ,
         \modmult_1/xin[200] , \modmult_1/xin[199] , \modmult_1/xin[198] ,
         \modmult_1/xin[197] , \modmult_1/xin[196] , \modmult_1/xin[195] ,
         \modmult_1/xin[194] , \modmult_1/xin[193] , \modmult_1/xin[192] ,
         \modmult_1/xin[191] , \modmult_1/xin[190] , \modmult_1/xin[189] ,
         \modmult_1/xin[188] , \modmult_1/xin[187] , \modmult_1/xin[186] ,
         \modmult_1/xin[185] , \modmult_1/xin[184] , \modmult_1/xin[183] ,
         \modmult_1/xin[182] , \modmult_1/xin[181] , \modmult_1/xin[180] ,
         \modmult_1/xin[179] , \modmult_1/xin[178] , \modmult_1/xin[177] ,
         \modmult_1/xin[176] , \modmult_1/xin[175] , \modmult_1/xin[174] ,
         \modmult_1/xin[173] , \modmult_1/xin[172] , \modmult_1/xin[171] ,
         \modmult_1/xin[170] , \modmult_1/xin[169] , \modmult_1/xin[168] ,
         \modmult_1/xin[167] , \modmult_1/xin[166] , \modmult_1/xin[165] ,
         \modmult_1/xin[164] , \modmult_1/xin[163] , \modmult_1/xin[162] ,
         \modmult_1/xin[161] , \modmult_1/xin[160] , \modmult_1/xin[159] ,
         \modmult_1/xin[158] , \modmult_1/xin[157] , \modmult_1/xin[156] ,
         \modmult_1/xin[155] , \modmult_1/xin[154] , \modmult_1/xin[153] ,
         \modmult_1/xin[152] , \modmult_1/xin[151] , \modmult_1/xin[150] ,
         \modmult_1/xin[149] , \modmult_1/xin[148] , \modmult_1/xin[147] ,
         \modmult_1/xin[146] , \modmult_1/xin[145] , \modmult_1/xin[144] ,
         \modmult_1/xin[143] , \modmult_1/xin[142] , \modmult_1/xin[141] ,
         \modmult_1/xin[140] , \modmult_1/xin[139] , \modmult_1/xin[138] ,
         \modmult_1/xin[137] , \modmult_1/xin[136] , \modmult_1/xin[135] ,
         \modmult_1/xin[134] , \modmult_1/xin[133] , \modmult_1/xin[132] ,
         \modmult_1/xin[131] , \modmult_1/xin[130] , \modmult_1/xin[129] ,
         \modmult_1/xin[128] , \modmult_1/xin[127] , \modmult_1/xin[126] ,
         \modmult_1/xin[125] , \modmult_1/xin[124] , \modmult_1/xin[123] ,
         \modmult_1/xin[122] , \modmult_1/xin[121] , \modmult_1/xin[120] ,
         \modmult_1/xin[119] , \modmult_1/xin[118] , \modmult_1/xin[117] ,
         \modmult_1/xin[116] , \modmult_1/xin[115] , \modmult_1/xin[114] ,
         \modmult_1/xin[113] , \modmult_1/xin[112] , \modmult_1/xin[111] ,
         \modmult_1/xin[110] , \modmult_1/xin[109] , \modmult_1/xin[108] ,
         \modmult_1/xin[107] , \modmult_1/xin[106] , \modmult_1/xin[105] ,
         \modmult_1/xin[104] , \modmult_1/xin[103] , \modmult_1/xin[102] ,
         \modmult_1/xin[101] , \modmult_1/xin[100] , \modmult_1/xin[99] ,
         \modmult_1/xin[98] , \modmult_1/xin[97] , \modmult_1/xin[96] ,
         \modmult_1/xin[95] , \modmult_1/xin[94] , \modmult_1/xin[93] ,
         \modmult_1/xin[92] , \modmult_1/xin[91] , \modmult_1/xin[90] ,
         \modmult_1/xin[89] , \modmult_1/xin[88] , \modmult_1/xin[87] ,
         \modmult_1/xin[86] , \modmult_1/xin[85] , \modmult_1/xin[84] ,
         \modmult_1/xin[83] , \modmult_1/xin[82] , \modmult_1/xin[81] ,
         \modmult_1/xin[80] , \modmult_1/xin[79] , \modmult_1/xin[78] ,
         \modmult_1/xin[77] , \modmult_1/xin[76] , \modmult_1/xin[75] ,
         \modmult_1/xin[74] , \modmult_1/xin[73] , \modmult_1/xin[72] ,
         \modmult_1/xin[71] , \modmult_1/xin[70] , \modmult_1/xin[69] ,
         \modmult_1/xin[68] , \modmult_1/xin[67] , \modmult_1/xin[66] ,
         \modmult_1/xin[65] , \modmult_1/xin[64] , \modmult_1/xin[63] ,
         \modmult_1/xin[62] , \modmult_1/xin[61] , \modmult_1/xin[60] ,
         \modmult_1/xin[59] , \modmult_1/xin[58] , \modmult_1/xin[57] ,
         \modmult_1/xin[56] , \modmult_1/xin[55] , \modmult_1/xin[54] ,
         \modmult_1/xin[53] , \modmult_1/xin[52] , \modmult_1/xin[51] ,
         \modmult_1/xin[50] , \modmult_1/xin[49] , \modmult_1/xin[48] ,
         \modmult_1/xin[47] , \modmult_1/xin[46] , \modmult_1/xin[45] ,
         \modmult_1/xin[44] , \modmult_1/xin[43] , \modmult_1/xin[42] ,
         \modmult_1/xin[41] , \modmult_1/xin[40] , \modmult_1/xin[39] ,
         \modmult_1/xin[38] , \modmult_1/xin[37] , \modmult_1/xin[36] ,
         \modmult_1/xin[35] , \modmult_1/xin[34] , \modmult_1/xin[33] ,
         \modmult_1/xin[32] , \modmult_1/xin[31] , \modmult_1/xin[30] ,
         \modmult_1/xin[29] , \modmult_1/xin[28] , \modmult_1/xin[27] ,
         \modmult_1/xin[26] , \modmult_1/xin[25] , \modmult_1/xin[24] ,
         \modmult_1/xin[23] , \modmult_1/xin[22] , \modmult_1/xin[21] ,
         \modmult_1/xin[20] , \modmult_1/xin[19] , \modmult_1/xin[18] ,
         \modmult_1/xin[17] , \modmult_1/xin[16] , \modmult_1/xin[15] ,
         \modmult_1/xin[14] , \modmult_1/xin[13] , \modmult_1/xin[12] ,
         \modmult_1/xin[11] , \modmult_1/xin[10] , \modmult_1/xin[9] ,
         \modmult_1/xin[8] , \modmult_1/xin[7] , \modmult_1/xin[6] ,
         \modmult_1/xin[5] , \modmult_1/xin[4] , \modmult_1/xin[3] ,
         \modmult_1/xin[2] , \modmult_1/xin[1] , \modmult_1/xin[0] ,
         \modmult_1/zin[0][1024] , \modmult_1/zin[0][1023] ,
         \modmult_1/zin[0][1022] , \modmult_1/zin[0][1021] ,
         \modmult_1/zin[0][1020] , \modmult_1/zin[0][1019] ,
         \modmult_1/zin[0][1018] , \modmult_1/zin[0][1017] ,
         \modmult_1/zin[0][1016] , \modmult_1/zin[0][1015] ,
         \modmult_1/zin[0][1014] , \modmult_1/zin[0][1013] ,
         \modmult_1/zin[0][1012] , \modmult_1/zin[0][1011] ,
         \modmult_1/zin[0][1010] , \modmult_1/zin[0][1009] ,
         \modmult_1/zin[0][1008] , \modmult_1/zin[0][1007] ,
         \modmult_1/zin[0][1006] , \modmult_1/zin[0][1005] ,
         \modmult_1/zin[0][1004] , \modmult_1/zin[0][1003] ,
         \modmult_1/zin[0][1002] , \modmult_1/zin[0][1001] ,
         \modmult_1/zin[0][1000] , \modmult_1/zin[0][999] ,
         \modmult_1/zin[0][998] , \modmult_1/zin[0][997] ,
         \modmult_1/zin[0][996] , \modmult_1/zin[0][995] ,
         \modmult_1/zin[0][994] , \modmult_1/zin[0][993] ,
         \modmult_1/zin[0][992] , \modmult_1/zin[0][991] ,
         \modmult_1/zin[0][990] , \modmult_1/zin[0][989] ,
         \modmult_1/zin[0][988] , \modmult_1/zin[0][987] ,
         \modmult_1/zin[0][986] , \modmult_1/zin[0][985] ,
         \modmult_1/zin[0][984] , \modmult_1/zin[0][983] ,
         \modmult_1/zin[0][982] , \modmult_1/zin[0][981] ,
         \modmult_1/zin[0][980] , \modmult_1/zin[0][979] ,
         \modmult_1/zin[0][978] , \modmult_1/zin[0][977] ,
         \modmult_1/zin[0][976] , \modmult_1/zin[0][975] ,
         \modmult_1/zin[0][974] , \modmult_1/zin[0][973] ,
         \modmult_1/zin[0][972] , \modmult_1/zin[0][971] ,
         \modmult_1/zin[0][970] , \modmult_1/zin[0][969] ,
         \modmult_1/zin[0][968] , \modmult_1/zin[0][967] ,
         \modmult_1/zin[0][966] , \modmult_1/zin[0][965] ,
         \modmult_1/zin[0][964] , \modmult_1/zin[0][963] ,
         \modmult_1/zin[0][962] , \modmult_1/zin[0][961] ,
         \modmult_1/zin[0][960] , \modmult_1/zin[0][959] ,
         \modmult_1/zin[0][958] , \modmult_1/zin[0][957] ,
         \modmult_1/zin[0][956] , \modmult_1/zin[0][955] ,
         \modmult_1/zin[0][954] , \modmult_1/zin[0][953] ,
         \modmult_1/zin[0][952] , \modmult_1/zin[0][951] ,
         \modmult_1/zin[0][950] , \modmult_1/zin[0][949] ,
         \modmult_1/zin[0][948] , \modmult_1/zin[0][947] ,
         \modmult_1/zin[0][946] , \modmult_1/zin[0][945] ,
         \modmult_1/zin[0][944] , \modmult_1/zin[0][943] ,
         \modmult_1/zin[0][942] , \modmult_1/zin[0][941] ,
         \modmult_1/zin[0][940] , \modmult_1/zin[0][939] ,
         \modmult_1/zin[0][938] , \modmult_1/zin[0][937] ,
         \modmult_1/zin[0][936] , \modmult_1/zin[0][935] ,
         \modmult_1/zin[0][934] , \modmult_1/zin[0][933] ,
         \modmult_1/zin[0][932] , \modmult_1/zin[0][931] ,
         \modmult_1/zin[0][930] , \modmult_1/zin[0][929] ,
         \modmult_1/zin[0][928] , \modmult_1/zin[0][927] ,
         \modmult_1/zin[0][926] , \modmult_1/zin[0][925] ,
         \modmult_1/zin[0][924] , \modmult_1/zin[0][923] ,
         \modmult_1/zin[0][922] , \modmult_1/zin[0][921] ,
         \modmult_1/zin[0][920] , \modmult_1/zin[0][919] ,
         \modmult_1/zin[0][918] , \modmult_1/zin[0][917] ,
         \modmult_1/zin[0][916] , \modmult_1/zin[0][915] ,
         \modmult_1/zin[0][914] , \modmult_1/zin[0][913] ,
         \modmult_1/zin[0][912] , \modmult_1/zin[0][911] ,
         \modmult_1/zin[0][910] , \modmult_1/zin[0][909] ,
         \modmult_1/zin[0][908] , \modmult_1/zin[0][907] ,
         \modmult_1/zin[0][906] , \modmult_1/zin[0][905] ,
         \modmult_1/zin[0][904] , \modmult_1/zin[0][903] ,
         \modmult_1/zin[0][902] , \modmult_1/zin[0][901] ,
         \modmult_1/zin[0][900] , \modmult_1/zin[0][899] ,
         \modmult_1/zin[0][898] , \modmult_1/zin[0][897] ,
         \modmult_1/zin[0][896] , \modmult_1/zin[0][895] ,
         \modmult_1/zin[0][894] , \modmult_1/zin[0][893] ,
         \modmult_1/zin[0][892] , \modmult_1/zin[0][891] ,
         \modmult_1/zin[0][890] , \modmult_1/zin[0][889] ,
         \modmult_1/zin[0][888] , \modmult_1/zin[0][887] ,
         \modmult_1/zin[0][886] , \modmult_1/zin[0][885] ,
         \modmult_1/zin[0][884] , \modmult_1/zin[0][883] ,
         \modmult_1/zin[0][882] , \modmult_1/zin[0][881] ,
         \modmult_1/zin[0][880] , \modmult_1/zin[0][879] ,
         \modmult_1/zin[0][878] , \modmult_1/zin[0][877] ,
         \modmult_1/zin[0][876] , \modmult_1/zin[0][875] ,
         \modmult_1/zin[0][874] , \modmult_1/zin[0][873] ,
         \modmult_1/zin[0][872] , \modmult_1/zin[0][871] ,
         \modmult_1/zin[0][870] , \modmult_1/zin[0][869] ,
         \modmult_1/zin[0][868] , \modmult_1/zin[0][867] ,
         \modmult_1/zin[0][866] , \modmult_1/zin[0][865] ,
         \modmult_1/zin[0][864] , \modmult_1/zin[0][863] ,
         \modmult_1/zin[0][862] , \modmult_1/zin[0][861] ,
         \modmult_1/zin[0][860] , \modmult_1/zin[0][859] ,
         \modmult_1/zin[0][858] , \modmult_1/zin[0][857] ,
         \modmult_1/zin[0][856] , \modmult_1/zin[0][855] ,
         \modmult_1/zin[0][854] , \modmult_1/zin[0][853] ,
         \modmult_1/zin[0][852] , \modmult_1/zin[0][851] ,
         \modmult_1/zin[0][850] , \modmult_1/zin[0][849] ,
         \modmult_1/zin[0][848] , \modmult_1/zin[0][847] ,
         \modmult_1/zin[0][846] , \modmult_1/zin[0][845] ,
         \modmult_1/zin[0][844] , \modmult_1/zin[0][843] ,
         \modmult_1/zin[0][842] , \modmult_1/zin[0][841] ,
         \modmult_1/zin[0][840] , \modmult_1/zin[0][839] ,
         \modmult_1/zin[0][838] , \modmult_1/zin[0][837] ,
         \modmult_1/zin[0][836] , \modmult_1/zin[0][835] ,
         \modmult_1/zin[0][834] , \modmult_1/zin[0][833] ,
         \modmult_1/zin[0][832] , \modmult_1/zin[0][831] ,
         \modmult_1/zin[0][830] , \modmult_1/zin[0][829] ,
         \modmult_1/zin[0][828] , \modmult_1/zin[0][827] ,
         \modmult_1/zin[0][826] , \modmult_1/zin[0][825] ,
         \modmult_1/zin[0][824] , \modmult_1/zin[0][823] ,
         \modmult_1/zin[0][822] , \modmult_1/zin[0][821] ,
         \modmult_1/zin[0][820] , \modmult_1/zin[0][819] ,
         \modmult_1/zin[0][818] , \modmult_1/zin[0][817] ,
         \modmult_1/zin[0][816] , \modmult_1/zin[0][815] ,
         \modmult_1/zin[0][814] , \modmult_1/zin[0][813] ,
         \modmult_1/zin[0][812] , \modmult_1/zin[0][811] ,
         \modmult_1/zin[0][810] , \modmult_1/zin[0][809] ,
         \modmult_1/zin[0][808] , \modmult_1/zin[0][807] ,
         \modmult_1/zin[0][806] , \modmult_1/zin[0][805] ,
         \modmult_1/zin[0][804] , \modmult_1/zin[0][803] ,
         \modmult_1/zin[0][802] , \modmult_1/zin[0][801] ,
         \modmult_1/zin[0][800] , \modmult_1/zin[0][799] ,
         \modmult_1/zin[0][798] , \modmult_1/zin[0][797] ,
         \modmult_1/zin[0][796] , \modmult_1/zin[0][795] ,
         \modmult_1/zin[0][794] , \modmult_1/zin[0][793] ,
         \modmult_1/zin[0][792] , \modmult_1/zin[0][791] ,
         \modmult_1/zin[0][790] , \modmult_1/zin[0][789] ,
         \modmult_1/zin[0][788] , \modmult_1/zin[0][787] ,
         \modmult_1/zin[0][786] , \modmult_1/zin[0][785] ,
         \modmult_1/zin[0][784] , \modmult_1/zin[0][783] ,
         \modmult_1/zin[0][782] , \modmult_1/zin[0][781] ,
         \modmult_1/zin[0][780] , \modmult_1/zin[0][779] ,
         \modmult_1/zin[0][778] , \modmult_1/zin[0][777] ,
         \modmult_1/zin[0][776] , \modmult_1/zin[0][775] ,
         \modmult_1/zin[0][774] , \modmult_1/zin[0][773] ,
         \modmult_1/zin[0][772] , \modmult_1/zin[0][771] ,
         \modmult_1/zin[0][770] , \modmult_1/zin[0][769] ,
         \modmult_1/zin[0][768] , \modmult_1/zin[0][767] ,
         \modmult_1/zin[0][766] , \modmult_1/zin[0][765] ,
         \modmult_1/zin[0][764] , \modmult_1/zin[0][763] ,
         \modmult_1/zin[0][762] , \modmult_1/zin[0][761] ,
         \modmult_1/zin[0][760] , \modmult_1/zin[0][759] ,
         \modmult_1/zin[0][758] , \modmult_1/zin[0][757] ,
         \modmult_1/zin[0][756] , \modmult_1/zin[0][755] ,
         \modmult_1/zin[0][754] , \modmult_1/zin[0][753] ,
         \modmult_1/zin[0][752] , \modmult_1/zin[0][751] ,
         \modmult_1/zin[0][750] , \modmult_1/zin[0][749] ,
         \modmult_1/zin[0][748] , \modmult_1/zin[0][747] ,
         \modmult_1/zin[0][746] , \modmult_1/zin[0][745] ,
         \modmult_1/zin[0][744] , \modmult_1/zin[0][743] ,
         \modmult_1/zin[0][742] , \modmult_1/zin[0][741] ,
         \modmult_1/zin[0][740] , \modmult_1/zin[0][739] ,
         \modmult_1/zin[0][738] , \modmult_1/zin[0][737] ,
         \modmult_1/zin[0][736] , \modmult_1/zin[0][735] ,
         \modmult_1/zin[0][734] , \modmult_1/zin[0][733] ,
         \modmult_1/zin[0][732] , \modmult_1/zin[0][731] ,
         \modmult_1/zin[0][730] , \modmult_1/zin[0][729] ,
         \modmult_1/zin[0][728] , \modmult_1/zin[0][727] ,
         \modmult_1/zin[0][726] , \modmult_1/zin[0][725] ,
         \modmult_1/zin[0][724] , \modmult_1/zin[0][723] ,
         \modmult_1/zin[0][722] , \modmult_1/zin[0][721] ,
         \modmult_1/zin[0][720] , \modmult_1/zin[0][719] ,
         \modmult_1/zin[0][718] , \modmult_1/zin[0][717] ,
         \modmult_1/zin[0][716] , \modmult_1/zin[0][715] ,
         \modmult_1/zin[0][714] , \modmult_1/zin[0][713] ,
         \modmult_1/zin[0][712] , \modmult_1/zin[0][711] ,
         \modmult_1/zin[0][710] , \modmult_1/zin[0][709] ,
         \modmult_1/zin[0][708] , \modmult_1/zin[0][707] ,
         \modmult_1/zin[0][706] , \modmult_1/zin[0][705] ,
         \modmult_1/zin[0][704] , \modmult_1/zin[0][703] ,
         \modmult_1/zin[0][702] , \modmult_1/zin[0][701] ,
         \modmult_1/zin[0][700] , \modmult_1/zin[0][699] ,
         \modmult_1/zin[0][698] , \modmult_1/zin[0][697] ,
         \modmult_1/zin[0][696] , \modmult_1/zin[0][695] ,
         \modmult_1/zin[0][694] , \modmult_1/zin[0][693] ,
         \modmult_1/zin[0][692] , \modmult_1/zin[0][691] ,
         \modmult_1/zin[0][690] , \modmult_1/zin[0][689] ,
         \modmult_1/zin[0][688] , \modmult_1/zin[0][687] ,
         \modmult_1/zin[0][686] , \modmult_1/zin[0][685] ,
         \modmult_1/zin[0][684] , \modmult_1/zin[0][683] ,
         \modmult_1/zin[0][682] , \modmult_1/zin[0][681] ,
         \modmult_1/zin[0][680] , \modmult_1/zin[0][679] ,
         \modmult_1/zin[0][678] , \modmult_1/zin[0][677] ,
         \modmult_1/zin[0][676] , \modmult_1/zin[0][675] ,
         \modmult_1/zin[0][674] , \modmult_1/zin[0][673] ,
         \modmult_1/zin[0][672] , \modmult_1/zin[0][671] ,
         \modmult_1/zin[0][670] , \modmult_1/zin[0][669] ,
         \modmult_1/zin[0][668] , \modmult_1/zin[0][667] ,
         \modmult_1/zin[0][666] , \modmult_1/zin[0][665] ,
         \modmult_1/zin[0][664] , \modmult_1/zin[0][663] ,
         \modmult_1/zin[0][662] , \modmult_1/zin[0][661] ,
         \modmult_1/zin[0][660] , \modmult_1/zin[0][659] ,
         \modmult_1/zin[0][658] , \modmult_1/zin[0][657] ,
         \modmult_1/zin[0][656] , \modmult_1/zin[0][655] ,
         \modmult_1/zin[0][654] , \modmult_1/zin[0][653] ,
         \modmult_1/zin[0][652] , \modmult_1/zin[0][651] ,
         \modmult_1/zin[0][650] , \modmult_1/zin[0][649] ,
         \modmult_1/zin[0][648] , \modmult_1/zin[0][647] ,
         \modmult_1/zin[0][646] , \modmult_1/zin[0][645] ,
         \modmult_1/zin[0][644] , \modmult_1/zin[0][643] ,
         \modmult_1/zin[0][642] , \modmult_1/zin[0][641] ,
         \modmult_1/zin[0][640] , \modmult_1/zin[0][639] ,
         \modmult_1/zin[0][638] , \modmult_1/zin[0][637] ,
         \modmult_1/zin[0][636] , \modmult_1/zin[0][635] ,
         \modmult_1/zin[0][634] , \modmult_1/zin[0][633] ,
         \modmult_1/zin[0][632] , \modmult_1/zin[0][631] ,
         \modmult_1/zin[0][630] , \modmult_1/zin[0][629] ,
         \modmult_1/zin[0][628] , \modmult_1/zin[0][627] ,
         \modmult_1/zin[0][626] , \modmult_1/zin[0][625] ,
         \modmult_1/zin[0][624] , \modmult_1/zin[0][623] ,
         \modmult_1/zin[0][622] , \modmult_1/zin[0][621] ,
         \modmult_1/zin[0][620] , \modmult_1/zin[0][619] ,
         \modmult_1/zin[0][618] , \modmult_1/zin[0][617] ,
         \modmult_1/zin[0][616] , \modmult_1/zin[0][615] ,
         \modmult_1/zin[0][614] , \modmult_1/zin[0][613] ,
         \modmult_1/zin[0][612] , \modmult_1/zin[0][611] ,
         \modmult_1/zin[0][610] , \modmult_1/zin[0][609] ,
         \modmult_1/zin[0][608] , \modmult_1/zin[0][607] ,
         \modmult_1/zin[0][606] , \modmult_1/zin[0][605] ,
         \modmult_1/zin[0][604] , \modmult_1/zin[0][603] ,
         \modmult_1/zin[0][602] , \modmult_1/zin[0][601] ,
         \modmult_1/zin[0][600] , \modmult_1/zin[0][599] ,
         \modmult_1/zin[0][598] , \modmult_1/zin[0][597] ,
         \modmult_1/zin[0][596] , \modmult_1/zin[0][595] ,
         \modmult_1/zin[0][594] , \modmult_1/zin[0][593] ,
         \modmult_1/zin[0][592] , \modmult_1/zin[0][591] ,
         \modmult_1/zin[0][590] , \modmult_1/zin[0][589] ,
         \modmult_1/zin[0][588] , \modmult_1/zin[0][587] ,
         \modmult_1/zin[0][586] , \modmult_1/zin[0][585] ,
         \modmult_1/zin[0][584] , \modmult_1/zin[0][583] ,
         \modmult_1/zin[0][582] , \modmult_1/zin[0][581] ,
         \modmult_1/zin[0][580] , \modmult_1/zin[0][579] ,
         \modmult_1/zin[0][578] , \modmult_1/zin[0][577] ,
         \modmult_1/zin[0][576] , \modmult_1/zin[0][575] ,
         \modmult_1/zin[0][574] , \modmult_1/zin[0][573] ,
         \modmult_1/zin[0][572] , \modmult_1/zin[0][571] ,
         \modmult_1/zin[0][570] , \modmult_1/zin[0][569] ,
         \modmult_1/zin[0][568] , \modmult_1/zin[0][567] ,
         \modmult_1/zin[0][566] , \modmult_1/zin[0][565] ,
         \modmult_1/zin[0][564] , \modmult_1/zin[0][563] ,
         \modmult_1/zin[0][562] , \modmult_1/zin[0][561] ,
         \modmult_1/zin[0][560] , \modmult_1/zin[0][559] ,
         \modmult_1/zin[0][558] , \modmult_1/zin[0][557] ,
         \modmult_1/zin[0][556] , \modmult_1/zin[0][555] ,
         \modmult_1/zin[0][554] , \modmult_1/zin[0][553] ,
         \modmult_1/zin[0][552] , \modmult_1/zin[0][551] ,
         \modmult_1/zin[0][550] , \modmult_1/zin[0][549] ,
         \modmult_1/zin[0][548] , \modmult_1/zin[0][547] ,
         \modmult_1/zin[0][546] , \modmult_1/zin[0][545] ,
         \modmult_1/zin[0][544] , \modmult_1/zin[0][543] ,
         \modmult_1/zin[0][542] , \modmult_1/zin[0][541] ,
         \modmult_1/zin[0][540] , \modmult_1/zin[0][539] ,
         \modmult_1/zin[0][538] , \modmult_1/zin[0][537] ,
         \modmult_1/zin[0][536] , \modmult_1/zin[0][535] ,
         \modmult_1/zin[0][534] , \modmult_1/zin[0][533] ,
         \modmult_1/zin[0][532] , \modmult_1/zin[0][531] ,
         \modmult_1/zin[0][530] , \modmult_1/zin[0][529] ,
         \modmult_1/zin[0][528] , \modmult_1/zin[0][527] ,
         \modmult_1/zin[0][526] , \modmult_1/zin[0][525] ,
         \modmult_1/zin[0][524] , \modmult_1/zin[0][523] ,
         \modmult_1/zin[0][522] , \modmult_1/zin[0][521] ,
         \modmult_1/zin[0][520] , \modmult_1/zin[0][519] ,
         \modmult_1/zin[0][518] , \modmult_1/zin[0][517] ,
         \modmult_1/zin[0][516] , \modmult_1/zin[0][515] ,
         \modmult_1/zin[0][514] , \modmult_1/zin[0][513] ,
         \modmult_1/zin[0][512] , \modmult_1/zin[0][511] ,
         \modmult_1/zin[0][510] , \modmult_1/zin[0][509] ,
         \modmult_1/zin[0][508] , \modmult_1/zin[0][507] ,
         \modmult_1/zin[0][506] , \modmult_1/zin[0][505] ,
         \modmult_1/zin[0][504] , \modmult_1/zin[0][503] ,
         \modmult_1/zin[0][502] , \modmult_1/zin[0][501] ,
         \modmult_1/zin[0][500] , \modmult_1/zin[0][499] ,
         \modmult_1/zin[0][498] , \modmult_1/zin[0][497] ,
         \modmult_1/zin[0][496] , \modmult_1/zin[0][495] ,
         \modmult_1/zin[0][494] , \modmult_1/zin[0][493] ,
         \modmult_1/zin[0][492] , \modmult_1/zin[0][491] ,
         \modmult_1/zin[0][490] , \modmult_1/zin[0][489] ,
         \modmult_1/zin[0][488] , \modmult_1/zin[0][487] ,
         \modmult_1/zin[0][486] , \modmult_1/zin[0][485] ,
         \modmult_1/zin[0][484] , \modmult_1/zin[0][483] ,
         \modmult_1/zin[0][482] , \modmult_1/zin[0][481] ,
         \modmult_1/zin[0][480] , \modmult_1/zin[0][479] ,
         \modmult_1/zin[0][478] , \modmult_1/zin[0][477] ,
         \modmult_1/zin[0][476] , \modmult_1/zin[0][475] ,
         \modmult_1/zin[0][474] , \modmult_1/zin[0][473] ,
         \modmult_1/zin[0][472] , \modmult_1/zin[0][471] ,
         \modmult_1/zin[0][470] , \modmult_1/zin[0][469] ,
         \modmult_1/zin[0][468] , \modmult_1/zin[0][467] ,
         \modmult_1/zin[0][466] , \modmult_1/zin[0][465] ,
         \modmult_1/zin[0][464] , \modmult_1/zin[0][463] ,
         \modmult_1/zin[0][462] , \modmult_1/zin[0][461] ,
         \modmult_1/zin[0][460] , \modmult_1/zin[0][459] ,
         \modmult_1/zin[0][458] , \modmult_1/zin[0][457] ,
         \modmult_1/zin[0][456] , \modmult_1/zin[0][455] ,
         \modmult_1/zin[0][454] , \modmult_1/zin[0][453] ,
         \modmult_1/zin[0][452] , \modmult_1/zin[0][451] ,
         \modmult_1/zin[0][450] , \modmult_1/zin[0][449] ,
         \modmult_1/zin[0][448] , \modmult_1/zin[0][447] ,
         \modmult_1/zin[0][446] , \modmult_1/zin[0][445] ,
         \modmult_1/zin[0][444] , \modmult_1/zin[0][443] ,
         \modmult_1/zin[0][442] , \modmult_1/zin[0][441] ,
         \modmult_1/zin[0][440] , \modmult_1/zin[0][439] ,
         \modmult_1/zin[0][438] , \modmult_1/zin[0][437] ,
         \modmult_1/zin[0][436] , \modmult_1/zin[0][435] ,
         \modmult_1/zin[0][434] , \modmult_1/zin[0][433] ,
         \modmult_1/zin[0][432] , \modmult_1/zin[0][431] ,
         \modmult_1/zin[0][430] , \modmult_1/zin[0][429] ,
         \modmult_1/zin[0][428] , \modmult_1/zin[0][427] ,
         \modmult_1/zin[0][426] , \modmult_1/zin[0][425] ,
         \modmult_1/zin[0][424] , \modmult_1/zin[0][423] ,
         \modmult_1/zin[0][422] , \modmult_1/zin[0][421] ,
         \modmult_1/zin[0][420] , \modmult_1/zin[0][419] ,
         \modmult_1/zin[0][418] , \modmult_1/zin[0][417] ,
         \modmult_1/zin[0][416] , \modmult_1/zin[0][415] ,
         \modmult_1/zin[0][414] , \modmult_1/zin[0][413] ,
         \modmult_1/zin[0][412] , \modmult_1/zin[0][411] ,
         \modmult_1/zin[0][410] , \modmult_1/zin[0][409] ,
         \modmult_1/zin[0][408] , \modmult_1/zin[0][407] ,
         \modmult_1/zin[0][406] , \modmult_1/zin[0][405] ,
         \modmult_1/zin[0][404] , \modmult_1/zin[0][403] ,
         \modmult_1/zin[0][402] , \modmult_1/zin[0][401] ,
         \modmult_1/zin[0][400] , \modmult_1/zin[0][399] ,
         \modmult_1/zin[0][398] , \modmult_1/zin[0][397] ,
         \modmult_1/zin[0][396] , \modmult_1/zin[0][395] ,
         \modmult_1/zin[0][394] , \modmult_1/zin[0][393] ,
         \modmult_1/zin[0][392] , \modmult_1/zin[0][391] ,
         \modmult_1/zin[0][390] , \modmult_1/zin[0][389] ,
         \modmult_1/zin[0][388] , \modmult_1/zin[0][387] ,
         \modmult_1/zin[0][386] , \modmult_1/zin[0][385] ,
         \modmult_1/zin[0][384] , \modmult_1/zin[0][383] ,
         \modmult_1/zin[0][382] , \modmult_1/zin[0][381] ,
         \modmult_1/zin[0][380] , \modmult_1/zin[0][379] ,
         \modmult_1/zin[0][378] , \modmult_1/zin[0][377] ,
         \modmult_1/zin[0][376] , \modmult_1/zin[0][375] ,
         \modmult_1/zin[0][374] , \modmult_1/zin[0][373] ,
         \modmult_1/zin[0][372] , \modmult_1/zin[0][371] ,
         \modmult_1/zin[0][370] , \modmult_1/zin[0][369] ,
         \modmult_1/zin[0][368] , \modmult_1/zin[0][367] ,
         \modmult_1/zin[0][366] , \modmult_1/zin[0][365] ,
         \modmult_1/zin[0][364] , \modmult_1/zin[0][363] ,
         \modmult_1/zin[0][362] , \modmult_1/zin[0][361] ,
         \modmult_1/zin[0][360] , \modmult_1/zin[0][359] ,
         \modmult_1/zin[0][358] , \modmult_1/zin[0][357] ,
         \modmult_1/zin[0][356] , \modmult_1/zin[0][355] ,
         \modmult_1/zin[0][354] , \modmult_1/zin[0][353] ,
         \modmult_1/zin[0][352] , \modmult_1/zin[0][351] ,
         \modmult_1/zin[0][350] , \modmult_1/zin[0][349] ,
         \modmult_1/zin[0][348] , \modmult_1/zin[0][347] ,
         \modmult_1/zin[0][346] , \modmult_1/zin[0][345] ,
         \modmult_1/zin[0][344] , \modmult_1/zin[0][343] ,
         \modmult_1/zin[0][342] , \modmult_1/zin[0][341] ,
         \modmult_1/zin[0][340] , \modmult_1/zin[0][339] ,
         \modmult_1/zin[0][338] , \modmult_1/zin[0][337] ,
         \modmult_1/zin[0][336] , \modmult_1/zin[0][335] ,
         \modmult_1/zin[0][334] , \modmult_1/zin[0][333] ,
         \modmult_1/zin[0][332] , \modmult_1/zin[0][331] ,
         \modmult_1/zin[0][330] , \modmult_1/zin[0][329] ,
         \modmult_1/zin[0][328] , \modmult_1/zin[0][327] ,
         \modmult_1/zin[0][326] , \modmult_1/zin[0][325] ,
         \modmult_1/zin[0][324] , \modmult_1/zin[0][323] ,
         \modmult_1/zin[0][322] , \modmult_1/zin[0][321] ,
         \modmult_1/zin[0][320] , \modmult_1/zin[0][319] ,
         \modmult_1/zin[0][318] , \modmult_1/zin[0][317] ,
         \modmult_1/zin[0][316] , \modmult_1/zin[0][315] ,
         \modmult_1/zin[0][314] , \modmult_1/zin[0][313] ,
         \modmult_1/zin[0][312] , \modmult_1/zin[0][311] ,
         \modmult_1/zin[0][310] , \modmult_1/zin[0][309] ,
         \modmult_1/zin[0][308] , \modmult_1/zin[0][307] ,
         \modmult_1/zin[0][306] , \modmult_1/zin[0][305] ,
         \modmult_1/zin[0][304] , \modmult_1/zin[0][303] ,
         \modmult_1/zin[0][302] , \modmult_1/zin[0][301] ,
         \modmult_1/zin[0][300] , \modmult_1/zin[0][299] ,
         \modmult_1/zin[0][298] , \modmult_1/zin[0][297] ,
         \modmult_1/zin[0][296] , \modmult_1/zin[0][295] ,
         \modmult_1/zin[0][294] , \modmult_1/zin[0][293] ,
         \modmult_1/zin[0][292] , \modmult_1/zin[0][291] ,
         \modmult_1/zin[0][290] , \modmult_1/zin[0][289] ,
         \modmult_1/zin[0][288] , \modmult_1/zin[0][287] ,
         \modmult_1/zin[0][286] , \modmult_1/zin[0][285] ,
         \modmult_1/zin[0][284] , \modmult_1/zin[0][283] ,
         \modmult_1/zin[0][282] , \modmult_1/zin[0][281] ,
         \modmult_1/zin[0][280] , \modmult_1/zin[0][279] ,
         \modmult_1/zin[0][278] , \modmult_1/zin[0][277] ,
         \modmult_1/zin[0][276] , \modmult_1/zin[0][275] ,
         \modmult_1/zin[0][274] , \modmult_1/zin[0][273] ,
         \modmult_1/zin[0][272] , \modmult_1/zin[0][271] ,
         \modmult_1/zin[0][270] , \modmult_1/zin[0][269] ,
         \modmult_1/zin[0][268] , \modmult_1/zin[0][267] ,
         \modmult_1/zin[0][266] , \modmult_1/zin[0][265] ,
         \modmult_1/zin[0][264] , \modmult_1/zin[0][263] ,
         \modmult_1/zin[0][262] , \modmult_1/zin[0][261] ,
         \modmult_1/zin[0][260] , \modmult_1/zin[0][259] ,
         \modmult_1/zin[0][258] , \modmult_1/zin[0][257] ,
         \modmult_1/zin[0][256] , \modmult_1/zin[0][255] ,
         \modmult_1/zin[0][254] , \modmult_1/zin[0][253] ,
         \modmult_1/zin[0][252] , \modmult_1/zin[0][251] ,
         \modmult_1/zin[0][250] , \modmult_1/zin[0][249] ,
         \modmult_1/zin[0][248] , \modmult_1/zin[0][247] ,
         \modmult_1/zin[0][246] , \modmult_1/zin[0][245] ,
         \modmult_1/zin[0][244] , \modmult_1/zin[0][243] ,
         \modmult_1/zin[0][242] , \modmult_1/zin[0][241] ,
         \modmult_1/zin[0][240] , \modmult_1/zin[0][239] ,
         \modmult_1/zin[0][238] , \modmult_1/zin[0][237] ,
         \modmult_1/zin[0][236] , \modmult_1/zin[0][235] ,
         \modmult_1/zin[0][234] , \modmult_1/zin[0][233] ,
         \modmult_1/zin[0][232] , \modmult_1/zin[0][231] ,
         \modmult_1/zin[0][230] , \modmult_1/zin[0][229] ,
         \modmult_1/zin[0][228] , \modmult_1/zin[0][227] ,
         \modmult_1/zin[0][226] , \modmult_1/zin[0][225] ,
         \modmult_1/zin[0][224] , \modmult_1/zin[0][223] ,
         \modmult_1/zin[0][222] , \modmult_1/zin[0][221] ,
         \modmult_1/zin[0][220] , \modmult_1/zin[0][219] ,
         \modmult_1/zin[0][218] , \modmult_1/zin[0][217] ,
         \modmult_1/zin[0][216] , \modmult_1/zin[0][215] ,
         \modmult_1/zin[0][214] , \modmult_1/zin[0][213] ,
         \modmult_1/zin[0][212] , \modmult_1/zin[0][211] ,
         \modmult_1/zin[0][210] , \modmult_1/zin[0][209] ,
         \modmult_1/zin[0][208] , \modmult_1/zin[0][207] ,
         \modmult_1/zin[0][206] , \modmult_1/zin[0][205] ,
         \modmult_1/zin[0][204] , \modmult_1/zin[0][203] ,
         \modmult_1/zin[0][202] , \modmult_1/zin[0][201] ,
         \modmult_1/zin[0][200] , \modmult_1/zin[0][199] ,
         \modmult_1/zin[0][198] , \modmult_1/zin[0][197] ,
         \modmult_1/zin[0][196] , \modmult_1/zin[0][195] ,
         \modmult_1/zin[0][194] , \modmult_1/zin[0][193] ,
         \modmult_1/zin[0][192] , \modmult_1/zin[0][191] ,
         \modmult_1/zin[0][190] , \modmult_1/zin[0][189] ,
         \modmult_1/zin[0][188] , \modmult_1/zin[0][187] ,
         \modmult_1/zin[0][186] , \modmult_1/zin[0][185] ,
         \modmult_1/zin[0][184] , \modmult_1/zin[0][183] ,
         \modmult_1/zin[0][182] , \modmult_1/zin[0][181] ,
         \modmult_1/zin[0][180] , \modmult_1/zin[0][179] ,
         \modmult_1/zin[0][178] , \modmult_1/zin[0][177] ,
         \modmult_1/zin[0][176] , \modmult_1/zin[0][175] ,
         \modmult_1/zin[0][174] , \modmult_1/zin[0][173] ,
         \modmult_1/zin[0][172] , \modmult_1/zin[0][171] ,
         \modmult_1/zin[0][170] , \modmult_1/zin[0][169] ,
         \modmult_1/zin[0][168] , \modmult_1/zin[0][167] ,
         \modmult_1/zin[0][166] , \modmult_1/zin[0][165] ,
         \modmult_1/zin[0][164] , \modmult_1/zin[0][163] ,
         \modmult_1/zin[0][162] , \modmult_1/zin[0][161] ,
         \modmult_1/zin[0][160] , \modmult_1/zin[0][159] ,
         \modmult_1/zin[0][158] , \modmult_1/zin[0][157] ,
         \modmult_1/zin[0][156] , \modmult_1/zin[0][155] ,
         \modmult_1/zin[0][154] , \modmult_1/zin[0][153] ,
         \modmult_1/zin[0][152] , \modmult_1/zin[0][151] ,
         \modmult_1/zin[0][150] , \modmult_1/zin[0][149] ,
         \modmult_1/zin[0][148] , \modmult_1/zin[0][147] ,
         \modmult_1/zin[0][146] , \modmult_1/zin[0][145] ,
         \modmult_1/zin[0][144] , \modmult_1/zin[0][143] ,
         \modmult_1/zin[0][142] , \modmult_1/zin[0][141] ,
         \modmult_1/zin[0][140] , \modmult_1/zin[0][139] ,
         \modmult_1/zin[0][138] , \modmult_1/zin[0][137] ,
         \modmult_1/zin[0][136] , \modmult_1/zin[0][135] ,
         \modmult_1/zin[0][134] , \modmult_1/zin[0][133] ,
         \modmult_1/zin[0][132] , \modmult_1/zin[0][131] ,
         \modmult_1/zin[0][130] , \modmult_1/zin[0][129] ,
         \modmult_1/zin[0][128] , \modmult_1/zin[0][127] ,
         \modmult_1/zin[0][126] , \modmult_1/zin[0][125] ,
         \modmult_1/zin[0][124] , \modmult_1/zin[0][123] ,
         \modmult_1/zin[0][122] , \modmult_1/zin[0][121] ,
         \modmult_1/zin[0][120] , \modmult_1/zin[0][119] ,
         \modmult_1/zin[0][118] , \modmult_1/zin[0][117] ,
         \modmult_1/zin[0][116] , \modmult_1/zin[0][115] ,
         \modmult_1/zin[0][114] , \modmult_1/zin[0][113] ,
         \modmult_1/zin[0][112] , \modmult_1/zin[0][111] ,
         \modmult_1/zin[0][110] , \modmult_1/zin[0][109] ,
         \modmult_1/zin[0][108] , \modmult_1/zin[0][107] ,
         \modmult_1/zin[0][106] , \modmult_1/zin[0][105] ,
         \modmult_1/zin[0][104] , \modmult_1/zin[0][103] ,
         \modmult_1/zin[0][102] , \modmult_1/zin[0][101] ,
         \modmult_1/zin[0][100] , \modmult_1/zin[0][99] ,
         \modmult_1/zin[0][98] , \modmult_1/zin[0][97] ,
         \modmult_1/zin[0][96] , \modmult_1/zin[0][95] ,
         \modmult_1/zin[0][94] , \modmult_1/zin[0][93] ,
         \modmult_1/zin[0][92] , \modmult_1/zin[0][91] ,
         \modmult_1/zin[0][90] , \modmult_1/zin[0][89] ,
         \modmult_1/zin[0][88] , \modmult_1/zin[0][87] ,
         \modmult_1/zin[0][86] , \modmult_1/zin[0][85] ,
         \modmult_1/zin[0][84] , \modmult_1/zin[0][83] ,
         \modmult_1/zin[0][82] , \modmult_1/zin[0][81] ,
         \modmult_1/zin[0][80] , \modmult_1/zin[0][79] ,
         \modmult_1/zin[0][78] , \modmult_1/zin[0][77] ,
         \modmult_1/zin[0][76] , \modmult_1/zin[0][75] ,
         \modmult_1/zin[0][74] , \modmult_1/zin[0][73] ,
         \modmult_1/zin[0][72] , \modmult_1/zin[0][71] ,
         \modmult_1/zin[0][70] , \modmult_1/zin[0][69] ,
         \modmult_1/zin[0][68] , \modmult_1/zin[0][67] ,
         \modmult_1/zin[0][66] , \modmult_1/zin[0][65] ,
         \modmult_1/zin[0][64] , \modmult_1/zin[0][63] ,
         \modmult_1/zin[0][62] , \modmult_1/zin[0][61] ,
         \modmult_1/zin[0][60] , \modmult_1/zin[0][59] ,
         \modmult_1/zin[0][58] , \modmult_1/zin[0][57] ,
         \modmult_1/zin[0][56] , \modmult_1/zin[0][55] ,
         \modmult_1/zin[0][54] , \modmult_1/zin[0][53] ,
         \modmult_1/zin[0][52] , \modmult_1/zin[0][51] ,
         \modmult_1/zin[0][50] , \modmult_1/zin[0][49] ,
         \modmult_1/zin[0][48] , \modmult_1/zin[0][47] ,
         \modmult_1/zin[0][46] , \modmult_1/zin[0][45] ,
         \modmult_1/zin[0][44] , \modmult_1/zin[0][43] ,
         \modmult_1/zin[0][42] , \modmult_1/zin[0][41] ,
         \modmult_1/zin[0][40] , \modmult_1/zin[0][39] ,
         \modmult_1/zin[0][38] , \modmult_1/zin[0][37] ,
         \modmult_1/zin[0][36] , \modmult_1/zin[0][35] ,
         \modmult_1/zin[0][34] , \modmult_1/zin[0][33] ,
         \modmult_1/zin[0][32] , \modmult_1/zin[0][31] ,
         \modmult_1/zin[0][30] , \modmult_1/zin[0][29] ,
         \modmult_1/zin[0][28] , \modmult_1/zin[0][27] ,
         \modmult_1/zin[0][26] , \modmult_1/zin[0][25] ,
         \modmult_1/zin[0][24] , \modmult_1/zin[0][23] ,
         \modmult_1/zin[0][22] , \modmult_1/zin[0][21] ,
         \modmult_1/zin[0][20] , \modmult_1/zin[0][19] ,
         \modmult_1/zin[0][18] , \modmult_1/zin[0][17] ,
         \modmult_1/zin[0][16] , \modmult_1/zin[0][15] ,
         \modmult_1/zin[0][14] , \modmult_1/zin[0][13] ,
         \modmult_1/zin[0][12] , \modmult_1/zin[0][11] ,
         \modmult_1/zin[0][10] , \modmult_1/zin[0][9] , \modmult_1/zin[0][8] ,
         \modmult_1/zin[0][7] , \modmult_1/zin[0][6] , \modmult_1/zin[0][5] ,
         \modmult_1/zin[0][4] , \modmult_1/zin[0][3] , \modmult_1/zin[0][2] ,
         \modmult_1/zin[0][1] , \modmult_1/zin[0][0] ,
         \modmult_1/zout[0][1024] , n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
         n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
         n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
         n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
         n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
         n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
         n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
         n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
         n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575,
         n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
         n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
         n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
         n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
         n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
         n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
         n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
         n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839,
         n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911,
         n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
         n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
         n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
         n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
         n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
         n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
         n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
         n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111,
         n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
         n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
         n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
         n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295,
         n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
         n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
         n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
         n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
         n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
         n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
         n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
         n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111,
         n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
         n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
         n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135,
         n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
         n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183,
         n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
         n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
         n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
         n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
         n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
         n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
         n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
         n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
         n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
         n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
         n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
         n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
         n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
         n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407,
         n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
         n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
         n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
         n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479,
         n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
         n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495,
         n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
         n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
         n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519,
         n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527,
         n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535,
         n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543,
         n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
         n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
         n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567,
         n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
         n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
         n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
         n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
         n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
         n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615,
         n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623,
         n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
         n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639,
         n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
         n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
         n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
         n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
         n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695,
         n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
         n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711,
         n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
         n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727,
         n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
         n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
         n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
         n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759,
         n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767,
         n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
         n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783,
         n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
         n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
         n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807,
         n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
         n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
         n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831,
         n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
         n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
         n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
         n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
         n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
         n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903,
         n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911,
         n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
         n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
         n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
         n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943,
         n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
         n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
         n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967,
         n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975,
         n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
         n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
         n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
         n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
         n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
         n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023,
         n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
         n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
         n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
         n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055,
         n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
         n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
         n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
         n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
         n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095,
         n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
         n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
         n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119,
         n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127,
         n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
         n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
         n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
         n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
         n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
         n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
         n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
         n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191,
         n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
         n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
         n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
         n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
         n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
         n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
         n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
         n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255,
         n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263,
         n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271,
         n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
         n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287,
         n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
         n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
         n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
         n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319,
         n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327,
         n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335,
         n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343,
         n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
         n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359,
         n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
         n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
         n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383,
         n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391,
         n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399,
         n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
         n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415,
         n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
         n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431,
         n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
         n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
         n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455,
         n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463,
         n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
         n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
         n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
         n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551,
         n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
         n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
         n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
         n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
         n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599,
         n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
         n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
         n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623,
         n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
         n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
         n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
         n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
         n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
         n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
         n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
         n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
         n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703,
         n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
         n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
         n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
         n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815,
         n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
         n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031,
         n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
         n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
         n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055,
         n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
         n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
         n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
         n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
         n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
         n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
         n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
         n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
         n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
         n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
         n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
         n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
         n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
         n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
         n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
         n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
         n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
         n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
         n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
         n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
         n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
         n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
         n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487,
         n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
         n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
         n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511,
         n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
         n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
         n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535,
         n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
         n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551,
         n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
         n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567,
         n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
         n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583,
         n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
         n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
         n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607,
         n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615,
         n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
         n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
         n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639,
         n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
         n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655,
         n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
         n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
         n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679,
         n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687,
         n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
         n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703,
         n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711,
         n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
         n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727,
         n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
         n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
         n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751,
         n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
         n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
         n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775,
         n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
         n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
         n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
         n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
         n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823,
         n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831,
         n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
         n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847,
         n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855,
         n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
         n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871,
         n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
         n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
         n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895,
         n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903,
         n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
         n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
         n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927,
         n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
         n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
         n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
         n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959,
         n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967,
         n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
         n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
         n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
         n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
         n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
         n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015,
         n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
         n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031,
         n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039,
         n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
         n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055,
         n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
         n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071,
         n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
         n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
         n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
         n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
         n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111,
         n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
         n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
         n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135,
         n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143,
         n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
         n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159,
         n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
         n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175,
         n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183,
         n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
         n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
         n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207,
         n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
         n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
         n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
         n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
         n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247,
         n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255,
         n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263,
         n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
         n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279,
         n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
         n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
         n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303,
         n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
         n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
         n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
         n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
         n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
         n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
         n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375,
         n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
         n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
         n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399,
         n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
         n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
         n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
         n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
         n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
         n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447,
         n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
         n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463,
         n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471,
         n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479,
         n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487,
         n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
         n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503,
         n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
         n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519,
         n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
         n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535,
         n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543,
         n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
         n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
         n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
         n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575,
         n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
         n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591,
         n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
         n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
         n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
         n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
         n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
         n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
         n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647,
         n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
         n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663,
         n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
         n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
         n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
         n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
         n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
         n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
         n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
         n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
         n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735,
         n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
         n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
         n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759,
         n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
         n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
         n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
         n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
         n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
         n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807,
         n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
         n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
         n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
         n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
         n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
         n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855,
         n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863,
         n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
         n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879,
         n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
         n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
         n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
         n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
         n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
         n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927,
         n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
         n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
         n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
         n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
         n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
         n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
         n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
         n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
         n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999,
         n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
         n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
         n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023,
         n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
         n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
         n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
         n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
         n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
         n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
         n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
         n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
         n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095,
         n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
         n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
         n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
         n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
         n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
         n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
         n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
         n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
         n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
         n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
         n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
         n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191,
         n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
         n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
         n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
         n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
         n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
         n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239,
         n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
         n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
         n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
         n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
         n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
         n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
         n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
         n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
         n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
         n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
         n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335,
         n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
         n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
         n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359,
         n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
         n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
         n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
         n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
         n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
         n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407,
         n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
         n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
         n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431,
         n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
         n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
         n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455,
         n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
         n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
         n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
         n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
         n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
         n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503,
         n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
         n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
         n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527,
         n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
         n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
         n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
         n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
         n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
         n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575,
         n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
         n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
         n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599,
         n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
         n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
         n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623,
         n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
         n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
         n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
         n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
         n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
         n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
         n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
         n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
         n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
         n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
         n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
         n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
         n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
         n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
         n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743,
         n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
         n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
         n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767,
         n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
         n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
         n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
         n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
         n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
         n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
         n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
         n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
         n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
         n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
         n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
         n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
         n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
         n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
         n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
         n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
         n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
         n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
         n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
         n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
         n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999,
         n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007,
         n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015,
         n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023,
         n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031,
         n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039,
         n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047,
         n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055,
         n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
         n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071,
         n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079,
         n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
         n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
         n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103,
         n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
         n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119,
         n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127,
         n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135,
         n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143,
         n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151,
         n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159,
         n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
         n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175,
         n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
         n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191,
         n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199,
         n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207,
         n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215,
         n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223,
         n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231,
         n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
         n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247,
         n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
         n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263,
         n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271,
         n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279,
         n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287,
         n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295,
         n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303,
         n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
         n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319,
         n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
         n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
         n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343,
         n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351,
         n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359,
         n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367,
         n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
         n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
         n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
         n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415,
         n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423,
         n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431,
         n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439,
         n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
         n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455,
         n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463,
         n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471,
         n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479,
         n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487,
         n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495,
         n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503,
         n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511,
         n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519,
         n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
         n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535,
         n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
         n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
         n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559,
         n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567,
         n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575,
         n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583,
         n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591,
         n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599,
         n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607,
         n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615,
         n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623,
         n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631,
         n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639,
         n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647,
         n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655,
         n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
         n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
         n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679,
         n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
         n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
         n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703,
         n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
         n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719,
         n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727,
         n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
         n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
         n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751,
         n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
         n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767,
         n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775,
         n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783,
         n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
         n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799,
         n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807,
         n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
         n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823,
         n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
         n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839,
         n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847,
         n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
         n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863,
         n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871,
         n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879,
         n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
         n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895,
         n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
         n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
         n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919,
         n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927,
         n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935,
         n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
         n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951,
         n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
         n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967,
         n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
         n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983,
         n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991,
         n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
         n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
         n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
         n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
         n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
         n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039,
         n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
         n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
         n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063,
         n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071,
         n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
         n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087,
         n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095,
         n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
         n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111,
         n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
         n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127,
         n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
         n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
         n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
         n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159,
         n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167,
         n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
         n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183,
         n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
         n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
         n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207,
         n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215,
         n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
         n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231,
         n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239,
         n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
         n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255,
         n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263,
         n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271,
         n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279,
         n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287,
         n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295,
         n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303,
         n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311,
         n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319,
         n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327,
         n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
         n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343,
         n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351,
         n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359,
         n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
         n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375,
         n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383,
         n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
         n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399,
         n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407,
         n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415,
         n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423,
         n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431,
         n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439,
         n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447,
         n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455,
         n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463,
         n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471,
         n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
         n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
         n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495,
         n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503,
         n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511,
         n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519,
         n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527,
         n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
         n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543,
         n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
         n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559,
         n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567,
         n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575,
         n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583,
         n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591,
         n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599,
         n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
         n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615,
         n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623,
         n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631,
         n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639,
         n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647,
         n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655,
         n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663,
         n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671,
         n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
         n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687,
         n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695,
         n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703,
         n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711,
         n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719,
         n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727,
         n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735,
         n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743,
         n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
         n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759,
         n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767,
         n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775,
         n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783,
         n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791,
         n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799,
         n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807,
         n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815,
         n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823,
         n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831,
         n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839,
         n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847,
         n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855,
         n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
         n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871,
         n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879,
         n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887,
         n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
         n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903,
         n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
         n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
         n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927,
         n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
         n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
         n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
         n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959,
         n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
         n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975,
         n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
         n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991,
         n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999,
         n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
         n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
         n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023,
         n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031,
         n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
         n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047,
         n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
         n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063,
         n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
         n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
         n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
         n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095,
         n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103,
         n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
         n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119,
         n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
         n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
         n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143,
         n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
         n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
         n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167,
         n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175,
         n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
         n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191,
         n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
         n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
         n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215,
         n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
         n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
         n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239,
         n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247,
         n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
         n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263,
         n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
         n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
         n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287,
         n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
         n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303,
         n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311,
         n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
         n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
         n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335,
         n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
         n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
         n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359,
         n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
         n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375,
         n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383,
         n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391,
         n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
         n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407,
         n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
         n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
         n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431,
         n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
         n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447,
         n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455,
         n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
         n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
         n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479,
         n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
         n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495,
         n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503,
         n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
         n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
         n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527,
         n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535,
         n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
         n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551,
         n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
         n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
         n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575,
         n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
         n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
         n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599,
         n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
         n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
         n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623,
         n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
         n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
         n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
         n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
         n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
         n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671,
         n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
         n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
         n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695,
         n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
         n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
         n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
         n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
         n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
         n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743,
         n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751,
         n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
         n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767,
         n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
         n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783,
         n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791,
         n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
         n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807,
         n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815,
         n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823,
         n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
         n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
         n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
         n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
         n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863,
         n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871,
         n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
         n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887,
         n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895,
         n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
         n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911,
         n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
         n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927,
         n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935,
         n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
         n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951,
         n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959,
         n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967,
         n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
         n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983,
         n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
         n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999,
         n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
         n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
         n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023,
         n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
         n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039,
         n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
         n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055,
         n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
         n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071,
         n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079,
         n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
         n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095,
         n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103,
         n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111,
         n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
         n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
         n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
         n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
         n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
         n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
         n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
         n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
         n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
         n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
         n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199,
         n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
         n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215,
         n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223,
         n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
         n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
         n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247,
         n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255,
         n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
         n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271,
         n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
         n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287,
         n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295,
         n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303,
         n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
         n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319,
         n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327,
         n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
         n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343,
         n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
         n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359,
         n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367,
         n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
         n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
         n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
         n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399,
         n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
         n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415,
         n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
         n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431,
         n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439,
         n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447,
         n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
         n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463,
         n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471,
         n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
         n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487,
         n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
         n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
         n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511,
         n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
         n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527,
         n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535,
         n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543,
         n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
         n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559,
         n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
         n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
         n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583,
         n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
         n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599,
         n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607,
         n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
         n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
         n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631,
         n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
         n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647,
         n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655,
         n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663,
         n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671,
         n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679,
         n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687,
         n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
         n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703,
         n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
         n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719,
         n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727,
         n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735,
         n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743,
         n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751,
         n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
         n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
         n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775,
         n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
         n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
         n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799,
         n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807,
         n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815,
         n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823,
         n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831,
         n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
         n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847,
         n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
         n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863,
         n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871,
         n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879,
         n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887,
         n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895,
         n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
         n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
         n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919,
         n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
         n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935,
         n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943,
         n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951,
         n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
         n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967,
         n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
         n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
         n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991,
         n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
         n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007,
         n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015,
         n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
         n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
         n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
         n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047,
         n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
         n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063,
         n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
         n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
         n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087,
         n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095,
         n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
         n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111,
         n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119,
         n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127,
         n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135,
         n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143,
         n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151,
         n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159,
         n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167,
         n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175,
         n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183,
         n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191,
         n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199,
         n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207,
         n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
         n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223,
         n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231,
         n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239,
         n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247,
         n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255,
         n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263,
         n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
         n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279,
         n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
         n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295,
         n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303,
         n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311,
         n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319,
         n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327,
         n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335,
         n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343,
         n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351,
         n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359,
         n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367,
         n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375,
         n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383,
         n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391,
         n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399,
         n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407,
         n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415,
         n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423,
         n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431,
         n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439,
         n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447,
         n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455,
         n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
         n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471,
         n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479,
         n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487,
         n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495,
         n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
         n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511,
         n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519,
         n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
         n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
         n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543,
         n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551,
         n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
         n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567,
         n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
         n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583,
         n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591,
         n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599,
         n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
         n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615,
         n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623,
         n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
         n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
         n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
         n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655,
         n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663,
         n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671,
         n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679,
         n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687,
         n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695,
         n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
         n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711,
         n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719,
         n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727,
         n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735,
         n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
         n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751,
         n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759,
         n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767,
         n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775,
         n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783,
         n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791,
         n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799,
         n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807,
         n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815,
         n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823,
         n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831,
         n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839,
         n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
         n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855,
         n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863,
         n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871,
         n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879,
         n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887,
         n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895,
         n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903,
         n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911,
         n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
         n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927,
         n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935,
         n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943,
         n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951,
         n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
         n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967,
         n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975,
         n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983,
         n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
         n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999,
         n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007,
         n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015,
         n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023,
         n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031,
         n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039,
         n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047,
         n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055,
         n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
         n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071,
         n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079,
         n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087,
         n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095,
         n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103,
         n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111,
         n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119,
         n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127,
         n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
         n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143,
         n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151,
         n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159,
         n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167,
         n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175,
         n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183,
         n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191,
         n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199,
         n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
         n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215,
         n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223,
         n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231,
         n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239,
         n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247,
         n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255,
         n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263,
         n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271,
         n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
         n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287,
         n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
         n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303,
         n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311,
         n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
         n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327,
         n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335,
         n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343,
         n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
         n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359,
         n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367,
         n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375,
         n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383,
         n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
         n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399,
         n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407,
         n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415,
         n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
         n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431,
         n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439,
         n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447,
         n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455,
         n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463,
         n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471,
         n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479,
         n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487,
         n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495,
         n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503,
         n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511,
         n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519,
         n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
         n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535,
         n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543,
         n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551,
         n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559,
         n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567,
         n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575,
         n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583,
         n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
         n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599,
         n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607,
         n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615,
         n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623,
         n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631,
         n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
         n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647,
         n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
         n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
         n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671,
         n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679,
         n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687,
         n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695,
         n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703,
         n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711,
         n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719,
         n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
         n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735,
         n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743,
         n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751,
         n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759,
         n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767,
         n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775,
         n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
         n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791,
         n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799,
         n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807,
         n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815,
         n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823,
         n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831,
         n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839,
         n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847,
         n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
         n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863,
         n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871,
         n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879,
         n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887,
         n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895,
         n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903,
         n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911,
         n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919,
         n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
         n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935,
         n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
         n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951,
         n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959,
         n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967,
         n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
         n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983,
         n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
         n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
         n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007,
         n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
         n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023,
         n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031,
         n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039,
         n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047,
         n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055,
         n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063,
         n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
         n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079,
         n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
         n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
         n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103,
         n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111,
         n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
         n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127,
         n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135,
         n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
         n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151,
         n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
         n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167,
         n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175,
         n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
         n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191,
         n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199,
         n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207,
         n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
         n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223,
         n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
         n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239,
         n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247,
         n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
         n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263,
         n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271,
         n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279,
         n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287,
         n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295,
         n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
         n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
         n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319,
         n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327,
         n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335,
         n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343,
         n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351,
         n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359,
         n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367,
         n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
         n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383,
         n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391,
         n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399,
         n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407,
         n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415,
         n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423,
         n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
         n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439,
         n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
         n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455,
         n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463,
         n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471,
         n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479,
         n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487,
         n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495,
         n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
         n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511,
         n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519,
         n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527,
         n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535,
         n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543,
         n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551,
         n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559,
         n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567,
         n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
         n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583,
         n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591,
         n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599,
         n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607,
         n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615,
         n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623,
         n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631,
         n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639,
         n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
         n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655,
         n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663,
         n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671,
         n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679,
         n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687,
         n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695,
         n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703,
         n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711,
         n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
         n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727,
         n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735,
         n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743,
         n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751,
         n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759,
         n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767,
         n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775,
         n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783,
         n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
         n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799,
         n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
         n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815,
         n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823,
         n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831,
         n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839,
         n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847,
         n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855,
         n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
         n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871,
         n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879,
         n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887,
         n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895,
         n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903,
         n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911,
         n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919,
         n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927,
         n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
         n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943,
         n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951,
         n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959,
         n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967,
         n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
         n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983,
         n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991,
         n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
         n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
         n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015,
         n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
         n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
         n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039,
         n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
         n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055,
         n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063,
         n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071,
         n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
         n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087,
         n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
         n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103,
         n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111,
         n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
         n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127,
         n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135,
         n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143,
         n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
         n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159,
         n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167,
         n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175,
         n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183,
         n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
         n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199,
         n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207,
         n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215,
         n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
         n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231,
         n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239,
         n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247,
         n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255,
         n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263,
         n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271,
         n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279,
         n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
         n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
         n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303,
         n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
         n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319,
         n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327,
         n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335,
         n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343,
         n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351,
         n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359,
         n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367,
         n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375,
         n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383,
         n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391,
         n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399,
         n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
         n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415,
         n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423,
         n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431,
         n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439,
         n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447,
         n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
         n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463,
         n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471,
         n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
         n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487,
         n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495,
         n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503,
         n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511,
         n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519,
         n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527,
         n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
         n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543,
         n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551,
         n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559,
         n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567,
         n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575,
         n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583,
         n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591,
         n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
         n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607,
         n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615,
         n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623,
         n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631,
         n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639,
         n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647,
         n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
         n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663,
         n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671,
         n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679,
         n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687,
         n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695,
         n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703,
         n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711,
         n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719,
         n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
         n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735,
         n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743,
         n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
         n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759,
         n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767,
         n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775,
         n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783,
         n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791,
         n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799,
         n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807,
         n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815,
         n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823,
         n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831,
         n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839,
         n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847,
         n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855,
         n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863,
         n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871,
         n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879,
         n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887,
         n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895,
         n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903,
         n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911,
         n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919,
         n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927,
         n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935,
         n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943,
         n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951,
         n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
         n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
         n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975,
         n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983,
         n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991,
         n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999,
         n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007,
         n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
         n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023,
         n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
         n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
         n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047,
         n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055,
         n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063,
         n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071,
         n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079,
         n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087,
         n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095,
         n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
         n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111,
         n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119,
         n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127,
         n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135,
         n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143,
         n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151,
         n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159,
         n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167,
         n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
         n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183,
         n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191,
         n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199,
         n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207,
         n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215,
         n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223,
         n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
         n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239,
         n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
         n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255,
         n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263,
         n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271,
         n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279,
         n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287,
         n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295,
         n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303,
         n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311,
         n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
         n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327,
         n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335,
         n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343,
         n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351,
         n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359,
         n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367,
         n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375,
         n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383,
         n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
         n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399,
         n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407,
         n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415,
         n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423,
         n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431,
         n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439,
         n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447,
         n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455,
         n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
         n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471,
         n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479,
         n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487,
         n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495,
         n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503,
         n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511,
         n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
         n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527,
         n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
         n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543,
         n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551,
         n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559,
         n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567,
         n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575,
         n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583,
         n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591,
         n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599,
         n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607,
         n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615,
         n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623,
         n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631,
         n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639,
         n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647,
         n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655,
         n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663,
         n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
         n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679,
         n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687,
         n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695,
         n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703,
         n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711,
         n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719,
         n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727,
         n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
         n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743,
         n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751,
         n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759,
         n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767,
         n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775,
         n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783,
         n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791,
         n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799,
         n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
         n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815,
         n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823,
         n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831,
         n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839,
         n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
         n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855,
         n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863,
         n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871,
         n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879,
         n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887,
         n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895,
         n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903,
         n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911,
         n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919,
         n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927,
         n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935,
         n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943,
         n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951,
         n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959,
         n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967,
         n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
         n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983,
         n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991,
         n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999,
         n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007,
         n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015,
         n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023,
         n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031,
         n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
         n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047,
         n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055,
         n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063,
         n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071,
         n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079,
         n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087,
         n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095,
         n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103,
         n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
         n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119,
         n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127,
         n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135,
         n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143,
         n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151,
         n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159,
         n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
         n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175,
         n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183,
         n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191,
         n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199,
         n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207,
         n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215,
         n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223,
         n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231,
         n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
         n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247,
         n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255,
         n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263,
         n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271,
         n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279,
         n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287,
         n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295,
         n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303,
         n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311,
         n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319,
         n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327,
         n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335,
         n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343,
         n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351,
         n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359,
         n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367,
         n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375,
         n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
         n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391,
         n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
         n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407,
         n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415,
         n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
         n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431,
         n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439,
         n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447,
         n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
         n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463,
         n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
         n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
         n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487,
         n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
         n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503,
         n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511,
         n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519,
         n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
         n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535,
         n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
         n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551,
         n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559,
         n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567,
         n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575,
         n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583,
         n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591,
         n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
         n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607,
         n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615,
         n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623,
         n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631,
         n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639,
         n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647,
         n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655,
         n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663,
         n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671,
         n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679,
         n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687,
         n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695,
         n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703,
         n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711,
         n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719,
         n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727,
         n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735,
         n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743,
         n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751,
         n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759,
         n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767,
         n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775,
         n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783,
         n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791,
         n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799,
         n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807,
         n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815,
         n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823,
         n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831,
         n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839,
         n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847,
         n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855,
         n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863,
         n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871,
         n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879,
         n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887,
         n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895,
         n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903,
         n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911,
         n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919,
         n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927,
         n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935,
         n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943,
         n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951,
         n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959,
         n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967,
         n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975,
         n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983,
         n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991;
  wire   [1023:0] start_in;
  wire   [1023:0] ein;
  wire   [1023:0] creg_next;
  wire   [1023:0] o;
  wire   [1023:0] ereg_next;

  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(start_in[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(start_in[1023]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(e[256]), 
        .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(e[257]), 
        .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(e[258]), 
        .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(e[259]), 
        .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(e[260]), 
        .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(e[261]), 
        .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(e[262]), 
        .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(e[263]), 
        .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(e[264]), 
        .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(e[265]), 
        .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(e[266]), 
        .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(e[267]), 
        .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(e[268]), 
        .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(e[269]), 
        .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(e[270]), 
        .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(e[271]), 
        .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(e[272]), 
        .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(e[273]), 
        .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(e[274]), 
        .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(e[275]), 
        .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(e[276]), 
        .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(e[277]), 
        .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(e[278]), 
        .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(e[279]), 
        .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(e[280]), 
        .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(e[281]), 
        .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(e[282]), 
        .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(e[283]), 
        .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(e[284]), 
        .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(e[285]), 
        .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(e[286]), 
        .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(e[287]), 
        .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(e[288]), 
        .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(e[289]), 
        .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(e[290]), 
        .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(e[291]), 
        .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(e[292]), 
        .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(e[293]), 
        .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(e[294]), 
        .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(e[295]), 
        .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(e[296]), 
        .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(e[297]), 
        .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(e[298]), 
        .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(e[299]), 
        .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(e[300]), 
        .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(e[301]), 
        .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(e[302]), 
        .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(e[303]), 
        .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(e[304]), 
        .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(e[305]), 
        .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(e[306]), 
        .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(e[307]), 
        .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(e[308]), 
        .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(e[309]), 
        .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(e[310]), 
        .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(e[311]), 
        .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(e[312]), 
        .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(e[313]), 
        .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(e[314]), 
        .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(e[315]), 
        .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(e[316]), 
        .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(e[317]), 
        .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(e[318]), 
        .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(e[319]), 
        .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(e[320]), 
        .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(e[321]), 
        .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(e[322]), 
        .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(e[323]), 
        .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(e[324]), 
        .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(e[325]), 
        .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(e[326]), 
        .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(e[327]), 
        .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(e[328]), 
        .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(e[329]), 
        .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(e[330]), 
        .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(e[331]), 
        .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(e[332]), 
        .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(e[333]), 
        .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(e[334]), 
        .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(e[335]), 
        .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(e[336]), 
        .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(e[337]), 
        .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(e[338]), 
        .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(e[339]), 
        .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(e[340]), 
        .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(e[341]), 
        .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(e[342]), 
        .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(e[343]), 
        .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(e[344]), 
        .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(e[345]), 
        .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(e[346]), 
        .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(e[347]), 
        .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(e[348]), 
        .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(e[349]), 
        .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(e[350]), 
        .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(e[351]), 
        .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(e[352]), 
        .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(e[353]), 
        .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(e[354]), 
        .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(e[355]), 
        .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(e[356]), 
        .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(e[357]), 
        .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(e[358]), 
        .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(e[359]), 
        .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(e[360]), 
        .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(e[361]), 
        .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(e[362]), 
        .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(e[363]), 
        .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(e[364]), 
        .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(e[365]), 
        .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(e[366]), 
        .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(e[367]), 
        .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(e[368]), 
        .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(e[369]), 
        .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(e[370]), 
        .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(e[371]), 
        .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(e[372]), 
        .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(e[373]), 
        .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(e[374]), 
        .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(e[375]), 
        .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(e[376]), 
        .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(e[377]), 
        .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(e[378]), 
        .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(e[379]), 
        .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(e[380]), 
        .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(e[381]), 
        .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(e[382]), 
        .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(e[383]), 
        .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(e[384]), 
        .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(e[385]), 
        .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(e[386]), 
        .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(e[387]), 
        .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(e[388]), 
        .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(e[389]), 
        .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(e[390]), 
        .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(e[391]), 
        .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(e[392]), 
        .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(e[393]), 
        .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(e[394]), 
        .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(e[395]), 
        .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(e[396]), 
        .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(e[397]), 
        .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(e[398]), 
        .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(e[399]), 
        .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(e[400]), 
        .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(e[401]), 
        .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(e[402]), 
        .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(e[403]), 
        .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(e[404]), 
        .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(e[405]), 
        .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(e[406]), 
        .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(e[407]), 
        .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(e[408]), 
        .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(e[409]), 
        .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(e[410]), 
        .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(e[411]), 
        .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(e[412]), 
        .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(e[413]), 
        .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(e[414]), 
        .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(e[415]), 
        .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(e[416]), 
        .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(e[417]), 
        .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(e[418]), 
        .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(e[419]), 
        .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(e[420]), 
        .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(e[421]), 
        .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(e[422]), 
        .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(e[423]), 
        .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(e[424]), 
        .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(e[425]), 
        .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(e[426]), 
        .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(e[427]), 
        .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(e[428]), 
        .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(e[429]), 
        .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(e[430]), 
        .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(e[431]), 
        .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(e[432]), 
        .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(e[433]), 
        .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(e[434]), 
        .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(e[435]), 
        .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(e[436]), 
        .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(e[437]), 
        .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(e[438]), 
        .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(e[439]), 
        .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(e[440]), 
        .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(e[441]), 
        .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(e[442]), 
        .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(e[443]), 
        .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(e[444]), 
        .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(e[445]), 
        .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(e[446]), 
        .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(e[447]), 
        .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(e[448]), 
        .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(e[449]), 
        .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(e[450]), 
        .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(e[451]), 
        .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(e[452]), 
        .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(e[453]), 
        .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(e[454]), 
        .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(e[455]), 
        .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(e[456]), 
        .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(e[457]), 
        .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(e[458]), 
        .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(e[459]), 
        .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(e[460]), 
        .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(e[461]), 
        .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(e[462]), 
        .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(e[463]), 
        .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(e[464]), 
        .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(e[465]), 
        .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(e[466]), 
        .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(e[467]), 
        .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(e[468]), 
        .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(e[469]), 
        .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(e[470]), 
        .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(e[471]), 
        .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(e[472]), 
        .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(e[473]), 
        .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(e[474]), 
        .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(e[475]), 
        .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(e[476]), 
        .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(e[477]), 
        .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(e[478]), 
        .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(e[479]), 
        .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(e[480]), 
        .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(e[481]), 
        .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(e[482]), 
        .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(e[483]), 
        .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(e[484]), 
        .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(e[485]), 
        .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(e[486]), 
        .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(e[487]), 
        .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(e[488]), 
        .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(e[489]), 
        .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(e[490]), 
        .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(e[491]), 
        .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(e[492]), 
        .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(e[493]), 
        .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(e[494]), 
        .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(e[495]), 
        .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(e[496]), 
        .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(e[497]), 
        .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(e[498]), 
        .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(e[499]), 
        .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(e[500]), 
        .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(e[501]), 
        .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(e[502]), 
        .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(e[503]), 
        .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(e[504]), 
        .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(e[505]), 
        .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(e[506]), 
        .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(e[507]), 
        .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(e[508]), 
        .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(e[509]), 
        .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(e[510]), 
        .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(e[511]), 
        .Q(ein[511]) );
  DFF \ereg_reg[512]  ( .D(ereg_next[512]), .CLK(clk), .RST(rst), .I(e[512]), 
        .Q(ein[512]) );
  DFF \ereg_reg[513]  ( .D(ereg_next[513]), .CLK(clk), .RST(rst), .I(e[513]), 
        .Q(ein[513]) );
  DFF \ereg_reg[514]  ( .D(ereg_next[514]), .CLK(clk), .RST(rst), .I(e[514]), 
        .Q(ein[514]) );
  DFF \ereg_reg[515]  ( .D(ereg_next[515]), .CLK(clk), .RST(rst), .I(e[515]), 
        .Q(ein[515]) );
  DFF \ereg_reg[516]  ( .D(ereg_next[516]), .CLK(clk), .RST(rst), .I(e[516]), 
        .Q(ein[516]) );
  DFF \ereg_reg[517]  ( .D(ereg_next[517]), .CLK(clk), .RST(rst), .I(e[517]), 
        .Q(ein[517]) );
  DFF \ereg_reg[518]  ( .D(ereg_next[518]), .CLK(clk), .RST(rst), .I(e[518]), 
        .Q(ein[518]) );
  DFF \ereg_reg[519]  ( .D(ereg_next[519]), .CLK(clk), .RST(rst), .I(e[519]), 
        .Q(ein[519]) );
  DFF \ereg_reg[520]  ( .D(ereg_next[520]), .CLK(clk), .RST(rst), .I(e[520]), 
        .Q(ein[520]) );
  DFF \ereg_reg[521]  ( .D(ereg_next[521]), .CLK(clk), .RST(rst), .I(e[521]), 
        .Q(ein[521]) );
  DFF \ereg_reg[522]  ( .D(ereg_next[522]), .CLK(clk), .RST(rst), .I(e[522]), 
        .Q(ein[522]) );
  DFF \ereg_reg[523]  ( .D(ereg_next[523]), .CLK(clk), .RST(rst), .I(e[523]), 
        .Q(ein[523]) );
  DFF \ereg_reg[524]  ( .D(ereg_next[524]), .CLK(clk), .RST(rst), .I(e[524]), 
        .Q(ein[524]) );
  DFF \ereg_reg[525]  ( .D(ereg_next[525]), .CLK(clk), .RST(rst), .I(e[525]), 
        .Q(ein[525]) );
  DFF \ereg_reg[526]  ( .D(ereg_next[526]), .CLK(clk), .RST(rst), .I(e[526]), 
        .Q(ein[526]) );
  DFF \ereg_reg[527]  ( .D(ereg_next[527]), .CLK(clk), .RST(rst), .I(e[527]), 
        .Q(ein[527]) );
  DFF \ereg_reg[528]  ( .D(ereg_next[528]), .CLK(clk), .RST(rst), .I(e[528]), 
        .Q(ein[528]) );
  DFF \ereg_reg[529]  ( .D(ereg_next[529]), .CLK(clk), .RST(rst), .I(e[529]), 
        .Q(ein[529]) );
  DFF \ereg_reg[530]  ( .D(ereg_next[530]), .CLK(clk), .RST(rst), .I(e[530]), 
        .Q(ein[530]) );
  DFF \ereg_reg[531]  ( .D(ereg_next[531]), .CLK(clk), .RST(rst), .I(e[531]), 
        .Q(ein[531]) );
  DFF \ereg_reg[532]  ( .D(ereg_next[532]), .CLK(clk), .RST(rst), .I(e[532]), 
        .Q(ein[532]) );
  DFF \ereg_reg[533]  ( .D(ereg_next[533]), .CLK(clk), .RST(rst), .I(e[533]), 
        .Q(ein[533]) );
  DFF \ereg_reg[534]  ( .D(ereg_next[534]), .CLK(clk), .RST(rst), .I(e[534]), 
        .Q(ein[534]) );
  DFF \ereg_reg[535]  ( .D(ereg_next[535]), .CLK(clk), .RST(rst), .I(e[535]), 
        .Q(ein[535]) );
  DFF \ereg_reg[536]  ( .D(ereg_next[536]), .CLK(clk), .RST(rst), .I(e[536]), 
        .Q(ein[536]) );
  DFF \ereg_reg[537]  ( .D(ereg_next[537]), .CLK(clk), .RST(rst), .I(e[537]), 
        .Q(ein[537]) );
  DFF \ereg_reg[538]  ( .D(ereg_next[538]), .CLK(clk), .RST(rst), .I(e[538]), 
        .Q(ein[538]) );
  DFF \ereg_reg[539]  ( .D(ereg_next[539]), .CLK(clk), .RST(rst), .I(e[539]), 
        .Q(ein[539]) );
  DFF \ereg_reg[540]  ( .D(ereg_next[540]), .CLK(clk), .RST(rst), .I(e[540]), 
        .Q(ein[540]) );
  DFF \ereg_reg[541]  ( .D(ereg_next[541]), .CLK(clk), .RST(rst), .I(e[541]), 
        .Q(ein[541]) );
  DFF \ereg_reg[542]  ( .D(ereg_next[542]), .CLK(clk), .RST(rst), .I(e[542]), 
        .Q(ein[542]) );
  DFF \ereg_reg[543]  ( .D(ereg_next[543]), .CLK(clk), .RST(rst), .I(e[543]), 
        .Q(ein[543]) );
  DFF \ereg_reg[544]  ( .D(ereg_next[544]), .CLK(clk), .RST(rst), .I(e[544]), 
        .Q(ein[544]) );
  DFF \ereg_reg[545]  ( .D(ereg_next[545]), .CLK(clk), .RST(rst), .I(e[545]), 
        .Q(ein[545]) );
  DFF \ereg_reg[546]  ( .D(ereg_next[546]), .CLK(clk), .RST(rst), .I(e[546]), 
        .Q(ein[546]) );
  DFF \ereg_reg[547]  ( .D(ereg_next[547]), .CLK(clk), .RST(rst), .I(e[547]), 
        .Q(ein[547]) );
  DFF \ereg_reg[548]  ( .D(ereg_next[548]), .CLK(clk), .RST(rst), .I(e[548]), 
        .Q(ein[548]) );
  DFF \ereg_reg[549]  ( .D(ereg_next[549]), .CLK(clk), .RST(rst), .I(e[549]), 
        .Q(ein[549]) );
  DFF \ereg_reg[550]  ( .D(ereg_next[550]), .CLK(clk), .RST(rst), .I(e[550]), 
        .Q(ein[550]) );
  DFF \ereg_reg[551]  ( .D(ereg_next[551]), .CLK(clk), .RST(rst), .I(e[551]), 
        .Q(ein[551]) );
  DFF \ereg_reg[552]  ( .D(ereg_next[552]), .CLK(clk), .RST(rst), .I(e[552]), 
        .Q(ein[552]) );
  DFF \ereg_reg[553]  ( .D(ereg_next[553]), .CLK(clk), .RST(rst), .I(e[553]), 
        .Q(ein[553]) );
  DFF \ereg_reg[554]  ( .D(ereg_next[554]), .CLK(clk), .RST(rst), .I(e[554]), 
        .Q(ein[554]) );
  DFF \ereg_reg[555]  ( .D(ereg_next[555]), .CLK(clk), .RST(rst), .I(e[555]), 
        .Q(ein[555]) );
  DFF \ereg_reg[556]  ( .D(ereg_next[556]), .CLK(clk), .RST(rst), .I(e[556]), 
        .Q(ein[556]) );
  DFF \ereg_reg[557]  ( .D(ereg_next[557]), .CLK(clk), .RST(rst), .I(e[557]), 
        .Q(ein[557]) );
  DFF \ereg_reg[558]  ( .D(ereg_next[558]), .CLK(clk), .RST(rst), .I(e[558]), 
        .Q(ein[558]) );
  DFF \ereg_reg[559]  ( .D(ereg_next[559]), .CLK(clk), .RST(rst), .I(e[559]), 
        .Q(ein[559]) );
  DFF \ereg_reg[560]  ( .D(ereg_next[560]), .CLK(clk), .RST(rst), .I(e[560]), 
        .Q(ein[560]) );
  DFF \ereg_reg[561]  ( .D(ereg_next[561]), .CLK(clk), .RST(rst), .I(e[561]), 
        .Q(ein[561]) );
  DFF \ereg_reg[562]  ( .D(ereg_next[562]), .CLK(clk), .RST(rst), .I(e[562]), 
        .Q(ein[562]) );
  DFF \ereg_reg[563]  ( .D(ereg_next[563]), .CLK(clk), .RST(rst), .I(e[563]), 
        .Q(ein[563]) );
  DFF \ereg_reg[564]  ( .D(ereg_next[564]), .CLK(clk), .RST(rst), .I(e[564]), 
        .Q(ein[564]) );
  DFF \ereg_reg[565]  ( .D(ereg_next[565]), .CLK(clk), .RST(rst), .I(e[565]), 
        .Q(ein[565]) );
  DFF \ereg_reg[566]  ( .D(ereg_next[566]), .CLK(clk), .RST(rst), .I(e[566]), 
        .Q(ein[566]) );
  DFF \ereg_reg[567]  ( .D(ereg_next[567]), .CLK(clk), .RST(rst), .I(e[567]), 
        .Q(ein[567]) );
  DFF \ereg_reg[568]  ( .D(ereg_next[568]), .CLK(clk), .RST(rst), .I(e[568]), 
        .Q(ein[568]) );
  DFF \ereg_reg[569]  ( .D(ereg_next[569]), .CLK(clk), .RST(rst), .I(e[569]), 
        .Q(ein[569]) );
  DFF \ereg_reg[570]  ( .D(ereg_next[570]), .CLK(clk), .RST(rst), .I(e[570]), 
        .Q(ein[570]) );
  DFF \ereg_reg[571]  ( .D(ereg_next[571]), .CLK(clk), .RST(rst), .I(e[571]), 
        .Q(ein[571]) );
  DFF \ereg_reg[572]  ( .D(ereg_next[572]), .CLK(clk), .RST(rst), .I(e[572]), 
        .Q(ein[572]) );
  DFF \ereg_reg[573]  ( .D(ereg_next[573]), .CLK(clk), .RST(rst), .I(e[573]), 
        .Q(ein[573]) );
  DFF \ereg_reg[574]  ( .D(ereg_next[574]), .CLK(clk), .RST(rst), .I(e[574]), 
        .Q(ein[574]) );
  DFF \ereg_reg[575]  ( .D(ereg_next[575]), .CLK(clk), .RST(rst), .I(e[575]), 
        .Q(ein[575]) );
  DFF \ereg_reg[576]  ( .D(ereg_next[576]), .CLK(clk), .RST(rst), .I(e[576]), 
        .Q(ein[576]) );
  DFF \ereg_reg[577]  ( .D(ereg_next[577]), .CLK(clk), .RST(rst), .I(e[577]), 
        .Q(ein[577]) );
  DFF \ereg_reg[578]  ( .D(ereg_next[578]), .CLK(clk), .RST(rst), .I(e[578]), 
        .Q(ein[578]) );
  DFF \ereg_reg[579]  ( .D(ereg_next[579]), .CLK(clk), .RST(rst), .I(e[579]), 
        .Q(ein[579]) );
  DFF \ereg_reg[580]  ( .D(ereg_next[580]), .CLK(clk), .RST(rst), .I(e[580]), 
        .Q(ein[580]) );
  DFF \ereg_reg[581]  ( .D(ereg_next[581]), .CLK(clk), .RST(rst), .I(e[581]), 
        .Q(ein[581]) );
  DFF \ereg_reg[582]  ( .D(ereg_next[582]), .CLK(clk), .RST(rst), .I(e[582]), 
        .Q(ein[582]) );
  DFF \ereg_reg[583]  ( .D(ereg_next[583]), .CLK(clk), .RST(rst), .I(e[583]), 
        .Q(ein[583]) );
  DFF \ereg_reg[584]  ( .D(ereg_next[584]), .CLK(clk), .RST(rst), .I(e[584]), 
        .Q(ein[584]) );
  DFF \ereg_reg[585]  ( .D(ereg_next[585]), .CLK(clk), .RST(rst), .I(e[585]), 
        .Q(ein[585]) );
  DFF \ereg_reg[586]  ( .D(ereg_next[586]), .CLK(clk), .RST(rst), .I(e[586]), 
        .Q(ein[586]) );
  DFF \ereg_reg[587]  ( .D(ereg_next[587]), .CLK(clk), .RST(rst), .I(e[587]), 
        .Q(ein[587]) );
  DFF \ereg_reg[588]  ( .D(ereg_next[588]), .CLK(clk), .RST(rst), .I(e[588]), 
        .Q(ein[588]) );
  DFF \ereg_reg[589]  ( .D(ereg_next[589]), .CLK(clk), .RST(rst), .I(e[589]), 
        .Q(ein[589]) );
  DFF \ereg_reg[590]  ( .D(ereg_next[590]), .CLK(clk), .RST(rst), .I(e[590]), 
        .Q(ein[590]) );
  DFF \ereg_reg[591]  ( .D(ereg_next[591]), .CLK(clk), .RST(rst), .I(e[591]), 
        .Q(ein[591]) );
  DFF \ereg_reg[592]  ( .D(ereg_next[592]), .CLK(clk), .RST(rst), .I(e[592]), 
        .Q(ein[592]) );
  DFF \ereg_reg[593]  ( .D(ereg_next[593]), .CLK(clk), .RST(rst), .I(e[593]), 
        .Q(ein[593]) );
  DFF \ereg_reg[594]  ( .D(ereg_next[594]), .CLK(clk), .RST(rst), .I(e[594]), 
        .Q(ein[594]) );
  DFF \ereg_reg[595]  ( .D(ereg_next[595]), .CLK(clk), .RST(rst), .I(e[595]), 
        .Q(ein[595]) );
  DFF \ereg_reg[596]  ( .D(ereg_next[596]), .CLK(clk), .RST(rst), .I(e[596]), 
        .Q(ein[596]) );
  DFF \ereg_reg[597]  ( .D(ereg_next[597]), .CLK(clk), .RST(rst), .I(e[597]), 
        .Q(ein[597]) );
  DFF \ereg_reg[598]  ( .D(ereg_next[598]), .CLK(clk), .RST(rst), .I(e[598]), 
        .Q(ein[598]) );
  DFF \ereg_reg[599]  ( .D(ereg_next[599]), .CLK(clk), .RST(rst), .I(e[599]), 
        .Q(ein[599]) );
  DFF \ereg_reg[600]  ( .D(ereg_next[600]), .CLK(clk), .RST(rst), .I(e[600]), 
        .Q(ein[600]) );
  DFF \ereg_reg[601]  ( .D(ereg_next[601]), .CLK(clk), .RST(rst), .I(e[601]), 
        .Q(ein[601]) );
  DFF \ereg_reg[602]  ( .D(ereg_next[602]), .CLK(clk), .RST(rst), .I(e[602]), 
        .Q(ein[602]) );
  DFF \ereg_reg[603]  ( .D(ereg_next[603]), .CLK(clk), .RST(rst), .I(e[603]), 
        .Q(ein[603]) );
  DFF \ereg_reg[604]  ( .D(ereg_next[604]), .CLK(clk), .RST(rst), .I(e[604]), 
        .Q(ein[604]) );
  DFF \ereg_reg[605]  ( .D(ereg_next[605]), .CLK(clk), .RST(rst), .I(e[605]), 
        .Q(ein[605]) );
  DFF \ereg_reg[606]  ( .D(ereg_next[606]), .CLK(clk), .RST(rst), .I(e[606]), 
        .Q(ein[606]) );
  DFF \ereg_reg[607]  ( .D(ereg_next[607]), .CLK(clk), .RST(rst), .I(e[607]), 
        .Q(ein[607]) );
  DFF \ereg_reg[608]  ( .D(ereg_next[608]), .CLK(clk), .RST(rst), .I(e[608]), 
        .Q(ein[608]) );
  DFF \ereg_reg[609]  ( .D(ereg_next[609]), .CLK(clk), .RST(rst), .I(e[609]), 
        .Q(ein[609]) );
  DFF \ereg_reg[610]  ( .D(ereg_next[610]), .CLK(clk), .RST(rst), .I(e[610]), 
        .Q(ein[610]) );
  DFF \ereg_reg[611]  ( .D(ereg_next[611]), .CLK(clk), .RST(rst), .I(e[611]), 
        .Q(ein[611]) );
  DFF \ereg_reg[612]  ( .D(ereg_next[612]), .CLK(clk), .RST(rst), .I(e[612]), 
        .Q(ein[612]) );
  DFF \ereg_reg[613]  ( .D(ereg_next[613]), .CLK(clk), .RST(rst), .I(e[613]), 
        .Q(ein[613]) );
  DFF \ereg_reg[614]  ( .D(ereg_next[614]), .CLK(clk), .RST(rst), .I(e[614]), 
        .Q(ein[614]) );
  DFF \ereg_reg[615]  ( .D(ereg_next[615]), .CLK(clk), .RST(rst), .I(e[615]), 
        .Q(ein[615]) );
  DFF \ereg_reg[616]  ( .D(ereg_next[616]), .CLK(clk), .RST(rst), .I(e[616]), 
        .Q(ein[616]) );
  DFF \ereg_reg[617]  ( .D(ereg_next[617]), .CLK(clk), .RST(rst), .I(e[617]), 
        .Q(ein[617]) );
  DFF \ereg_reg[618]  ( .D(ereg_next[618]), .CLK(clk), .RST(rst), .I(e[618]), 
        .Q(ein[618]) );
  DFF \ereg_reg[619]  ( .D(ereg_next[619]), .CLK(clk), .RST(rst), .I(e[619]), 
        .Q(ein[619]) );
  DFF \ereg_reg[620]  ( .D(ereg_next[620]), .CLK(clk), .RST(rst), .I(e[620]), 
        .Q(ein[620]) );
  DFF \ereg_reg[621]  ( .D(ereg_next[621]), .CLK(clk), .RST(rst), .I(e[621]), 
        .Q(ein[621]) );
  DFF \ereg_reg[622]  ( .D(ereg_next[622]), .CLK(clk), .RST(rst), .I(e[622]), 
        .Q(ein[622]) );
  DFF \ereg_reg[623]  ( .D(ereg_next[623]), .CLK(clk), .RST(rst), .I(e[623]), 
        .Q(ein[623]) );
  DFF \ereg_reg[624]  ( .D(ereg_next[624]), .CLK(clk), .RST(rst), .I(e[624]), 
        .Q(ein[624]) );
  DFF \ereg_reg[625]  ( .D(ereg_next[625]), .CLK(clk), .RST(rst), .I(e[625]), 
        .Q(ein[625]) );
  DFF \ereg_reg[626]  ( .D(ereg_next[626]), .CLK(clk), .RST(rst), .I(e[626]), 
        .Q(ein[626]) );
  DFF \ereg_reg[627]  ( .D(ereg_next[627]), .CLK(clk), .RST(rst), .I(e[627]), 
        .Q(ein[627]) );
  DFF \ereg_reg[628]  ( .D(ereg_next[628]), .CLK(clk), .RST(rst), .I(e[628]), 
        .Q(ein[628]) );
  DFF \ereg_reg[629]  ( .D(ereg_next[629]), .CLK(clk), .RST(rst), .I(e[629]), 
        .Q(ein[629]) );
  DFF \ereg_reg[630]  ( .D(ereg_next[630]), .CLK(clk), .RST(rst), .I(e[630]), 
        .Q(ein[630]) );
  DFF \ereg_reg[631]  ( .D(ereg_next[631]), .CLK(clk), .RST(rst), .I(e[631]), 
        .Q(ein[631]) );
  DFF \ereg_reg[632]  ( .D(ereg_next[632]), .CLK(clk), .RST(rst), .I(e[632]), 
        .Q(ein[632]) );
  DFF \ereg_reg[633]  ( .D(ereg_next[633]), .CLK(clk), .RST(rst), .I(e[633]), 
        .Q(ein[633]) );
  DFF \ereg_reg[634]  ( .D(ereg_next[634]), .CLK(clk), .RST(rst), .I(e[634]), 
        .Q(ein[634]) );
  DFF \ereg_reg[635]  ( .D(ereg_next[635]), .CLK(clk), .RST(rst), .I(e[635]), 
        .Q(ein[635]) );
  DFF \ereg_reg[636]  ( .D(ereg_next[636]), .CLK(clk), .RST(rst), .I(e[636]), 
        .Q(ein[636]) );
  DFF \ereg_reg[637]  ( .D(ereg_next[637]), .CLK(clk), .RST(rst), .I(e[637]), 
        .Q(ein[637]) );
  DFF \ereg_reg[638]  ( .D(ereg_next[638]), .CLK(clk), .RST(rst), .I(e[638]), 
        .Q(ein[638]) );
  DFF \ereg_reg[639]  ( .D(ereg_next[639]), .CLK(clk), .RST(rst), .I(e[639]), 
        .Q(ein[639]) );
  DFF \ereg_reg[640]  ( .D(ereg_next[640]), .CLK(clk), .RST(rst), .I(e[640]), 
        .Q(ein[640]) );
  DFF \ereg_reg[641]  ( .D(ereg_next[641]), .CLK(clk), .RST(rst), .I(e[641]), 
        .Q(ein[641]) );
  DFF \ereg_reg[642]  ( .D(ereg_next[642]), .CLK(clk), .RST(rst), .I(e[642]), 
        .Q(ein[642]) );
  DFF \ereg_reg[643]  ( .D(ereg_next[643]), .CLK(clk), .RST(rst), .I(e[643]), 
        .Q(ein[643]) );
  DFF \ereg_reg[644]  ( .D(ereg_next[644]), .CLK(clk), .RST(rst), .I(e[644]), 
        .Q(ein[644]) );
  DFF \ereg_reg[645]  ( .D(ereg_next[645]), .CLK(clk), .RST(rst), .I(e[645]), 
        .Q(ein[645]) );
  DFF \ereg_reg[646]  ( .D(ereg_next[646]), .CLK(clk), .RST(rst), .I(e[646]), 
        .Q(ein[646]) );
  DFF \ereg_reg[647]  ( .D(ereg_next[647]), .CLK(clk), .RST(rst), .I(e[647]), 
        .Q(ein[647]) );
  DFF \ereg_reg[648]  ( .D(ereg_next[648]), .CLK(clk), .RST(rst), .I(e[648]), 
        .Q(ein[648]) );
  DFF \ereg_reg[649]  ( .D(ereg_next[649]), .CLK(clk), .RST(rst), .I(e[649]), 
        .Q(ein[649]) );
  DFF \ereg_reg[650]  ( .D(ereg_next[650]), .CLK(clk), .RST(rst), .I(e[650]), 
        .Q(ein[650]) );
  DFF \ereg_reg[651]  ( .D(ereg_next[651]), .CLK(clk), .RST(rst), .I(e[651]), 
        .Q(ein[651]) );
  DFF \ereg_reg[652]  ( .D(ereg_next[652]), .CLK(clk), .RST(rst), .I(e[652]), 
        .Q(ein[652]) );
  DFF \ereg_reg[653]  ( .D(ereg_next[653]), .CLK(clk), .RST(rst), .I(e[653]), 
        .Q(ein[653]) );
  DFF \ereg_reg[654]  ( .D(ereg_next[654]), .CLK(clk), .RST(rst), .I(e[654]), 
        .Q(ein[654]) );
  DFF \ereg_reg[655]  ( .D(ereg_next[655]), .CLK(clk), .RST(rst), .I(e[655]), 
        .Q(ein[655]) );
  DFF \ereg_reg[656]  ( .D(ereg_next[656]), .CLK(clk), .RST(rst), .I(e[656]), 
        .Q(ein[656]) );
  DFF \ereg_reg[657]  ( .D(ereg_next[657]), .CLK(clk), .RST(rst), .I(e[657]), 
        .Q(ein[657]) );
  DFF \ereg_reg[658]  ( .D(ereg_next[658]), .CLK(clk), .RST(rst), .I(e[658]), 
        .Q(ein[658]) );
  DFF \ereg_reg[659]  ( .D(ereg_next[659]), .CLK(clk), .RST(rst), .I(e[659]), 
        .Q(ein[659]) );
  DFF \ereg_reg[660]  ( .D(ereg_next[660]), .CLK(clk), .RST(rst), .I(e[660]), 
        .Q(ein[660]) );
  DFF \ereg_reg[661]  ( .D(ereg_next[661]), .CLK(clk), .RST(rst), .I(e[661]), 
        .Q(ein[661]) );
  DFF \ereg_reg[662]  ( .D(ereg_next[662]), .CLK(clk), .RST(rst), .I(e[662]), 
        .Q(ein[662]) );
  DFF \ereg_reg[663]  ( .D(ereg_next[663]), .CLK(clk), .RST(rst), .I(e[663]), 
        .Q(ein[663]) );
  DFF \ereg_reg[664]  ( .D(ereg_next[664]), .CLK(clk), .RST(rst), .I(e[664]), 
        .Q(ein[664]) );
  DFF \ereg_reg[665]  ( .D(ereg_next[665]), .CLK(clk), .RST(rst), .I(e[665]), 
        .Q(ein[665]) );
  DFF \ereg_reg[666]  ( .D(ereg_next[666]), .CLK(clk), .RST(rst), .I(e[666]), 
        .Q(ein[666]) );
  DFF \ereg_reg[667]  ( .D(ereg_next[667]), .CLK(clk), .RST(rst), .I(e[667]), 
        .Q(ein[667]) );
  DFF \ereg_reg[668]  ( .D(ereg_next[668]), .CLK(clk), .RST(rst), .I(e[668]), 
        .Q(ein[668]) );
  DFF \ereg_reg[669]  ( .D(ereg_next[669]), .CLK(clk), .RST(rst), .I(e[669]), 
        .Q(ein[669]) );
  DFF \ereg_reg[670]  ( .D(ereg_next[670]), .CLK(clk), .RST(rst), .I(e[670]), 
        .Q(ein[670]) );
  DFF \ereg_reg[671]  ( .D(ereg_next[671]), .CLK(clk), .RST(rst), .I(e[671]), 
        .Q(ein[671]) );
  DFF \ereg_reg[672]  ( .D(ereg_next[672]), .CLK(clk), .RST(rst), .I(e[672]), 
        .Q(ein[672]) );
  DFF \ereg_reg[673]  ( .D(ereg_next[673]), .CLK(clk), .RST(rst), .I(e[673]), 
        .Q(ein[673]) );
  DFF \ereg_reg[674]  ( .D(ereg_next[674]), .CLK(clk), .RST(rst), .I(e[674]), 
        .Q(ein[674]) );
  DFF \ereg_reg[675]  ( .D(ereg_next[675]), .CLK(clk), .RST(rst), .I(e[675]), 
        .Q(ein[675]) );
  DFF \ereg_reg[676]  ( .D(ereg_next[676]), .CLK(clk), .RST(rst), .I(e[676]), 
        .Q(ein[676]) );
  DFF \ereg_reg[677]  ( .D(ereg_next[677]), .CLK(clk), .RST(rst), .I(e[677]), 
        .Q(ein[677]) );
  DFF \ereg_reg[678]  ( .D(ereg_next[678]), .CLK(clk), .RST(rst), .I(e[678]), 
        .Q(ein[678]) );
  DFF \ereg_reg[679]  ( .D(ereg_next[679]), .CLK(clk), .RST(rst), .I(e[679]), 
        .Q(ein[679]) );
  DFF \ereg_reg[680]  ( .D(ereg_next[680]), .CLK(clk), .RST(rst), .I(e[680]), 
        .Q(ein[680]) );
  DFF \ereg_reg[681]  ( .D(ereg_next[681]), .CLK(clk), .RST(rst), .I(e[681]), 
        .Q(ein[681]) );
  DFF \ereg_reg[682]  ( .D(ereg_next[682]), .CLK(clk), .RST(rst), .I(e[682]), 
        .Q(ein[682]) );
  DFF \ereg_reg[683]  ( .D(ereg_next[683]), .CLK(clk), .RST(rst), .I(e[683]), 
        .Q(ein[683]) );
  DFF \ereg_reg[684]  ( .D(ereg_next[684]), .CLK(clk), .RST(rst), .I(e[684]), 
        .Q(ein[684]) );
  DFF \ereg_reg[685]  ( .D(ereg_next[685]), .CLK(clk), .RST(rst), .I(e[685]), 
        .Q(ein[685]) );
  DFF \ereg_reg[686]  ( .D(ereg_next[686]), .CLK(clk), .RST(rst), .I(e[686]), 
        .Q(ein[686]) );
  DFF \ereg_reg[687]  ( .D(ereg_next[687]), .CLK(clk), .RST(rst), .I(e[687]), 
        .Q(ein[687]) );
  DFF \ereg_reg[688]  ( .D(ereg_next[688]), .CLK(clk), .RST(rst), .I(e[688]), 
        .Q(ein[688]) );
  DFF \ereg_reg[689]  ( .D(ereg_next[689]), .CLK(clk), .RST(rst), .I(e[689]), 
        .Q(ein[689]) );
  DFF \ereg_reg[690]  ( .D(ereg_next[690]), .CLK(clk), .RST(rst), .I(e[690]), 
        .Q(ein[690]) );
  DFF \ereg_reg[691]  ( .D(ereg_next[691]), .CLK(clk), .RST(rst), .I(e[691]), 
        .Q(ein[691]) );
  DFF \ereg_reg[692]  ( .D(ereg_next[692]), .CLK(clk), .RST(rst), .I(e[692]), 
        .Q(ein[692]) );
  DFF \ereg_reg[693]  ( .D(ereg_next[693]), .CLK(clk), .RST(rst), .I(e[693]), 
        .Q(ein[693]) );
  DFF \ereg_reg[694]  ( .D(ereg_next[694]), .CLK(clk), .RST(rst), .I(e[694]), 
        .Q(ein[694]) );
  DFF \ereg_reg[695]  ( .D(ereg_next[695]), .CLK(clk), .RST(rst), .I(e[695]), 
        .Q(ein[695]) );
  DFF \ereg_reg[696]  ( .D(ereg_next[696]), .CLK(clk), .RST(rst), .I(e[696]), 
        .Q(ein[696]) );
  DFF \ereg_reg[697]  ( .D(ereg_next[697]), .CLK(clk), .RST(rst), .I(e[697]), 
        .Q(ein[697]) );
  DFF \ereg_reg[698]  ( .D(ereg_next[698]), .CLK(clk), .RST(rst), .I(e[698]), 
        .Q(ein[698]) );
  DFF \ereg_reg[699]  ( .D(ereg_next[699]), .CLK(clk), .RST(rst), .I(e[699]), 
        .Q(ein[699]) );
  DFF \ereg_reg[700]  ( .D(ereg_next[700]), .CLK(clk), .RST(rst), .I(e[700]), 
        .Q(ein[700]) );
  DFF \ereg_reg[701]  ( .D(ereg_next[701]), .CLK(clk), .RST(rst), .I(e[701]), 
        .Q(ein[701]) );
  DFF \ereg_reg[702]  ( .D(ereg_next[702]), .CLK(clk), .RST(rst), .I(e[702]), 
        .Q(ein[702]) );
  DFF \ereg_reg[703]  ( .D(ereg_next[703]), .CLK(clk), .RST(rst), .I(e[703]), 
        .Q(ein[703]) );
  DFF \ereg_reg[704]  ( .D(ereg_next[704]), .CLK(clk), .RST(rst), .I(e[704]), 
        .Q(ein[704]) );
  DFF \ereg_reg[705]  ( .D(ereg_next[705]), .CLK(clk), .RST(rst), .I(e[705]), 
        .Q(ein[705]) );
  DFF \ereg_reg[706]  ( .D(ereg_next[706]), .CLK(clk), .RST(rst), .I(e[706]), 
        .Q(ein[706]) );
  DFF \ereg_reg[707]  ( .D(ereg_next[707]), .CLK(clk), .RST(rst), .I(e[707]), 
        .Q(ein[707]) );
  DFF \ereg_reg[708]  ( .D(ereg_next[708]), .CLK(clk), .RST(rst), .I(e[708]), 
        .Q(ein[708]) );
  DFF \ereg_reg[709]  ( .D(ereg_next[709]), .CLK(clk), .RST(rst), .I(e[709]), 
        .Q(ein[709]) );
  DFF \ereg_reg[710]  ( .D(ereg_next[710]), .CLK(clk), .RST(rst), .I(e[710]), 
        .Q(ein[710]) );
  DFF \ereg_reg[711]  ( .D(ereg_next[711]), .CLK(clk), .RST(rst), .I(e[711]), 
        .Q(ein[711]) );
  DFF \ereg_reg[712]  ( .D(ereg_next[712]), .CLK(clk), .RST(rst), .I(e[712]), 
        .Q(ein[712]) );
  DFF \ereg_reg[713]  ( .D(ereg_next[713]), .CLK(clk), .RST(rst), .I(e[713]), 
        .Q(ein[713]) );
  DFF \ereg_reg[714]  ( .D(ereg_next[714]), .CLK(clk), .RST(rst), .I(e[714]), 
        .Q(ein[714]) );
  DFF \ereg_reg[715]  ( .D(ereg_next[715]), .CLK(clk), .RST(rst), .I(e[715]), 
        .Q(ein[715]) );
  DFF \ereg_reg[716]  ( .D(ereg_next[716]), .CLK(clk), .RST(rst), .I(e[716]), 
        .Q(ein[716]) );
  DFF \ereg_reg[717]  ( .D(ereg_next[717]), .CLK(clk), .RST(rst), .I(e[717]), 
        .Q(ein[717]) );
  DFF \ereg_reg[718]  ( .D(ereg_next[718]), .CLK(clk), .RST(rst), .I(e[718]), 
        .Q(ein[718]) );
  DFF \ereg_reg[719]  ( .D(ereg_next[719]), .CLK(clk), .RST(rst), .I(e[719]), 
        .Q(ein[719]) );
  DFF \ereg_reg[720]  ( .D(ereg_next[720]), .CLK(clk), .RST(rst), .I(e[720]), 
        .Q(ein[720]) );
  DFF \ereg_reg[721]  ( .D(ereg_next[721]), .CLK(clk), .RST(rst), .I(e[721]), 
        .Q(ein[721]) );
  DFF \ereg_reg[722]  ( .D(ereg_next[722]), .CLK(clk), .RST(rst), .I(e[722]), 
        .Q(ein[722]) );
  DFF \ereg_reg[723]  ( .D(ereg_next[723]), .CLK(clk), .RST(rst), .I(e[723]), 
        .Q(ein[723]) );
  DFF \ereg_reg[724]  ( .D(ereg_next[724]), .CLK(clk), .RST(rst), .I(e[724]), 
        .Q(ein[724]) );
  DFF \ereg_reg[725]  ( .D(ereg_next[725]), .CLK(clk), .RST(rst), .I(e[725]), 
        .Q(ein[725]) );
  DFF \ereg_reg[726]  ( .D(ereg_next[726]), .CLK(clk), .RST(rst), .I(e[726]), 
        .Q(ein[726]) );
  DFF \ereg_reg[727]  ( .D(ereg_next[727]), .CLK(clk), .RST(rst), .I(e[727]), 
        .Q(ein[727]) );
  DFF \ereg_reg[728]  ( .D(ereg_next[728]), .CLK(clk), .RST(rst), .I(e[728]), 
        .Q(ein[728]) );
  DFF \ereg_reg[729]  ( .D(ereg_next[729]), .CLK(clk), .RST(rst), .I(e[729]), 
        .Q(ein[729]) );
  DFF \ereg_reg[730]  ( .D(ereg_next[730]), .CLK(clk), .RST(rst), .I(e[730]), 
        .Q(ein[730]) );
  DFF \ereg_reg[731]  ( .D(ereg_next[731]), .CLK(clk), .RST(rst), .I(e[731]), 
        .Q(ein[731]) );
  DFF \ereg_reg[732]  ( .D(ereg_next[732]), .CLK(clk), .RST(rst), .I(e[732]), 
        .Q(ein[732]) );
  DFF \ereg_reg[733]  ( .D(ereg_next[733]), .CLK(clk), .RST(rst), .I(e[733]), 
        .Q(ein[733]) );
  DFF \ereg_reg[734]  ( .D(ereg_next[734]), .CLK(clk), .RST(rst), .I(e[734]), 
        .Q(ein[734]) );
  DFF \ereg_reg[735]  ( .D(ereg_next[735]), .CLK(clk), .RST(rst), .I(e[735]), 
        .Q(ein[735]) );
  DFF \ereg_reg[736]  ( .D(ereg_next[736]), .CLK(clk), .RST(rst), .I(e[736]), 
        .Q(ein[736]) );
  DFF \ereg_reg[737]  ( .D(ereg_next[737]), .CLK(clk), .RST(rst), .I(e[737]), 
        .Q(ein[737]) );
  DFF \ereg_reg[738]  ( .D(ereg_next[738]), .CLK(clk), .RST(rst), .I(e[738]), 
        .Q(ein[738]) );
  DFF \ereg_reg[739]  ( .D(ereg_next[739]), .CLK(clk), .RST(rst), .I(e[739]), 
        .Q(ein[739]) );
  DFF \ereg_reg[740]  ( .D(ereg_next[740]), .CLK(clk), .RST(rst), .I(e[740]), 
        .Q(ein[740]) );
  DFF \ereg_reg[741]  ( .D(ereg_next[741]), .CLK(clk), .RST(rst), .I(e[741]), 
        .Q(ein[741]) );
  DFF \ereg_reg[742]  ( .D(ereg_next[742]), .CLK(clk), .RST(rst), .I(e[742]), 
        .Q(ein[742]) );
  DFF \ereg_reg[743]  ( .D(ereg_next[743]), .CLK(clk), .RST(rst), .I(e[743]), 
        .Q(ein[743]) );
  DFF \ereg_reg[744]  ( .D(ereg_next[744]), .CLK(clk), .RST(rst), .I(e[744]), 
        .Q(ein[744]) );
  DFF \ereg_reg[745]  ( .D(ereg_next[745]), .CLK(clk), .RST(rst), .I(e[745]), 
        .Q(ein[745]) );
  DFF \ereg_reg[746]  ( .D(ereg_next[746]), .CLK(clk), .RST(rst), .I(e[746]), 
        .Q(ein[746]) );
  DFF \ereg_reg[747]  ( .D(ereg_next[747]), .CLK(clk), .RST(rst), .I(e[747]), 
        .Q(ein[747]) );
  DFF \ereg_reg[748]  ( .D(ereg_next[748]), .CLK(clk), .RST(rst), .I(e[748]), 
        .Q(ein[748]) );
  DFF \ereg_reg[749]  ( .D(ereg_next[749]), .CLK(clk), .RST(rst), .I(e[749]), 
        .Q(ein[749]) );
  DFF \ereg_reg[750]  ( .D(ereg_next[750]), .CLK(clk), .RST(rst), .I(e[750]), 
        .Q(ein[750]) );
  DFF \ereg_reg[751]  ( .D(ereg_next[751]), .CLK(clk), .RST(rst), .I(e[751]), 
        .Q(ein[751]) );
  DFF \ereg_reg[752]  ( .D(ereg_next[752]), .CLK(clk), .RST(rst), .I(e[752]), 
        .Q(ein[752]) );
  DFF \ereg_reg[753]  ( .D(ereg_next[753]), .CLK(clk), .RST(rst), .I(e[753]), 
        .Q(ein[753]) );
  DFF \ereg_reg[754]  ( .D(ereg_next[754]), .CLK(clk), .RST(rst), .I(e[754]), 
        .Q(ein[754]) );
  DFF \ereg_reg[755]  ( .D(ereg_next[755]), .CLK(clk), .RST(rst), .I(e[755]), 
        .Q(ein[755]) );
  DFF \ereg_reg[756]  ( .D(ereg_next[756]), .CLK(clk), .RST(rst), .I(e[756]), 
        .Q(ein[756]) );
  DFF \ereg_reg[757]  ( .D(ereg_next[757]), .CLK(clk), .RST(rst), .I(e[757]), 
        .Q(ein[757]) );
  DFF \ereg_reg[758]  ( .D(ereg_next[758]), .CLK(clk), .RST(rst), .I(e[758]), 
        .Q(ein[758]) );
  DFF \ereg_reg[759]  ( .D(ereg_next[759]), .CLK(clk), .RST(rst), .I(e[759]), 
        .Q(ein[759]) );
  DFF \ereg_reg[760]  ( .D(ereg_next[760]), .CLK(clk), .RST(rst), .I(e[760]), 
        .Q(ein[760]) );
  DFF \ereg_reg[761]  ( .D(ereg_next[761]), .CLK(clk), .RST(rst), .I(e[761]), 
        .Q(ein[761]) );
  DFF \ereg_reg[762]  ( .D(ereg_next[762]), .CLK(clk), .RST(rst), .I(e[762]), 
        .Q(ein[762]) );
  DFF \ereg_reg[763]  ( .D(ereg_next[763]), .CLK(clk), .RST(rst), .I(e[763]), 
        .Q(ein[763]) );
  DFF \ereg_reg[764]  ( .D(ereg_next[764]), .CLK(clk), .RST(rst), .I(e[764]), 
        .Q(ein[764]) );
  DFF \ereg_reg[765]  ( .D(ereg_next[765]), .CLK(clk), .RST(rst), .I(e[765]), 
        .Q(ein[765]) );
  DFF \ereg_reg[766]  ( .D(ereg_next[766]), .CLK(clk), .RST(rst), .I(e[766]), 
        .Q(ein[766]) );
  DFF \ereg_reg[767]  ( .D(ereg_next[767]), .CLK(clk), .RST(rst), .I(e[767]), 
        .Q(ein[767]) );
  DFF \ereg_reg[768]  ( .D(ereg_next[768]), .CLK(clk), .RST(rst), .I(e[768]), 
        .Q(ein[768]) );
  DFF \ereg_reg[769]  ( .D(ereg_next[769]), .CLK(clk), .RST(rst), .I(e[769]), 
        .Q(ein[769]) );
  DFF \ereg_reg[770]  ( .D(ereg_next[770]), .CLK(clk), .RST(rst), .I(e[770]), 
        .Q(ein[770]) );
  DFF \ereg_reg[771]  ( .D(ereg_next[771]), .CLK(clk), .RST(rst), .I(e[771]), 
        .Q(ein[771]) );
  DFF \ereg_reg[772]  ( .D(ereg_next[772]), .CLK(clk), .RST(rst), .I(e[772]), 
        .Q(ein[772]) );
  DFF \ereg_reg[773]  ( .D(ereg_next[773]), .CLK(clk), .RST(rst), .I(e[773]), 
        .Q(ein[773]) );
  DFF \ereg_reg[774]  ( .D(ereg_next[774]), .CLK(clk), .RST(rst), .I(e[774]), 
        .Q(ein[774]) );
  DFF \ereg_reg[775]  ( .D(ereg_next[775]), .CLK(clk), .RST(rst), .I(e[775]), 
        .Q(ein[775]) );
  DFF \ereg_reg[776]  ( .D(ereg_next[776]), .CLK(clk), .RST(rst), .I(e[776]), 
        .Q(ein[776]) );
  DFF \ereg_reg[777]  ( .D(ereg_next[777]), .CLK(clk), .RST(rst), .I(e[777]), 
        .Q(ein[777]) );
  DFF \ereg_reg[778]  ( .D(ereg_next[778]), .CLK(clk), .RST(rst), .I(e[778]), 
        .Q(ein[778]) );
  DFF \ereg_reg[779]  ( .D(ereg_next[779]), .CLK(clk), .RST(rst), .I(e[779]), 
        .Q(ein[779]) );
  DFF \ereg_reg[780]  ( .D(ereg_next[780]), .CLK(clk), .RST(rst), .I(e[780]), 
        .Q(ein[780]) );
  DFF \ereg_reg[781]  ( .D(ereg_next[781]), .CLK(clk), .RST(rst), .I(e[781]), 
        .Q(ein[781]) );
  DFF \ereg_reg[782]  ( .D(ereg_next[782]), .CLK(clk), .RST(rst), .I(e[782]), 
        .Q(ein[782]) );
  DFF \ereg_reg[783]  ( .D(ereg_next[783]), .CLK(clk), .RST(rst), .I(e[783]), 
        .Q(ein[783]) );
  DFF \ereg_reg[784]  ( .D(ereg_next[784]), .CLK(clk), .RST(rst), .I(e[784]), 
        .Q(ein[784]) );
  DFF \ereg_reg[785]  ( .D(ereg_next[785]), .CLK(clk), .RST(rst), .I(e[785]), 
        .Q(ein[785]) );
  DFF \ereg_reg[786]  ( .D(ereg_next[786]), .CLK(clk), .RST(rst), .I(e[786]), 
        .Q(ein[786]) );
  DFF \ereg_reg[787]  ( .D(ereg_next[787]), .CLK(clk), .RST(rst), .I(e[787]), 
        .Q(ein[787]) );
  DFF \ereg_reg[788]  ( .D(ereg_next[788]), .CLK(clk), .RST(rst), .I(e[788]), 
        .Q(ein[788]) );
  DFF \ereg_reg[789]  ( .D(ereg_next[789]), .CLK(clk), .RST(rst), .I(e[789]), 
        .Q(ein[789]) );
  DFF \ereg_reg[790]  ( .D(ereg_next[790]), .CLK(clk), .RST(rst), .I(e[790]), 
        .Q(ein[790]) );
  DFF \ereg_reg[791]  ( .D(ereg_next[791]), .CLK(clk), .RST(rst), .I(e[791]), 
        .Q(ein[791]) );
  DFF \ereg_reg[792]  ( .D(ereg_next[792]), .CLK(clk), .RST(rst), .I(e[792]), 
        .Q(ein[792]) );
  DFF \ereg_reg[793]  ( .D(ereg_next[793]), .CLK(clk), .RST(rst), .I(e[793]), 
        .Q(ein[793]) );
  DFF \ereg_reg[794]  ( .D(ereg_next[794]), .CLK(clk), .RST(rst), .I(e[794]), 
        .Q(ein[794]) );
  DFF \ereg_reg[795]  ( .D(ereg_next[795]), .CLK(clk), .RST(rst), .I(e[795]), 
        .Q(ein[795]) );
  DFF \ereg_reg[796]  ( .D(ereg_next[796]), .CLK(clk), .RST(rst), .I(e[796]), 
        .Q(ein[796]) );
  DFF \ereg_reg[797]  ( .D(ereg_next[797]), .CLK(clk), .RST(rst), .I(e[797]), 
        .Q(ein[797]) );
  DFF \ereg_reg[798]  ( .D(ereg_next[798]), .CLK(clk), .RST(rst), .I(e[798]), 
        .Q(ein[798]) );
  DFF \ereg_reg[799]  ( .D(ereg_next[799]), .CLK(clk), .RST(rst), .I(e[799]), 
        .Q(ein[799]) );
  DFF \ereg_reg[800]  ( .D(ereg_next[800]), .CLK(clk), .RST(rst), .I(e[800]), 
        .Q(ein[800]) );
  DFF \ereg_reg[801]  ( .D(ereg_next[801]), .CLK(clk), .RST(rst), .I(e[801]), 
        .Q(ein[801]) );
  DFF \ereg_reg[802]  ( .D(ereg_next[802]), .CLK(clk), .RST(rst), .I(e[802]), 
        .Q(ein[802]) );
  DFF \ereg_reg[803]  ( .D(ereg_next[803]), .CLK(clk), .RST(rst), .I(e[803]), 
        .Q(ein[803]) );
  DFF \ereg_reg[804]  ( .D(ereg_next[804]), .CLK(clk), .RST(rst), .I(e[804]), 
        .Q(ein[804]) );
  DFF \ereg_reg[805]  ( .D(ereg_next[805]), .CLK(clk), .RST(rst), .I(e[805]), 
        .Q(ein[805]) );
  DFF \ereg_reg[806]  ( .D(ereg_next[806]), .CLK(clk), .RST(rst), .I(e[806]), 
        .Q(ein[806]) );
  DFF \ereg_reg[807]  ( .D(ereg_next[807]), .CLK(clk), .RST(rst), .I(e[807]), 
        .Q(ein[807]) );
  DFF \ereg_reg[808]  ( .D(ereg_next[808]), .CLK(clk), .RST(rst), .I(e[808]), 
        .Q(ein[808]) );
  DFF \ereg_reg[809]  ( .D(ereg_next[809]), .CLK(clk), .RST(rst), .I(e[809]), 
        .Q(ein[809]) );
  DFF \ereg_reg[810]  ( .D(ereg_next[810]), .CLK(clk), .RST(rst), .I(e[810]), 
        .Q(ein[810]) );
  DFF \ereg_reg[811]  ( .D(ereg_next[811]), .CLK(clk), .RST(rst), .I(e[811]), 
        .Q(ein[811]) );
  DFF \ereg_reg[812]  ( .D(ereg_next[812]), .CLK(clk), .RST(rst), .I(e[812]), 
        .Q(ein[812]) );
  DFF \ereg_reg[813]  ( .D(ereg_next[813]), .CLK(clk), .RST(rst), .I(e[813]), 
        .Q(ein[813]) );
  DFF \ereg_reg[814]  ( .D(ereg_next[814]), .CLK(clk), .RST(rst), .I(e[814]), 
        .Q(ein[814]) );
  DFF \ereg_reg[815]  ( .D(ereg_next[815]), .CLK(clk), .RST(rst), .I(e[815]), 
        .Q(ein[815]) );
  DFF \ereg_reg[816]  ( .D(ereg_next[816]), .CLK(clk), .RST(rst), .I(e[816]), 
        .Q(ein[816]) );
  DFF \ereg_reg[817]  ( .D(ereg_next[817]), .CLK(clk), .RST(rst), .I(e[817]), 
        .Q(ein[817]) );
  DFF \ereg_reg[818]  ( .D(ereg_next[818]), .CLK(clk), .RST(rst), .I(e[818]), 
        .Q(ein[818]) );
  DFF \ereg_reg[819]  ( .D(ereg_next[819]), .CLK(clk), .RST(rst), .I(e[819]), 
        .Q(ein[819]) );
  DFF \ereg_reg[820]  ( .D(ereg_next[820]), .CLK(clk), .RST(rst), .I(e[820]), 
        .Q(ein[820]) );
  DFF \ereg_reg[821]  ( .D(ereg_next[821]), .CLK(clk), .RST(rst), .I(e[821]), 
        .Q(ein[821]) );
  DFF \ereg_reg[822]  ( .D(ereg_next[822]), .CLK(clk), .RST(rst), .I(e[822]), 
        .Q(ein[822]) );
  DFF \ereg_reg[823]  ( .D(ereg_next[823]), .CLK(clk), .RST(rst), .I(e[823]), 
        .Q(ein[823]) );
  DFF \ereg_reg[824]  ( .D(ereg_next[824]), .CLK(clk), .RST(rst), .I(e[824]), 
        .Q(ein[824]) );
  DFF \ereg_reg[825]  ( .D(ereg_next[825]), .CLK(clk), .RST(rst), .I(e[825]), 
        .Q(ein[825]) );
  DFF \ereg_reg[826]  ( .D(ereg_next[826]), .CLK(clk), .RST(rst), .I(e[826]), 
        .Q(ein[826]) );
  DFF \ereg_reg[827]  ( .D(ereg_next[827]), .CLK(clk), .RST(rst), .I(e[827]), 
        .Q(ein[827]) );
  DFF \ereg_reg[828]  ( .D(ereg_next[828]), .CLK(clk), .RST(rst), .I(e[828]), 
        .Q(ein[828]) );
  DFF \ereg_reg[829]  ( .D(ereg_next[829]), .CLK(clk), .RST(rst), .I(e[829]), 
        .Q(ein[829]) );
  DFF \ereg_reg[830]  ( .D(ereg_next[830]), .CLK(clk), .RST(rst), .I(e[830]), 
        .Q(ein[830]) );
  DFF \ereg_reg[831]  ( .D(ereg_next[831]), .CLK(clk), .RST(rst), .I(e[831]), 
        .Q(ein[831]) );
  DFF \ereg_reg[832]  ( .D(ereg_next[832]), .CLK(clk), .RST(rst), .I(e[832]), 
        .Q(ein[832]) );
  DFF \ereg_reg[833]  ( .D(ereg_next[833]), .CLK(clk), .RST(rst), .I(e[833]), 
        .Q(ein[833]) );
  DFF \ereg_reg[834]  ( .D(ereg_next[834]), .CLK(clk), .RST(rst), .I(e[834]), 
        .Q(ein[834]) );
  DFF \ereg_reg[835]  ( .D(ereg_next[835]), .CLK(clk), .RST(rst), .I(e[835]), 
        .Q(ein[835]) );
  DFF \ereg_reg[836]  ( .D(ereg_next[836]), .CLK(clk), .RST(rst), .I(e[836]), 
        .Q(ein[836]) );
  DFF \ereg_reg[837]  ( .D(ereg_next[837]), .CLK(clk), .RST(rst), .I(e[837]), 
        .Q(ein[837]) );
  DFF \ereg_reg[838]  ( .D(ereg_next[838]), .CLK(clk), .RST(rst), .I(e[838]), 
        .Q(ein[838]) );
  DFF \ereg_reg[839]  ( .D(ereg_next[839]), .CLK(clk), .RST(rst), .I(e[839]), 
        .Q(ein[839]) );
  DFF \ereg_reg[840]  ( .D(ereg_next[840]), .CLK(clk), .RST(rst), .I(e[840]), 
        .Q(ein[840]) );
  DFF \ereg_reg[841]  ( .D(ereg_next[841]), .CLK(clk), .RST(rst), .I(e[841]), 
        .Q(ein[841]) );
  DFF \ereg_reg[842]  ( .D(ereg_next[842]), .CLK(clk), .RST(rst), .I(e[842]), 
        .Q(ein[842]) );
  DFF \ereg_reg[843]  ( .D(ereg_next[843]), .CLK(clk), .RST(rst), .I(e[843]), 
        .Q(ein[843]) );
  DFF \ereg_reg[844]  ( .D(ereg_next[844]), .CLK(clk), .RST(rst), .I(e[844]), 
        .Q(ein[844]) );
  DFF \ereg_reg[845]  ( .D(ereg_next[845]), .CLK(clk), .RST(rst), .I(e[845]), 
        .Q(ein[845]) );
  DFF \ereg_reg[846]  ( .D(ereg_next[846]), .CLK(clk), .RST(rst), .I(e[846]), 
        .Q(ein[846]) );
  DFF \ereg_reg[847]  ( .D(ereg_next[847]), .CLK(clk), .RST(rst), .I(e[847]), 
        .Q(ein[847]) );
  DFF \ereg_reg[848]  ( .D(ereg_next[848]), .CLK(clk), .RST(rst), .I(e[848]), 
        .Q(ein[848]) );
  DFF \ereg_reg[849]  ( .D(ereg_next[849]), .CLK(clk), .RST(rst), .I(e[849]), 
        .Q(ein[849]) );
  DFF \ereg_reg[850]  ( .D(ereg_next[850]), .CLK(clk), .RST(rst), .I(e[850]), 
        .Q(ein[850]) );
  DFF \ereg_reg[851]  ( .D(ereg_next[851]), .CLK(clk), .RST(rst), .I(e[851]), 
        .Q(ein[851]) );
  DFF \ereg_reg[852]  ( .D(ereg_next[852]), .CLK(clk), .RST(rst), .I(e[852]), 
        .Q(ein[852]) );
  DFF \ereg_reg[853]  ( .D(ereg_next[853]), .CLK(clk), .RST(rst), .I(e[853]), 
        .Q(ein[853]) );
  DFF \ereg_reg[854]  ( .D(ereg_next[854]), .CLK(clk), .RST(rst), .I(e[854]), 
        .Q(ein[854]) );
  DFF \ereg_reg[855]  ( .D(ereg_next[855]), .CLK(clk), .RST(rst), .I(e[855]), 
        .Q(ein[855]) );
  DFF \ereg_reg[856]  ( .D(ereg_next[856]), .CLK(clk), .RST(rst), .I(e[856]), 
        .Q(ein[856]) );
  DFF \ereg_reg[857]  ( .D(ereg_next[857]), .CLK(clk), .RST(rst), .I(e[857]), 
        .Q(ein[857]) );
  DFF \ereg_reg[858]  ( .D(ereg_next[858]), .CLK(clk), .RST(rst), .I(e[858]), 
        .Q(ein[858]) );
  DFF \ereg_reg[859]  ( .D(ereg_next[859]), .CLK(clk), .RST(rst), .I(e[859]), 
        .Q(ein[859]) );
  DFF \ereg_reg[860]  ( .D(ereg_next[860]), .CLK(clk), .RST(rst), .I(e[860]), 
        .Q(ein[860]) );
  DFF \ereg_reg[861]  ( .D(ereg_next[861]), .CLK(clk), .RST(rst), .I(e[861]), 
        .Q(ein[861]) );
  DFF \ereg_reg[862]  ( .D(ereg_next[862]), .CLK(clk), .RST(rst), .I(e[862]), 
        .Q(ein[862]) );
  DFF \ereg_reg[863]  ( .D(ereg_next[863]), .CLK(clk), .RST(rst), .I(e[863]), 
        .Q(ein[863]) );
  DFF \ereg_reg[864]  ( .D(ereg_next[864]), .CLK(clk), .RST(rst), .I(e[864]), 
        .Q(ein[864]) );
  DFF \ereg_reg[865]  ( .D(ereg_next[865]), .CLK(clk), .RST(rst), .I(e[865]), 
        .Q(ein[865]) );
  DFF \ereg_reg[866]  ( .D(ereg_next[866]), .CLK(clk), .RST(rst), .I(e[866]), 
        .Q(ein[866]) );
  DFF \ereg_reg[867]  ( .D(ereg_next[867]), .CLK(clk), .RST(rst), .I(e[867]), 
        .Q(ein[867]) );
  DFF \ereg_reg[868]  ( .D(ereg_next[868]), .CLK(clk), .RST(rst), .I(e[868]), 
        .Q(ein[868]) );
  DFF \ereg_reg[869]  ( .D(ereg_next[869]), .CLK(clk), .RST(rst), .I(e[869]), 
        .Q(ein[869]) );
  DFF \ereg_reg[870]  ( .D(ereg_next[870]), .CLK(clk), .RST(rst), .I(e[870]), 
        .Q(ein[870]) );
  DFF \ereg_reg[871]  ( .D(ereg_next[871]), .CLK(clk), .RST(rst), .I(e[871]), 
        .Q(ein[871]) );
  DFF \ereg_reg[872]  ( .D(ereg_next[872]), .CLK(clk), .RST(rst), .I(e[872]), 
        .Q(ein[872]) );
  DFF \ereg_reg[873]  ( .D(ereg_next[873]), .CLK(clk), .RST(rst), .I(e[873]), 
        .Q(ein[873]) );
  DFF \ereg_reg[874]  ( .D(ereg_next[874]), .CLK(clk), .RST(rst), .I(e[874]), 
        .Q(ein[874]) );
  DFF \ereg_reg[875]  ( .D(ereg_next[875]), .CLK(clk), .RST(rst), .I(e[875]), 
        .Q(ein[875]) );
  DFF \ereg_reg[876]  ( .D(ereg_next[876]), .CLK(clk), .RST(rst), .I(e[876]), 
        .Q(ein[876]) );
  DFF \ereg_reg[877]  ( .D(ereg_next[877]), .CLK(clk), .RST(rst), .I(e[877]), 
        .Q(ein[877]) );
  DFF \ereg_reg[878]  ( .D(ereg_next[878]), .CLK(clk), .RST(rst), .I(e[878]), 
        .Q(ein[878]) );
  DFF \ereg_reg[879]  ( .D(ereg_next[879]), .CLK(clk), .RST(rst), .I(e[879]), 
        .Q(ein[879]) );
  DFF \ereg_reg[880]  ( .D(ereg_next[880]), .CLK(clk), .RST(rst), .I(e[880]), 
        .Q(ein[880]) );
  DFF \ereg_reg[881]  ( .D(ereg_next[881]), .CLK(clk), .RST(rst), .I(e[881]), 
        .Q(ein[881]) );
  DFF \ereg_reg[882]  ( .D(ereg_next[882]), .CLK(clk), .RST(rst), .I(e[882]), 
        .Q(ein[882]) );
  DFF \ereg_reg[883]  ( .D(ereg_next[883]), .CLK(clk), .RST(rst), .I(e[883]), 
        .Q(ein[883]) );
  DFF \ereg_reg[884]  ( .D(ereg_next[884]), .CLK(clk), .RST(rst), .I(e[884]), 
        .Q(ein[884]) );
  DFF \ereg_reg[885]  ( .D(ereg_next[885]), .CLK(clk), .RST(rst), .I(e[885]), 
        .Q(ein[885]) );
  DFF \ereg_reg[886]  ( .D(ereg_next[886]), .CLK(clk), .RST(rst), .I(e[886]), 
        .Q(ein[886]) );
  DFF \ereg_reg[887]  ( .D(ereg_next[887]), .CLK(clk), .RST(rst), .I(e[887]), 
        .Q(ein[887]) );
  DFF \ereg_reg[888]  ( .D(ereg_next[888]), .CLK(clk), .RST(rst), .I(e[888]), 
        .Q(ein[888]) );
  DFF \ereg_reg[889]  ( .D(ereg_next[889]), .CLK(clk), .RST(rst), .I(e[889]), 
        .Q(ein[889]) );
  DFF \ereg_reg[890]  ( .D(ereg_next[890]), .CLK(clk), .RST(rst), .I(e[890]), 
        .Q(ein[890]) );
  DFF \ereg_reg[891]  ( .D(ereg_next[891]), .CLK(clk), .RST(rst), .I(e[891]), 
        .Q(ein[891]) );
  DFF \ereg_reg[892]  ( .D(ereg_next[892]), .CLK(clk), .RST(rst), .I(e[892]), 
        .Q(ein[892]) );
  DFF \ereg_reg[893]  ( .D(ereg_next[893]), .CLK(clk), .RST(rst), .I(e[893]), 
        .Q(ein[893]) );
  DFF \ereg_reg[894]  ( .D(ereg_next[894]), .CLK(clk), .RST(rst), .I(e[894]), 
        .Q(ein[894]) );
  DFF \ereg_reg[895]  ( .D(ereg_next[895]), .CLK(clk), .RST(rst), .I(e[895]), 
        .Q(ein[895]) );
  DFF \ereg_reg[896]  ( .D(ereg_next[896]), .CLK(clk), .RST(rst), .I(e[896]), 
        .Q(ein[896]) );
  DFF \ereg_reg[897]  ( .D(ereg_next[897]), .CLK(clk), .RST(rst), .I(e[897]), 
        .Q(ein[897]) );
  DFF \ereg_reg[898]  ( .D(ereg_next[898]), .CLK(clk), .RST(rst), .I(e[898]), 
        .Q(ein[898]) );
  DFF \ereg_reg[899]  ( .D(ereg_next[899]), .CLK(clk), .RST(rst), .I(e[899]), 
        .Q(ein[899]) );
  DFF \ereg_reg[900]  ( .D(ereg_next[900]), .CLK(clk), .RST(rst), .I(e[900]), 
        .Q(ein[900]) );
  DFF \ereg_reg[901]  ( .D(ereg_next[901]), .CLK(clk), .RST(rst), .I(e[901]), 
        .Q(ein[901]) );
  DFF \ereg_reg[902]  ( .D(ereg_next[902]), .CLK(clk), .RST(rst), .I(e[902]), 
        .Q(ein[902]) );
  DFF \ereg_reg[903]  ( .D(ereg_next[903]), .CLK(clk), .RST(rst), .I(e[903]), 
        .Q(ein[903]) );
  DFF \ereg_reg[904]  ( .D(ereg_next[904]), .CLK(clk), .RST(rst), .I(e[904]), 
        .Q(ein[904]) );
  DFF \ereg_reg[905]  ( .D(ereg_next[905]), .CLK(clk), .RST(rst), .I(e[905]), 
        .Q(ein[905]) );
  DFF \ereg_reg[906]  ( .D(ereg_next[906]), .CLK(clk), .RST(rst), .I(e[906]), 
        .Q(ein[906]) );
  DFF \ereg_reg[907]  ( .D(ereg_next[907]), .CLK(clk), .RST(rst), .I(e[907]), 
        .Q(ein[907]) );
  DFF \ereg_reg[908]  ( .D(ereg_next[908]), .CLK(clk), .RST(rst), .I(e[908]), 
        .Q(ein[908]) );
  DFF \ereg_reg[909]  ( .D(ereg_next[909]), .CLK(clk), .RST(rst), .I(e[909]), 
        .Q(ein[909]) );
  DFF \ereg_reg[910]  ( .D(ereg_next[910]), .CLK(clk), .RST(rst), .I(e[910]), 
        .Q(ein[910]) );
  DFF \ereg_reg[911]  ( .D(ereg_next[911]), .CLK(clk), .RST(rst), .I(e[911]), 
        .Q(ein[911]) );
  DFF \ereg_reg[912]  ( .D(ereg_next[912]), .CLK(clk), .RST(rst), .I(e[912]), 
        .Q(ein[912]) );
  DFF \ereg_reg[913]  ( .D(ereg_next[913]), .CLK(clk), .RST(rst), .I(e[913]), 
        .Q(ein[913]) );
  DFF \ereg_reg[914]  ( .D(ereg_next[914]), .CLK(clk), .RST(rst), .I(e[914]), 
        .Q(ein[914]) );
  DFF \ereg_reg[915]  ( .D(ereg_next[915]), .CLK(clk), .RST(rst), .I(e[915]), 
        .Q(ein[915]) );
  DFF \ereg_reg[916]  ( .D(ereg_next[916]), .CLK(clk), .RST(rst), .I(e[916]), 
        .Q(ein[916]) );
  DFF \ereg_reg[917]  ( .D(ereg_next[917]), .CLK(clk), .RST(rst), .I(e[917]), 
        .Q(ein[917]) );
  DFF \ereg_reg[918]  ( .D(ereg_next[918]), .CLK(clk), .RST(rst), .I(e[918]), 
        .Q(ein[918]) );
  DFF \ereg_reg[919]  ( .D(ereg_next[919]), .CLK(clk), .RST(rst), .I(e[919]), 
        .Q(ein[919]) );
  DFF \ereg_reg[920]  ( .D(ereg_next[920]), .CLK(clk), .RST(rst), .I(e[920]), 
        .Q(ein[920]) );
  DFF \ereg_reg[921]  ( .D(ereg_next[921]), .CLK(clk), .RST(rst), .I(e[921]), 
        .Q(ein[921]) );
  DFF \ereg_reg[922]  ( .D(ereg_next[922]), .CLK(clk), .RST(rst), .I(e[922]), 
        .Q(ein[922]) );
  DFF \ereg_reg[923]  ( .D(ereg_next[923]), .CLK(clk), .RST(rst), .I(e[923]), 
        .Q(ein[923]) );
  DFF \ereg_reg[924]  ( .D(ereg_next[924]), .CLK(clk), .RST(rst), .I(e[924]), 
        .Q(ein[924]) );
  DFF \ereg_reg[925]  ( .D(ereg_next[925]), .CLK(clk), .RST(rst), .I(e[925]), 
        .Q(ein[925]) );
  DFF \ereg_reg[926]  ( .D(ereg_next[926]), .CLK(clk), .RST(rst), .I(e[926]), 
        .Q(ein[926]) );
  DFF \ereg_reg[927]  ( .D(ereg_next[927]), .CLK(clk), .RST(rst), .I(e[927]), 
        .Q(ein[927]) );
  DFF \ereg_reg[928]  ( .D(ereg_next[928]), .CLK(clk), .RST(rst), .I(e[928]), 
        .Q(ein[928]) );
  DFF \ereg_reg[929]  ( .D(ereg_next[929]), .CLK(clk), .RST(rst), .I(e[929]), 
        .Q(ein[929]) );
  DFF \ereg_reg[930]  ( .D(ereg_next[930]), .CLK(clk), .RST(rst), .I(e[930]), 
        .Q(ein[930]) );
  DFF \ereg_reg[931]  ( .D(ereg_next[931]), .CLK(clk), .RST(rst), .I(e[931]), 
        .Q(ein[931]) );
  DFF \ereg_reg[932]  ( .D(ereg_next[932]), .CLK(clk), .RST(rst), .I(e[932]), 
        .Q(ein[932]) );
  DFF \ereg_reg[933]  ( .D(ereg_next[933]), .CLK(clk), .RST(rst), .I(e[933]), 
        .Q(ein[933]) );
  DFF \ereg_reg[934]  ( .D(ereg_next[934]), .CLK(clk), .RST(rst), .I(e[934]), 
        .Q(ein[934]) );
  DFF \ereg_reg[935]  ( .D(ereg_next[935]), .CLK(clk), .RST(rst), .I(e[935]), 
        .Q(ein[935]) );
  DFF \ereg_reg[936]  ( .D(ereg_next[936]), .CLK(clk), .RST(rst), .I(e[936]), 
        .Q(ein[936]) );
  DFF \ereg_reg[937]  ( .D(ereg_next[937]), .CLK(clk), .RST(rst), .I(e[937]), 
        .Q(ein[937]) );
  DFF \ereg_reg[938]  ( .D(ereg_next[938]), .CLK(clk), .RST(rst), .I(e[938]), 
        .Q(ein[938]) );
  DFF \ereg_reg[939]  ( .D(ereg_next[939]), .CLK(clk), .RST(rst), .I(e[939]), 
        .Q(ein[939]) );
  DFF \ereg_reg[940]  ( .D(ereg_next[940]), .CLK(clk), .RST(rst), .I(e[940]), 
        .Q(ein[940]) );
  DFF \ereg_reg[941]  ( .D(ereg_next[941]), .CLK(clk), .RST(rst), .I(e[941]), 
        .Q(ein[941]) );
  DFF \ereg_reg[942]  ( .D(ereg_next[942]), .CLK(clk), .RST(rst), .I(e[942]), 
        .Q(ein[942]) );
  DFF \ereg_reg[943]  ( .D(ereg_next[943]), .CLK(clk), .RST(rst), .I(e[943]), 
        .Q(ein[943]) );
  DFF \ereg_reg[944]  ( .D(ereg_next[944]), .CLK(clk), .RST(rst), .I(e[944]), 
        .Q(ein[944]) );
  DFF \ereg_reg[945]  ( .D(ereg_next[945]), .CLK(clk), .RST(rst), .I(e[945]), 
        .Q(ein[945]) );
  DFF \ereg_reg[946]  ( .D(ereg_next[946]), .CLK(clk), .RST(rst), .I(e[946]), 
        .Q(ein[946]) );
  DFF \ereg_reg[947]  ( .D(ereg_next[947]), .CLK(clk), .RST(rst), .I(e[947]), 
        .Q(ein[947]) );
  DFF \ereg_reg[948]  ( .D(ereg_next[948]), .CLK(clk), .RST(rst), .I(e[948]), 
        .Q(ein[948]) );
  DFF \ereg_reg[949]  ( .D(ereg_next[949]), .CLK(clk), .RST(rst), .I(e[949]), 
        .Q(ein[949]) );
  DFF \ereg_reg[950]  ( .D(ereg_next[950]), .CLK(clk), .RST(rst), .I(e[950]), 
        .Q(ein[950]) );
  DFF \ereg_reg[951]  ( .D(ereg_next[951]), .CLK(clk), .RST(rst), .I(e[951]), 
        .Q(ein[951]) );
  DFF \ereg_reg[952]  ( .D(ereg_next[952]), .CLK(clk), .RST(rst), .I(e[952]), 
        .Q(ein[952]) );
  DFF \ereg_reg[953]  ( .D(ereg_next[953]), .CLK(clk), .RST(rst), .I(e[953]), 
        .Q(ein[953]) );
  DFF \ereg_reg[954]  ( .D(ereg_next[954]), .CLK(clk), .RST(rst), .I(e[954]), 
        .Q(ein[954]) );
  DFF \ereg_reg[955]  ( .D(ereg_next[955]), .CLK(clk), .RST(rst), .I(e[955]), 
        .Q(ein[955]) );
  DFF \ereg_reg[956]  ( .D(ereg_next[956]), .CLK(clk), .RST(rst), .I(e[956]), 
        .Q(ein[956]) );
  DFF \ereg_reg[957]  ( .D(ereg_next[957]), .CLK(clk), .RST(rst), .I(e[957]), 
        .Q(ein[957]) );
  DFF \ereg_reg[958]  ( .D(ereg_next[958]), .CLK(clk), .RST(rst), .I(e[958]), 
        .Q(ein[958]) );
  DFF \ereg_reg[959]  ( .D(ereg_next[959]), .CLK(clk), .RST(rst), .I(e[959]), 
        .Q(ein[959]) );
  DFF \ereg_reg[960]  ( .D(ereg_next[960]), .CLK(clk), .RST(rst), .I(e[960]), 
        .Q(ein[960]) );
  DFF \ereg_reg[961]  ( .D(ereg_next[961]), .CLK(clk), .RST(rst), .I(e[961]), 
        .Q(ein[961]) );
  DFF \ereg_reg[962]  ( .D(ereg_next[962]), .CLK(clk), .RST(rst), .I(e[962]), 
        .Q(ein[962]) );
  DFF \ereg_reg[963]  ( .D(ereg_next[963]), .CLK(clk), .RST(rst), .I(e[963]), 
        .Q(ein[963]) );
  DFF \ereg_reg[964]  ( .D(ereg_next[964]), .CLK(clk), .RST(rst), .I(e[964]), 
        .Q(ein[964]) );
  DFF \ereg_reg[965]  ( .D(ereg_next[965]), .CLK(clk), .RST(rst), .I(e[965]), 
        .Q(ein[965]) );
  DFF \ereg_reg[966]  ( .D(ereg_next[966]), .CLK(clk), .RST(rst), .I(e[966]), 
        .Q(ein[966]) );
  DFF \ereg_reg[967]  ( .D(ereg_next[967]), .CLK(clk), .RST(rst), .I(e[967]), 
        .Q(ein[967]) );
  DFF \ereg_reg[968]  ( .D(ereg_next[968]), .CLK(clk), .RST(rst), .I(e[968]), 
        .Q(ein[968]) );
  DFF \ereg_reg[969]  ( .D(ereg_next[969]), .CLK(clk), .RST(rst), .I(e[969]), 
        .Q(ein[969]) );
  DFF \ereg_reg[970]  ( .D(ereg_next[970]), .CLK(clk), .RST(rst), .I(e[970]), 
        .Q(ein[970]) );
  DFF \ereg_reg[971]  ( .D(ereg_next[971]), .CLK(clk), .RST(rst), .I(e[971]), 
        .Q(ein[971]) );
  DFF \ereg_reg[972]  ( .D(ereg_next[972]), .CLK(clk), .RST(rst), .I(e[972]), 
        .Q(ein[972]) );
  DFF \ereg_reg[973]  ( .D(ereg_next[973]), .CLK(clk), .RST(rst), .I(e[973]), 
        .Q(ein[973]) );
  DFF \ereg_reg[974]  ( .D(ereg_next[974]), .CLK(clk), .RST(rst), .I(e[974]), 
        .Q(ein[974]) );
  DFF \ereg_reg[975]  ( .D(ereg_next[975]), .CLK(clk), .RST(rst), .I(e[975]), 
        .Q(ein[975]) );
  DFF \ereg_reg[976]  ( .D(ereg_next[976]), .CLK(clk), .RST(rst), .I(e[976]), 
        .Q(ein[976]) );
  DFF \ereg_reg[977]  ( .D(ereg_next[977]), .CLK(clk), .RST(rst), .I(e[977]), 
        .Q(ein[977]) );
  DFF \ereg_reg[978]  ( .D(ereg_next[978]), .CLK(clk), .RST(rst), .I(e[978]), 
        .Q(ein[978]) );
  DFF \ereg_reg[979]  ( .D(ereg_next[979]), .CLK(clk), .RST(rst), .I(e[979]), 
        .Q(ein[979]) );
  DFF \ereg_reg[980]  ( .D(ereg_next[980]), .CLK(clk), .RST(rst), .I(e[980]), 
        .Q(ein[980]) );
  DFF \ereg_reg[981]  ( .D(ereg_next[981]), .CLK(clk), .RST(rst), .I(e[981]), 
        .Q(ein[981]) );
  DFF \ereg_reg[982]  ( .D(ereg_next[982]), .CLK(clk), .RST(rst), .I(e[982]), 
        .Q(ein[982]) );
  DFF \ereg_reg[983]  ( .D(ereg_next[983]), .CLK(clk), .RST(rst), .I(e[983]), 
        .Q(ein[983]) );
  DFF \ereg_reg[984]  ( .D(ereg_next[984]), .CLK(clk), .RST(rst), .I(e[984]), 
        .Q(ein[984]) );
  DFF \ereg_reg[985]  ( .D(ereg_next[985]), .CLK(clk), .RST(rst), .I(e[985]), 
        .Q(ein[985]) );
  DFF \ereg_reg[986]  ( .D(ereg_next[986]), .CLK(clk), .RST(rst), .I(e[986]), 
        .Q(ein[986]) );
  DFF \ereg_reg[987]  ( .D(ereg_next[987]), .CLK(clk), .RST(rst), .I(e[987]), 
        .Q(ein[987]) );
  DFF \ereg_reg[988]  ( .D(ereg_next[988]), .CLK(clk), .RST(rst), .I(e[988]), 
        .Q(ein[988]) );
  DFF \ereg_reg[989]  ( .D(ereg_next[989]), .CLK(clk), .RST(rst), .I(e[989]), 
        .Q(ein[989]) );
  DFF \ereg_reg[990]  ( .D(ereg_next[990]), .CLK(clk), .RST(rst), .I(e[990]), 
        .Q(ein[990]) );
  DFF \ereg_reg[991]  ( .D(ereg_next[991]), .CLK(clk), .RST(rst), .I(e[991]), 
        .Q(ein[991]) );
  DFF \ereg_reg[992]  ( .D(ereg_next[992]), .CLK(clk), .RST(rst), .I(e[992]), 
        .Q(ein[992]) );
  DFF \ereg_reg[993]  ( .D(ereg_next[993]), .CLK(clk), .RST(rst), .I(e[993]), 
        .Q(ein[993]) );
  DFF \ereg_reg[994]  ( .D(ereg_next[994]), .CLK(clk), .RST(rst), .I(e[994]), 
        .Q(ein[994]) );
  DFF \ereg_reg[995]  ( .D(ereg_next[995]), .CLK(clk), .RST(rst), .I(e[995]), 
        .Q(ein[995]) );
  DFF \ereg_reg[996]  ( .D(ereg_next[996]), .CLK(clk), .RST(rst), .I(e[996]), 
        .Q(ein[996]) );
  DFF \ereg_reg[997]  ( .D(ereg_next[997]), .CLK(clk), .RST(rst), .I(e[997]), 
        .Q(ein[997]) );
  DFF \ereg_reg[998]  ( .D(ereg_next[998]), .CLK(clk), .RST(rst), .I(e[998]), 
        .Q(ein[998]) );
  DFF \ereg_reg[999]  ( .D(ereg_next[999]), .CLK(clk), .RST(rst), .I(e[999]), 
        .Q(ein[999]) );
  DFF \ereg_reg[1000]  ( .D(ereg_next[1000]), .CLK(clk), .RST(rst), .I(e[1000]), .Q(ein[1000]) );
  DFF \ereg_reg[1001]  ( .D(ereg_next[1001]), .CLK(clk), .RST(rst), .I(e[1001]), .Q(ein[1001]) );
  DFF \ereg_reg[1002]  ( .D(ereg_next[1002]), .CLK(clk), .RST(rst), .I(e[1002]), .Q(ein[1002]) );
  DFF \ereg_reg[1003]  ( .D(ereg_next[1003]), .CLK(clk), .RST(rst), .I(e[1003]), .Q(ein[1003]) );
  DFF \ereg_reg[1004]  ( .D(ereg_next[1004]), .CLK(clk), .RST(rst), .I(e[1004]), .Q(ein[1004]) );
  DFF \ereg_reg[1005]  ( .D(ereg_next[1005]), .CLK(clk), .RST(rst), .I(e[1005]), .Q(ein[1005]) );
  DFF \ereg_reg[1006]  ( .D(ereg_next[1006]), .CLK(clk), .RST(rst), .I(e[1006]), .Q(ein[1006]) );
  DFF \ereg_reg[1007]  ( .D(ereg_next[1007]), .CLK(clk), .RST(rst), .I(e[1007]), .Q(ein[1007]) );
  DFF \ereg_reg[1008]  ( .D(ereg_next[1008]), .CLK(clk), .RST(rst), .I(e[1008]), .Q(ein[1008]) );
  DFF \ereg_reg[1009]  ( .D(ereg_next[1009]), .CLK(clk), .RST(rst), .I(e[1009]), .Q(ein[1009]) );
  DFF \ereg_reg[1010]  ( .D(ereg_next[1010]), .CLK(clk), .RST(rst), .I(e[1010]), .Q(ein[1010]) );
  DFF \ereg_reg[1011]  ( .D(ereg_next[1011]), .CLK(clk), .RST(rst), .I(e[1011]), .Q(ein[1011]) );
  DFF \ereg_reg[1012]  ( .D(ereg_next[1012]), .CLK(clk), .RST(rst), .I(e[1012]), .Q(ein[1012]) );
  DFF \ereg_reg[1013]  ( .D(ereg_next[1013]), .CLK(clk), .RST(rst), .I(e[1013]), .Q(ein[1013]) );
  DFF \ereg_reg[1014]  ( .D(ereg_next[1014]), .CLK(clk), .RST(rst), .I(e[1014]), .Q(ein[1014]) );
  DFF \ereg_reg[1015]  ( .D(ereg_next[1015]), .CLK(clk), .RST(rst), .I(e[1015]), .Q(ein[1015]) );
  DFF \ereg_reg[1016]  ( .D(ereg_next[1016]), .CLK(clk), .RST(rst), .I(e[1016]), .Q(ein[1016]) );
  DFF \ereg_reg[1017]  ( .D(ereg_next[1017]), .CLK(clk), .RST(rst), .I(e[1017]), .Q(ein[1017]) );
  DFF \ereg_reg[1018]  ( .D(ereg_next[1018]), .CLK(clk), .RST(rst), .I(e[1018]), .Q(ein[1018]) );
  DFF \ereg_reg[1019]  ( .D(ereg_next[1019]), .CLK(clk), .RST(rst), .I(e[1019]), .Q(ein[1019]) );
  DFF \ereg_reg[1020]  ( .D(ereg_next[1020]), .CLK(clk), .RST(rst), .I(e[1020]), .Q(ein[1020]) );
  DFF \ereg_reg[1021]  ( .D(ereg_next[1021]), .CLK(clk), .RST(rst), .I(e[1021]), .Q(ein[1021]) );
  DFF \ereg_reg[1022]  ( .D(ereg_next[1022]), .CLK(clk), .RST(rst), .I(e[1022]), .Q(ein[1022]) );
  DFF \ereg_reg[1023]  ( .D(ereg_next[1023]), .CLK(clk), .RST(rst), .I(e[1023]), .Q(ein[1023]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  DFF \creg_reg[256]  ( .D(creg_next[256]), .CLK(clk), .RST(rst), .I(m[256]), 
        .Q(c[256]) );
  DFF \creg_reg[257]  ( .D(creg_next[257]), .CLK(clk), .RST(rst), .I(m[257]), 
        .Q(c[257]) );
  DFF \creg_reg[258]  ( .D(creg_next[258]), .CLK(clk), .RST(rst), .I(m[258]), 
        .Q(c[258]) );
  DFF \creg_reg[259]  ( .D(creg_next[259]), .CLK(clk), .RST(rst), .I(m[259]), 
        .Q(c[259]) );
  DFF \creg_reg[260]  ( .D(creg_next[260]), .CLK(clk), .RST(rst), .I(m[260]), 
        .Q(c[260]) );
  DFF \creg_reg[261]  ( .D(creg_next[261]), .CLK(clk), .RST(rst), .I(m[261]), 
        .Q(c[261]) );
  DFF \creg_reg[262]  ( .D(creg_next[262]), .CLK(clk), .RST(rst), .I(m[262]), 
        .Q(c[262]) );
  DFF \creg_reg[263]  ( .D(creg_next[263]), .CLK(clk), .RST(rst), .I(m[263]), 
        .Q(c[263]) );
  DFF \creg_reg[264]  ( .D(creg_next[264]), .CLK(clk), .RST(rst), .I(m[264]), 
        .Q(c[264]) );
  DFF \creg_reg[265]  ( .D(creg_next[265]), .CLK(clk), .RST(rst), .I(m[265]), 
        .Q(c[265]) );
  DFF \creg_reg[266]  ( .D(creg_next[266]), .CLK(clk), .RST(rst), .I(m[266]), 
        .Q(c[266]) );
  DFF \creg_reg[267]  ( .D(creg_next[267]), .CLK(clk), .RST(rst), .I(m[267]), 
        .Q(c[267]) );
  DFF \creg_reg[268]  ( .D(creg_next[268]), .CLK(clk), .RST(rst), .I(m[268]), 
        .Q(c[268]) );
  DFF \creg_reg[269]  ( .D(creg_next[269]), .CLK(clk), .RST(rst), .I(m[269]), 
        .Q(c[269]) );
  DFF \creg_reg[270]  ( .D(creg_next[270]), .CLK(clk), .RST(rst), .I(m[270]), 
        .Q(c[270]) );
  DFF \creg_reg[271]  ( .D(creg_next[271]), .CLK(clk), .RST(rst), .I(m[271]), 
        .Q(c[271]) );
  DFF \creg_reg[272]  ( .D(creg_next[272]), .CLK(clk), .RST(rst), .I(m[272]), 
        .Q(c[272]) );
  DFF \creg_reg[273]  ( .D(creg_next[273]), .CLK(clk), .RST(rst), .I(m[273]), 
        .Q(c[273]) );
  DFF \creg_reg[274]  ( .D(creg_next[274]), .CLK(clk), .RST(rst), .I(m[274]), 
        .Q(c[274]) );
  DFF \creg_reg[275]  ( .D(creg_next[275]), .CLK(clk), .RST(rst), .I(m[275]), 
        .Q(c[275]) );
  DFF \creg_reg[276]  ( .D(creg_next[276]), .CLK(clk), .RST(rst), .I(m[276]), 
        .Q(c[276]) );
  DFF \creg_reg[277]  ( .D(creg_next[277]), .CLK(clk), .RST(rst), .I(m[277]), 
        .Q(c[277]) );
  DFF \creg_reg[278]  ( .D(creg_next[278]), .CLK(clk), .RST(rst), .I(m[278]), 
        .Q(c[278]) );
  DFF \creg_reg[279]  ( .D(creg_next[279]), .CLK(clk), .RST(rst), .I(m[279]), 
        .Q(c[279]) );
  DFF \creg_reg[280]  ( .D(creg_next[280]), .CLK(clk), .RST(rst), .I(m[280]), 
        .Q(c[280]) );
  DFF \creg_reg[281]  ( .D(creg_next[281]), .CLK(clk), .RST(rst), .I(m[281]), 
        .Q(c[281]) );
  DFF \creg_reg[282]  ( .D(creg_next[282]), .CLK(clk), .RST(rst), .I(m[282]), 
        .Q(c[282]) );
  DFF \creg_reg[283]  ( .D(creg_next[283]), .CLK(clk), .RST(rst), .I(m[283]), 
        .Q(c[283]) );
  DFF \creg_reg[284]  ( .D(creg_next[284]), .CLK(clk), .RST(rst), .I(m[284]), 
        .Q(c[284]) );
  DFF \creg_reg[285]  ( .D(creg_next[285]), .CLK(clk), .RST(rst), .I(m[285]), 
        .Q(c[285]) );
  DFF \creg_reg[286]  ( .D(creg_next[286]), .CLK(clk), .RST(rst), .I(m[286]), 
        .Q(c[286]) );
  DFF \creg_reg[287]  ( .D(creg_next[287]), .CLK(clk), .RST(rst), .I(m[287]), 
        .Q(c[287]) );
  DFF \creg_reg[288]  ( .D(creg_next[288]), .CLK(clk), .RST(rst), .I(m[288]), 
        .Q(c[288]) );
  DFF \creg_reg[289]  ( .D(creg_next[289]), .CLK(clk), .RST(rst), .I(m[289]), 
        .Q(c[289]) );
  DFF \creg_reg[290]  ( .D(creg_next[290]), .CLK(clk), .RST(rst), .I(m[290]), 
        .Q(c[290]) );
  DFF \creg_reg[291]  ( .D(creg_next[291]), .CLK(clk), .RST(rst), .I(m[291]), 
        .Q(c[291]) );
  DFF \creg_reg[292]  ( .D(creg_next[292]), .CLK(clk), .RST(rst), .I(m[292]), 
        .Q(c[292]) );
  DFF \creg_reg[293]  ( .D(creg_next[293]), .CLK(clk), .RST(rst), .I(m[293]), 
        .Q(c[293]) );
  DFF \creg_reg[294]  ( .D(creg_next[294]), .CLK(clk), .RST(rst), .I(m[294]), 
        .Q(c[294]) );
  DFF \creg_reg[295]  ( .D(creg_next[295]), .CLK(clk), .RST(rst), .I(m[295]), 
        .Q(c[295]) );
  DFF \creg_reg[296]  ( .D(creg_next[296]), .CLK(clk), .RST(rst), .I(m[296]), 
        .Q(c[296]) );
  DFF \creg_reg[297]  ( .D(creg_next[297]), .CLK(clk), .RST(rst), .I(m[297]), 
        .Q(c[297]) );
  DFF \creg_reg[298]  ( .D(creg_next[298]), .CLK(clk), .RST(rst), .I(m[298]), 
        .Q(c[298]) );
  DFF \creg_reg[299]  ( .D(creg_next[299]), .CLK(clk), .RST(rst), .I(m[299]), 
        .Q(c[299]) );
  DFF \creg_reg[300]  ( .D(creg_next[300]), .CLK(clk), .RST(rst), .I(m[300]), 
        .Q(c[300]) );
  DFF \creg_reg[301]  ( .D(creg_next[301]), .CLK(clk), .RST(rst), .I(m[301]), 
        .Q(c[301]) );
  DFF \creg_reg[302]  ( .D(creg_next[302]), .CLK(clk), .RST(rst), .I(m[302]), 
        .Q(c[302]) );
  DFF \creg_reg[303]  ( .D(creg_next[303]), .CLK(clk), .RST(rst), .I(m[303]), 
        .Q(c[303]) );
  DFF \creg_reg[304]  ( .D(creg_next[304]), .CLK(clk), .RST(rst), .I(m[304]), 
        .Q(c[304]) );
  DFF \creg_reg[305]  ( .D(creg_next[305]), .CLK(clk), .RST(rst), .I(m[305]), 
        .Q(c[305]) );
  DFF \creg_reg[306]  ( .D(creg_next[306]), .CLK(clk), .RST(rst), .I(m[306]), 
        .Q(c[306]) );
  DFF \creg_reg[307]  ( .D(creg_next[307]), .CLK(clk), .RST(rst), .I(m[307]), 
        .Q(c[307]) );
  DFF \creg_reg[308]  ( .D(creg_next[308]), .CLK(clk), .RST(rst), .I(m[308]), 
        .Q(c[308]) );
  DFF \creg_reg[309]  ( .D(creg_next[309]), .CLK(clk), .RST(rst), .I(m[309]), 
        .Q(c[309]) );
  DFF \creg_reg[310]  ( .D(creg_next[310]), .CLK(clk), .RST(rst), .I(m[310]), 
        .Q(c[310]) );
  DFF \creg_reg[311]  ( .D(creg_next[311]), .CLK(clk), .RST(rst), .I(m[311]), 
        .Q(c[311]) );
  DFF \creg_reg[312]  ( .D(creg_next[312]), .CLK(clk), .RST(rst), .I(m[312]), 
        .Q(c[312]) );
  DFF \creg_reg[313]  ( .D(creg_next[313]), .CLK(clk), .RST(rst), .I(m[313]), 
        .Q(c[313]) );
  DFF \creg_reg[314]  ( .D(creg_next[314]), .CLK(clk), .RST(rst), .I(m[314]), 
        .Q(c[314]) );
  DFF \creg_reg[315]  ( .D(creg_next[315]), .CLK(clk), .RST(rst), .I(m[315]), 
        .Q(c[315]) );
  DFF \creg_reg[316]  ( .D(creg_next[316]), .CLK(clk), .RST(rst), .I(m[316]), 
        .Q(c[316]) );
  DFF \creg_reg[317]  ( .D(creg_next[317]), .CLK(clk), .RST(rst), .I(m[317]), 
        .Q(c[317]) );
  DFF \creg_reg[318]  ( .D(creg_next[318]), .CLK(clk), .RST(rst), .I(m[318]), 
        .Q(c[318]) );
  DFF \creg_reg[319]  ( .D(creg_next[319]), .CLK(clk), .RST(rst), .I(m[319]), 
        .Q(c[319]) );
  DFF \creg_reg[320]  ( .D(creg_next[320]), .CLK(clk), .RST(rst), .I(m[320]), 
        .Q(c[320]) );
  DFF \creg_reg[321]  ( .D(creg_next[321]), .CLK(clk), .RST(rst), .I(m[321]), 
        .Q(c[321]) );
  DFF \creg_reg[322]  ( .D(creg_next[322]), .CLK(clk), .RST(rst), .I(m[322]), 
        .Q(c[322]) );
  DFF \creg_reg[323]  ( .D(creg_next[323]), .CLK(clk), .RST(rst), .I(m[323]), 
        .Q(c[323]) );
  DFF \creg_reg[324]  ( .D(creg_next[324]), .CLK(clk), .RST(rst), .I(m[324]), 
        .Q(c[324]) );
  DFF \creg_reg[325]  ( .D(creg_next[325]), .CLK(clk), .RST(rst), .I(m[325]), 
        .Q(c[325]) );
  DFF \creg_reg[326]  ( .D(creg_next[326]), .CLK(clk), .RST(rst), .I(m[326]), 
        .Q(c[326]) );
  DFF \creg_reg[327]  ( .D(creg_next[327]), .CLK(clk), .RST(rst), .I(m[327]), 
        .Q(c[327]) );
  DFF \creg_reg[328]  ( .D(creg_next[328]), .CLK(clk), .RST(rst), .I(m[328]), 
        .Q(c[328]) );
  DFF \creg_reg[329]  ( .D(creg_next[329]), .CLK(clk), .RST(rst), .I(m[329]), 
        .Q(c[329]) );
  DFF \creg_reg[330]  ( .D(creg_next[330]), .CLK(clk), .RST(rst), .I(m[330]), 
        .Q(c[330]) );
  DFF \creg_reg[331]  ( .D(creg_next[331]), .CLK(clk), .RST(rst), .I(m[331]), 
        .Q(c[331]) );
  DFF \creg_reg[332]  ( .D(creg_next[332]), .CLK(clk), .RST(rst), .I(m[332]), 
        .Q(c[332]) );
  DFF \creg_reg[333]  ( .D(creg_next[333]), .CLK(clk), .RST(rst), .I(m[333]), 
        .Q(c[333]) );
  DFF \creg_reg[334]  ( .D(creg_next[334]), .CLK(clk), .RST(rst), .I(m[334]), 
        .Q(c[334]) );
  DFF \creg_reg[335]  ( .D(creg_next[335]), .CLK(clk), .RST(rst), .I(m[335]), 
        .Q(c[335]) );
  DFF \creg_reg[336]  ( .D(creg_next[336]), .CLK(clk), .RST(rst), .I(m[336]), 
        .Q(c[336]) );
  DFF \creg_reg[337]  ( .D(creg_next[337]), .CLK(clk), .RST(rst), .I(m[337]), 
        .Q(c[337]) );
  DFF \creg_reg[338]  ( .D(creg_next[338]), .CLK(clk), .RST(rst), .I(m[338]), 
        .Q(c[338]) );
  DFF \creg_reg[339]  ( .D(creg_next[339]), .CLK(clk), .RST(rst), .I(m[339]), 
        .Q(c[339]) );
  DFF \creg_reg[340]  ( .D(creg_next[340]), .CLK(clk), .RST(rst), .I(m[340]), 
        .Q(c[340]) );
  DFF \creg_reg[341]  ( .D(creg_next[341]), .CLK(clk), .RST(rst), .I(m[341]), 
        .Q(c[341]) );
  DFF \creg_reg[342]  ( .D(creg_next[342]), .CLK(clk), .RST(rst), .I(m[342]), 
        .Q(c[342]) );
  DFF \creg_reg[343]  ( .D(creg_next[343]), .CLK(clk), .RST(rst), .I(m[343]), 
        .Q(c[343]) );
  DFF \creg_reg[344]  ( .D(creg_next[344]), .CLK(clk), .RST(rst), .I(m[344]), 
        .Q(c[344]) );
  DFF \creg_reg[345]  ( .D(creg_next[345]), .CLK(clk), .RST(rst), .I(m[345]), 
        .Q(c[345]) );
  DFF \creg_reg[346]  ( .D(creg_next[346]), .CLK(clk), .RST(rst), .I(m[346]), 
        .Q(c[346]) );
  DFF \creg_reg[347]  ( .D(creg_next[347]), .CLK(clk), .RST(rst), .I(m[347]), 
        .Q(c[347]) );
  DFF \creg_reg[348]  ( .D(creg_next[348]), .CLK(clk), .RST(rst), .I(m[348]), 
        .Q(c[348]) );
  DFF \creg_reg[349]  ( .D(creg_next[349]), .CLK(clk), .RST(rst), .I(m[349]), 
        .Q(c[349]) );
  DFF \creg_reg[350]  ( .D(creg_next[350]), .CLK(clk), .RST(rst), .I(m[350]), 
        .Q(c[350]) );
  DFF \creg_reg[351]  ( .D(creg_next[351]), .CLK(clk), .RST(rst), .I(m[351]), 
        .Q(c[351]) );
  DFF \creg_reg[352]  ( .D(creg_next[352]), .CLK(clk), .RST(rst), .I(m[352]), 
        .Q(c[352]) );
  DFF \creg_reg[353]  ( .D(creg_next[353]), .CLK(clk), .RST(rst), .I(m[353]), 
        .Q(c[353]) );
  DFF \creg_reg[354]  ( .D(creg_next[354]), .CLK(clk), .RST(rst), .I(m[354]), 
        .Q(c[354]) );
  DFF \creg_reg[355]  ( .D(creg_next[355]), .CLK(clk), .RST(rst), .I(m[355]), 
        .Q(c[355]) );
  DFF \creg_reg[356]  ( .D(creg_next[356]), .CLK(clk), .RST(rst), .I(m[356]), 
        .Q(c[356]) );
  DFF \creg_reg[357]  ( .D(creg_next[357]), .CLK(clk), .RST(rst), .I(m[357]), 
        .Q(c[357]) );
  DFF \creg_reg[358]  ( .D(creg_next[358]), .CLK(clk), .RST(rst), .I(m[358]), 
        .Q(c[358]) );
  DFF \creg_reg[359]  ( .D(creg_next[359]), .CLK(clk), .RST(rst), .I(m[359]), 
        .Q(c[359]) );
  DFF \creg_reg[360]  ( .D(creg_next[360]), .CLK(clk), .RST(rst), .I(m[360]), 
        .Q(c[360]) );
  DFF \creg_reg[361]  ( .D(creg_next[361]), .CLK(clk), .RST(rst), .I(m[361]), 
        .Q(c[361]) );
  DFF \creg_reg[362]  ( .D(creg_next[362]), .CLK(clk), .RST(rst), .I(m[362]), 
        .Q(c[362]) );
  DFF \creg_reg[363]  ( .D(creg_next[363]), .CLK(clk), .RST(rst), .I(m[363]), 
        .Q(c[363]) );
  DFF \creg_reg[364]  ( .D(creg_next[364]), .CLK(clk), .RST(rst), .I(m[364]), 
        .Q(c[364]) );
  DFF \creg_reg[365]  ( .D(creg_next[365]), .CLK(clk), .RST(rst), .I(m[365]), 
        .Q(c[365]) );
  DFF \creg_reg[366]  ( .D(creg_next[366]), .CLK(clk), .RST(rst), .I(m[366]), 
        .Q(c[366]) );
  DFF \creg_reg[367]  ( .D(creg_next[367]), .CLK(clk), .RST(rst), .I(m[367]), 
        .Q(c[367]) );
  DFF \creg_reg[368]  ( .D(creg_next[368]), .CLK(clk), .RST(rst), .I(m[368]), 
        .Q(c[368]) );
  DFF \creg_reg[369]  ( .D(creg_next[369]), .CLK(clk), .RST(rst), .I(m[369]), 
        .Q(c[369]) );
  DFF \creg_reg[370]  ( .D(creg_next[370]), .CLK(clk), .RST(rst), .I(m[370]), 
        .Q(c[370]) );
  DFF \creg_reg[371]  ( .D(creg_next[371]), .CLK(clk), .RST(rst), .I(m[371]), 
        .Q(c[371]) );
  DFF \creg_reg[372]  ( .D(creg_next[372]), .CLK(clk), .RST(rst), .I(m[372]), 
        .Q(c[372]) );
  DFF \creg_reg[373]  ( .D(creg_next[373]), .CLK(clk), .RST(rst), .I(m[373]), 
        .Q(c[373]) );
  DFF \creg_reg[374]  ( .D(creg_next[374]), .CLK(clk), .RST(rst), .I(m[374]), 
        .Q(c[374]) );
  DFF \creg_reg[375]  ( .D(creg_next[375]), .CLK(clk), .RST(rst), .I(m[375]), 
        .Q(c[375]) );
  DFF \creg_reg[376]  ( .D(creg_next[376]), .CLK(clk), .RST(rst), .I(m[376]), 
        .Q(c[376]) );
  DFF \creg_reg[377]  ( .D(creg_next[377]), .CLK(clk), .RST(rst), .I(m[377]), 
        .Q(c[377]) );
  DFF \creg_reg[378]  ( .D(creg_next[378]), .CLK(clk), .RST(rst), .I(m[378]), 
        .Q(c[378]) );
  DFF \creg_reg[379]  ( .D(creg_next[379]), .CLK(clk), .RST(rst), .I(m[379]), 
        .Q(c[379]) );
  DFF \creg_reg[380]  ( .D(creg_next[380]), .CLK(clk), .RST(rst), .I(m[380]), 
        .Q(c[380]) );
  DFF \creg_reg[381]  ( .D(creg_next[381]), .CLK(clk), .RST(rst), .I(m[381]), 
        .Q(c[381]) );
  DFF \creg_reg[382]  ( .D(creg_next[382]), .CLK(clk), .RST(rst), .I(m[382]), 
        .Q(c[382]) );
  DFF \creg_reg[383]  ( .D(creg_next[383]), .CLK(clk), .RST(rst), .I(m[383]), 
        .Q(c[383]) );
  DFF \creg_reg[384]  ( .D(creg_next[384]), .CLK(clk), .RST(rst), .I(m[384]), 
        .Q(c[384]) );
  DFF \creg_reg[385]  ( .D(creg_next[385]), .CLK(clk), .RST(rst), .I(m[385]), 
        .Q(c[385]) );
  DFF \creg_reg[386]  ( .D(creg_next[386]), .CLK(clk), .RST(rst), .I(m[386]), 
        .Q(c[386]) );
  DFF \creg_reg[387]  ( .D(creg_next[387]), .CLK(clk), .RST(rst), .I(m[387]), 
        .Q(c[387]) );
  DFF \creg_reg[388]  ( .D(creg_next[388]), .CLK(clk), .RST(rst), .I(m[388]), 
        .Q(c[388]) );
  DFF \creg_reg[389]  ( .D(creg_next[389]), .CLK(clk), .RST(rst), .I(m[389]), 
        .Q(c[389]) );
  DFF \creg_reg[390]  ( .D(creg_next[390]), .CLK(clk), .RST(rst), .I(m[390]), 
        .Q(c[390]) );
  DFF \creg_reg[391]  ( .D(creg_next[391]), .CLK(clk), .RST(rst), .I(m[391]), 
        .Q(c[391]) );
  DFF \creg_reg[392]  ( .D(creg_next[392]), .CLK(clk), .RST(rst), .I(m[392]), 
        .Q(c[392]) );
  DFF \creg_reg[393]  ( .D(creg_next[393]), .CLK(clk), .RST(rst), .I(m[393]), 
        .Q(c[393]) );
  DFF \creg_reg[394]  ( .D(creg_next[394]), .CLK(clk), .RST(rst), .I(m[394]), 
        .Q(c[394]) );
  DFF \creg_reg[395]  ( .D(creg_next[395]), .CLK(clk), .RST(rst), .I(m[395]), 
        .Q(c[395]) );
  DFF \creg_reg[396]  ( .D(creg_next[396]), .CLK(clk), .RST(rst), .I(m[396]), 
        .Q(c[396]) );
  DFF \creg_reg[397]  ( .D(creg_next[397]), .CLK(clk), .RST(rst), .I(m[397]), 
        .Q(c[397]) );
  DFF \creg_reg[398]  ( .D(creg_next[398]), .CLK(clk), .RST(rst), .I(m[398]), 
        .Q(c[398]) );
  DFF \creg_reg[399]  ( .D(creg_next[399]), .CLK(clk), .RST(rst), .I(m[399]), 
        .Q(c[399]) );
  DFF \creg_reg[400]  ( .D(creg_next[400]), .CLK(clk), .RST(rst), .I(m[400]), 
        .Q(c[400]) );
  DFF \creg_reg[401]  ( .D(creg_next[401]), .CLK(clk), .RST(rst), .I(m[401]), 
        .Q(c[401]) );
  DFF \creg_reg[402]  ( .D(creg_next[402]), .CLK(clk), .RST(rst), .I(m[402]), 
        .Q(c[402]) );
  DFF \creg_reg[403]  ( .D(creg_next[403]), .CLK(clk), .RST(rst), .I(m[403]), 
        .Q(c[403]) );
  DFF \creg_reg[404]  ( .D(creg_next[404]), .CLK(clk), .RST(rst), .I(m[404]), 
        .Q(c[404]) );
  DFF \creg_reg[405]  ( .D(creg_next[405]), .CLK(clk), .RST(rst), .I(m[405]), 
        .Q(c[405]) );
  DFF \creg_reg[406]  ( .D(creg_next[406]), .CLK(clk), .RST(rst), .I(m[406]), 
        .Q(c[406]) );
  DFF \creg_reg[407]  ( .D(creg_next[407]), .CLK(clk), .RST(rst), .I(m[407]), 
        .Q(c[407]) );
  DFF \creg_reg[408]  ( .D(creg_next[408]), .CLK(clk), .RST(rst), .I(m[408]), 
        .Q(c[408]) );
  DFF \creg_reg[409]  ( .D(creg_next[409]), .CLK(clk), .RST(rst), .I(m[409]), 
        .Q(c[409]) );
  DFF \creg_reg[410]  ( .D(creg_next[410]), .CLK(clk), .RST(rst), .I(m[410]), 
        .Q(c[410]) );
  DFF \creg_reg[411]  ( .D(creg_next[411]), .CLK(clk), .RST(rst), .I(m[411]), 
        .Q(c[411]) );
  DFF \creg_reg[412]  ( .D(creg_next[412]), .CLK(clk), .RST(rst), .I(m[412]), 
        .Q(c[412]) );
  DFF \creg_reg[413]  ( .D(creg_next[413]), .CLK(clk), .RST(rst), .I(m[413]), 
        .Q(c[413]) );
  DFF \creg_reg[414]  ( .D(creg_next[414]), .CLK(clk), .RST(rst), .I(m[414]), 
        .Q(c[414]) );
  DFF \creg_reg[415]  ( .D(creg_next[415]), .CLK(clk), .RST(rst), .I(m[415]), 
        .Q(c[415]) );
  DFF \creg_reg[416]  ( .D(creg_next[416]), .CLK(clk), .RST(rst), .I(m[416]), 
        .Q(c[416]) );
  DFF \creg_reg[417]  ( .D(creg_next[417]), .CLK(clk), .RST(rst), .I(m[417]), 
        .Q(c[417]) );
  DFF \creg_reg[418]  ( .D(creg_next[418]), .CLK(clk), .RST(rst), .I(m[418]), 
        .Q(c[418]) );
  DFF \creg_reg[419]  ( .D(creg_next[419]), .CLK(clk), .RST(rst), .I(m[419]), 
        .Q(c[419]) );
  DFF \creg_reg[420]  ( .D(creg_next[420]), .CLK(clk), .RST(rst), .I(m[420]), 
        .Q(c[420]) );
  DFF \creg_reg[421]  ( .D(creg_next[421]), .CLK(clk), .RST(rst), .I(m[421]), 
        .Q(c[421]) );
  DFF \creg_reg[422]  ( .D(creg_next[422]), .CLK(clk), .RST(rst), .I(m[422]), 
        .Q(c[422]) );
  DFF \creg_reg[423]  ( .D(creg_next[423]), .CLK(clk), .RST(rst), .I(m[423]), 
        .Q(c[423]) );
  DFF \creg_reg[424]  ( .D(creg_next[424]), .CLK(clk), .RST(rst), .I(m[424]), 
        .Q(c[424]) );
  DFF \creg_reg[425]  ( .D(creg_next[425]), .CLK(clk), .RST(rst), .I(m[425]), 
        .Q(c[425]) );
  DFF \creg_reg[426]  ( .D(creg_next[426]), .CLK(clk), .RST(rst), .I(m[426]), 
        .Q(c[426]) );
  DFF \creg_reg[427]  ( .D(creg_next[427]), .CLK(clk), .RST(rst), .I(m[427]), 
        .Q(c[427]) );
  DFF \creg_reg[428]  ( .D(creg_next[428]), .CLK(clk), .RST(rst), .I(m[428]), 
        .Q(c[428]) );
  DFF \creg_reg[429]  ( .D(creg_next[429]), .CLK(clk), .RST(rst), .I(m[429]), 
        .Q(c[429]) );
  DFF \creg_reg[430]  ( .D(creg_next[430]), .CLK(clk), .RST(rst), .I(m[430]), 
        .Q(c[430]) );
  DFF \creg_reg[431]  ( .D(creg_next[431]), .CLK(clk), .RST(rst), .I(m[431]), 
        .Q(c[431]) );
  DFF \creg_reg[432]  ( .D(creg_next[432]), .CLK(clk), .RST(rst), .I(m[432]), 
        .Q(c[432]) );
  DFF \creg_reg[433]  ( .D(creg_next[433]), .CLK(clk), .RST(rst), .I(m[433]), 
        .Q(c[433]) );
  DFF \creg_reg[434]  ( .D(creg_next[434]), .CLK(clk), .RST(rst), .I(m[434]), 
        .Q(c[434]) );
  DFF \creg_reg[435]  ( .D(creg_next[435]), .CLK(clk), .RST(rst), .I(m[435]), 
        .Q(c[435]) );
  DFF \creg_reg[436]  ( .D(creg_next[436]), .CLK(clk), .RST(rst), .I(m[436]), 
        .Q(c[436]) );
  DFF \creg_reg[437]  ( .D(creg_next[437]), .CLK(clk), .RST(rst), .I(m[437]), 
        .Q(c[437]) );
  DFF \creg_reg[438]  ( .D(creg_next[438]), .CLK(clk), .RST(rst), .I(m[438]), 
        .Q(c[438]) );
  DFF \creg_reg[439]  ( .D(creg_next[439]), .CLK(clk), .RST(rst), .I(m[439]), 
        .Q(c[439]) );
  DFF \creg_reg[440]  ( .D(creg_next[440]), .CLK(clk), .RST(rst), .I(m[440]), 
        .Q(c[440]) );
  DFF \creg_reg[441]  ( .D(creg_next[441]), .CLK(clk), .RST(rst), .I(m[441]), 
        .Q(c[441]) );
  DFF \creg_reg[442]  ( .D(creg_next[442]), .CLK(clk), .RST(rst), .I(m[442]), 
        .Q(c[442]) );
  DFF \creg_reg[443]  ( .D(creg_next[443]), .CLK(clk), .RST(rst), .I(m[443]), 
        .Q(c[443]) );
  DFF \creg_reg[444]  ( .D(creg_next[444]), .CLK(clk), .RST(rst), .I(m[444]), 
        .Q(c[444]) );
  DFF \creg_reg[445]  ( .D(creg_next[445]), .CLK(clk), .RST(rst), .I(m[445]), 
        .Q(c[445]) );
  DFF \creg_reg[446]  ( .D(creg_next[446]), .CLK(clk), .RST(rst), .I(m[446]), 
        .Q(c[446]) );
  DFF \creg_reg[447]  ( .D(creg_next[447]), .CLK(clk), .RST(rst), .I(m[447]), 
        .Q(c[447]) );
  DFF \creg_reg[448]  ( .D(creg_next[448]), .CLK(clk), .RST(rst), .I(m[448]), 
        .Q(c[448]) );
  DFF \creg_reg[449]  ( .D(creg_next[449]), .CLK(clk), .RST(rst), .I(m[449]), 
        .Q(c[449]) );
  DFF \creg_reg[450]  ( .D(creg_next[450]), .CLK(clk), .RST(rst), .I(m[450]), 
        .Q(c[450]) );
  DFF \creg_reg[451]  ( .D(creg_next[451]), .CLK(clk), .RST(rst), .I(m[451]), 
        .Q(c[451]) );
  DFF \creg_reg[452]  ( .D(creg_next[452]), .CLK(clk), .RST(rst), .I(m[452]), 
        .Q(c[452]) );
  DFF \creg_reg[453]  ( .D(creg_next[453]), .CLK(clk), .RST(rst), .I(m[453]), 
        .Q(c[453]) );
  DFF \creg_reg[454]  ( .D(creg_next[454]), .CLK(clk), .RST(rst), .I(m[454]), 
        .Q(c[454]) );
  DFF \creg_reg[455]  ( .D(creg_next[455]), .CLK(clk), .RST(rst), .I(m[455]), 
        .Q(c[455]) );
  DFF \creg_reg[456]  ( .D(creg_next[456]), .CLK(clk), .RST(rst), .I(m[456]), 
        .Q(c[456]) );
  DFF \creg_reg[457]  ( .D(creg_next[457]), .CLK(clk), .RST(rst), .I(m[457]), 
        .Q(c[457]) );
  DFF \creg_reg[458]  ( .D(creg_next[458]), .CLK(clk), .RST(rst), .I(m[458]), 
        .Q(c[458]) );
  DFF \creg_reg[459]  ( .D(creg_next[459]), .CLK(clk), .RST(rst), .I(m[459]), 
        .Q(c[459]) );
  DFF \creg_reg[460]  ( .D(creg_next[460]), .CLK(clk), .RST(rst), .I(m[460]), 
        .Q(c[460]) );
  DFF \creg_reg[461]  ( .D(creg_next[461]), .CLK(clk), .RST(rst), .I(m[461]), 
        .Q(c[461]) );
  DFF \creg_reg[462]  ( .D(creg_next[462]), .CLK(clk), .RST(rst), .I(m[462]), 
        .Q(c[462]) );
  DFF \creg_reg[463]  ( .D(creg_next[463]), .CLK(clk), .RST(rst), .I(m[463]), 
        .Q(c[463]) );
  DFF \creg_reg[464]  ( .D(creg_next[464]), .CLK(clk), .RST(rst), .I(m[464]), 
        .Q(c[464]) );
  DFF \creg_reg[465]  ( .D(creg_next[465]), .CLK(clk), .RST(rst), .I(m[465]), 
        .Q(c[465]) );
  DFF \creg_reg[466]  ( .D(creg_next[466]), .CLK(clk), .RST(rst), .I(m[466]), 
        .Q(c[466]) );
  DFF \creg_reg[467]  ( .D(creg_next[467]), .CLK(clk), .RST(rst), .I(m[467]), 
        .Q(c[467]) );
  DFF \creg_reg[468]  ( .D(creg_next[468]), .CLK(clk), .RST(rst), .I(m[468]), 
        .Q(c[468]) );
  DFF \creg_reg[469]  ( .D(creg_next[469]), .CLK(clk), .RST(rst), .I(m[469]), 
        .Q(c[469]) );
  DFF \creg_reg[470]  ( .D(creg_next[470]), .CLK(clk), .RST(rst), .I(m[470]), 
        .Q(c[470]) );
  DFF \creg_reg[471]  ( .D(creg_next[471]), .CLK(clk), .RST(rst), .I(m[471]), 
        .Q(c[471]) );
  DFF \creg_reg[472]  ( .D(creg_next[472]), .CLK(clk), .RST(rst), .I(m[472]), 
        .Q(c[472]) );
  DFF \creg_reg[473]  ( .D(creg_next[473]), .CLK(clk), .RST(rst), .I(m[473]), 
        .Q(c[473]) );
  DFF \creg_reg[474]  ( .D(creg_next[474]), .CLK(clk), .RST(rst), .I(m[474]), 
        .Q(c[474]) );
  DFF \creg_reg[475]  ( .D(creg_next[475]), .CLK(clk), .RST(rst), .I(m[475]), 
        .Q(c[475]) );
  DFF \creg_reg[476]  ( .D(creg_next[476]), .CLK(clk), .RST(rst), .I(m[476]), 
        .Q(c[476]) );
  DFF \creg_reg[477]  ( .D(creg_next[477]), .CLK(clk), .RST(rst), .I(m[477]), 
        .Q(c[477]) );
  DFF \creg_reg[478]  ( .D(creg_next[478]), .CLK(clk), .RST(rst), .I(m[478]), 
        .Q(c[478]) );
  DFF \creg_reg[479]  ( .D(creg_next[479]), .CLK(clk), .RST(rst), .I(m[479]), 
        .Q(c[479]) );
  DFF \creg_reg[480]  ( .D(creg_next[480]), .CLK(clk), .RST(rst), .I(m[480]), 
        .Q(c[480]) );
  DFF \creg_reg[481]  ( .D(creg_next[481]), .CLK(clk), .RST(rst), .I(m[481]), 
        .Q(c[481]) );
  DFF \creg_reg[482]  ( .D(creg_next[482]), .CLK(clk), .RST(rst), .I(m[482]), 
        .Q(c[482]) );
  DFF \creg_reg[483]  ( .D(creg_next[483]), .CLK(clk), .RST(rst), .I(m[483]), 
        .Q(c[483]) );
  DFF \creg_reg[484]  ( .D(creg_next[484]), .CLK(clk), .RST(rst), .I(m[484]), 
        .Q(c[484]) );
  DFF \creg_reg[485]  ( .D(creg_next[485]), .CLK(clk), .RST(rst), .I(m[485]), 
        .Q(c[485]) );
  DFF \creg_reg[486]  ( .D(creg_next[486]), .CLK(clk), .RST(rst), .I(m[486]), 
        .Q(c[486]) );
  DFF \creg_reg[487]  ( .D(creg_next[487]), .CLK(clk), .RST(rst), .I(m[487]), 
        .Q(c[487]) );
  DFF \creg_reg[488]  ( .D(creg_next[488]), .CLK(clk), .RST(rst), .I(m[488]), 
        .Q(c[488]) );
  DFF \creg_reg[489]  ( .D(creg_next[489]), .CLK(clk), .RST(rst), .I(m[489]), 
        .Q(c[489]) );
  DFF \creg_reg[490]  ( .D(creg_next[490]), .CLK(clk), .RST(rst), .I(m[490]), 
        .Q(c[490]) );
  DFF \creg_reg[491]  ( .D(creg_next[491]), .CLK(clk), .RST(rst), .I(m[491]), 
        .Q(c[491]) );
  DFF \creg_reg[492]  ( .D(creg_next[492]), .CLK(clk), .RST(rst), .I(m[492]), 
        .Q(c[492]) );
  DFF \creg_reg[493]  ( .D(creg_next[493]), .CLK(clk), .RST(rst), .I(m[493]), 
        .Q(c[493]) );
  DFF \creg_reg[494]  ( .D(creg_next[494]), .CLK(clk), .RST(rst), .I(m[494]), 
        .Q(c[494]) );
  DFF \creg_reg[495]  ( .D(creg_next[495]), .CLK(clk), .RST(rst), .I(m[495]), 
        .Q(c[495]) );
  DFF \creg_reg[496]  ( .D(creg_next[496]), .CLK(clk), .RST(rst), .I(m[496]), 
        .Q(c[496]) );
  DFF \creg_reg[497]  ( .D(creg_next[497]), .CLK(clk), .RST(rst), .I(m[497]), 
        .Q(c[497]) );
  DFF \creg_reg[498]  ( .D(creg_next[498]), .CLK(clk), .RST(rst), .I(m[498]), 
        .Q(c[498]) );
  DFF \creg_reg[499]  ( .D(creg_next[499]), .CLK(clk), .RST(rst), .I(m[499]), 
        .Q(c[499]) );
  DFF \creg_reg[500]  ( .D(creg_next[500]), .CLK(clk), .RST(rst), .I(m[500]), 
        .Q(c[500]) );
  DFF \creg_reg[501]  ( .D(creg_next[501]), .CLK(clk), .RST(rst), .I(m[501]), 
        .Q(c[501]) );
  DFF \creg_reg[502]  ( .D(creg_next[502]), .CLK(clk), .RST(rst), .I(m[502]), 
        .Q(c[502]) );
  DFF \creg_reg[503]  ( .D(creg_next[503]), .CLK(clk), .RST(rst), .I(m[503]), 
        .Q(c[503]) );
  DFF \creg_reg[504]  ( .D(creg_next[504]), .CLK(clk), .RST(rst), .I(m[504]), 
        .Q(c[504]) );
  DFF \creg_reg[505]  ( .D(creg_next[505]), .CLK(clk), .RST(rst), .I(m[505]), 
        .Q(c[505]) );
  DFF \creg_reg[506]  ( .D(creg_next[506]), .CLK(clk), .RST(rst), .I(m[506]), 
        .Q(c[506]) );
  DFF \creg_reg[507]  ( .D(creg_next[507]), .CLK(clk), .RST(rst), .I(m[507]), 
        .Q(c[507]) );
  DFF \creg_reg[508]  ( .D(creg_next[508]), .CLK(clk), .RST(rst), .I(m[508]), 
        .Q(c[508]) );
  DFF \creg_reg[509]  ( .D(creg_next[509]), .CLK(clk), .RST(rst), .I(m[509]), 
        .Q(c[509]) );
  DFF \creg_reg[510]  ( .D(creg_next[510]), .CLK(clk), .RST(rst), .I(m[510]), 
        .Q(c[510]) );
  DFF \creg_reg[511]  ( .D(creg_next[511]), .CLK(clk), .RST(rst), .I(m[511]), 
        .Q(c[511]) );
  DFF \creg_reg[512]  ( .D(creg_next[512]), .CLK(clk), .RST(rst), .I(m[512]), 
        .Q(c[512]) );
  DFF \creg_reg[513]  ( .D(creg_next[513]), .CLK(clk), .RST(rst), .I(m[513]), 
        .Q(c[513]) );
  DFF \creg_reg[514]  ( .D(creg_next[514]), .CLK(clk), .RST(rst), .I(m[514]), 
        .Q(c[514]) );
  DFF \creg_reg[515]  ( .D(creg_next[515]), .CLK(clk), .RST(rst), .I(m[515]), 
        .Q(c[515]) );
  DFF \creg_reg[516]  ( .D(creg_next[516]), .CLK(clk), .RST(rst), .I(m[516]), 
        .Q(c[516]) );
  DFF \creg_reg[517]  ( .D(creg_next[517]), .CLK(clk), .RST(rst), .I(m[517]), 
        .Q(c[517]) );
  DFF \creg_reg[518]  ( .D(creg_next[518]), .CLK(clk), .RST(rst), .I(m[518]), 
        .Q(c[518]) );
  DFF \creg_reg[519]  ( .D(creg_next[519]), .CLK(clk), .RST(rst), .I(m[519]), 
        .Q(c[519]) );
  DFF \creg_reg[520]  ( .D(creg_next[520]), .CLK(clk), .RST(rst), .I(m[520]), 
        .Q(c[520]) );
  DFF \creg_reg[521]  ( .D(creg_next[521]), .CLK(clk), .RST(rst), .I(m[521]), 
        .Q(c[521]) );
  DFF \creg_reg[522]  ( .D(creg_next[522]), .CLK(clk), .RST(rst), .I(m[522]), 
        .Q(c[522]) );
  DFF \creg_reg[523]  ( .D(creg_next[523]), .CLK(clk), .RST(rst), .I(m[523]), 
        .Q(c[523]) );
  DFF \creg_reg[524]  ( .D(creg_next[524]), .CLK(clk), .RST(rst), .I(m[524]), 
        .Q(c[524]) );
  DFF \creg_reg[525]  ( .D(creg_next[525]), .CLK(clk), .RST(rst), .I(m[525]), 
        .Q(c[525]) );
  DFF \creg_reg[526]  ( .D(creg_next[526]), .CLK(clk), .RST(rst), .I(m[526]), 
        .Q(c[526]) );
  DFF \creg_reg[527]  ( .D(creg_next[527]), .CLK(clk), .RST(rst), .I(m[527]), 
        .Q(c[527]) );
  DFF \creg_reg[528]  ( .D(creg_next[528]), .CLK(clk), .RST(rst), .I(m[528]), 
        .Q(c[528]) );
  DFF \creg_reg[529]  ( .D(creg_next[529]), .CLK(clk), .RST(rst), .I(m[529]), 
        .Q(c[529]) );
  DFF \creg_reg[530]  ( .D(creg_next[530]), .CLK(clk), .RST(rst), .I(m[530]), 
        .Q(c[530]) );
  DFF \creg_reg[531]  ( .D(creg_next[531]), .CLK(clk), .RST(rst), .I(m[531]), 
        .Q(c[531]) );
  DFF \creg_reg[532]  ( .D(creg_next[532]), .CLK(clk), .RST(rst), .I(m[532]), 
        .Q(c[532]) );
  DFF \creg_reg[533]  ( .D(creg_next[533]), .CLK(clk), .RST(rst), .I(m[533]), 
        .Q(c[533]) );
  DFF \creg_reg[534]  ( .D(creg_next[534]), .CLK(clk), .RST(rst), .I(m[534]), 
        .Q(c[534]) );
  DFF \creg_reg[535]  ( .D(creg_next[535]), .CLK(clk), .RST(rst), .I(m[535]), 
        .Q(c[535]) );
  DFF \creg_reg[536]  ( .D(creg_next[536]), .CLK(clk), .RST(rst), .I(m[536]), 
        .Q(c[536]) );
  DFF \creg_reg[537]  ( .D(creg_next[537]), .CLK(clk), .RST(rst), .I(m[537]), 
        .Q(c[537]) );
  DFF \creg_reg[538]  ( .D(creg_next[538]), .CLK(clk), .RST(rst), .I(m[538]), 
        .Q(c[538]) );
  DFF \creg_reg[539]  ( .D(creg_next[539]), .CLK(clk), .RST(rst), .I(m[539]), 
        .Q(c[539]) );
  DFF \creg_reg[540]  ( .D(creg_next[540]), .CLK(clk), .RST(rst), .I(m[540]), 
        .Q(c[540]) );
  DFF \creg_reg[541]  ( .D(creg_next[541]), .CLK(clk), .RST(rst), .I(m[541]), 
        .Q(c[541]) );
  DFF \creg_reg[542]  ( .D(creg_next[542]), .CLK(clk), .RST(rst), .I(m[542]), 
        .Q(c[542]) );
  DFF \creg_reg[543]  ( .D(creg_next[543]), .CLK(clk), .RST(rst), .I(m[543]), 
        .Q(c[543]) );
  DFF \creg_reg[544]  ( .D(creg_next[544]), .CLK(clk), .RST(rst), .I(m[544]), 
        .Q(c[544]) );
  DFF \creg_reg[545]  ( .D(creg_next[545]), .CLK(clk), .RST(rst), .I(m[545]), 
        .Q(c[545]) );
  DFF \creg_reg[546]  ( .D(creg_next[546]), .CLK(clk), .RST(rst), .I(m[546]), 
        .Q(c[546]) );
  DFF \creg_reg[547]  ( .D(creg_next[547]), .CLK(clk), .RST(rst), .I(m[547]), 
        .Q(c[547]) );
  DFF \creg_reg[548]  ( .D(creg_next[548]), .CLK(clk), .RST(rst), .I(m[548]), 
        .Q(c[548]) );
  DFF \creg_reg[549]  ( .D(creg_next[549]), .CLK(clk), .RST(rst), .I(m[549]), 
        .Q(c[549]) );
  DFF \creg_reg[550]  ( .D(creg_next[550]), .CLK(clk), .RST(rst), .I(m[550]), 
        .Q(c[550]) );
  DFF \creg_reg[551]  ( .D(creg_next[551]), .CLK(clk), .RST(rst), .I(m[551]), 
        .Q(c[551]) );
  DFF \creg_reg[552]  ( .D(creg_next[552]), .CLK(clk), .RST(rst), .I(m[552]), 
        .Q(c[552]) );
  DFF \creg_reg[553]  ( .D(creg_next[553]), .CLK(clk), .RST(rst), .I(m[553]), 
        .Q(c[553]) );
  DFF \creg_reg[554]  ( .D(creg_next[554]), .CLK(clk), .RST(rst), .I(m[554]), 
        .Q(c[554]) );
  DFF \creg_reg[555]  ( .D(creg_next[555]), .CLK(clk), .RST(rst), .I(m[555]), 
        .Q(c[555]) );
  DFF \creg_reg[556]  ( .D(creg_next[556]), .CLK(clk), .RST(rst), .I(m[556]), 
        .Q(c[556]) );
  DFF \creg_reg[557]  ( .D(creg_next[557]), .CLK(clk), .RST(rst), .I(m[557]), 
        .Q(c[557]) );
  DFF \creg_reg[558]  ( .D(creg_next[558]), .CLK(clk), .RST(rst), .I(m[558]), 
        .Q(c[558]) );
  DFF \creg_reg[559]  ( .D(creg_next[559]), .CLK(clk), .RST(rst), .I(m[559]), 
        .Q(c[559]) );
  DFF \creg_reg[560]  ( .D(creg_next[560]), .CLK(clk), .RST(rst), .I(m[560]), 
        .Q(c[560]) );
  DFF \creg_reg[561]  ( .D(creg_next[561]), .CLK(clk), .RST(rst), .I(m[561]), 
        .Q(c[561]) );
  DFF \creg_reg[562]  ( .D(creg_next[562]), .CLK(clk), .RST(rst), .I(m[562]), 
        .Q(c[562]) );
  DFF \creg_reg[563]  ( .D(creg_next[563]), .CLK(clk), .RST(rst), .I(m[563]), 
        .Q(c[563]) );
  DFF \creg_reg[564]  ( .D(creg_next[564]), .CLK(clk), .RST(rst), .I(m[564]), 
        .Q(c[564]) );
  DFF \creg_reg[565]  ( .D(creg_next[565]), .CLK(clk), .RST(rst), .I(m[565]), 
        .Q(c[565]) );
  DFF \creg_reg[566]  ( .D(creg_next[566]), .CLK(clk), .RST(rst), .I(m[566]), 
        .Q(c[566]) );
  DFF \creg_reg[567]  ( .D(creg_next[567]), .CLK(clk), .RST(rst), .I(m[567]), 
        .Q(c[567]) );
  DFF \creg_reg[568]  ( .D(creg_next[568]), .CLK(clk), .RST(rst), .I(m[568]), 
        .Q(c[568]) );
  DFF \creg_reg[569]  ( .D(creg_next[569]), .CLK(clk), .RST(rst), .I(m[569]), 
        .Q(c[569]) );
  DFF \creg_reg[570]  ( .D(creg_next[570]), .CLK(clk), .RST(rst), .I(m[570]), 
        .Q(c[570]) );
  DFF \creg_reg[571]  ( .D(creg_next[571]), .CLK(clk), .RST(rst), .I(m[571]), 
        .Q(c[571]) );
  DFF \creg_reg[572]  ( .D(creg_next[572]), .CLK(clk), .RST(rst), .I(m[572]), 
        .Q(c[572]) );
  DFF \creg_reg[573]  ( .D(creg_next[573]), .CLK(clk), .RST(rst), .I(m[573]), 
        .Q(c[573]) );
  DFF \creg_reg[574]  ( .D(creg_next[574]), .CLK(clk), .RST(rst), .I(m[574]), 
        .Q(c[574]) );
  DFF \creg_reg[575]  ( .D(creg_next[575]), .CLK(clk), .RST(rst), .I(m[575]), 
        .Q(c[575]) );
  DFF \creg_reg[576]  ( .D(creg_next[576]), .CLK(clk), .RST(rst), .I(m[576]), 
        .Q(c[576]) );
  DFF \creg_reg[577]  ( .D(creg_next[577]), .CLK(clk), .RST(rst), .I(m[577]), 
        .Q(c[577]) );
  DFF \creg_reg[578]  ( .D(creg_next[578]), .CLK(clk), .RST(rst), .I(m[578]), 
        .Q(c[578]) );
  DFF \creg_reg[579]  ( .D(creg_next[579]), .CLK(clk), .RST(rst), .I(m[579]), 
        .Q(c[579]) );
  DFF \creg_reg[580]  ( .D(creg_next[580]), .CLK(clk), .RST(rst), .I(m[580]), 
        .Q(c[580]) );
  DFF \creg_reg[581]  ( .D(creg_next[581]), .CLK(clk), .RST(rst), .I(m[581]), 
        .Q(c[581]) );
  DFF \creg_reg[582]  ( .D(creg_next[582]), .CLK(clk), .RST(rst), .I(m[582]), 
        .Q(c[582]) );
  DFF \creg_reg[583]  ( .D(creg_next[583]), .CLK(clk), .RST(rst), .I(m[583]), 
        .Q(c[583]) );
  DFF \creg_reg[584]  ( .D(creg_next[584]), .CLK(clk), .RST(rst), .I(m[584]), 
        .Q(c[584]) );
  DFF \creg_reg[585]  ( .D(creg_next[585]), .CLK(clk), .RST(rst), .I(m[585]), 
        .Q(c[585]) );
  DFF \creg_reg[586]  ( .D(creg_next[586]), .CLK(clk), .RST(rst), .I(m[586]), 
        .Q(c[586]) );
  DFF \creg_reg[587]  ( .D(creg_next[587]), .CLK(clk), .RST(rst), .I(m[587]), 
        .Q(c[587]) );
  DFF \creg_reg[588]  ( .D(creg_next[588]), .CLK(clk), .RST(rst), .I(m[588]), 
        .Q(c[588]) );
  DFF \creg_reg[589]  ( .D(creg_next[589]), .CLK(clk), .RST(rst), .I(m[589]), 
        .Q(c[589]) );
  DFF \creg_reg[590]  ( .D(creg_next[590]), .CLK(clk), .RST(rst), .I(m[590]), 
        .Q(c[590]) );
  DFF \creg_reg[591]  ( .D(creg_next[591]), .CLK(clk), .RST(rst), .I(m[591]), 
        .Q(c[591]) );
  DFF \creg_reg[592]  ( .D(creg_next[592]), .CLK(clk), .RST(rst), .I(m[592]), 
        .Q(c[592]) );
  DFF \creg_reg[593]  ( .D(creg_next[593]), .CLK(clk), .RST(rst), .I(m[593]), 
        .Q(c[593]) );
  DFF \creg_reg[594]  ( .D(creg_next[594]), .CLK(clk), .RST(rst), .I(m[594]), 
        .Q(c[594]) );
  DFF \creg_reg[595]  ( .D(creg_next[595]), .CLK(clk), .RST(rst), .I(m[595]), 
        .Q(c[595]) );
  DFF \creg_reg[596]  ( .D(creg_next[596]), .CLK(clk), .RST(rst), .I(m[596]), 
        .Q(c[596]) );
  DFF \creg_reg[597]  ( .D(creg_next[597]), .CLK(clk), .RST(rst), .I(m[597]), 
        .Q(c[597]) );
  DFF \creg_reg[598]  ( .D(creg_next[598]), .CLK(clk), .RST(rst), .I(m[598]), 
        .Q(c[598]) );
  DFF \creg_reg[599]  ( .D(creg_next[599]), .CLK(clk), .RST(rst), .I(m[599]), 
        .Q(c[599]) );
  DFF \creg_reg[600]  ( .D(creg_next[600]), .CLK(clk), .RST(rst), .I(m[600]), 
        .Q(c[600]) );
  DFF \creg_reg[601]  ( .D(creg_next[601]), .CLK(clk), .RST(rst), .I(m[601]), 
        .Q(c[601]) );
  DFF \creg_reg[602]  ( .D(creg_next[602]), .CLK(clk), .RST(rst), .I(m[602]), 
        .Q(c[602]) );
  DFF \creg_reg[603]  ( .D(creg_next[603]), .CLK(clk), .RST(rst), .I(m[603]), 
        .Q(c[603]) );
  DFF \creg_reg[604]  ( .D(creg_next[604]), .CLK(clk), .RST(rst), .I(m[604]), 
        .Q(c[604]) );
  DFF \creg_reg[605]  ( .D(creg_next[605]), .CLK(clk), .RST(rst), .I(m[605]), 
        .Q(c[605]) );
  DFF \creg_reg[606]  ( .D(creg_next[606]), .CLK(clk), .RST(rst), .I(m[606]), 
        .Q(c[606]) );
  DFF \creg_reg[607]  ( .D(creg_next[607]), .CLK(clk), .RST(rst), .I(m[607]), 
        .Q(c[607]) );
  DFF \creg_reg[608]  ( .D(creg_next[608]), .CLK(clk), .RST(rst), .I(m[608]), 
        .Q(c[608]) );
  DFF \creg_reg[609]  ( .D(creg_next[609]), .CLK(clk), .RST(rst), .I(m[609]), 
        .Q(c[609]) );
  DFF \creg_reg[610]  ( .D(creg_next[610]), .CLK(clk), .RST(rst), .I(m[610]), 
        .Q(c[610]) );
  DFF \creg_reg[611]  ( .D(creg_next[611]), .CLK(clk), .RST(rst), .I(m[611]), 
        .Q(c[611]) );
  DFF \creg_reg[612]  ( .D(creg_next[612]), .CLK(clk), .RST(rst), .I(m[612]), 
        .Q(c[612]) );
  DFF \creg_reg[613]  ( .D(creg_next[613]), .CLK(clk), .RST(rst), .I(m[613]), 
        .Q(c[613]) );
  DFF \creg_reg[614]  ( .D(creg_next[614]), .CLK(clk), .RST(rst), .I(m[614]), 
        .Q(c[614]) );
  DFF \creg_reg[615]  ( .D(creg_next[615]), .CLK(clk), .RST(rst), .I(m[615]), 
        .Q(c[615]) );
  DFF \creg_reg[616]  ( .D(creg_next[616]), .CLK(clk), .RST(rst), .I(m[616]), 
        .Q(c[616]) );
  DFF \creg_reg[617]  ( .D(creg_next[617]), .CLK(clk), .RST(rst), .I(m[617]), 
        .Q(c[617]) );
  DFF \creg_reg[618]  ( .D(creg_next[618]), .CLK(clk), .RST(rst), .I(m[618]), 
        .Q(c[618]) );
  DFF \creg_reg[619]  ( .D(creg_next[619]), .CLK(clk), .RST(rst), .I(m[619]), 
        .Q(c[619]) );
  DFF \creg_reg[620]  ( .D(creg_next[620]), .CLK(clk), .RST(rst), .I(m[620]), 
        .Q(c[620]) );
  DFF \creg_reg[621]  ( .D(creg_next[621]), .CLK(clk), .RST(rst), .I(m[621]), 
        .Q(c[621]) );
  DFF \creg_reg[622]  ( .D(creg_next[622]), .CLK(clk), .RST(rst), .I(m[622]), 
        .Q(c[622]) );
  DFF \creg_reg[623]  ( .D(creg_next[623]), .CLK(clk), .RST(rst), .I(m[623]), 
        .Q(c[623]) );
  DFF \creg_reg[624]  ( .D(creg_next[624]), .CLK(clk), .RST(rst), .I(m[624]), 
        .Q(c[624]) );
  DFF \creg_reg[625]  ( .D(creg_next[625]), .CLK(clk), .RST(rst), .I(m[625]), 
        .Q(c[625]) );
  DFF \creg_reg[626]  ( .D(creg_next[626]), .CLK(clk), .RST(rst), .I(m[626]), 
        .Q(c[626]) );
  DFF \creg_reg[627]  ( .D(creg_next[627]), .CLK(clk), .RST(rst), .I(m[627]), 
        .Q(c[627]) );
  DFF \creg_reg[628]  ( .D(creg_next[628]), .CLK(clk), .RST(rst), .I(m[628]), 
        .Q(c[628]) );
  DFF \creg_reg[629]  ( .D(creg_next[629]), .CLK(clk), .RST(rst), .I(m[629]), 
        .Q(c[629]) );
  DFF \creg_reg[630]  ( .D(creg_next[630]), .CLK(clk), .RST(rst), .I(m[630]), 
        .Q(c[630]) );
  DFF \creg_reg[631]  ( .D(creg_next[631]), .CLK(clk), .RST(rst), .I(m[631]), 
        .Q(c[631]) );
  DFF \creg_reg[632]  ( .D(creg_next[632]), .CLK(clk), .RST(rst), .I(m[632]), 
        .Q(c[632]) );
  DFF \creg_reg[633]  ( .D(creg_next[633]), .CLK(clk), .RST(rst), .I(m[633]), 
        .Q(c[633]) );
  DFF \creg_reg[634]  ( .D(creg_next[634]), .CLK(clk), .RST(rst), .I(m[634]), 
        .Q(c[634]) );
  DFF \creg_reg[635]  ( .D(creg_next[635]), .CLK(clk), .RST(rst), .I(m[635]), 
        .Q(c[635]) );
  DFF \creg_reg[636]  ( .D(creg_next[636]), .CLK(clk), .RST(rst), .I(m[636]), 
        .Q(c[636]) );
  DFF \creg_reg[637]  ( .D(creg_next[637]), .CLK(clk), .RST(rst), .I(m[637]), 
        .Q(c[637]) );
  DFF \creg_reg[638]  ( .D(creg_next[638]), .CLK(clk), .RST(rst), .I(m[638]), 
        .Q(c[638]) );
  DFF \creg_reg[639]  ( .D(creg_next[639]), .CLK(clk), .RST(rst), .I(m[639]), 
        .Q(c[639]) );
  DFF \creg_reg[640]  ( .D(creg_next[640]), .CLK(clk), .RST(rst), .I(m[640]), 
        .Q(c[640]) );
  DFF \creg_reg[641]  ( .D(creg_next[641]), .CLK(clk), .RST(rst), .I(m[641]), 
        .Q(c[641]) );
  DFF \creg_reg[642]  ( .D(creg_next[642]), .CLK(clk), .RST(rst), .I(m[642]), 
        .Q(c[642]) );
  DFF \creg_reg[643]  ( .D(creg_next[643]), .CLK(clk), .RST(rst), .I(m[643]), 
        .Q(c[643]) );
  DFF \creg_reg[644]  ( .D(creg_next[644]), .CLK(clk), .RST(rst), .I(m[644]), 
        .Q(c[644]) );
  DFF \creg_reg[645]  ( .D(creg_next[645]), .CLK(clk), .RST(rst), .I(m[645]), 
        .Q(c[645]) );
  DFF \creg_reg[646]  ( .D(creg_next[646]), .CLK(clk), .RST(rst), .I(m[646]), 
        .Q(c[646]) );
  DFF \creg_reg[647]  ( .D(creg_next[647]), .CLK(clk), .RST(rst), .I(m[647]), 
        .Q(c[647]) );
  DFF \creg_reg[648]  ( .D(creg_next[648]), .CLK(clk), .RST(rst), .I(m[648]), 
        .Q(c[648]) );
  DFF \creg_reg[649]  ( .D(creg_next[649]), .CLK(clk), .RST(rst), .I(m[649]), 
        .Q(c[649]) );
  DFF \creg_reg[650]  ( .D(creg_next[650]), .CLK(clk), .RST(rst), .I(m[650]), 
        .Q(c[650]) );
  DFF \creg_reg[651]  ( .D(creg_next[651]), .CLK(clk), .RST(rst), .I(m[651]), 
        .Q(c[651]) );
  DFF \creg_reg[652]  ( .D(creg_next[652]), .CLK(clk), .RST(rst), .I(m[652]), 
        .Q(c[652]) );
  DFF \creg_reg[653]  ( .D(creg_next[653]), .CLK(clk), .RST(rst), .I(m[653]), 
        .Q(c[653]) );
  DFF \creg_reg[654]  ( .D(creg_next[654]), .CLK(clk), .RST(rst), .I(m[654]), 
        .Q(c[654]) );
  DFF \creg_reg[655]  ( .D(creg_next[655]), .CLK(clk), .RST(rst), .I(m[655]), 
        .Q(c[655]) );
  DFF \creg_reg[656]  ( .D(creg_next[656]), .CLK(clk), .RST(rst), .I(m[656]), 
        .Q(c[656]) );
  DFF \creg_reg[657]  ( .D(creg_next[657]), .CLK(clk), .RST(rst), .I(m[657]), 
        .Q(c[657]) );
  DFF \creg_reg[658]  ( .D(creg_next[658]), .CLK(clk), .RST(rst), .I(m[658]), 
        .Q(c[658]) );
  DFF \creg_reg[659]  ( .D(creg_next[659]), .CLK(clk), .RST(rst), .I(m[659]), 
        .Q(c[659]) );
  DFF \creg_reg[660]  ( .D(creg_next[660]), .CLK(clk), .RST(rst), .I(m[660]), 
        .Q(c[660]) );
  DFF \creg_reg[661]  ( .D(creg_next[661]), .CLK(clk), .RST(rst), .I(m[661]), 
        .Q(c[661]) );
  DFF \creg_reg[662]  ( .D(creg_next[662]), .CLK(clk), .RST(rst), .I(m[662]), 
        .Q(c[662]) );
  DFF \creg_reg[663]  ( .D(creg_next[663]), .CLK(clk), .RST(rst), .I(m[663]), 
        .Q(c[663]) );
  DFF \creg_reg[664]  ( .D(creg_next[664]), .CLK(clk), .RST(rst), .I(m[664]), 
        .Q(c[664]) );
  DFF \creg_reg[665]  ( .D(creg_next[665]), .CLK(clk), .RST(rst), .I(m[665]), 
        .Q(c[665]) );
  DFF \creg_reg[666]  ( .D(creg_next[666]), .CLK(clk), .RST(rst), .I(m[666]), 
        .Q(c[666]) );
  DFF \creg_reg[667]  ( .D(creg_next[667]), .CLK(clk), .RST(rst), .I(m[667]), 
        .Q(c[667]) );
  DFF \creg_reg[668]  ( .D(creg_next[668]), .CLK(clk), .RST(rst), .I(m[668]), 
        .Q(c[668]) );
  DFF \creg_reg[669]  ( .D(creg_next[669]), .CLK(clk), .RST(rst), .I(m[669]), 
        .Q(c[669]) );
  DFF \creg_reg[670]  ( .D(creg_next[670]), .CLK(clk), .RST(rst), .I(m[670]), 
        .Q(c[670]) );
  DFF \creg_reg[671]  ( .D(creg_next[671]), .CLK(clk), .RST(rst), .I(m[671]), 
        .Q(c[671]) );
  DFF \creg_reg[672]  ( .D(creg_next[672]), .CLK(clk), .RST(rst), .I(m[672]), 
        .Q(c[672]) );
  DFF \creg_reg[673]  ( .D(creg_next[673]), .CLK(clk), .RST(rst), .I(m[673]), 
        .Q(c[673]) );
  DFF \creg_reg[674]  ( .D(creg_next[674]), .CLK(clk), .RST(rst), .I(m[674]), 
        .Q(c[674]) );
  DFF \creg_reg[675]  ( .D(creg_next[675]), .CLK(clk), .RST(rst), .I(m[675]), 
        .Q(c[675]) );
  DFF \creg_reg[676]  ( .D(creg_next[676]), .CLK(clk), .RST(rst), .I(m[676]), 
        .Q(c[676]) );
  DFF \creg_reg[677]  ( .D(creg_next[677]), .CLK(clk), .RST(rst), .I(m[677]), 
        .Q(c[677]) );
  DFF \creg_reg[678]  ( .D(creg_next[678]), .CLK(clk), .RST(rst), .I(m[678]), 
        .Q(c[678]) );
  DFF \creg_reg[679]  ( .D(creg_next[679]), .CLK(clk), .RST(rst), .I(m[679]), 
        .Q(c[679]) );
  DFF \creg_reg[680]  ( .D(creg_next[680]), .CLK(clk), .RST(rst), .I(m[680]), 
        .Q(c[680]) );
  DFF \creg_reg[681]  ( .D(creg_next[681]), .CLK(clk), .RST(rst), .I(m[681]), 
        .Q(c[681]) );
  DFF \creg_reg[682]  ( .D(creg_next[682]), .CLK(clk), .RST(rst), .I(m[682]), 
        .Q(c[682]) );
  DFF \creg_reg[683]  ( .D(creg_next[683]), .CLK(clk), .RST(rst), .I(m[683]), 
        .Q(c[683]) );
  DFF \creg_reg[684]  ( .D(creg_next[684]), .CLK(clk), .RST(rst), .I(m[684]), 
        .Q(c[684]) );
  DFF \creg_reg[685]  ( .D(creg_next[685]), .CLK(clk), .RST(rst), .I(m[685]), 
        .Q(c[685]) );
  DFF \creg_reg[686]  ( .D(creg_next[686]), .CLK(clk), .RST(rst), .I(m[686]), 
        .Q(c[686]) );
  DFF \creg_reg[687]  ( .D(creg_next[687]), .CLK(clk), .RST(rst), .I(m[687]), 
        .Q(c[687]) );
  DFF \creg_reg[688]  ( .D(creg_next[688]), .CLK(clk), .RST(rst), .I(m[688]), 
        .Q(c[688]) );
  DFF \creg_reg[689]  ( .D(creg_next[689]), .CLK(clk), .RST(rst), .I(m[689]), 
        .Q(c[689]) );
  DFF \creg_reg[690]  ( .D(creg_next[690]), .CLK(clk), .RST(rst), .I(m[690]), 
        .Q(c[690]) );
  DFF \creg_reg[691]  ( .D(creg_next[691]), .CLK(clk), .RST(rst), .I(m[691]), 
        .Q(c[691]) );
  DFF \creg_reg[692]  ( .D(creg_next[692]), .CLK(clk), .RST(rst), .I(m[692]), 
        .Q(c[692]) );
  DFF \creg_reg[693]  ( .D(creg_next[693]), .CLK(clk), .RST(rst), .I(m[693]), 
        .Q(c[693]) );
  DFF \creg_reg[694]  ( .D(creg_next[694]), .CLK(clk), .RST(rst), .I(m[694]), 
        .Q(c[694]) );
  DFF \creg_reg[695]  ( .D(creg_next[695]), .CLK(clk), .RST(rst), .I(m[695]), 
        .Q(c[695]) );
  DFF \creg_reg[696]  ( .D(creg_next[696]), .CLK(clk), .RST(rst), .I(m[696]), 
        .Q(c[696]) );
  DFF \creg_reg[697]  ( .D(creg_next[697]), .CLK(clk), .RST(rst), .I(m[697]), 
        .Q(c[697]) );
  DFF \creg_reg[698]  ( .D(creg_next[698]), .CLK(clk), .RST(rst), .I(m[698]), 
        .Q(c[698]) );
  DFF \creg_reg[699]  ( .D(creg_next[699]), .CLK(clk), .RST(rst), .I(m[699]), 
        .Q(c[699]) );
  DFF \creg_reg[700]  ( .D(creg_next[700]), .CLK(clk), .RST(rst), .I(m[700]), 
        .Q(c[700]) );
  DFF \creg_reg[701]  ( .D(creg_next[701]), .CLK(clk), .RST(rst), .I(m[701]), 
        .Q(c[701]) );
  DFF \creg_reg[702]  ( .D(creg_next[702]), .CLK(clk), .RST(rst), .I(m[702]), 
        .Q(c[702]) );
  DFF \creg_reg[703]  ( .D(creg_next[703]), .CLK(clk), .RST(rst), .I(m[703]), 
        .Q(c[703]) );
  DFF \creg_reg[704]  ( .D(creg_next[704]), .CLK(clk), .RST(rst), .I(m[704]), 
        .Q(c[704]) );
  DFF \creg_reg[705]  ( .D(creg_next[705]), .CLK(clk), .RST(rst), .I(m[705]), 
        .Q(c[705]) );
  DFF \creg_reg[706]  ( .D(creg_next[706]), .CLK(clk), .RST(rst), .I(m[706]), 
        .Q(c[706]) );
  DFF \creg_reg[707]  ( .D(creg_next[707]), .CLK(clk), .RST(rst), .I(m[707]), 
        .Q(c[707]) );
  DFF \creg_reg[708]  ( .D(creg_next[708]), .CLK(clk), .RST(rst), .I(m[708]), 
        .Q(c[708]) );
  DFF \creg_reg[709]  ( .D(creg_next[709]), .CLK(clk), .RST(rst), .I(m[709]), 
        .Q(c[709]) );
  DFF \creg_reg[710]  ( .D(creg_next[710]), .CLK(clk), .RST(rst), .I(m[710]), 
        .Q(c[710]) );
  DFF \creg_reg[711]  ( .D(creg_next[711]), .CLK(clk), .RST(rst), .I(m[711]), 
        .Q(c[711]) );
  DFF \creg_reg[712]  ( .D(creg_next[712]), .CLK(clk), .RST(rst), .I(m[712]), 
        .Q(c[712]) );
  DFF \creg_reg[713]  ( .D(creg_next[713]), .CLK(clk), .RST(rst), .I(m[713]), 
        .Q(c[713]) );
  DFF \creg_reg[714]  ( .D(creg_next[714]), .CLK(clk), .RST(rst), .I(m[714]), 
        .Q(c[714]) );
  DFF \creg_reg[715]  ( .D(creg_next[715]), .CLK(clk), .RST(rst), .I(m[715]), 
        .Q(c[715]) );
  DFF \creg_reg[716]  ( .D(creg_next[716]), .CLK(clk), .RST(rst), .I(m[716]), 
        .Q(c[716]) );
  DFF \creg_reg[717]  ( .D(creg_next[717]), .CLK(clk), .RST(rst), .I(m[717]), 
        .Q(c[717]) );
  DFF \creg_reg[718]  ( .D(creg_next[718]), .CLK(clk), .RST(rst), .I(m[718]), 
        .Q(c[718]) );
  DFF \creg_reg[719]  ( .D(creg_next[719]), .CLK(clk), .RST(rst), .I(m[719]), 
        .Q(c[719]) );
  DFF \creg_reg[720]  ( .D(creg_next[720]), .CLK(clk), .RST(rst), .I(m[720]), 
        .Q(c[720]) );
  DFF \creg_reg[721]  ( .D(creg_next[721]), .CLK(clk), .RST(rst), .I(m[721]), 
        .Q(c[721]) );
  DFF \creg_reg[722]  ( .D(creg_next[722]), .CLK(clk), .RST(rst), .I(m[722]), 
        .Q(c[722]) );
  DFF \creg_reg[723]  ( .D(creg_next[723]), .CLK(clk), .RST(rst), .I(m[723]), 
        .Q(c[723]) );
  DFF \creg_reg[724]  ( .D(creg_next[724]), .CLK(clk), .RST(rst), .I(m[724]), 
        .Q(c[724]) );
  DFF \creg_reg[725]  ( .D(creg_next[725]), .CLK(clk), .RST(rst), .I(m[725]), 
        .Q(c[725]) );
  DFF \creg_reg[726]  ( .D(creg_next[726]), .CLK(clk), .RST(rst), .I(m[726]), 
        .Q(c[726]) );
  DFF \creg_reg[727]  ( .D(creg_next[727]), .CLK(clk), .RST(rst), .I(m[727]), 
        .Q(c[727]) );
  DFF \creg_reg[728]  ( .D(creg_next[728]), .CLK(clk), .RST(rst), .I(m[728]), 
        .Q(c[728]) );
  DFF \creg_reg[729]  ( .D(creg_next[729]), .CLK(clk), .RST(rst), .I(m[729]), 
        .Q(c[729]) );
  DFF \creg_reg[730]  ( .D(creg_next[730]), .CLK(clk), .RST(rst), .I(m[730]), 
        .Q(c[730]) );
  DFF \creg_reg[731]  ( .D(creg_next[731]), .CLK(clk), .RST(rst), .I(m[731]), 
        .Q(c[731]) );
  DFF \creg_reg[732]  ( .D(creg_next[732]), .CLK(clk), .RST(rst), .I(m[732]), 
        .Q(c[732]) );
  DFF \creg_reg[733]  ( .D(creg_next[733]), .CLK(clk), .RST(rst), .I(m[733]), 
        .Q(c[733]) );
  DFF \creg_reg[734]  ( .D(creg_next[734]), .CLK(clk), .RST(rst), .I(m[734]), 
        .Q(c[734]) );
  DFF \creg_reg[735]  ( .D(creg_next[735]), .CLK(clk), .RST(rst), .I(m[735]), 
        .Q(c[735]) );
  DFF \creg_reg[736]  ( .D(creg_next[736]), .CLK(clk), .RST(rst), .I(m[736]), 
        .Q(c[736]) );
  DFF \creg_reg[737]  ( .D(creg_next[737]), .CLK(clk), .RST(rst), .I(m[737]), 
        .Q(c[737]) );
  DFF \creg_reg[738]  ( .D(creg_next[738]), .CLK(clk), .RST(rst), .I(m[738]), 
        .Q(c[738]) );
  DFF \creg_reg[739]  ( .D(creg_next[739]), .CLK(clk), .RST(rst), .I(m[739]), 
        .Q(c[739]) );
  DFF \creg_reg[740]  ( .D(creg_next[740]), .CLK(clk), .RST(rst), .I(m[740]), 
        .Q(c[740]) );
  DFF \creg_reg[741]  ( .D(creg_next[741]), .CLK(clk), .RST(rst), .I(m[741]), 
        .Q(c[741]) );
  DFF \creg_reg[742]  ( .D(creg_next[742]), .CLK(clk), .RST(rst), .I(m[742]), 
        .Q(c[742]) );
  DFF \creg_reg[743]  ( .D(creg_next[743]), .CLK(clk), .RST(rst), .I(m[743]), 
        .Q(c[743]) );
  DFF \creg_reg[744]  ( .D(creg_next[744]), .CLK(clk), .RST(rst), .I(m[744]), 
        .Q(c[744]) );
  DFF \creg_reg[745]  ( .D(creg_next[745]), .CLK(clk), .RST(rst), .I(m[745]), 
        .Q(c[745]) );
  DFF \creg_reg[746]  ( .D(creg_next[746]), .CLK(clk), .RST(rst), .I(m[746]), 
        .Q(c[746]) );
  DFF \creg_reg[747]  ( .D(creg_next[747]), .CLK(clk), .RST(rst), .I(m[747]), 
        .Q(c[747]) );
  DFF \creg_reg[748]  ( .D(creg_next[748]), .CLK(clk), .RST(rst), .I(m[748]), 
        .Q(c[748]) );
  DFF \creg_reg[749]  ( .D(creg_next[749]), .CLK(clk), .RST(rst), .I(m[749]), 
        .Q(c[749]) );
  DFF \creg_reg[750]  ( .D(creg_next[750]), .CLK(clk), .RST(rst), .I(m[750]), 
        .Q(c[750]) );
  DFF \creg_reg[751]  ( .D(creg_next[751]), .CLK(clk), .RST(rst), .I(m[751]), 
        .Q(c[751]) );
  DFF \creg_reg[752]  ( .D(creg_next[752]), .CLK(clk), .RST(rst), .I(m[752]), 
        .Q(c[752]) );
  DFF \creg_reg[753]  ( .D(creg_next[753]), .CLK(clk), .RST(rst), .I(m[753]), 
        .Q(c[753]) );
  DFF \creg_reg[754]  ( .D(creg_next[754]), .CLK(clk), .RST(rst), .I(m[754]), 
        .Q(c[754]) );
  DFF \creg_reg[755]  ( .D(creg_next[755]), .CLK(clk), .RST(rst), .I(m[755]), 
        .Q(c[755]) );
  DFF \creg_reg[756]  ( .D(creg_next[756]), .CLK(clk), .RST(rst), .I(m[756]), 
        .Q(c[756]) );
  DFF \creg_reg[757]  ( .D(creg_next[757]), .CLK(clk), .RST(rst), .I(m[757]), 
        .Q(c[757]) );
  DFF \creg_reg[758]  ( .D(creg_next[758]), .CLK(clk), .RST(rst), .I(m[758]), 
        .Q(c[758]) );
  DFF \creg_reg[759]  ( .D(creg_next[759]), .CLK(clk), .RST(rst), .I(m[759]), 
        .Q(c[759]) );
  DFF \creg_reg[760]  ( .D(creg_next[760]), .CLK(clk), .RST(rst), .I(m[760]), 
        .Q(c[760]) );
  DFF \creg_reg[761]  ( .D(creg_next[761]), .CLK(clk), .RST(rst), .I(m[761]), 
        .Q(c[761]) );
  DFF \creg_reg[762]  ( .D(creg_next[762]), .CLK(clk), .RST(rst), .I(m[762]), 
        .Q(c[762]) );
  DFF \creg_reg[763]  ( .D(creg_next[763]), .CLK(clk), .RST(rst), .I(m[763]), 
        .Q(c[763]) );
  DFF \creg_reg[764]  ( .D(creg_next[764]), .CLK(clk), .RST(rst), .I(m[764]), 
        .Q(c[764]) );
  DFF \creg_reg[765]  ( .D(creg_next[765]), .CLK(clk), .RST(rst), .I(m[765]), 
        .Q(c[765]) );
  DFF \creg_reg[766]  ( .D(creg_next[766]), .CLK(clk), .RST(rst), .I(m[766]), 
        .Q(c[766]) );
  DFF \creg_reg[767]  ( .D(creg_next[767]), .CLK(clk), .RST(rst), .I(m[767]), 
        .Q(c[767]) );
  DFF \creg_reg[768]  ( .D(creg_next[768]), .CLK(clk), .RST(rst), .I(m[768]), 
        .Q(c[768]) );
  DFF \creg_reg[769]  ( .D(creg_next[769]), .CLK(clk), .RST(rst), .I(m[769]), 
        .Q(c[769]) );
  DFF \creg_reg[770]  ( .D(creg_next[770]), .CLK(clk), .RST(rst), .I(m[770]), 
        .Q(c[770]) );
  DFF \creg_reg[771]  ( .D(creg_next[771]), .CLK(clk), .RST(rst), .I(m[771]), 
        .Q(c[771]) );
  DFF \creg_reg[772]  ( .D(creg_next[772]), .CLK(clk), .RST(rst), .I(m[772]), 
        .Q(c[772]) );
  DFF \creg_reg[773]  ( .D(creg_next[773]), .CLK(clk), .RST(rst), .I(m[773]), 
        .Q(c[773]) );
  DFF \creg_reg[774]  ( .D(creg_next[774]), .CLK(clk), .RST(rst), .I(m[774]), 
        .Q(c[774]) );
  DFF \creg_reg[775]  ( .D(creg_next[775]), .CLK(clk), .RST(rst), .I(m[775]), 
        .Q(c[775]) );
  DFF \creg_reg[776]  ( .D(creg_next[776]), .CLK(clk), .RST(rst), .I(m[776]), 
        .Q(c[776]) );
  DFF \creg_reg[777]  ( .D(creg_next[777]), .CLK(clk), .RST(rst), .I(m[777]), 
        .Q(c[777]) );
  DFF \creg_reg[778]  ( .D(creg_next[778]), .CLK(clk), .RST(rst), .I(m[778]), 
        .Q(c[778]) );
  DFF \creg_reg[779]  ( .D(creg_next[779]), .CLK(clk), .RST(rst), .I(m[779]), 
        .Q(c[779]) );
  DFF \creg_reg[780]  ( .D(creg_next[780]), .CLK(clk), .RST(rst), .I(m[780]), 
        .Q(c[780]) );
  DFF \creg_reg[781]  ( .D(creg_next[781]), .CLK(clk), .RST(rst), .I(m[781]), 
        .Q(c[781]) );
  DFF \creg_reg[782]  ( .D(creg_next[782]), .CLK(clk), .RST(rst), .I(m[782]), 
        .Q(c[782]) );
  DFF \creg_reg[783]  ( .D(creg_next[783]), .CLK(clk), .RST(rst), .I(m[783]), 
        .Q(c[783]) );
  DFF \creg_reg[784]  ( .D(creg_next[784]), .CLK(clk), .RST(rst), .I(m[784]), 
        .Q(c[784]) );
  DFF \creg_reg[785]  ( .D(creg_next[785]), .CLK(clk), .RST(rst), .I(m[785]), 
        .Q(c[785]) );
  DFF \creg_reg[786]  ( .D(creg_next[786]), .CLK(clk), .RST(rst), .I(m[786]), 
        .Q(c[786]) );
  DFF \creg_reg[787]  ( .D(creg_next[787]), .CLK(clk), .RST(rst), .I(m[787]), 
        .Q(c[787]) );
  DFF \creg_reg[788]  ( .D(creg_next[788]), .CLK(clk), .RST(rst), .I(m[788]), 
        .Q(c[788]) );
  DFF \creg_reg[789]  ( .D(creg_next[789]), .CLK(clk), .RST(rst), .I(m[789]), 
        .Q(c[789]) );
  DFF \creg_reg[790]  ( .D(creg_next[790]), .CLK(clk), .RST(rst), .I(m[790]), 
        .Q(c[790]) );
  DFF \creg_reg[791]  ( .D(creg_next[791]), .CLK(clk), .RST(rst), .I(m[791]), 
        .Q(c[791]) );
  DFF \creg_reg[792]  ( .D(creg_next[792]), .CLK(clk), .RST(rst), .I(m[792]), 
        .Q(c[792]) );
  DFF \creg_reg[793]  ( .D(creg_next[793]), .CLK(clk), .RST(rst), .I(m[793]), 
        .Q(c[793]) );
  DFF \creg_reg[794]  ( .D(creg_next[794]), .CLK(clk), .RST(rst), .I(m[794]), 
        .Q(c[794]) );
  DFF \creg_reg[795]  ( .D(creg_next[795]), .CLK(clk), .RST(rst), .I(m[795]), 
        .Q(c[795]) );
  DFF \creg_reg[796]  ( .D(creg_next[796]), .CLK(clk), .RST(rst), .I(m[796]), 
        .Q(c[796]) );
  DFF \creg_reg[797]  ( .D(creg_next[797]), .CLK(clk), .RST(rst), .I(m[797]), 
        .Q(c[797]) );
  DFF \creg_reg[798]  ( .D(creg_next[798]), .CLK(clk), .RST(rst), .I(m[798]), 
        .Q(c[798]) );
  DFF \creg_reg[799]  ( .D(creg_next[799]), .CLK(clk), .RST(rst), .I(m[799]), 
        .Q(c[799]) );
  DFF \creg_reg[800]  ( .D(creg_next[800]), .CLK(clk), .RST(rst), .I(m[800]), 
        .Q(c[800]) );
  DFF \creg_reg[801]  ( .D(creg_next[801]), .CLK(clk), .RST(rst), .I(m[801]), 
        .Q(c[801]) );
  DFF \creg_reg[802]  ( .D(creg_next[802]), .CLK(clk), .RST(rst), .I(m[802]), 
        .Q(c[802]) );
  DFF \creg_reg[803]  ( .D(creg_next[803]), .CLK(clk), .RST(rst), .I(m[803]), 
        .Q(c[803]) );
  DFF \creg_reg[804]  ( .D(creg_next[804]), .CLK(clk), .RST(rst), .I(m[804]), 
        .Q(c[804]) );
  DFF \creg_reg[805]  ( .D(creg_next[805]), .CLK(clk), .RST(rst), .I(m[805]), 
        .Q(c[805]) );
  DFF \creg_reg[806]  ( .D(creg_next[806]), .CLK(clk), .RST(rst), .I(m[806]), 
        .Q(c[806]) );
  DFF \creg_reg[807]  ( .D(creg_next[807]), .CLK(clk), .RST(rst), .I(m[807]), 
        .Q(c[807]) );
  DFF \creg_reg[808]  ( .D(creg_next[808]), .CLK(clk), .RST(rst), .I(m[808]), 
        .Q(c[808]) );
  DFF \creg_reg[809]  ( .D(creg_next[809]), .CLK(clk), .RST(rst), .I(m[809]), 
        .Q(c[809]) );
  DFF \creg_reg[810]  ( .D(creg_next[810]), .CLK(clk), .RST(rst), .I(m[810]), 
        .Q(c[810]) );
  DFF \creg_reg[811]  ( .D(creg_next[811]), .CLK(clk), .RST(rst), .I(m[811]), 
        .Q(c[811]) );
  DFF \creg_reg[812]  ( .D(creg_next[812]), .CLK(clk), .RST(rst), .I(m[812]), 
        .Q(c[812]) );
  DFF \creg_reg[813]  ( .D(creg_next[813]), .CLK(clk), .RST(rst), .I(m[813]), 
        .Q(c[813]) );
  DFF \creg_reg[814]  ( .D(creg_next[814]), .CLK(clk), .RST(rst), .I(m[814]), 
        .Q(c[814]) );
  DFF \creg_reg[815]  ( .D(creg_next[815]), .CLK(clk), .RST(rst), .I(m[815]), 
        .Q(c[815]) );
  DFF \creg_reg[816]  ( .D(creg_next[816]), .CLK(clk), .RST(rst), .I(m[816]), 
        .Q(c[816]) );
  DFF \creg_reg[817]  ( .D(creg_next[817]), .CLK(clk), .RST(rst), .I(m[817]), 
        .Q(c[817]) );
  DFF \creg_reg[818]  ( .D(creg_next[818]), .CLK(clk), .RST(rst), .I(m[818]), 
        .Q(c[818]) );
  DFF \creg_reg[819]  ( .D(creg_next[819]), .CLK(clk), .RST(rst), .I(m[819]), 
        .Q(c[819]) );
  DFF \creg_reg[820]  ( .D(creg_next[820]), .CLK(clk), .RST(rst), .I(m[820]), 
        .Q(c[820]) );
  DFF \creg_reg[821]  ( .D(creg_next[821]), .CLK(clk), .RST(rst), .I(m[821]), 
        .Q(c[821]) );
  DFF \creg_reg[822]  ( .D(creg_next[822]), .CLK(clk), .RST(rst), .I(m[822]), 
        .Q(c[822]) );
  DFF \creg_reg[823]  ( .D(creg_next[823]), .CLK(clk), .RST(rst), .I(m[823]), 
        .Q(c[823]) );
  DFF \creg_reg[824]  ( .D(creg_next[824]), .CLK(clk), .RST(rst), .I(m[824]), 
        .Q(c[824]) );
  DFF \creg_reg[825]  ( .D(creg_next[825]), .CLK(clk), .RST(rst), .I(m[825]), 
        .Q(c[825]) );
  DFF \creg_reg[826]  ( .D(creg_next[826]), .CLK(clk), .RST(rst), .I(m[826]), 
        .Q(c[826]) );
  DFF \creg_reg[827]  ( .D(creg_next[827]), .CLK(clk), .RST(rst), .I(m[827]), 
        .Q(c[827]) );
  DFF \creg_reg[828]  ( .D(creg_next[828]), .CLK(clk), .RST(rst), .I(m[828]), 
        .Q(c[828]) );
  DFF \creg_reg[829]  ( .D(creg_next[829]), .CLK(clk), .RST(rst), .I(m[829]), 
        .Q(c[829]) );
  DFF \creg_reg[830]  ( .D(creg_next[830]), .CLK(clk), .RST(rst), .I(m[830]), 
        .Q(c[830]) );
  DFF \creg_reg[831]  ( .D(creg_next[831]), .CLK(clk), .RST(rst), .I(m[831]), 
        .Q(c[831]) );
  DFF \creg_reg[832]  ( .D(creg_next[832]), .CLK(clk), .RST(rst), .I(m[832]), 
        .Q(c[832]) );
  DFF \creg_reg[833]  ( .D(creg_next[833]), .CLK(clk), .RST(rst), .I(m[833]), 
        .Q(c[833]) );
  DFF \creg_reg[834]  ( .D(creg_next[834]), .CLK(clk), .RST(rst), .I(m[834]), 
        .Q(c[834]) );
  DFF \creg_reg[835]  ( .D(creg_next[835]), .CLK(clk), .RST(rst), .I(m[835]), 
        .Q(c[835]) );
  DFF \creg_reg[836]  ( .D(creg_next[836]), .CLK(clk), .RST(rst), .I(m[836]), 
        .Q(c[836]) );
  DFF \creg_reg[837]  ( .D(creg_next[837]), .CLK(clk), .RST(rst), .I(m[837]), 
        .Q(c[837]) );
  DFF \creg_reg[838]  ( .D(creg_next[838]), .CLK(clk), .RST(rst), .I(m[838]), 
        .Q(c[838]) );
  DFF \creg_reg[839]  ( .D(creg_next[839]), .CLK(clk), .RST(rst), .I(m[839]), 
        .Q(c[839]) );
  DFF \creg_reg[840]  ( .D(creg_next[840]), .CLK(clk), .RST(rst), .I(m[840]), 
        .Q(c[840]) );
  DFF \creg_reg[841]  ( .D(creg_next[841]), .CLK(clk), .RST(rst), .I(m[841]), 
        .Q(c[841]) );
  DFF \creg_reg[842]  ( .D(creg_next[842]), .CLK(clk), .RST(rst), .I(m[842]), 
        .Q(c[842]) );
  DFF \creg_reg[843]  ( .D(creg_next[843]), .CLK(clk), .RST(rst), .I(m[843]), 
        .Q(c[843]) );
  DFF \creg_reg[844]  ( .D(creg_next[844]), .CLK(clk), .RST(rst), .I(m[844]), 
        .Q(c[844]) );
  DFF \creg_reg[845]  ( .D(creg_next[845]), .CLK(clk), .RST(rst), .I(m[845]), 
        .Q(c[845]) );
  DFF \creg_reg[846]  ( .D(creg_next[846]), .CLK(clk), .RST(rst), .I(m[846]), 
        .Q(c[846]) );
  DFF \creg_reg[847]  ( .D(creg_next[847]), .CLK(clk), .RST(rst), .I(m[847]), 
        .Q(c[847]) );
  DFF \creg_reg[848]  ( .D(creg_next[848]), .CLK(clk), .RST(rst), .I(m[848]), 
        .Q(c[848]) );
  DFF \creg_reg[849]  ( .D(creg_next[849]), .CLK(clk), .RST(rst), .I(m[849]), 
        .Q(c[849]) );
  DFF \creg_reg[850]  ( .D(creg_next[850]), .CLK(clk), .RST(rst), .I(m[850]), 
        .Q(c[850]) );
  DFF \creg_reg[851]  ( .D(creg_next[851]), .CLK(clk), .RST(rst), .I(m[851]), 
        .Q(c[851]) );
  DFF \creg_reg[852]  ( .D(creg_next[852]), .CLK(clk), .RST(rst), .I(m[852]), 
        .Q(c[852]) );
  DFF \creg_reg[853]  ( .D(creg_next[853]), .CLK(clk), .RST(rst), .I(m[853]), 
        .Q(c[853]) );
  DFF \creg_reg[854]  ( .D(creg_next[854]), .CLK(clk), .RST(rst), .I(m[854]), 
        .Q(c[854]) );
  DFF \creg_reg[855]  ( .D(creg_next[855]), .CLK(clk), .RST(rst), .I(m[855]), 
        .Q(c[855]) );
  DFF \creg_reg[856]  ( .D(creg_next[856]), .CLK(clk), .RST(rst), .I(m[856]), 
        .Q(c[856]) );
  DFF \creg_reg[857]  ( .D(creg_next[857]), .CLK(clk), .RST(rst), .I(m[857]), 
        .Q(c[857]) );
  DFF \creg_reg[858]  ( .D(creg_next[858]), .CLK(clk), .RST(rst), .I(m[858]), 
        .Q(c[858]) );
  DFF \creg_reg[859]  ( .D(creg_next[859]), .CLK(clk), .RST(rst), .I(m[859]), 
        .Q(c[859]) );
  DFF \creg_reg[860]  ( .D(creg_next[860]), .CLK(clk), .RST(rst), .I(m[860]), 
        .Q(c[860]) );
  DFF \creg_reg[861]  ( .D(creg_next[861]), .CLK(clk), .RST(rst), .I(m[861]), 
        .Q(c[861]) );
  DFF \creg_reg[862]  ( .D(creg_next[862]), .CLK(clk), .RST(rst), .I(m[862]), 
        .Q(c[862]) );
  DFF \creg_reg[863]  ( .D(creg_next[863]), .CLK(clk), .RST(rst), .I(m[863]), 
        .Q(c[863]) );
  DFF \creg_reg[864]  ( .D(creg_next[864]), .CLK(clk), .RST(rst), .I(m[864]), 
        .Q(c[864]) );
  DFF \creg_reg[865]  ( .D(creg_next[865]), .CLK(clk), .RST(rst), .I(m[865]), 
        .Q(c[865]) );
  DFF \creg_reg[866]  ( .D(creg_next[866]), .CLK(clk), .RST(rst), .I(m[866]), 
        .Q(c[866]) );
  DFF \creg_reg[867]  ( .D(creg_next[867]), .CLK(clk), .RST(rst), .I(m[867]), 
        .Q(c[867]) );
  DFF \creg_reg[868]  ( .D(creg_next[868]), .CLK(clk), .RST(rst), .I(m[868]), 
        .Q(c[868]) );
  DFF \creg_reg[869]  ( .D(creg_next[869]), .CLK(clk), .RST(rst), .I(m[869]), 
        .Q(c[869]) );
  DFF \creg_reg[870]  ( .D(creg_next[870]), .CLK(clk), .RST(rst), .I(m[870]), 
        .Q(c[870]) );
  DFF \creg_reg[871]  ( .D(creg_next[871]), .CLK(clk), .RST(rst), .I(m[871]), 
        .Q(c[871]) );
  DFF \creg_reg[872]  ( .D(creg_next[872]), .CLK(clk), .RST(rst), .I(m[872]), 
        .Q(c[872]) );
  DFF \creg_reg[873]  ( .D(creg_next[873]), .CLK(clk), .RST(rst), .I(m[873]), 
        .Q(c[873]) );
  DFF \creg_reg[874]  ( .D(creg_next[874]), .CLK(clk), .RST(rst), .I(m[874]), 
        .Q(c[874]) );
  DFF \creg_reg[875]  ( .D(creg_next[875]), .CLK(clk), .RST(rst), .I(m[875]), 
        .Q(c[875]) );
  DFF \creg_reg[876]  ( .D(creg_next[876]), .CLK(clk), .RST(rst), .I(m[876]), 
        .Q(c[876]) );
  DFF \creg_reg[877]  ( .D(creg_next[877]), .CLK(clk), .RST(rst), .I(m[877]), 
        .Q(c[877]) );
  DFF \creg_reg[878]  ( .D(creg_next[878]), .CLK(clk), .RST(rst), .I(m[878]), 
        .Q(c[878]) );
  DFF \creg_reg[879]  ( .D(creg_next[879]), .CLK(clk), .RST(rst), .I(m[879]), 
        .Q(c[879]) );
  DFF \creg_reg[880]  ( .D(creg_next[880]), .CLK(clk), .RST(rst), .I(m[880]), 
        .Q(c[880]) );
  DFF \creg_reg[881]  ( .D(creg_next[881]), .CLK(clk), .RST(rst), .I(m[881]), 
        .Q(c[881]) );
  DFF \creg_reg[882]  ( .D(creg_next[882]), .CLK(clk), .RST(rst), .I(m[882]), 
        .Q(c[882]) );
  DFF \creg_reg[883]  ( .D(creg_next[883]), .CLK(clk), .RST(rst), .I(m[883]), 
        .Q(c[883]) );
  DFF \creg_reg[884]  ( .D(creg_next[884]), .CLK(clk), .RST(rst), .I(m[884]), 
        .Q(c[884]) );
  DFF \creg_reg[885]  ( .D(creg_next[885]), .CLK(clk), .RST(rst), .I(m[885]), 
        .Q(c[885]) );
  DFF \creg_reg[886]  ( .D(creg_next[886]), .CLK(clk), .RST(rst), .I(m[886]), 
        .Q(c[886]) );
  DFF \creg_reg[887]  ( .D(creg_next[887]), .CLK(clk), .RST(rst), .I(m[887]), 
        .Q(c[887]) );
  DFF \creg_reg[888]  ( .D(creg_next[888]), .CLK(clk), .RST(rst), .I(m[888]), 
        .Q(c[888]) );
  DFF \creg_reg[889]  ( .D(creg_next[889]), .CLK(clk), .RST(rst), .I(m[889]), 
        .Q(c[889]) );
  DFF \creg_reg[890]  ( .D(creg_next[890]), .CLK(clk), .RST(rst), .I(m[890]), 
        .Q(c[890]) );
  DFF \creg_reg[891]  ( .D(creg_next[891]), .CLK(clk), .RST(rst), .I(m[891]), 
        .Q(c[891]) );
  DFF \creg_reg[892]  ( .D(creg_next[892]), .CLK(clk), .RST(rst), .I(m[892]), 
        .Q(c[892]) );
  DFF \creg_reg[893]  ( .D(creg_next[893]), .CLK(clk), .RST(rst), .I(m[893]), 
        .Q(c[893]) );
  DFF \creg_reg[894]  ( .D(creg_next[894]), .CLK(clk), .RST(rst), .I(m[894]), 
        .Q(c[894]) );
  DFF \creg_reg[895]  ( .D(creg_next[895]), .CLK(clk), .RST(rst), .I(m[895]), 
        .Q(c[895]) );
  DFF \creg_reg[896]  ( .D(creg_next[896]), .CLK(clk), .RST(rst), .I(m[896]), 
        .Q(c[896]) );
  DFF \creg_reg[897]  ( .D(creg_next[897]), .CLK(clk), .RST(rst), .I(m[897]), 
        .Q(c[897]) );
  DFF \creg_reg[898]  ( .D(creg_next[898]), .CLK(clk), .RST(rst), .I(m[898]), 
        .Q(c[898]) );
  DFF \creg_reg[899]  ( .D(creg_next[899]), .CLK(clk), .RST(rst), .I(m[899]), 
        .Q(c[899]) );
  DFF \creg_reg[900]  ( .D(creg_next[900]), .CLK(clk), .RST(rst), .I(m[900]), 
        .Q(c[900]) );
  DFF \creg_reg[901]  ( .D(creg_next[901]), .CLK(clk), .RST(rst), .I(m[901]), 
        .Q(c[901]) );
  DFF \creg_reg[902]  ( .D(creg_next[902]), .CLK(clk), .RST(rst), .I(m[902]), 
        .Q(c[902]) );
  DFF \creg_reg[903]  ( .D(creg_next[903]), .CLK(clk), .RST(rst), .I(m[903]), 
        .Q(c[903]) );
  DFF \creg_reg[904]  ( .D(creg_next[904]), .CLK(clk), .RST(rst), .I(m[904]), 
        .Q(c[904]) );
  DFF \creg_reg[905]  ( .D(creg_next[905]), .CLK(clk), .RST(rst), .I(m[905]), 
        .Q(c[905]) );
  DFF \creg_reg[906]  ( .D(creg_next[906]), .CLK(clk), .RST(rst), .I(m[906]), 
        .Q(c[906]) );
  DFF \creg_reg[907]  ( .D(creg_next[907]), .CLK(clk), .RST(rst), .I(m[907]), 
        .Q(c[907]) );
  DFF \creg_reg[908]  ( .D(creg_next[908]), .CLK(clk), .RST(rst), .I(m[908]), 
        .Q(c[908]) );
  DFF \creg_reg[909]  ( .D(creg_next[909]), .CLK(clk), .RST(rst), .I(m[909]), 
        .Q(c[909]) );
  DFF \creg_reg[910]  ( .D(creg_next[910]), .CLK(clk), .RST(rst), .I(m[910]), 
        .Q(c[910]) );
  DFF \creg_reg[911]  ( .D(creg_next[911]), .CLK(clk), .RST(rst), .I(m[911]), 
        .Q(c[911]) );
  DFF \creg_reg[912]  ( .D(creg_next[912]), .CLK(clk), .RST(rst), .I(m[912]), 
        .Q(c[912]) );
  DFF \creg_reg[913]  ( .D(creg_next[913]), .CLK(clk), .RST(rst), .I(m[913]), 
        .Q(c[913]) );
  DFF \creg_reg[914]  ( .D(creg_next[914]), .CLK(clk), .RST(rst), .I(m[914]), 
        .Q(c[914]) );
  DFF \creg_reg[915]  ( .D(creg_next[915]), .CLK(clk), .RST(rst), .I(m[915]), 
        .Q(c[915]) );
  DFF \creg_reg[916]  ( .D(creg_next[916]), .CLK(clk), .RST(rst), .I(m[916]), 
        .Q(c[916]) );
  DFF \creg_reg[917]  ( .D(creg_next[917]), .CLK(clk), .RST(rst), .I(m[917]), 
        .Q(c[917]) );
  DFF \creg_reg[918]  ( .D(creg_next[918]), .CLK(clk), .RST(rst), .I(m[918]), 
        .Q(c[918]) );
  DFF \creg_reg[919]  ( .D(creg_next[919]), .CLK(clk), .RST(rst), .I(m[919]), 
        .Q(c[919]) );
  DFF \creg_reg[920]  ( .D(creg_next[920]), .CLK(clk), .RST(rst), .I(m[920]), 
        .Q(c[920]) );
  DFF \creg_reg[921]  ( .D(creg_next[921]), .CLK(clk), .RST(rst), .I(m[921]), 
        .Q(c[921]) );
  DFF \creg_reg[922]  ( .D(creg_next[922]), .CLK(clk), .RST(rst), .I(m[922]), 
        .Q(c[922]) );
  DFF \creg_reg[923]  ( .D(creg_next[923]), .CLK(clk), .RST(rst), .I(m[923]), 
        .Q(c[923]) );
  DFF \creg_reg[924]  ( .D(creg_next[924]), .CLK(clk), .RST(rst), .I(m[924]), 
        .Q(c[924]) );
  DFF \creg_reg[925]  ( .D(creg_next[925]), .CLK(clk), .RST(rst), .I(m[925]), 
        .Q(c[925]) );
  DFF \creg_reg[926]  ( .D(creg_next[926]), .CLK(clk), .RST(rst), .I(m[926]), 
        .Q(c[926]) );
  DFF \creg_reg[927]  ( .D(creg_next[927]), .CLK(clk), .RST(rst), .I(m[927]), 
        .Q(c[927]) );
  DFF \creg_reg[928]  ( .D(creg_next[928]), .CLK(clk), .RST(rst), .I(m[928]), 
        .Q(c[928]) );
  DFF \creg_reg[929]  ( .D(creg_next[929]), .CLK(clk), .RST(rst), .I(m[929]), 
        .Q(c[929]) );
  DFF \creg_reg[930]  ( .D(creg_next[930]), .CLK(clk), .RST(rst), .I(m[930]), 
        .Q(c[930]) );
  DFF \creg_reg[931]  ( .D(creg_next[931]), .CLK(clk), .RST(rst), .I(m[931]), 
        .Q(c[931]) );
  DFF \creg_reg[932]  ( .D(creg_next[932]), .CLK(clk), .RST(rst), .I(m[932]), 
        .Q(c[932]) );
  DFF \creg_reg[933]  ( .D(creg_next[933]), .CLK(clk), .RST(rst), .I(m[933]), 
        .Q(c[933]) );
  DFF \creg_reg[934]  ( .D(creg_next[934]), .CLK(clk), .RST(rst), .I(m[934]), 
        .Q(c[934]) );
  DFF \creg_reg[935]  ( .D(creg_next[935]), .CLK(clk), .RST(rst), .I(m[935]), 
        .Q(c[935]) );
  DFF \creg_reg[936]  ( .D(creg_next[936]), .CLK(clk), .RST(rst), .I(m[936]), 
        .Q(c[936]) );
  DFF \creg_reg[937]  ( .D(creg_next[937]), .CLK(clk), .RST(rst), .I(m[937]), 
        .Q(c[937]) );
  DFF \creg_reg[938]  ( .D(creg_next[938]), .CLK(clk), .RST(rst), .I(m[938]), 
        .Q(c[938]) );
  DFF \creg_reg[939]  ( .D(creg_next[939]), .CLK(clk), .RST(rst), .I(m[939]), 
        .Q(c[939]) );
  DFF \creg_reg[940]  ( .D(creg_next[940]), .CLK(clk), .RST(rst), .I(m[940]), 
        .Q(c[940]) );
  DFF \creg_reg[941]  ( .D(creg_next[941]), .CLK(clk), .RST(rst), .I(m[941]), 
        .Q(c[941]) );
  DFF \creg_reg[942]  ( .D(creg_next[942]), .CLK(clk), .RST(rst), .I(m[942]), 
        .Q(c[942]) );
  DFF \creg_reg[943]  ( .D(creg_next[943]), .CLK(clk), .RST(rst), .I(m[943]), 
        .Q(c[943]) );
  DFF \creg_reg[944]  ( .D(creg_next[944]), .CLK(clk), .RST(rst), .I(m[944]), 
        .Q(c[944]) );
  DFF \creg_reg[945]  ( .D(creg_next[945]), .CLK(clk), .RST(rst), .I(m[945]), 
        .Q(c[945]) );
  DFF \creg_reg[946]  ( .D(creg_next[946]), .CLK(clk), .RST(rst), .I(m[946]), 
        .Q(c[946]) );
  DFF \creg_reg[947]  ( .D(creg_next[947]), .CLK(clk), .RST(rst), .I(m[947]), 
        .Q(c[947]) );
  DFF \creg_reg[948]  ( .D(creg_next[948]), .CLK(clk), .RST(rst), .I(m[948]), 
        .Q(c[948]) );
  DFF \creg_reg[949]  ( .D(creg_next[949]), .CLK(clk), .RST(rst), .I(m[949]), 
        .Q(c[949]) );
  DFF \creg_reg[950]  ( .D(creg_next[950]), .CLK(clk), .RST(rst), .I(m[950]), 
        .Q(c[950]) );
  DFF \creg_reg[951]  ( .D(creg_next[951]), .CLK(clk), .RST(rst), .I(m[951]), 
        .Q(c[951]) );
  DFF \creg_reg[952]  ( .D(creg_next[952]), .CLK(clk), .RST(rst), .I(m[952]), 
        .Q(c[952]) );
  DFF \creg_reg[953]  ( .D(creg_next[953]), .CLK(clk), .RST(rst), .I(m[953]), 
        .Q(c[953]) );
  DFF \creg_reg[954]  ( .D(creg_next[954]), .CLK(clk), .RST(rst), .I(m[954]), 
        .Q(c[954]) );
  DFF \creg_reg[955]  ( .D(creg_next[955]), .CLK(clk), .RST(rst), .I(m[955]), 
        .Q(c[955]) );
  DFF \creg_reg[956]  ( .D(creg_next[956]), .CLK(clk), .RST(rst), .I(m[956]), 
        .Q(c[956]) );
  DFF \creg_reg[957]  ( .D(creg_next[957]), .CLK(clk), .RST(rst), .I(m[957]), 
        .Q(c[957]) );
  DFF \creg_reg[958]  ( .D(creg_next[958]), .CLK(clk), .RST(rst), .I(m[958]), 
        .Q(c[958]) );
  DFF \creg_reg[959]  ( .D(creg_next[959]), .CLK(clk), .RST(rst), .I(m[959]), 
        .Q(c[959]) );
  DFF \creg_reg[960]  ( .D(creg_next[960]), .CLK(clk), .RST(rst), .I(m[960]), 
        .Q(c[960]) );
  DFF \creg_reg[961]  ( .D(creg_next[961]), .CLK(clk), .RST(rst), .I(m[961]), 
        .Q(c[961]) );
  DFF \creg_reg[962]  ( .D(creg_next[962]), .CLK(clk), .RST(rst), .I(m[962]), 
        .Q(c[962]) );
  DFF \creg_reg[963]  ( .D(creg_next[963]), .CLK(clk), .RST(rst), .I(m[963]), 
        .Q(c[963]) );
  DFF \creg_reg[964]  ( .D(creg_next[964]), .CLK(clk), .RST(rst), .I(m[964]), 
        .Q(c[964]) );
  DFF \creg_reg[965]  ( .D(creg_next[965]), .CLK(clk), .RST(rst), .I(m[965]), 
        .Q(c[965]) );
  DFF \creg_reg[966]  ( .D(creg_next[966]), .CLK(clk), .RST(rst), .I(m[966]), 
        .Q(c[966]) );
  DFF \creg_reg[967]  ( .D(creg_next[967]), .CLK(clk), .RST(rst), .I(m[967]), 
        .Q(c[967]) );
  DFF \creg_reg[968]  ( .D(creg_next[968]), .CLK(clk), .RST(rst), .I(m[968]), 
        .Q(c[968]) );
  DFF \creg_reg[969]  ( .D(creg_next[969]), .CLK(clk), .RST(rst), .I(m[969]), 
        .Q(c[969]) );
  DFF \creg_reg[970]  ( .D(creg_next[970]), .CLK(clk), .RST(rst), .I(m[970]), 
        .Q(c[970]) );
  DFF \creg_reg[971]  ( .D(creg_next[971]), .CLK(clk), .RST(rst), .I(m[971]), 
        .Q(c[971]) );
  DFF \creg_reg[972]  ( .D(creg_next[972]), .CLK(clk), .RST(rst), .I(m[972]), 
        .Q(c[972]) );
  DFF \creg_reg[973]  ( .D(creg_next[973]), .CLK(clk), .RST(rst), .I(m[973]), 
        .Q(c[973]) );
  DFF \creg_reg[974]  ( .D(creg_next[974]), .CLK(clk), .RST(rst), .I(m[974]), 
        .Q(c[974]) );
  DFF \creg_reg[975]  ( .D(creg_next[975]), .CLK(clk), .RST(rst), .I(m[975]), 
        .Q(c[975]) );
  DFF \creg_reg[976]  ( .D(creg_next[976]), .CLK(clk), .RST(rst), .I(m[976]), 
        .Q(c[976]) );
  DFF \creg_reg[977]  ( .D(creg_next[977]), .CLK(clk), .RST(rst), .I(m[977]), 
        .Q(c[977]) );
  DFF \creg_reg[978]  ( .D(creg_next[978]), .CLK(clk), .RST(rst), .I(m[978]), 
        .Q(c[978]) );
  DFF \creg_reg[979]  ( .D(creg_next[979]), .CLK(clk), .RST(rst), .I(m[979]), 
        .Q(c[979]) );
  DFF \creg_reg[980]  ( .D(creg_next[980]), .CLK(clk), .RST(rst), .I(m[980]), 
        .Q(c[980]) );
  DFF \creg_reg[981]  ( .D(creg_next[981]), .CLK(clk), .RST(rst), .I(m[981]), 
        .Q(c[981]) );
  DFF \creg_reg[982]  ( .D(creg_next[982]), .CLK(clk), .RST(rst), .I(m[982]), 
        .Q(c[982]) );
  DFF \creg_reg[983]  ( .D(creg_next[983]), .CLK(clk), .RST(rst), .I(m[983]), 
        .Q(c[983]) );
  DFF \creg_reg[984]  ( .D(creg_next[984]), .CLK(clk), .RST(rst), .I(m[984]), 
        .Q(c[984]) );
  DFF \creg_reg[985]  ( .D(creg_next[985]), .CLK(clk), .RST(rst), .I(m[985]), 
        .Q(c[985]) );
  DFF \creg_reg[986]  ( .D(creg_next[986]), .CLK(clk), .RST(rst), .I(m[986]), 
        .Q(c[986]) );
  DFF \creg_reg[987]  ( .D(creg_next[987]), .CLK(clk), .RST(rst), .I(m[987]), 
        .Q(c[987]) );
  DFF \creg_reg[988]  ( .D(creg_next[988]), .CLK(clk), .RST(rst), .I(m[988]), 
        .Q(c[988]) );
  DFF \creg_reg[989]  ( .D(creg_next[989]), .CLK(clk), .RST(rst), .I(m[989]), 
        .Q(c[989]) );
  DFF \creg_reg[990]  ( .D(creg_next[990]), .CLK(clk), .RST(rst), .I(m[990]), 
        .Q(c[990]) );
  DFF \creg_reg[991]  ( .D(creg_next[991]), .CLK(clk), .RST(rst), .I(m[991]), 
        .Q(c[991]) );
  DFF \creg_reg[992]  ( .D(creg_next[992]), .CLK(clk), .RST(rst), .I(m[992]), 
        .Q(c[992]) );
  DFF \creg_reg[993]  ( .D(creg_next[993]), .CLK(clk), .RST(rst), .I(m[993]), 
        .Q(c[993]) );
  DFF \creg_reg[994]  ( .D(creg_next[994]), .CLK(clk), .RST(rst), .I(m[994]), 
        .Q(c[994]) );
  DFF \creg_reg[995]  ( .D(creg_next[995]), .CLK(clk), .RST(rst), .I(m[995]), 
        .Q(c[995]) );
  DFF \creg_reg[996]  ( .D(creg_next[996]), .CLK(clk), .RST(rst), .I(m[996]), 
        .Q(c[996]) );
  DFF \creg_reg[997]  ( .D(creg_next[997]), .CLK(clk), .RST(rst), .I(m[997]), 
        .Q(c[997]) );
  DFF \creg_reg[998]  ( .D(creg_next[998]), .CLK(clk), .RST(rst), .I(m[998]), 
        .Q(c[998]) );
  DFF \creg_reg[999]  ( .D(creg_next[999]), .CLK(clk), .RST(rst), .I(m[999]), 
        .Q(c[999]) );
  DFF \creg_reg[1000]  ( .D(creg_next[1000]), .CLK(clk), .RST(rst), .I(m[1000]), .Q(c[1000]) );
  DFF \creg_reg[1001]  ( .D(creg_next[1001]), .CLK(clk), .RST(rst), .I(m[1001]), .Q(c[1001]) );
  DFF \creg_reg[1002]  ( .D(creg_next[1002]), .CLK(clk), .RST(rst), .I(m[1002]), .Q(c[1002]) );
  DFF \creg_reg[1003]  ( .D(creg_next[1003]), .CLK(clk), .RST(rst), .I(m[1003]), .Q(c[1003]) );
  DFF \creg_reg[1004]  ( .D(creg_next[1004]), .CLK(clk), .RST(rst), .I(m[1004]), .Q(c[1004]) );
  DFF \creg_reg[1005]  ( .D(creg_next[1005]), .CLK(clk), .RST(rst), .I(m[1005]), .Q(c[1005]) );
  DFF \creg_reg[1006]  ( .D(creg_next[1006]), .CLK(clk), .RST(rst), .I(m[1006]), .Q(c[1006]) );
  DFF \creg_reg[1007]  ( .D(creg_next[1007]), .CLK(clk), .RST(rst), .I(m[1007]), .Q(c[1007]) );
  DFF \creg_reg[1008]  ( .D(creg_next[1008]), .CLK(clk), .RST(rst), .I(m[1008]), .Q(c[1008]) );
  DFF \creg_reg[1009]  ( .D(creg_next[1009]), .CLK(clk), .RST(rst), .I(m[1009]), .Q(c[1009]) );
  DFF \creg_reg[1010]  ( .D(creg_next[1010]), .CLK(clk), .RST(rst), .I(m[1010]), .Q(c[1010]) );
  DFF \creg_reg[1011]  ( .D(creg_next[1011]), .CLK(clk), .RST(rst), .I(m[1011]), .Q(c[1011]) );
  DFF \creg_reg[1012]  ( .D(creg_next[1012]), .CLK(clk), .RST(rst), .I(m[1012]), .Q(c[1012]) );
  DFF \creg_reg[1013]  ( .D(creg_next[1013]), .CLK(clk), .RST(rst), .I(m[1013]), .Q(c[1013]) );
  DFF \creg_reg[1014]  ( .D(creg_next[1014]), .CLK(clk), .RST(rst), .I(m[1014]), .Q(c[1014]) );
  DFF \creg_reg[1015]  ( .D(creg_next[1015]), .CLK(clk), .RST(rst), .I(m[1015]), .Q(c[1015]) );
  DFF \creg_reg[1016]  ( .D(creg_next[1016]), .CLK(clk), .RST(rst), .I(m[1016]), .Q(c[1016]) );
  DFF \creg_reg[1017]  ( .D(creg_next[1017]), .CLK(clk), .RST(rst), .I(m[1017]), .Q(c[1017]) );
  DFF \creg_reg[1018]  ( .D(creg_next[1018]), .CLK(clk), .RST(rst), .I(m[1018]), .Q(c[1018]) );
  DFF \creg_reg[1019]  ( .D(creg_next[1019]), .CLK(clk), .RST(rst), .I(m[1019]), .Q(c[1019]) );
  DFF \creg_reg[1020]  ( .D(creg_next[1020]), .CLK(clk), .RST(rst), .I(m[1020]), .Q(c[1020]) );
  DFF \creg_reg[1021]  ( .D(creg_next[1021]), .CLK(clk), .RST(rst), .I(m[1021]), .Q(c[1021]) );
  DFF \creg_reg[1022]  ( .D(creg_next[1022]), .CLK(clk), .RST(rst), .I(m[1022]), .Q(c[1022]) );
  DFF \creg_reg[1023]  ( .D(creg_next[1023]), .CLK(clk), .RST(rst), .I(m[1023]), .Q(c[1023]) );
  DFF \modmult_1/zreg_reg[1024]  ( .D(\modmult_1/zout[0][1024] ), .CLK(clk), 
        .RST(start_in[0]), .I(1'b0), .Q(\modmult_1/zin[0][1024] ) );
  DFF \modmult_1/zreg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1023] ) );
  DFF \modmult_1/zreg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1022] ) );
  DFF \modmult_1/zreg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1021] ) );
  DFF \modmult_1/zreg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1020] ) );
  DFF \modmult_1/zreg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1019] ) );
  DFF \modmult_1/zreg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1018] ) );
  DFF \modmult_1/zreg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1017] ) );
  DFF \modmult_1/zreg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1016] ) );
  DFF \modmult_1/zreg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1015] ) );
  DFF \modmult_1/zreg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1014] ) );
  DFF \modmult_1/zreg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1013] ) );
  DFF \modmult_1/zreg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1012] ) );
  DFF \modmult_1/zreg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1011] ) );
  DFF \modmult_1/zreg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1010] ) );
  DFF \modmult_1/zreg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1009] ) );
  DFF \modmult_1/zreg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1008] ) );
  DFF \modmult_1/zreg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1007] ) );
  DFF \modmult_1/zreg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1006] ) );
  DFF \modmult_1/zreg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1005] ) );
  DFF \modmult_1/zreg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1004] ) );
  DFF \modmult_1/zreg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1003] ) );
  DFF \modmult_1/zreg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1002] ) );
  DFF \modmult_1/zreg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1001] ) );
  DFF \modmult_1/zreg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][1000] ) );
  DFF \modmult_1/zreg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][999] ) );
  DFF \modmult_1/zreg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][998] ) );
  DFF \modmult_1/zreg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][997] ) );
  DFF \modmult_1/zreg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][996] ) );
  DFF \modmult_1/zreg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][995] ) );
  DFF \modmult_1/zreg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][994] ) );
  DFF \modmult_1/zreg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][993] ) );
  DFF \modmult_1/zreg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][992] ) );
  DFF \modmult_1/zreg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][991] ) );
  DFF \modmult_1/zreg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][990] ) );
  DFF \modmult_1/zreg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][989] ) );
  DFF \modmult_1/zreg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][988] ) );
  DFF \modmult_1/zreg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][987] ) );
  DFF \modmult_1/zreg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][986] ) );
  DFF \modmult_1/zreg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][985] ) );
  DFF \modmult_1/zreg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][984] ) );
  DFF \modmult_1/zreg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][983] ) );
  DFF \modmult_1/zreg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][982] ) );
  DFF \modmult_1/zreg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][981] ) );
  DFF \modmult_1/zreg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][980] ) );
  DFF \modmult_1/zreg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][979] ) );
  DFF \modmult_1/zreg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][978] ) );
  DFF \modmult_1/zreg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][977] ) );
  DFF \modmult_1/zreg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][976] ) );
  DFF \modmult_1/zreg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][975] ) );
  DFF \modmult_1/zreg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][974] ) );
  DFF \modmult_1/zreg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][973] ) );
  DFF \modmult_1/zreg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][972] ) );
  DFF \modmult_1/zreg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][971] ) );
  DFF \modmult_1/zreg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][970] ) );
  DFF \modmult_1/zreg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][969] ) );
  DFF \modmult_1/zreg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][968] ) );
  DFF \modmult_1/zreg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][967] ) );
  DFF \modmult_1/zreg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][966] ) );
  DFF \modmult_1/zreg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][965] ) );
  DFF \modmult_1/zreg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][964] ) );
  DFF \modmult_1/zreg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][963] ) );
  DFF \modmult_1/zreg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][962] ) );
  DFF \modmult_1/zreg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][961] ) );
  DFF \modmult_1/zreg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][960] ) );
  DFF \modmult_1/zreg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][959] ) );
  DFF \modmult_1/zreg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][958] ) );
  DFF \modmult_1/zreg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][957] ) );
  DFF \modmult_1/zreg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][956] ) );
  DFF \modmult_1/zreg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][955] ) );
  DFF \modmult_1/zreg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][954] ) );
  DFF \modmult_1/zreg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][953] ) );
  DFF \modmult_1/zreg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][952] ) );
  DFF \modmult_1/zreg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][951] ) );
  DFF \modmult_1/zreg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][950] ) );
  DFF \modmult_1/zreg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][949] ) );
  DFF \modmult_1/zreg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][948] ) );
  DFF \modmult_1/zreg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][947] ) );
  DFF \modmult_1/zreg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][946] ) );
  DFF \modmult_1/zreg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][945] ) );
  DFF \modmult_1/zreg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][944] ) );
  DFF \modmult_1/zreg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][943] ) );
  DFF \modmult_1/zreg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][942] ) );
  DFF \modmult_1/zreg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][941] ) );
  DFF \modmult_1/zreg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][940] ) );
  DFF \modmult_1/zreg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][939] ) );
  DFF \modmult_1/zreg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][938] ) );
  DFF \modmult_1/zreg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][937] ) );
  DFF \modmult_1/zreg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][936] ) );
  DFF \modmult_1/zreg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][935] ) );
  DFF \modmult_1/zreg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][934] ) );
  DFF \modmult_1/zreg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][933] ) );
  DFF \modmult_1/zreg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][932] ) );
  DFF \modmult_1/zreg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][931] ) );
  DFF \modmult_1/zreg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][930] ) );
  DFF \modmult_1/zreg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][929] ) );
  DFF \modmult_1/zreg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][928] ) );
  DFF \modmult_1/zreg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][927] ) );
  DFF \modmult_1/zreg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][926] ) );
  DFF \modmult_1/zreg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][925] ) );
  DFF \modmult_1/zreg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][924] ) );
  DFF \modmult_1/zreg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][923] ) );
  DFF \modmult_1/zreg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][922] ) );
  DFF \modmult_1/zreg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][921] ) );
  DFF \modmult_1/zreg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][920] ) );
  DFF \modmult_1/zreg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][919] ) );
  DFF \modmult_1/zreg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][918] ) );
  DFF \modmult_1/zreg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][917] ) );
  DFF \modmult_1/zreg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][916] ) );
  DFF \modmult_1/zreg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][915] ) );
  DFF \modmult_1/zreg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][914] ) );
  DFF \modmult_1/zreg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][913] ) );
  DFF \modmult_1/zreg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][912] ) );
  DFF \modmult_1/zreg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][911] ) );
  DFF \modmult_1/zreg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][910] ) );
  DFF \modmult_1/zreg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][909] ) );
  DFF \modmult_1/zreg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][908] ) );
  DFF \modmult_1/zreg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][907] ) );
  DFF \modmult_1/zreg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][906] ) );
  DFF \modmult_1/zreg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][905] ) );
  DFF \modmult_1/zreg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][904] ) );
  DFF \modmult_1/zreg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][903] ) );
  DFF \modmult_1/zreg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][902] ) );
  DFF \modmult_1/zreg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][901] ) );
  DFF \modmult_1/zreg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][900] ) );
  DFF \modmult_1/zreg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][899] ) );
  DFF \modmult_1/zreg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][898] ) );
  DFF \modmult_1/zreg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][897] ) );
  DFF \modmult_1/zreg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][896] ) );
  DFF \modmult_1/zreg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][895] ) );
  DFF \modmult_1/zreg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][894] ) );
  DFF \modmult_1/zreg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][893] ) );
  DFF \modmult_1/zreg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][892] ) );
  DFF \modmult_1/zreg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][891] ) );
  DFF \modmult_1/zreg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][890] ) );
  DFF \modmult_1/zreg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][889] ) );
  DFF \modmult_1/zreg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][888] ) );
  DFF \modmult_1/zreg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][887] ) );
  DFF \modmult_1/zreg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][886] ) );
  DFF \modmult_1/zreg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][885] ) );
  DFF \modmult_1/zreg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][884] ) );
  DFF \modmult_1/zreg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][883] ) );
  DFF \modmult_1/zreg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][882] ) );
  DFF \modmult_1/zreg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][881] ) );
  DFF \modmult_1/zreg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][880] ) );
  DFF \modmult_1/zreg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][879] ) );
  DFF \modmult_1/zreg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][878] ) );
  DFF \modmult_1/zreg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][877] ) );
  DFF \modmult_1/zreg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][876] ) );
  DFF \modmult_1/zreg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][875] ) );
  DFF \modmult_1/zreg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][874] ) );
  DFF \modmult_1/zreg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][873] ) );
  DFF \modmult_1/zreg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][872] ) );
  DFF \modmult_1/zreg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][871] ) );
  DFF \modmult_1/zreg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][870] ) );
  DFF \modmult_1/zreg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][869] ) );
  DFF \modmult_1/zreg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][868] ) );
  DFF \modmult_1/zreg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][867] ) );
  DFF \modmult_1/zreg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][866] ) );
  DFF \modmult_1/zreg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][865] ) );
  DFF \modmult_1/zreg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][864] ) );
  DFF \modmult_1/zreg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][863] ) );
  DFF \modmult_1/zreg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][862] ) );
  DFF \modmult_1/zreg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][861] ) );
  DFF \modmult_1/zreg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][860] ) );
  DFF \modmult_1/zreg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][859] ) );
  DFF \modmult_1/zreg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][858] ) );
  DFF \modmult_1/zreg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][857] ) );
  DFF \modmult_1/zreg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][856] ) );
  DFF \modmult_1/zreg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][855] ) );
  DFF \modmult_1/zreg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][854] ) );
  DFF \modmult_1/zreg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][853] ) );
  DFF \modmult_1/zreg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][852] ) );
  DFF \modmult_1/zreg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][851] ) );
  DFF \modmult_1/zreg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][850] ) );
  DFF \modmult_1/zreg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][849] ) );
  DFF \modmult_1/zreg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][848] ) );
  DFF \modmult_1/zreg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][847] ) );
  DFF \modmult_1/zreg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][846] ) );
  DFF \modmult_1/zreg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][845] ) );
  DFF \modmult_1/zreg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][844] ) );
  DFF \modmult_1/zreg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][843] ) );
  DFF \modmult_1/zreg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][842] ) );
  DFF \modmult_1/zreg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][841] ) );
  DFF \modmult_1/zreg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][840] ) );
  DFF \modmult_1/zreg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][839] ) );
  DFF \modmult_1/zreg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][838] ) );
  DFF \modmult_1/zreg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][837] ) );
  DFF \modmult_1/zreg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][836] ) );
  DFF \modmult_1/zreg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][835] ) );
  DFF \modmult_1/zreg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][834] ) );
  DFF \modmult_1/zreg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][833] ) );
  DFF \modmult_1/zreg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][832] ) );
  DFF \modmult_1/zreg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][831] ) );
  DFF \modmult_1/zreg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][830] ) );
  DFF \modmult_1/zreg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][829] ) );
  DFF \modmult_1/zreg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][828] ) );
  DFF \modmult_1/zreg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][827] ) );
  DFF \modmult_1/zreg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][826] ) );
  DFF \modmult_1/zreg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][825] ) );
  DFF \modmult_1/zreg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][824] ) );
  DFF \modmult_1/zreg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][823] ) );
  DFF \modmult_1/zreg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][822] ) );
  DFF \modmult_1/zreg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][821] ) );
  DFF \modmult_1/zreg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][820] ) );
  DFF \modmult_1/zreg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][819] ) );
  DFF \modmult_1/zreg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][818] ) );
  DFF \modmult_1/zreg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][817] ) );
  DFF \modmult_1/zreg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][816] ) );
  DFF \modmult_1/zreg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][815] ) );
  DFF \modmult_1/zreg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][814] ) );
  DFF \modmult_1/zreg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][813] ) );
  DFF \modmult_1/zreg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][812] ) );
  DFF \modmult_1/zreg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][811] ) );
  DFF \modmult_1/zreg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][810] ) );
  DFF \modmult_1/zreg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][809] ) );
  DFF \modmult_1/zreg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][808] ) );
  DFF \modmult_1/zreg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][807] ) );
  DFF \modmult_1/zreg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][806] ) );
  DFF \modmult_1/zreg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][805] ) );
  DFF \modmult_1/zreg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][804] ) );
  DFF \modmult_1/zreg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][803] ) );
  DFF \modmult_1/zreg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][802] ) );
  DFF \modmult_1/zreg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][801] ) );
  DFF \modmult_1/zreg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][800] ) );
  DFF \modmult_1/zreg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][799] ) );
  DFF \modmult_1/zreg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][798] ) );
  DFF \modmult_1/zreg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][797] ) );
  DFF \modmult_1/zreg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][796] ) );
  DFF \modmult_1/zreg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][795] ) );
  DFF \modmult_1/zreg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][794] ) );
  DFF \modmult_1/zreg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][793] ) );
  DFF \modmult_1/zreg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][792] ) );
  DFF \modmult_1/zreg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][791] ) );
  DFF \modmult_1/zreg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][790] ) );
  DFF \modmult_1/zreg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][789] ) );
  DFF \modmult_1/zreg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][788] ) );
  DFF \modmult_1/zreg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][787] ) );
  DFF \modmult_1/zreg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][786] ) );
  DFF \modmult_1/zreg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][785] ) );
  DFF \modmult_1/zreg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][784] ) );
  DFF \modmult_1/zreg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][783] ) );
  DFF \modmult_1/zreg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][782] ) );
  DFF \modmult_1/zreg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][781] ) );
  DFF \modmult_1/zreg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][780] ) );
  DFF \modmult_1/zreg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][779] ) );
  DFF \modmult_1/zreg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][778] ) );
  DFF \modmult_1/zreg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][777] ) );
  DFF \modmult_1/zreg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][776] ) );
  DFF \modmult_1/zreg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][775] ) );
  DFF \modmult_1/zreg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][774] ) );
  DFF \modmult_1/zreg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][773] ) );
  DFF \modmult_1/zreg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][772] ) );
  DFF \modmult_1/zreg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][771] ) );
  DFF \modmult_1/zreg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][770] ) );
  DFF \modmult_1/zreg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][769] ) );
  DFF \modmult_1/zreg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][768] ) );
  DFF \modmult_1/zreg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][767] ) );
  DFF \modmult_1/zreg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][766] ) );
  DFF \modmult_1/zreg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][765] ) );
  DFF \modmult_1/zreg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][764] ) );
  DFF \modmult_1/zreg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][763] ) );
  DFF \modmult_1/zreg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][762] ) );
  DFF \modmult_1/zreg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][761] ) );
  DFF \modmult_1/zreg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][760] ) );
  DFF \modmult_1/zreg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][759] ) );
  DFF \modmult_1/zreg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][758] ) );
  DFF \modmult_1/zreg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][757] ) );
  DFF \modmult_1/zreg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][756] ) );
  DFF \modmult_1/zreg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][755] ) );
  DFF \modmult_1/zreg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][754] ) );
  DFF \modmult_1/zreg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][753] ) );
  DFF \modmult_1/zreg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][752] ) );
  DFF \modmult_1/zreg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][751] ) );
  DFF \modmult_1/zreg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][750] ) );
  DFF \modmult_1/zreg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][749] ) );
  DFF \modmult_1/zreg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][748] ) );
  DFF \modmult_1/zreg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][747] ) );
  DFF \modmult_1/zreg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][746] ) );
  DFF \modmult_1/zreg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][745] ) );
  DFF \modmult_1/zreg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][744] ) );
  DFF \modmult_1/zreg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][743] ) );
  DFF \modmult_1/zreg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][742] ) );
  DFF \modmult_1/zreg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][741] ) );
  DFF \modmult_1/zreg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][740] ) );
  DFF \modmult_1/zreg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][739] ) );
  DFF \modmult_1/zreg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][738] ) );
  DFF \modmult_1/zreg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][737] ) );
  DFF \modmult_1/zreg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][736] ) );
  DFF \modmult_1/zreg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][735] ) );
  DFF \modmult_1/zreg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][734] ) );
  DFF \modmult_1/zreg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][733] ) );
  DFF \modmult_1/zreg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][732] ) );
  DFF \modmult_1/zreg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][731] ) );
  DFF \modmult_1/zreg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][730] ) );
  DFF \modmult_1/zreg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][729] ) );
  DFF \modmult_1/zreg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][728] ) );
  DFF \modmult_1/zreg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][727] ) );
  DFF \modmult_1/zreg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][726] ) );
  DFF \modmult_1/zreg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][725] ) );
  DFF \modmult_1/zreg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][724] ) );
  DFF \modmult_1/zreg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][723] ) );
  DFF \modmult_1/zreg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][722] ) );
  DFF \modmult_1/zreg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][721] ) );
  DFF \modmult_1/zreg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][720] ) );
  DFF \modmult_1/zreg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][719] ) );
  DFF \modmult_1/zreg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][718] ) );
  DFF \modmult_1/zreg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][717] ) );
  DFF \modmult_1/zreg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][716] ) );
  DFF \modmult_1/zreg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][715] ) );
  DFF \modmult_1/zreg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][714] ) );
  DFF \modmult_1/zreg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][713] ) );
  DFF \modmult_1/zreg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][712] ) );
  DFF \modmult_1/zreg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][711] ) );
  DFF \modmult_1/zreg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][710] ) );
  DFF \modmult_1/zreg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][709] ) );
  DFF \modmult_1/zreg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][708] ) );
  DFF \modmult_1/zreg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][707] ) );
  DFF \modmult_1/zreg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][706] ) );
  DFF \modmult_1/zreg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][705] ) );
  DFF \modmult_1/zreg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][704] ) );
  DFF \modmult_1/zreg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][703] ) );
  DFF \modmult_1/zreg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][702] ) );
  DFF \modmult_1/zreg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][701] ) );
  DFF \modmult_1/zreg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][700] ) );
  DFF \modmult_1/zreg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][699] ) );
  DFF \modmult_1/zreg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][698] ) );
  DFF \modmult_1/zreg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][697] ) );
  DFF \modmult_1/zreg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][696] ) );
  DFF \modmult_1/zreg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][695] ) );
  DFF \modmult_1/zreg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][694] ) );
  DFF \modmult_1/zreg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][693] ) );
  DFF \modmult_1/zreg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][692] ) );
  DFF \modmult_1/zreg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][691] ) );
  DFF \modmult_1/zreg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][690] ) );
  DFF \modmult_1/zreg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][689] ) );
  DFF \modmult_1/zreg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][688] ) );
  DFF \modmult_1/zreg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][687] ) );
  DFF \modmult_1/zreg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][686] ) );
  DFF \modmult_1/zreg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][685] ) );
  DFF \modmult_1/zreg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][684] ) );
  DFF \modmult_1/zreg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][683] ) );
  DFF \modmult_1/zreg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][682] ) );
  DFF \modmult_1/zreg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][681] ) );
  DFF \modmult_1/zreg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][680] ) );
  DFF \modmult_1/zreg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][679] ) );
  DFF \modmult_1/zreg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][678] ) );
  DFF \modmult_1/zreg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][677] ) );
  DFF \modmult_1/zreg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][676] ) );
  DFF \modmult_1/zreg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][675] ) );
  DFF \modmult_1/zreg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][674] ) );
  DFF \modmult_1/zreg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][673] ) );
  DFF \modmult_1/zreg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][672] ) );
  DFF \modmult_1/zreg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][671] ) );
  DFF \modmult_1/zreg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][670] ) );
  DFF \modmult_1/zreg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][669] ) );
  DFF \modmult_1/zreg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][668] ) );
  DFF \modmult_1/zreg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][667] ) );
  DFF \modmult_1/zreg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][666] ) );
  DFF \modmult_1/zreg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][665] ) );
  DFF \modmult_1/zreg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][664] ) );
  DFF \modmult_1/zreg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][663] ) );
  DFF \modmult_1/zreg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][662] ) );
  DFF \modmult_1/zreg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][661] ) );
  DFF \modmult_1/zreg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][660] ) );
  DFF \modmult_1/zreg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][659] ) );
  DFF \modmult_1/zreg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][658] ) );
  DFF \modmult_1/zreg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][657] ) );
  DFF \modmult_1/zreg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][656] ) );
  DFF \modmult_1/zreg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][655] ) );
  DFF \modmult_1/zreg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][654] ) );
  DFF \modmult_1/zreg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][653] ) );
  DFF \modmult_1/zreg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][652] ) );
  DFF \modmult_1/zreg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][651] ) );
  DFF \modmult_1/zreg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][650] ) );
  DFF \modmult_1/zreg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][649] ) );
  DFF \modmult_1/zreg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][648] ) );
  DFF \modmult_1/zreg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][647] ) );
  DFF \modmult_1/zreg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][646] ) );
  DFF \modmult_1/zreg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][645] ) );
  DFF \modmult_1/zreg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][644] ) );
  DFF \modmult_1/zreg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][643] ) );
  DFF \modmult_1/zreg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][642] ) );
  DFF \modmult_1/zreg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][641] ) );
  DFF \modmult_1/zreg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][640] ) );
  DFF \modmult_1/zreg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][639] ) );
  DFF \modmult_1/zreg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][638] ) );
  DFF \modmult_1/zreg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][637] ) );
  DFF \modmult_1/zreg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][636] ) );
  DFF \modmult_1/zreg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][635] ) );
  DFF \modmult_1/zreg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][634] ) );
  DFF \modmult_1/zreg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][633] ) );
  DFF \modmult_1/zreg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][632] ) );
  DFF \modmult_1/zreg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][631] ) );
  DFF \modmult_1/zreg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][630] ) );
  DFF \modmult_1/zreg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][629] ) );
  DFF \modmult_1/zreg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][628] ) );
  DFF \modmult_1/zreg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][627] ) );
  DFF \modmult_1/zreg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][626] ) );
  DFF \modmult_1/zreg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][625] ) );
  DFF \modmult_1/zreg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][624] ) );
  DFF \modmult_1/zreg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][623] ) );
  DFF \modmult_1/zreg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][622] ) );
  DFF \modmult_1/zreg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][621] ) );
  DFF \modmult_1/zreg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][620] ) );
  DFF \modmult_1/zreg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][619] ) );
  DFF \modmult_1/zreg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][618] ) );
  DFF \modmult_1/zreg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][617] ) );
  DFF \modmult_1/zreg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][616] ) );
  DFF \modmult_1/zreg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][615] ) );
  DFF \modmult_1/zreg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][614] ) );
  DFF \modmult_1/zreg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][613] ) );
  DFF \modmult_1/zreg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][612] ) );
  DFF \modmult_1/zreg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][611] ) );
  DFF \modmult_1/zreg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][610] ) );
  DFF \modmult_1/zreg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][609] ) );
  DFF \modmult_1/zreg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][608] ) );
  DFF \modmult_1/zreg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][607] ) );
  DFF \modmult_1/zreg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][606] ) );
  DFF \modmult_1/zreg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][605] ) );
  DFF \modmult_1/zreg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][604] ) );
  DFF \modmult_1/zreg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][603] ) );
  DFF \modmult_1/zreg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][602] ) );
  DFF \modmult_1/zreg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][601] ) );
  DFF \modmult_1/zreg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][600] ) );
  DFF \modmult_1/zreg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][599] ) );
  DFF \modmult_1/zreg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][598] ) );
  DFF \modmult_1/zreg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][597] ) );
  DFF \modmult_1/zreg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][596] ) );
  DFF \modmult_1/zreg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][595] ) );
  DFF \modmult_1/zreg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][594] ) );
  DFF \modmult_1/zreg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][593] ) );
  DFF \modmult_1/zreg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][592] ) );
  DFF \modmult_1/zreg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][591] ) );
  DFF \modmult_1/zreg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][590] ) );
  DFF \modmult_1/zreg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][589] ) );
  DFF \modmult_1/zreg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][588] ) );
  DFF \modmult_1/zreg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][587] ) );
  DFF \modmult_1/zreg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][586] ) );
  DFF \modmult_1/zreg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][585] ) );
  DFF \modmult_1/zreg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][584] ) );
  DFF \modmult_1/zreg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][583] ) );
  DFF \modmult_1/zreg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][582] ) );
  DFF \modmult_1/zreg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][581] ) );
  DFF \modmult_1/zreg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][580] ) );
  DFF \modmult_1/zreg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][579] ) );
  DFF \modmult_1/zreg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][578] ) );
  DFF \modmult_1/zreg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][577] ) );
  DFF \modmult_1/zreg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][576] ) );
  DFF \modmult_1/zreg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][575] ) );
  DFF \modmult_1/zreg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][574] ) );
  DFF \modmult_1/zreg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][573] ) );
  DFF \modmult_1/zreg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][572] ) );
  DFF \modmult_1/zreg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][571] ) );
  DFF \modmult_1/zreg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][570] ) );
  DFF \modmult_1/zreg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][569] ) );
  DFF \modmult_1/zreg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][568] ) );
  DFF \modmult_1/zreg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][567] ) );
  DFF \modmult_1/zreg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][566] ) );
  DFF \modmult_1/zreg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][565] ) );
  DFF \modmult_1/zreg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][564] ) );
  DFF \modmult_1/zreg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][563] ) );
  DFF \modmult_1/zreg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][562] ) );
  DFF \modmult_1/zreg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][561] ) );
  DFF \modmult_1/zreg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][560] ) );
  DFF \modmult_1/zreg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][559] ) );
  DFF \modmult_1/zreg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][558] ) );
  DFF \modmult_1/zreg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][557] ) );
  DFF \modmult_1/zreg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][556] ) );
  DFF \modmult_1/zreg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][555] ) );
  DFF \modmult_1/zreg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][554] ) );
  DFF \modmult_1/zreg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][553] ) );
  DFF \modmult_1/zreg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][552] ) );
  DFF \modmult_1/zreg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][551] ) );
  DFF \modmult_1/zreg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][550] ) );
  DFF \modmult_1/zreg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][549] ) );
  DFF \modmult_1/zreg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][548] ) );
  DFF \modmult_1/zreg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][547] ) );
  DFF \modmult_1/zreg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][546] ) );
  DFF \modmult_1/zreg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][545] ) );
  DFF \modmult_1/zreg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][544] ) );
  DFF \modmult_1/zreg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][543] ) );
  DFF \modmult_1/zreg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][542] ) );
  DFF \modmult_1/zreg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][541] ) );
  DFF \modmult_1/zreg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][540] ) );
  DFF \modmult_1/zreg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][539] ) );
  DFF \modmult_1/zreg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][538] ) );
  DFF \modmult_1/zreg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][537] ) );
  DFF \modmult_1/zreg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][536] ) );
  DFF \modmult_1/zreg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][535] ) );
  DFF \modmult_1/zreg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][534] ) );
  DFF \modmult_1/zreg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][533] ) );
  DFF \modmult_1/zreg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][532] ) );
  DFF \modmult_1/zreg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][531] ) );
  DFF \modmult_1/zreg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][530] ) );
  DFF \modmult_1/zreg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][529] ) );
  DFF \modmult_1/zreg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][528] ) );
  DFF \modmult_1/zreg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][527] ) );
  DFF \modmult_1/zreg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][526] ) );
  DFF \modmult_1/zreg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][525] ) );
  DFF \modmult_1/zreg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][524] ) );
  DFF \modmult_1/zreg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][523] ) );
  DFF \modmult_1/zreg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][522] ) );
  DFF \modmult_1/zreg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][521] ) );
  DFF \modmult_1/zreg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][520] ) );
  DFF \modmult_1/zreg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][519] ) );
  DFF \modmult_1/zreg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][518] ) );
  DFF \modmult_1/zreg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][517] ) );
  DFF \modmult_1/zreg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][516] ) );
  DFF \modmult_1/zreg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][515] ) );
  DFF \modmult_1/zreg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][514] ) );
  DFF \modmult_1/zreg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][513] ) );
  DFF \modmult_1/zreg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][512] ) );
  DFF \modmult_1/zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][511] ) );
  DFF \modmult_1/zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][510] ) );
  DFF \modmult_1/zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][509] ) );
  DFF \modmult_1/zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][508] ) );
  DFF \modmult_1/zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][507] ) );
  DFF \modmult_1/zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][506] ) );
  DFF \modmult_1/zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][505] ) );
  DFF \modmult_1/zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][504] ) );
  DFF \modmult_1/zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][503] ) );
  DFF \modmult_1/zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][502] ) );
  DFF \modmult_1/zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][501] ) );
  DFF \modmult_1/zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][500] ) );
  DFF \modmult_1/zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][499] ) );
  DFF \modmult_1/zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][498] ) );
  DFF \modmult_1/zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][497] ) );
  DFF \modmult_1/zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][496] ) );
  DFF \modmult_1/zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][495] ) );
  DFF \modmult_1/zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][494] ) );
  DFF \modmult_1/zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][493] ) );
  DFF \modmult_1/zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][492] ) );
  DFF \modmult_1/zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][491] ) );
  DFF \modmult_1/zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][490] ) );
  DFF \modmult_1/zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][489] ) );
  DFF \modmult_1/zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][488] ) );
  DFF \modmult_1/zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][487] ) );
  DFF \modmult_1/zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][486] ) );
  DFF \modmult_1/zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][485] ) );
  DFF \modmult_1/zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][484] ) );
  DFF \modmult_1/zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][483] ) );
  DFF \modmult_1/zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][482] ) );
  DFF \modmult_1/zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][481] ) );
  DFF \modmult_1/zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][480] ) );
  DFF \modmult_1/zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][479] ) );
  DFF \modmult_1/zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][478] ) );
  DFF \modmult_1/zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][477] ) );
  DFF \modmult_1/zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][476] ) );
  DFF \modmult_1/zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][475] ) );
  DFF \modmult_1/zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][474] ) );
  DFF \modmult_1/zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][473] ) );
  DFF \modmult_1/zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][472] ) );
  DFF \modmult_1/zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][471] ) );
  DFF \modmult_1/zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][470] ) );
  DFF \modmult_1/zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][469] ) );
  DFF \modmult_1/zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][468] ) );
  DFF \modmult_1/zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][467] ) );
  DFF \modmult_1/zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][466] ) );
  DFF \modmult_1/zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][465] ) );
  DFF \modmult_1/zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][464] ) );
  DFF \modmult_1/zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][463] ) );
  DFF \modmult_1/zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][462] ) );
  DFF \modmult_1/zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][461] ) );
  DFF \modmult_1/zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][460] ) );
  DFF \modmult_1/zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][459] ) );
  DFF \modmult_1/zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][458] ) );
  DFF \modmult_1/zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][457] ) );
  DFF \modmult_1/zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][456] ) );
  DFF \modmult_1/zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][455] ) );
  DFF \modmult_1/zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][454] ) );
  DFF \modmult_1/zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][453] ) );
  DFF \modmult_1/zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][452] ) );
  DFF \modmult_1/zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][451] ) );
  DFF \modmult_1/zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][450] ) );
  DFF \modmult_1/zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][449] ) );
  DFF \modmult_1/zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][448] ) );
  DFF \modmult_1/zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][447] ) );
  DFF \modmult_1/zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][446] ) );
  DFF \modmult_1/zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][445] ) );
  DFF \modmult_1/zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][444] ) );
  DFF \modmult_1/zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][443] ) );
  DFF \modmult_1/zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][442] ) );
  DFF \modmult_1/zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][441] ) );
  DFF \modmult_1/zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][440] ) );
  DFF \modmult_1/zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][439] ) );
  DFF \modmult_1/zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][438] ) );
  DFF \modmult_1/zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][437] ) );
  DFF \modmult_1/zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][436] ) );
  DFF \modmult_1/zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][435] ) );
  DFF \modmult_1/zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][434] ) );
  DFF \modmult_1/zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][433] ) );
  DFF \modmult_1/zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][432] ) );
  DFF \modmult_1/zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][431] ) );
  DFF \modmult_1/zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][430] ) );
  DFF \modmult_1/zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][429] ) );
  DFF \modmult_1/zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][428] ) );
  DFF \modmult_1/zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][427] ) );
  DFF \modmult_1/zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][426] ) );
  DFF \modmult_1/zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][425] ) );
  DFF \modmult_1/zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][424] ) );
  DFF \modmult_1/zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][423] ) );
  DFF \modmult_1/zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][422] ) );
  DFF \modmult_1/zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][421] ) );
  DFF \modmult_1/zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][420] ) );
  DFF \modmult_1/zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][419] ) );
  DFF \modmult_1/zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][418] ) );
  DFF \modmult_1/zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][417] ) );
  DFF \modmult_1/zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][416] ) );
  DFF \modmult_1/zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][415] ) );
  DFF \modmult_1/zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][414] ) );
  DFF \modmult_1/zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][413] ) );
  DFF \modmult_1/zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][412] ) );
  DFF \modmult_1/zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][411] ) );
  DFF \modmult_1/zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][410] ) );
  DFF \modmult_1/zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][409] ) );
  DFF \modmult_1/zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][408] ) );
  DFF \modmult_1/zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][407] ) );
  DFF \modmult_1/zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][406] ) );
  DFF \modmult_1/zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][405] ) );
  DFF \modmult_1/zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][404] ) );
  DFF \modmult_1/zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][403] ) );
  DFF \modmult_1/zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][402] ) );
  DFF \modmult_1/zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][401] ) );
  DFF \modmult_1/zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][400] ) );
  DFF \modmult_1/zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][399] ) );
  DFF \modmult_1/zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][398] ) );
  DFF \modmult_1/zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][397] ) );
  DFF \modmult_1/zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][396] ) );
  DFF \modmult_1/zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][395] ) );
  DFF \modmult_1/zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][394] ) );
  DFF \modmult_1/zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][393] ) );
  DFF \modmult_1/zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][392] ) );
  DFF \modmult_1/zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][391] ) );
  DFF \modmult_1/zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][390] ) );
  DFF \modmult_1/zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][389] ) );
  DFF \modmult_1/zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][388] ) );
  DFF \modmult_1/zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][387] ) );
  DFF \modmult_1/zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][386] ) );
  DFF \modmult_1/zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][385] ) );
  DFF \modmult_1/zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][384] ) );
  DFF \modmult_1/zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][383] ) );
  DFF \modmult_1/zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][382] ) );
  DFF \modmult_1/zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][381] ) );
  DFF \modmult_1/zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][380] ) );
  DFF \modmult_1/zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][379] ) );
  DFF \modmult_1/zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][378] ) );
  DFF \modmult_1/zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][377] ) );
  DFF \modmult_1/zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][376] ) );
  DFF \modmult_1/zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][375] ) );
  DFF \modmult_1/zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][374] ) );
  DFF \modmult_1/zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][373] ) );
  DFF \modmult_1/zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][372] ) );
  DFF \modmult_1/zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][371] ) );
  DFF \modmult_1/zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][370] ) );
  DFF \modmult_1/zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][369] ) );
  DFF \modmult_1/zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][368] ) );
  DFF \modmult_1/zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][367] ) );
  DFF \modmult_1/zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][366] ) );
  DFF \modmult_1/zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][365] ) );
  DFF \modmult_1/zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][364] ) );
  DFF \modmult_1/zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][363] ) );
  DFF \modmult_1/zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][362] ) );
  DFF \modmult_1/zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][361] ) );
  DFF \modmult_1/zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][360] ) );
  DFF \modmult_1/zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][359] ) );
  DFF \modmult_1/zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][358] ) );
  DFF \modmult_1/zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][357] ) );
  DFF \modmult_1/zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][356] ) );
  DFF \modmult_1/zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][355] ) );
  DFF \modmult_1/zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][354] ) );
  DFF \modmult_1/zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][353] ) );
  DFF \modmult_1/zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][352] ) );
  DFF \modmult_1/zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][351] ) );
  DFF \modmult_1/zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][350] ) );
  DFF \modmult_1/zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][349] ) );
  DFF \modmult_1/zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][348] ) );
  DFF \modmult_1/zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][347] ) );
  DFF \modmult_1/zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][346] ) );
  DFF \modmult_1/zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][345] ) );
  DFF \modmult_1/zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][344] ) );
  DFF \modmult_1/zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][343] ) );
  DFF \modmult_1/zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][342] ) );
  DFF \modmult_1/zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][341] ) );
  DFF \modmult_1/zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][340] ) );
  DFF \modmult_1/zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][339] ) );
  DFF \modmult_1/zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][338] ) );
  DFF \modmult_1/zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][337] ) );
  DFF \modmult_1/zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][336] ) );
  DFF \modmult_1/zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][335] ) );
  DFF \modmult_1/zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][334] ) );
  DFF \modmult_1/zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][333] ) );
  DFF \modmult_1/zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][332] ) );
  DFF \modmult_1/zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][331] ) );
  DFF \modmult_1/zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][330] ) );
  DFF \modmult_1/zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][329] ) );
  DFF \modmult_1/zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][328] ) );
  DFF \modmult_1/zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][327] ) );
  DFF \modmult_1/zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][326] ) );
  DFF \modmult_1/zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][325] ) );
  DFF \modmult_1/zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][324] ) );
  DFF \modmult_1/zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][323] ) );
  DFF \modmult_1/zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][322] ) );
  DFF \modmult_1/zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][321] ) );
  DFF \modmult_1/zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][320] ) );
  DFF \modmult_1/zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][319] ) );
  DFF \modmult_1/zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][318] ) );
  DFF \modmult_1/zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][317] ) );
  DFF \modmult_1/zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][316] ) );
  DFF \modmult_1/zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][315] ) );
  DFF \modmult_1/zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][314] ) );
  DFF \modmult_1/zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][313] ) );
  DFF \modmult_1/zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][312] ) );
  DFF \modmult_1/zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][311] ) );
  DFF \modmult_1/zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][310] ) );
  DFF \modmult_1/zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][309] ) );
  DFF \modmult_1/zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][308] ) );
  DFF \modmult_1/zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][307] ) );
  DFF \modmult_1/zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][306] ) );
  DFF \modmult_1/zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][305] ) );
  DFF \modmult_1/zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][304] ) );
  DFF \modmult_1/zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][303] ) );
  DFF \modmult_1/zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][302] ) );
  DFF \modmult_1/zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][301] ) );
  DFF \modmult_1/zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][300] ) );
  DFF \modmult_1/zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][299] ) );
  DFF \modmult_1/zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][298] ) );
  DFF \modmult_1/zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][297] ) );
  DFF \modmult_1/zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][296] ) );
  DFF \modmult_1/zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][295] ) );
  DFF \modmult_1/zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][294] ) );
  DFF \modmult_1/zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][293] ) );
  DFF \modmult_1/zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][292] ) );
  DFF \modmult_1/zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][291] ) );
  DFF \modmult_1/zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][290] ) );
  DFF \modmult_1/zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][289] ) );
  DFF \modmult_1/zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][288] ) );
  DFF \modmult_1/zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][287] ) );
  DFF \modmult_1/zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][286] ) );
  DFF \modmult_1/zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][285] ) );
  DFF \modmult_1/zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][284] ) );
  DFF \modmult_1/zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][283] ) );
  DFF \modmult_1/zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][282] ) );
  DFF \modmult_1/zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][281] ) );
  DFF \modmult_1/zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][280] ) );
  DFF \modmult_1/zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][279] ) );
  DFF \modmult_1/zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][278] ) );
  DFF \modmult_1/zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][277] ) );
  DFF \modmult_1/zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][276] ) );
  DFF \modmult_1/zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][275] ) );
  DFF \modmult_1/zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][274] ) );
  DFF \modmult_1/zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][273] ) );
  DFF \modmult_1/zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][272] ) );
  DFF \modmult_1/zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][271] ) );
  DFF \modmult_1/zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][270] ) );
  DFF \modmult_1/zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][269] ) );
  DFF \modmult_1/zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][268] ) );
  DFF \modmult_1/zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][267] ) );
  DFF \modmult_1/zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][266] ) );
  DFF \modmult_1/zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][265] ) );
  DFF \modmult_1/zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][264] ) );
  DFF \modmult_1/zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][263] ) );
  DFF \modmult_1/zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][262] ) );
  DFF \modmult_1/zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][261] ) );
  DFF \modmult_1/zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][260] ) );
  DFF \modmult_1/zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][259] ) );
  DFF \modmult_1/zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][258] ) );
  DFF \modmult_1/zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][257] ) );
  DFF \modmult_1/zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][256] ) );
  DFF \modmult_1/zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][255] ) );
  DFF \modmult_1/zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][254] ) );
  DFF \modmult_1/zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][253] ) );
  DFF \modmult_1/zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][252] ) );
  DFF \modmult_1/zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][251] ) );
  DFF \modmult_1/zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][250] ) );
  DFF \modmult_1/zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][249] ) );
  DFF \modmult_1/zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][248] ) );
  DFF \modmult_1/zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][247] ) );
  DFF \modmult_1/zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][246] ) );
  DFF \modmult_1/zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][245] ) );
  DFF \modmult_1/zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][244] ) );
  DFF \modmult_1/zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][243] ) );
  DFF \modmult_1/zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][242] ) );
  DFF \modmult_1/zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][241] ) );
  DFF \modmult_1/zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][240] ) );
  DFF \modmult_1/zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][239] ) );
  DFF \modmult_1/zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][238] ) );
  DFF \modmult_1/zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][237] ) );
  DFF \modmult_1/zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][236] ) );
  DFF \modmult_1/zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][235] ) );
  DFF \modmult_1/zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][234] ) );
  DFF \modmult_1/zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][233] ) );
  DFF \modmult_1/zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][232] ) );
  DFF \modmult_1/zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][231] ) );
  DFF \modmult_1/zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][230] ) );
  DFF \modmult_1/zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][229] ) );
  DFF \modmult_1/zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][228] ) );
  DFF \modmult_1/zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][227] ) );
  DFF \modmult_1/zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][226] ) );
  DFF \modmult_1/zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][225] ) );
  DFF \modmult_1/zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][224] ) );
  DFF \modmult_1/zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][223] ) );
  DFF \modmult_1/zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][222] ) );
  DFF \modmult_1/zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][221] ) );
  DFF \modmult_1/zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][220] ) );
  DFF \modmult_1/zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][219] ) );
  DFF \modmult_1/zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][218] ) );
  DFF \modmult_1/zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][217] ) );
  DFF \modmult_1/zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][216] ) );
  DFF \modmult_1/zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][215] ) );
  DFF \modmult_1/zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][214] ) );
  DFF \modmult_1/zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][213] ) );
  DFF \modmult_1/zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][212] ) );
  DFF \modmult_1/zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][211] ) );
  DFF \modmult_1/zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][210] ) );
  DFF \modmult_1/zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][209] ) );
  DFF \modmult_1/zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][208] ) );
  DFF \modmult_1/zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][207] ) );
  DFF \modmult_1/zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][206] ) );
  DFF \modmult_1/zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][205] ) );
  DFF \modmult_1/zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][204] ) );
  DFF \modmult_1/zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][203] ) );
  DFF \modmult_1/zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][202] ) );
  DFF \modmult_1/zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][201] ) );
  DFF \modmult_1/zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][200] ) );
  DFF \modmult_1/zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][199] ) );
  DFF \modmult_1/zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][198] ) );
  DFF \modmult_1/zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][197] ) );
  DFF \modmult_1/zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][196] ) );
  DFF \modmult_1/zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][195] ) );
  DFF \modmult_1/zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][194] ) );
  DFF \modmult_1/zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][193] ) );
  DFF \modmult_1/zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][192] ) );
  DFF \modmult_1/zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][191] ) );
  DFF \modmult_1/zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][190] ) );
  DFF \modmult_1/zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][189] ) );
  DFF \modmult_1/zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][188] ) );
  DFF \modmult_1/zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][187] ) );
  DFF \modmult_1/zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][186] ) );
  DFF \modmult_1/zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][185] ) );
  DFF \modmult_1/zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][184] ) );
  DFF \modmult_1/zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][183] ) );
  DFF \modmult_1/zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][182] ) );
  DFF \modmult_1/zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][181] ) );
  DFF \modmult_1/zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][180] ) );
  DFF \modmult_1/zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][179] ) );
  DFF \modmult_1/zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][178] ) );
  DFF \modmult_1/zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][177] ) );
  DFF \modmult_1/zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][176] ) );
  DFF \modmult_1/zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][175] ) );
  DFF \modmult_1/zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][174] ) );
  DFF \modmult_1/zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][173] ) );
  DFF \modmult_1/zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][172] ) );
  DFF \modmult_1/zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][171] ) );
  DFF \modmult_1/zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][170] ) );
  DFF \modmult_1/zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][169] ) );
  DFF \modmult_1/zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][168] ) );
  DFF \modmult_1/zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][167] ) );
  DFF \modmult_1/zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][166] ) );
  DFF \modmult_1/zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][165] ) );
  DFF \modmult_1/zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][164] ) );
  DFF \modmult_1/zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][163] ) );
  DFF \modmult_1/zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][162] ) );
  DFF \modmult_1/zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][161] ) );
  DFF \modmult_1/zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][160] ) );
  DFF \modmult_1/zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][159] ) );
  DFF \modmult_1/zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][158] ) );
  DFF \modmult_1/zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][157] ) );
  DFF \modmult_1/zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][156] ) );
  DFF \modmult_1/zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][155] ) );
  DFF \modmult_1/zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][154] ) );
  DFF \modmult_1/zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][153] ) );
  DFF \modmult_1/zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][152] ) );
  DFF \modmult_1/zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][151] ) );
  DFF \modmult_1/zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][150] ) );
  DFF \modmult_1/zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][149] ) );
  DFF \modmult_1/zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][148] ) );
  DFF \modmult_1/zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][147] ) );
  DFF \modmult_1/zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][146] ) );
  DFF \modmult_1/zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][145] ) );
  DFF \modmult_1/zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][144] ) );
  DFF \modmult_1/zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][143] ) );
  DFF \modmult_1/zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][142] ) );
  DFF \modmult_1/zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][141] ) );
  DFF \modmult_1/zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][140] ) );
  DFF \modmult_1/zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][139] ) );
  DFF \modmult_1/zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][138] ) );
  DFF \modmult_1/zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][137] ) );
  DFF \modmult_1/zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][136] ) );
  DFF \modmult_1/zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][135] ) );
  DFF \modmult_1/zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][134] ) );
  DFF \modmult_1/zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][133] ) );
  DFF \modmult_1/zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][132] ) );
  DFF \modmult_1/zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][131] ) );
  DFF \modmult_1/zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][130] ) );
  DFF \modmult_1/zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][129] ) );
  DFF \modmult_1/zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][128] ) );
  DFF \modmult_1/zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][127] ) );
  DFF \modmult_1/zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][126] ) );
  DFF \modmult_1/zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][125] ) );
  DFF \modmult_1/zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][124] ) );
  DFF \modmult_1/zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][123] ) );
  DFF \modmult_1/zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][122] ) );
  DFF \modmult_1/zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][121] ) );
  DFF \modmult_1/zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][120] ) );
  DFF \modmult_1/zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][119] ) );
  DFF \modmult_1/zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][118] ) );
  DFF \modmult_1/zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][117] ) );
  DFF \modmult_1/zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][116] ) );
  DFF \modmult_1/zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][115] ) );
  DFF \modmult_1/zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][114] ) );
  DFF \modmult_1/zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][113] ) );
  DFF \modmult_1/zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][112] ) );
  DFF \modmult_1/zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][111] ) );
  DFF \modmult_1/zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][110] ) );
  DFF \modmult_1/zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][109] ) );
  DFF \modmult_1/zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][108] ) );
  DFF \modmult_1/zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][107] ) );
  DFF \modmult_1/zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][106] ) );
  DFF \modmult_1/zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][105] ) );
  DFF \modmult_1/zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][104] ) );
  DFF \modmult_1/zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][103] ) );
  DFF \modmult_1/zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][102] ) );
  DFF \modmult_1/zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][101] ) );
  DFF \modmult_1/zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start_in[0]), 
        .I(1'b0), .Q(\modmult_1/zin[0][100] ) );
  DFF \modmult_1/zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][99] ) );
  DFF \modmult_1/zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][98] ) );
  DFF \modmult_1/zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][97] ) );
  DFF \modmult_1/zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][96] ) );
  DFF \modmult_1/zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][95] ) );
  DFF \modmult_1/zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][94] ) );
  DFF \modmult_1/zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][93] ) );
  DFF \modmult_1/zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][92] ) );
  DFF \modmult_1/zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][91] ) );
  DFF \modmult_1/zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][90] ) );
  DFF \modmult_1/zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][89] ) );
  DFF \modmult_1/zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][88] ) );
  DFF \modmult_1/zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][87] ) );
  DFF \modmult_1/zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][86] ) );
  DFF \modmult_1/zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][85] ) );
  DFF \modmult_1/zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][84] ) );
  DFF \modmult_1/zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][83] ) );
  DFF \modmult_1/zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][82] ) );
  DFF \modmult_1/zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][81] ) );
  DFF \modmult_1/zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][80] ) );
  DFF \modmult_1/zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][79] ) );
  DFF \modmult_1/zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][78] ) );
  DFF \modmult_1/zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][77] ) );
  DFF \modmult_1/zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][76] ) );
  DFF \modmult_1/zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][75] ) );
  DFF \modmult_1/zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][74] ) );
  DFF \modmult_1/zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][73] ) );
  DFF \modmult_1/zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][72] ) );
  DFF \modmult_1/zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][71] ) );
  DFF \modmult_1/zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][70] ) );
  DFF \modmult_1/zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][69] ) );
  DFF \modmult_1/zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][68] ) );
  DFF \modmult_1/zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][67] ) );
  DFF \modmult_1/zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][66] ) );
  DFF \modmult_1/zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][65] ) );
  DFF \modmult_1/zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][64] ) );
  DFF \modmult_1/zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][63] ) );
  DFF \modmult_1/zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][62] ) );
  DFF \modmult_1/zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][61] ) );
  DFF \modmult_1/zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][60] ) );
  DFF \modmult_1/zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][59] ) );
  DFF \modmult_1/zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][58] ) );
  DFF \modmult_1/zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][57] ) );
  DFF \modmult_1/zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][56] ) );
  DFF \modmult_1/zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][55] ) );
  DFF \modmult_1/zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][54] ) );
  DFF \modmult_1/zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][53] ) );
  DFF \modmult_1/zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][52] ) );
  DFF \modmult_1/zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][51] ) );
  DFF \modmult_1/zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][50] ) );
  DFF \modmult_1/zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][49] ) );
  DFF \modmult_1/zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][48] ) );
  DFF \modmult_1/zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][47] ) );
  DFF \modmult_1/zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][46] ) );
  DFF \modmult_1/zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][45] ) );
  DFF \modmult_1/zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][44] ) );
  DFF \modmult_1/zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][43] ) );
  DFF \modmult_1/zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][42] ) );
  DFF \modmult_1/zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][41] ) );
  DFF \modmult_1/zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][40] ) );
  DFF \modmult_1/zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][39] ) );
  DFF \modmult_1/zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][38] ) );
  DFF \modmult_1/zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][37] ) );
  DFF \modmult_1/zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][36] ) );
  DFF \modmult_1/zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][35] ) );
  DFF \modmult_1/zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][34] ) );
  DFF \modmult_1/zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][33] ) );
  DFF \modmult_1/zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][32] ) );
  DFF \modmult_1/zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][31] ) );
  DFF \modmult_1/zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][30] ) );
  DFF \modmult_1/zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][29] ) );
  DFF \modmult_1/zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][28] ) );
  DFF \modmult_1/zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][27] ) );
  DFF \modmult_1/zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][26] ) );
  DFF \modmult_1/zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][25] ) );
  DFF \modmult_1/zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][24] ) );
  DFF \modmult_1/zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][23] ) );
  DFF \modmult_1/zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][22] ) );
  DFF \modmult_1/zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][21] ) );
  DFF \modmult_1/zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][20] ) );
  DFF \modmult_1/zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][19] ) );
  DFF \modmult_1/zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][18] ) );
  DFF \modmult_1/zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][17] ) );
  DFF \modmult_1/zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][16] ) );
  DFF \modmult_1/zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][15] ) );
  DFF \modmult_1/zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][14] ) );
  DFF \modmult_1/zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][13] ) );
  DFF \modmult_1/zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][12] ) );
  DFF \modmult_1/zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][11] ) );
  DFF \modmult_1/zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][10] ) );
  DFF \modmult_1/zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][9] ) );
  DFF \modmult_1/zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][8] ) );
  DFF \modmult_1/zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][7] ) );
  DFF \modmult_1/zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][6] ) );
  DFF \modmult_1/zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][5] ) );
  DFF \modmult_1/zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][4] ) );
  DFF \modmult_1/zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][3] ) );
  DFF \modmult_1/zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][2] ) );
  DFF \modmult_1/zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][1] ) );
  DFF \modmult_1/zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start_in[0]), .I(
        1'b0), .Q(\modmult_1/zin[0][0] ) );
  DFF \modmult_1/xreg_reg[1023]  ( .D(\modmult_1/xin[1022] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1023]), .Q(\modmult_1/xin[1023] ) );
  DFF \modmult_1/xreg_reg[1022]  ( .D(\modmult_1/xin[1021] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1022]), .Q(\modmult_1/xin[1022] ) );
  DFF \modmult_1/xreg_reg[1021]  ( .D(\modmult_1/xin[1020] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1021]), .Q(\modmult_1/xin[1021] ) );
  DFF \modmult_1/xreg_reg[1020]  ( .D(\modmult_1/xin[1019] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1020]), .Q(\modmult_1/xin[1020] ) );
  DFF \modmult_1/xreg_reg[1019]  ( .D(\modmult_1/xin[1018] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1019]), .Q(\modmult_1/xin[1019] ) );
  DFF \modmult_1/xreg_reg[1018]  ( .D(\modmult_1/xin[1017] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1018]), .Q(\modmult_1/xin[1018] ) );
  DFF \modmult_1/xreg_reg[1017]  ( .D(\modmult_1/xin[1016] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1017]), .Q(\modmult_1/xin[1017] ) );
  DFF \modmult_1/xreg_reg[1016]  ( .D(\modmult_1/xin[1015] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1016]), .Q(\modmult_1/xin[1016] ) );
  DFF \modmult_1/xreg_reg[1015]  ( .D(\modmult_1/xin[1014] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1015]), .Q(\modmult_1/xin[1015] ) );
  DFF \modmult_1/xreg_reg[1014]  ( .D(\modmult_1/xin[1013] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1014]), .Q(\modmult_1/xin[1014] ) );
  DFF \modmult_1/xreg_reg[1013]  ( .D(\modmult_1/xin[1012] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1013]), .Q(\modmult_1/xin[1013] ) );
  DFF \modmult_1/xreg_reg[1012]  ( .D(\modmult_1/xin[1011] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1012]), .Q(\modmult_1/xin[1012] ) );
  DFF \modmult_1/xreg_reg[1011]  ( .D(\modmult_1/xin[1010] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1011]), .Q(\modmult_1/xin[1011] ) );
  DFF \modmult_1/xreg_reg[1010]  ( .D(\modmult_1/xin[1009] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1010]), .Q(\modmult_1/xin[1010] ) );
  DFF \modmult_1/xreg_reg[1009]  ( .D(\modmult_1/xin[1008] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1009]), .Q(\modmult_1/xin[1009] ) );
  DFF \modmult_1/xreg_reg[1008]  ( .D(\modmult_1/xin[1007] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1008]), .Q(\modmult_1/xin[1008] ) );
  DFF \modmult_1/xreg_reg[1007]  ( .D(\modmult_1/xin[1006] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1007]), .Q(\modmult_1/xin[1007] ) );
  DFF \modmult_1/xreg_reg[1006]  ( .D(\modmult_1/xin[1005] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1006]), .Q(\modmult_1/xin[1006] ) );
  DFF \modmult_1/xreg_reg[1005]  ( .D(\modmult_1/xin[1004] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1005]), .Q(\modmult_1/xin[1005] ) );
  DFF \modmult_1/xreg_reg[1004]  ( .D(\modmult_1/xin[1003] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1004]), .Q(\modmult_1/xin[1004] ) );
  DFF \modmult_1/xreg_reg[1003]  ( .D(\modmult_1/xin[1002] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1003]), .Q(\modmult_1/xin[1003] ) );
  DFF \modmult_1/xreg_reg[1002]  ( .D(\modmult_1/xin[1001] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1002]), .Q(\modmult_1/xin[1002] ) );
  DFF \modmult_1/xreg_reg[1001]  ( .D(\modmult_1/xin[1000] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1001]), .Q(\modmult_1/xin[1001] ) );
  DFF \modmult_1/xreg_reg[1000]  ( .D(\modmult_1/xin[999] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1000]), .Q(\modmult_1/xin[1000] ) );
  DFF \modmult_1/xreg_reg[999]  ( .D(\modmult_1/xin[998] ), .CLK(clk), .RST(
        start_in[0]), .I(c[999]), .Q(\modmult_1/xin[999] ) );
  DFF \modmult_1/xreg_reg[998]  ( .D(\modmult_1/xin[997] ), .CLK(clk), .RST(
        start_in[0]), .I(c[998]), .Q(\modmult_1/xin[998] ) );
  DFF \modmult_1/xreg_reg[997]  ( .D(\modmult_1/xin[996] ), .CLK(clk), .RST(
        start_in[0]), .I(c[997]), .Q(\modmult_1/xin[997] ) );
  DFF \modmult_1/xreg_reg[996]  ( .D(\modmult_1/xin[995] ), .CLK(clk), .RST(
        start_in[0]), .I(c[996]), .Q(\modmult_1/xin[996] ) );
  DFF \modmult_1/xreg_reg[995]  ( .D(\modmult_1/xin[994] ), .CLK(clk), .RST(
        start_in[0]), .I(c[995]), .Q(\modmult_1/xin[995] ) );
  DFF \modmult_1/xreg_reg[994]  ( .D(\modmult_1/xin[993] ), .CLK(clk), .RST(
        start_in[0]), .I(c[994]), .Q(\modmult_1/xin[994] ) );
  DFF \modmult_1/xreg_reg[993]  ( .D(\modmult_1/xin[992] ), .CLK(clk), .RST(
        start_in[0]), .I(c[993]), .Q(\modmult_1/xin[993] ) );
  DFF \modmult_1/xreg_reg[992]  ( .D(\modmult_1/xin[991] ), .CLK(clk), .RST(
        start_in[0]), .I(c[992]), .Q(\modmult_1/xin[992] ) );
  DFF \modmult_1/xreg_reg[991]  ( .D(\modmult_1/xin[990] ), .CLK(clk), .RST(
        start_in[0]), .I(c[991]), .Q(\modmult_1/xin[991] ) );
  DFF \modmult_1/xreg_reg[990]  ( .D(\modmult_1/xin[989] ), .CLK(clk), .RST(
        start_in[0]), .I(c[990]), .Q(\modmult_1/xin[990] ) );
  DFF \modmult_1/xreg_reg[989]  ( .D(\modmult_1/xin[988] ), .CLK(clk), .RST(
        start_in[0]), .I(c[989]), .Q(\modmult_1/xin[989] ) );
  DFF \modmult_1/xreg_reg[988]  ( .D(\modmult_1/xin[987] ), .CLK(clk), .RST(
        start_in[0]), .I(c[988]), .Q(\modmult_1/xin[988] ) );
  DFF \modmult_1/xreg_reg[987]  ( .D(\modmult_1/xin[986] ), .CLK(clk), .RST(
        start_in[0]), .I(c[987]), .Q(\modmult_1/xin[987] ) );
  DFF \modmult_1/xreg_reg[986]  ( .D(\modmult_1/xin[985] ), .CLK(clk), .RST(
        start_in[0]), .I(c[986]), .Q(\modmult_1/xin[986] ) );
  DFF \modmult_1/xreg_reg[985]  ( .D(\modmult_1/xin[984] ), .CLK(clk), .RST(
        start_in[0]), .I(c[985]), .Q(\modmult_1/xin[985] ) );
  DFF \modmult_1/xreg_reg[984]  ( .D(\modmult_1/xin[983] ), .CLK(clk), .RST(
        start_in[0]), .I(c[984]), .Q(\modmult_1/xin[984] ) );
  DFF \modmult_1/xreg_reg[983]  ( .D(\modmult_1/xin[982] ), .CLK(clk), .RST(
        start_in[0]), .I(c[983]), .Q(\modmult_1/xin[983] ) );
  DFF \modmult_1/xreg_reg[982]  ( .D(\modmult_1/xin[981] ), .CLK(clk), .RST(
        start_in[0]), .I(c[982]), .Q(\modmult_1/xin[982] ) );
  DFF \modmult_1/xreg_reg[981]  ( .D(\modmult_1/xin[980] ), .CLK(clk), .RST(
        start_in[0]), .I(c[981]), .Q(\modmult_1/xin[981] ) );
  DFF \modmult_1/xreg_reg[980]  ( .D(\modmult_1/xin[979] ), .CLK(clk), .RST(
        start_in[0]), .I(c[980]), .Q(\modmult_1/xin[980] ) );
  DFF \modmult_1/xreg_reg[979]  ( .D(\modmult_1/xin[978] ), .CLK(clk), .RST(
        start_in[0]), .I(c[979]), .Q(\modmult_1/xin[979] ) );
  DFF \modmult_1/xreg_reg[978]  ( .D(\modmult_1/xin[977] ), .CLK(clk), .RST(
        start_in[0]), .I(c[978]), .Q(\modmult_1/xin[978] ) );
  DFF \modmult_1/xreg_reg[977]  ( .D(\modmult_1/xin[976] ), .CLK(clk), .RST(
        start_in[0]), .I(c[977]), .Q(\modmult_1/xin[977] ) );
  DFF \modmult_1/xreg_reg[976]  ( .D(\modmult_1/xin[975] ), .CLK(clk), .RST(
        start_in[0]), .I(c[976]), .Q(\modmult_1/xin[976] ) );
  DFF \modmult_1/xreg_reg[975]  ( .D(\modmult_1/xin[974] ), .CLK(clk), .RST(
        start_in[0]), .I(c[975]), .Q(\modmult_1/xin[975] ) );
  DFF \modmult_1/xreg_reg[974]  ( .D(\modmult_1/xin[973] ), .CLK(clk), .RST(
        start_in[0]), .I(c[974]), .Q(\modmult_1/xin[974] ) );
  DFF \modmult_1/xreg_reg[973]  ( .D(\modmult_1/xin[972] ), .CLK(clk), .RST(
        start_in[0]), .I(c[973]), .Q(\modmult_1/xin[973] ) );
  DFF \modmult_1/xreg_reg[972]  ( .D(\modmult_1/xin[971] ), .CLK(clk), .RST(
        start_in[0]), .I(c[972]), .Q(\modmult_1/xin[972] ) );
  DFF \modmult_1/xreg_reg[971]  ( .D(\modmult_1/xin[970] ), .CLK(clk), .RST(
        start_in[0]), .I(c[971]), .Q(\modmult_1/xin[971] ) );
  DFF \modmult_1/xreg_reg[970]  ( .D(\modmult_1/xin[969] ), .CLK(clk), .RST(
        start_in[0]), .I(c[970]), .Q(\modmult_1/xin[970] ) );
  DFF \modmult_1/xreg_reg[969]  ( .D(\modmult_1/xin[968] ), .CLK(clk), .RST(
        start_in[0]), .I(c[969]), .Q(\modmult_1/xin[969] ) );
  DFF \modmult_1/xreg_reg[968]  ( .D(\modmult_1/xin[967] ), .CLK(clk), .RST(
        start_in[0]), .I(c[968]), .Q(\modmult_1/xin[968] ) );
  DFF \modmult_1/xreg_reg[967]  ( .D(\modmult_1/xin[966] ), .CLK(clk), .RST(
        start_in[0]), .I(c[967]), .Q(\modmult_1/xin[967] ) );
  DFF \modmult_1/xreg_reg[966]  ( .D(\modmult_1/xin[965] ), .CLK(clk), .RST(
        start_in[0]), .I(c[966]), .Q(\modmult_1/xin[966] ) );
  DFF \modmult_1/xreg_reg[965]  ( .D(\modmult_1/xin[964] ), .CLK(clk), .RST(
        start_in[0]), .I(c[965]), .Q(\modmult_1/xin[965] ) );
  DFF \modmult_1/xreg_reg[964]  ( .D(\modmult_1/xin[963] ), .CLK(clk), .RST(
        start_in[0]), .I(c[964]), .Q(\modmult_1/xin[964] ) );
  DFF \modmult_1/xreg_reg[963]  ( .D(\modmult_1/xin[962] ), .CLK(clk), .RST(
        start_in[0]), .I(c[963]), .Q(\modmult_1/xin[963] ) );
  DFF \modmult_1/xreg_reg[962]  ( .D(\modmult_1/xin[961] ), .CLK(clk), .RST(
        start_in[0]), .I(c[962]), .Q(\modmult_1/xin[962] ) );
  DFF \modmult_1/xreg_reg[961]  ( .D(\modmult_1/xin[960] ), .CLK(clk), .RST(
        start_in[0]), .I(c[961]), .Q(\modmult_1/xin[961] ) );
  DFF \modmult_1/xreg_reg[960]  ( .D(\modmult_1/xin[959] ), .CLK(clk), .RST(
        start_in[0]), .I(c[960]), .Q(\modmult_1/xin[960] ) );
  DFF \modmult_1/xreg_reg[959]  ( .D(\modmult_1/xin[958] ), .CLK(clk), .RST(
        start_in[0]), .I(c[959]), .Q(\modmult_1/xin[959] ) );
  DFF \modmult_1/xreg_reg[958]  ( .D(\modmult_1/xin[957] ), .CLK(clk), .RST(
        start_in[0]), .I(c[958]), .Q(\modmult_1/xin[958] ) );
  DFF \modmult_1/xreg_reg[957]  ( .D(\modmult_1/xin[956] ), .CLK(clk), .RST(
        start_in[0]), .I(c[957]), .Q(\modmult_1/xin[957] ) );
  DFF \modmult_1/xreg_reg[956]  ( .D(\modmult_1/xin[955] ), .CLK(clk), .RST(
        start_in[0]), .I(c[956]), .Q(\modmult_1/xin[956] ) );
  DFF \modmult_1/xreg_reg[955]  ( .D(\modmult_1/xin[954] ), .CLK(clk), .RST(
        start_in[0]), .I(c[955]), .Q(\modmult_1/xin[955] ) );
  DFF \modmult_1/xreg_reg[954]  ( .D(\modmult_1/xin[953] ), .CLK(clk), .RST(
        start_in[0]), .I(c[954]), .Q(\modmult_1/xin[954] ) );
  DFF \modmult_1/xreg_reg[953]  ( .D(\modmult_1/xin[952] ), .CLK(clk), .RST(
        start_in[0]), .I(c[953]), .Q(\modmult_1/xin[953] ) );
  DFF \modmult_1/xreg_reg[952]  ( .D(\modmult_1/xin[951] ), .CLK(clk), .RST(
        start_in[0]), .I(c[952]), .Q(\modmult_1/xin[952] ) );
  DFF \modmult_1/xreg_reg[951]  ( .D(\modmult_1/xin[950] ), .CLK(clk), .RST(
        start_in[0]), .I(c[951]), .Q(\modmult_1/xin[951] ) );
  DFF \modmult_1/xreg_reg[950]  ( .D(\modmult_1/xin[949] ), .CLK(clk), .RST(
        start_in[0]), .I(c[950]), .Q(\modmult_1/xin[950] ) );
  DFF \modmult_1/xreg_reg[949]  ( .D(\modmult_1/xin[948] ), .CLK(clk), .RST(
        start_in[0]), .I(c[949]), .Q(\modmult_1/xin[949] ) );
  DFF \modmult_1/xreg_reg[948]  ( .D(\modmult_1/xin[947] ), .CLK(clk), .RST(
        start_in[0]), .I(c[948]), .Q(\modmult_1/xin[948] ) );
  DFF \modmult_1/xreg_reg[947]  ( .D(\modmult_1/xin[946] ), .CLK(clk), .RST(
        start_in[0]), .I(c[947]), .Q(\modmult_1/xin[947] ) );
  DFF \modmult_1/xreg_reg[946]  ( .D(\modmult_1/xin[945] ), .CLK(clk), .RST(
        start_in[0]), .I(c[946]), .Q(\modmult_1/xin[946] ) );
  DFF \modmult_1/xreg_reg[945]  ( .D(\modmult_1/xin[944] ), .CLK(clk), .RST(
        start_in[0]), .I(c[945]), .Q(\modmult_1/xin[945] ) );
  DFF \modmult_1/xreg_reg[944]  ( .D(\modmult_1/xin[943] ), .CLK(clk), .RST(
        start_in[0]), .I(c[944]), .Q(\modmult_1/xin[944] ) );
  DFF \modmult_1/xreg_reg[943]  ( .D(\modmult_1/xin[942] ), .CLK(clk), .RST(
        start_in[0]), .I(c[943]), .Q(\modmult_1/xin[943] ) );
  DFF \modmult_1/xreg_reg[942]  ( .D(\modmult_1/xin[941] ), .CLK(clk), .RST(
        start_in[0]), .I(c[942]), .Q(\modmult_1/xin[942] ) );
  DFF \modmult_1/xreg_reg[941]  ( .D(\modmult_1/xin[940] ), .CLK(clk), .RST(
        start_in[0]), .I(c[941]), .Q(\modmult_1/xin[941] ) );
  DFF \modmult_1/xreg_reg[940]  ( .D(\modmult_1/xin[939] ), .CLK(clk), .RST(
        start_in[0]), .I(c[940]), .Q(\modmult_1/xin[940] ) );
  DFF \modmult_1/xreg_reg[939]  ( .D(\modmult_1/xin[938] ), .CLK(clk), .RST(
        start_in[0]), .I(c[939]), .Q(\modmult_1/xin[939] ) );
  DFF \modmult_1/xreg_reg[938]  ( .D(\modmult_1/xin[937] ), .CLK(clk), .RST(
        start_in[0]), .I(c[938]), .Q(\modmult_1/xin[938] ) );
  DFF \modmult_1/xreg_reg[937]  ( .D(\modmult_1/xin[936] ), .CLK(clk), .RST(
        start_in[0]), .I(c[937]), .Q(\modmult_1/xin[937] ) );
  DFF \modmult_1/xreg_reg[936]  ( .D(\modmult_1/xin[935] ), .CLK(clk), .RST(
        start_in[0]), .I(c[936]), .Q(\modmult_1/xin[936] ) );
  DFF \modmult_1/xreg_reg[935]  ( .D(\modmult_1/xin[934] ), .CLK(clk), .RST(
        start_in[0]), .I(c[935]), .Q(\modmult_1/xin[935] ) );
  DFF \modmult_1/xreg_reg[934]  ( .D(\modmult_1/xin[933] ), .CLK(clk), .RST(
        start_in[0]), .I(c[934]), .Q(\modmult_1/xin[934] ) );
  DFF \modmult_1/xreg_reg[933]  ( .D(\modmult_1/xin[932] ), .CLK(clk), .RST(
        start_in[0]), .I(c[933]), .Q(\modmult_1/xin[933] ) );
  DFF \modmult_1/xreg_reg[932]  ( .D(\modmult_1/xin[931] ), .CLK(clk), .RST(
        start_in[0]), .I(c[932]), .Q(\modmult_1/xin[932] ) );
  DFF \modmult_1/xreg_reg[931]  ( .D(\modmult_1/xin[930] ), .CLK(clk), .RST(
        start_in[0]), .I(c[931]), .Q(\modmult_1/xin[931] ) );
  DFF \modmult_1/xreg_reg[930]  ( .D(\modmult_1/xin[929] ), .CLK(clk), .RST(
        start_in[0]), .I(c[930]), .Q(\modmult_1/xin[930] ) );
  DFF \modmult_1/xreg_reg[929]  ( .D(\modmult_1/xin[928] ), .CLK(clk), .RST(
        start_in[0]), .I(c[929]), .Q(\modmult_1/xin[929] ) );
  DFF \modmult_1/xreg_reg[928]  ( .D(\modmult_1/xin[927] ), .CLK(clk), .RST(
        start_in[0]), .I(c[928]), .Q(\modmult_1/xin[928] ) );
  DFF \modmult_1/xreg_reg[927]  ( .D(\modmult_1/xin[926] ), .CLK(clk), .RST(
        start_in[0]), .I(c[927]), .Q(\modmult_1/xin[927] ) );
  DFF \modmult_1/xreg_reg[926]  ( .D(\modmult_1/xin[925] ), .CLK(clk), .RST(
        start_in[0]), .I(c[926]), .Q(\modmult_1/xin[926] ) );
  DFF \modmult_1/xreg_reg[925]  ( .D(\modmult_1/xin[924] ), .CLK(clk), .RST(
        start_in[0]), .I(c[925]), .Q(\modmult_1/xin[925] ) );
  DFF \modmult_1/xreg_reg[924]  ( .D(\modmult_1/xin[923] ), .CLK(clk), .RST(
        start_in[0]), .I(c[924]), .Q(\modmult_1/xin[924] ) );
  DFF \modmult_1/xreg_reg[923]  ( .D(\modmult_1/xin[922] ), .CLK(clk), .RST(
        start_in[0]), .I(c[923]), .Q(\modmult_1/xin[923] ) );
  DFF \modmult_1/xreg_reg[922]  ( .D(\modmult_1/xin[921] ), .CLK(clk), .RST(
        start_in[0]), .I(c[922]), .Q(\modmult_1/xin[922] ) );
  DFF \modmult_1/xreg_reg[921]  ( .D(\modmult_1/xin[920] ), .CLK(clk), .RST(
        start_in[0]), .I(c[921]), .Q(\modmult_1/xin[921] ) );
  DFF \modmult_1/xreg_reg[920]  ( .D(\modmult_1/xin[919] ), .CLK(clk), .RST(
        start_in[0]), .I(c[920]), .Q(\modmult_1/xin[920] ) );
  DFF \modmult_1/xreg_reg[919]  ( .D(\modmult_1/xin[918] ), .CLK(clk), .RST(
        start_in[0]), .I(c[919]), .Q(\modmult_1/xin[919] ) );
  DFF \modmult_1/xreg_reg[918]  ( .D(\modmult_1/xin[917] ), .CLK(clk), .RST(
        start_in[0]), .I(c[918]), .Q(\modmult_1/xin[918] ) );
  DFF \modmult_1/xreg_reg[917]  ( .D(\modmult_1/xin[916] ), .CLK(clk), .RST(
        start_in[0]), .I(c[917]), .Q(\modmult_1/xin[917] ) );
  DFF \modmult_1/xreg_reg[916]  ( .D(\modmult_1/xin[915] ), .CLK(clk), .RST(
        start_in[0]), .I(c[916]), .Q(\modmult_1/xin[916] ) );
  DFF \modmult_1/xreg_reg[915]  ( .D(\modmult_1/xin[914] ), .CLK(clk), .RST(
        start_in[0]), .I(c[915]), .Q(\modmult_1/xin[915] ) );
  DFF \modmult_1/xreg_reg[914]  ( .D(\modmult_1/xin[913] ), .CLK(clk), .RST(
        start_in[0]), .I(c[914]), .Q(\modmult_1/xin[914] ) );
  DFF \modmult_1/xreg_reg[913]  ( .D(\modmult_1/xin[912] ), .CLK(clk), .RST(
        start_in[0]), .I(c[913]), .Q(\modmult_1/xin[913] ) );
  DFF \modmult_1/xreg_reg[912]  ( .D(\modmult_1/xin[911] ), .CLK(clk), .RST(
        start_in[0]), .I(c[912]), .Q(\modmult_1/xin[912] ) );
  DFF \modmult_1/xreg_reg[911]  ( .D(\modmult_1/xin[910] ), .CLK(clk), .RST(
        start_in[0]), .I(c[911]), .Q(\modmult_1/xin[911] ) );
  DFF \modmult_1/xreg_reg[910]  ( .D(\modmult_1/xin[909] ), .CLK(clk), .RST(
        start_in[0]), .I(c[910]), .Q(\modmult_1/xin[910] ) );
  DFF \modmult_1/xreg_reg[909]  ( .D(\modmult_1/xin[908] ), .CLK(clk), .RST(
        start_in[0]), .I(c[909]), .Q(\modmult_1/xin[909] ) );
  DFF \modmult_1/xreg_reg[908]  ( .D(\modmult_1/xin[907] ), .CLK(clk), .RST(
        start_in[0]), .I(c[908]), .Q(\modmult_1/xin[908] ) );
  DFF \modmult_1/xreg_reg[907]  ( .D(\modmult_1/xin[906] ), .CLK(clk), .RST(
        start_in[0]), .I(c[907]), .Q(\modmult_1/xin[907] ) );
  DFF \modmult_1/xreg_reg[906]  ( .D(\modmult_1/xin[905] ), .CLK(clk), .RST(
        start_in[0]), .I(c[906]), .Q(\modmult_1/xin[906] ) );
  DFF \modmult_1/xreg_reg[905]  ( .D(\modmult_1/xin[904] ), .CLK(clk), .RST(
        start_in[0]), .I(c[905]), .Q(\modmult_1/xin[905] ) );
  DFF \modmult_1/xreg_reg[904]  ( .D(\modmult_1/xin[903] ), .CLK(clk), .RST(
        start_in[0]), .I(c[904]), .Q(\modmult_1/xin[904] ) );
  DFF \modmult_1/xreg_reg[903]  ( .D(\modmult_1/xin[902] ), .CLK(clk), .RST(
        start_in[0]), .I(c[903]), .Q(\modmult_1/xin[903] ) );
  DFF \modmult_1/xreg_reg[902]  ( .D(\modmult_1/xin[901] ), .CLK(clk), .RST(
        start_in[0]), .I(c[902]), .Q(\modmult_1/xin[902] ) );
  DFF \modmult_1/xreg_reg[901]  ( .D(\modmult_1/xin[900] ), .CLK(clk), .RST(
        start_in[0]), .I(c[901]), .Q(\modmult_1/xin[901] ) );
  DFF \modmult_1/xreg_reg[900]  ( .D(\modmult_1/xin[899] ), .CLK(clk), .RST(
        start_in[0]), .I(c[900]), .Q(\modmult_1/xin[900] ) );
  DFF \modmult_1/xreg_reg[899]  ( .D(\modmult_1/xin[898] ), .CLK(clk), .RST(
        start_in[0]), .I(c[899]), .Q(\modmult_1/xin[899] ) );
  DFF \modmult_1/xreg_reg[898]  ( .D(\modmult_1/xin[897] ), .CLK(clk), .RST(
        start_in[0]), .I(c[898]), .Q(\modmult_1/xin[898] ) );
  DFF \modmult_1/xreg_reg[897]  ( .D(\modmult_1/xin[896] ), .CLK(clk), .RST(
        start_in[0]), .I(c[897]), .Q(\modmult_1/xin[897] ) );
  DFF \modmult_1/xreg_reg[896]  ( .D(\modmult_1/xin[895] ), .CLK(clk), .RST(
        start_in[0]), .I(c[896]), .Q(\modmult_1/xin[896] ) );
  DFF \modmult_1/xreg_reg[895]  ( .D(\modmult_1/xin[894] ), .CLK(clk), .RST(
        start_in[0]), .I(c[895]), .Q(\modmult_1/xin[895] ) );
  DFF \modmult_1/xreg_reg[894]  ( .D(\modmult_1/xin[893] ), .CLK(clk), .RST(
        start_in[0]), .I(c[894]), .Q(\modmult_1/xin[894] ) );
  DFF \modmult_1/xreg_reg[893]  ( .D(\modmult_1/xin[892] ), .CLK(clk), .RST(
        start_in[0]), .I(c[893]), .Q(\modmult_1/xin[893] ) );
  DFF \modmult_1/xreg_reg[892]  ( .D(\modmult_1/xin[891] ), .CLK(clk), .RST(
        start_in[0]), .I(c[892]), .Q(\modmult_1/xin[892] ) );
  DFF \modmult_1/xreg_reg[891]  ( .D(\modmult_1/xin[890] ), .CLK(clk), .RST(
        start_in[0]), .I(c[891]), .Q(\modmult_1/xin[891] ) );
  DFF \modmult_1/xreg_reg[890]  ( .D(\modmult_1/xin[889] ), .CLK(clk), .RST(
        start_in[0]), .I(c[890]), .Q(\modmult_1/xin[890] ) );
  DFF \modmult_1/xreg_reg[889]  ( .D(\modmult_1/xin[888] ), .CLK(clk), .RST(
        start_in[0]), .I(c[889]), .Q(\modmult_1/xin[889] ) );
  DFF \modmult_1/xreg_reg[888]  ( .D(\modmult_1/xin[887] ), .CLK(clk), .RST(
        start_in[0]), .I(c[888]), .Q(\modmult_1/xin[888] ) );
  DFF \modmult_1/xreg_reg[887]  ( .D(\modmult_1/xin[886] ), .CLK(clk), .RST(
        start_in[0]), .I(c[887]), .Q(\modmult_1/xin[887] ) );
  DFF \modmult_1/xreg_reg[886]  ( .D(\modmult_1/xin[885] ), .CLK(clk), .RST(
        start_in[0]), .I(c[886]), .Q(\modmult_1/xin[886] ) );
  DFF \modmult_1/xreg_reg[885]  ( .D(\modmult_1/xin[884] ), .CLK(clk), .RST(
        start_in[0]), .I(c[885]), .Q(\modmult_1/xin[885] ) );
  DFF \modmult_1/xreg_reg[884]  ( .D(\modmult_1/xin[883] ), .CLK(clk), .RST(
        start_in[0]), .I(c[884]), .Q(\modmult_1/xin[884] ) );
  DFF \modmult_1/xreg_reg[883]  ( .D(\modmult_1/xin[882] ), .CLK(clk), .RST(
        start_in[0]), .I(c[883]), .Q(\modmult_1/xin[883] ) );
  DFF \modmult_1/xreg_reg[882]  ( .D(\modmult_1/xin[881] ), .CLK(clk), .RST(
        start_in[0]), .I(c[882]), .Q(\modmult_1/xin[882] ) );
  DFF \modmult_1/xreg_reg[881]  ( .D(\modmult_1/xin[880] ), .CLK(clk), .RST(
        start_in[0]), .I(c[881]), .Q(\modmult_1/xin[881] ) );
  DFF \modmult_1/xreg_reg[880]  ( .D(\modmult_1/xin[879] ), .CLK(clk), .RST(
        start_in[0]), .I(c[880]), .Q(\modmult_1/xin[880] ) );
  DFF \modmult_1/xreg_reg[879]  ( .D(\modmult_1/xin[878] ), .CLK(clk), .RST(
        start_in[0]), .I(c[879]), .Q(\modmult_1/xin[879] ) );
  DFF \modmult_1/xreg_reg[878]  ( .D(\modmult_1/xin[877] ), .CLK(clk), .RST(
        start_in[0]), .I(c[878]), .Q(\modmult_1/xin[878] ) );
  DFF \modmult_1/xreg_reg[877]  ( .D(\modmult_1/xin[876] ), .CLK(clk), .RST(
        start_in[0]), .I(c[877]), .Q(\modmult_1/xin[877] ) );
  DFF \modmult_1/xreg_reg[876]  ( .D(\modmult_1/xin[875] ), .CLK(clk), .RST(
        start_in[0]), .I(c[876]), .Q(\modmult_1/xin[876] ) );
  DFF \modmult_1/xreg_reg[875]  ( .D(\modmult_1/xin[874] ), .CLK(clk), .RST(
        start_in[0]), .I(c[875]), .Q(\modmult_1/xin[875] ) );
  DFF \modmult_1/xreg_reg[874]  ( .D(\modmult_1/xin[873] ), .CLK(clk), .RST(
        start_in[0]), .I(c[874]), .Q(\modmult_1/xin[874] ) );
  DFF \modmult_1/xreg_reg[873]  ( .D(\modmult_1/xin[872] ), .CLK(clk), .RST(
        start_in[0]), .I(c[873]), .Q(\modmult_1/xin[873] ) );
  DFF \modmult_1/xreg_reg[872]  ( .D(\modmult_1/xin[871] ), .CLK(clk), .RST(
        start_in[0]), .I(c[872]), .Q(\modmult_1/xin[872] ) );
  DFF \modmult_1/xreg_reg[871]  ( .D(\modmult_1/xin[870] ), .CLK(clk), .RST(
        start_in[0]), .I(c[871]), .Q(\modmult_1/xin[871] ) );
  DFF \modmult_1/xreg_reg[870]  ( .D(\modmult_1/xin[869] ), .CLK(clk), .RST(
        start_in[0]), .I(c[870]), .Q(\modmult_1/xin[870] ) );
  DFF \modmult_1/xreg_reg[869]  ( .D(\modmult_1/xin[868] ), .CLK(clk), .RST(
        start_in[0]), .I(c[869]), .Q(\modmult_1/xin[869] ) );
  DFF \modmult_1/xreg_reg[868]  ( .D(\modmult_1/xin[867] ), .CLK(clk), .RST(
        start_in[0]), .I(c[868]), .Q(\modmult_1/xin[868] ) );
  DFF \modmult_1/xreg_reg[867]  ( .D(\modmult_1/xin[866] ), .CLK(clk), .RST(
        start_in[0]), .I(c[867]), .Q(\modmult_1/xin[867] ) );
  DFF \modmult_1/xreg_reg[866]  ( .D(\modmult_1/xin[865] ), .CLK(clk), .RST(
        start_in[0]), .I(c[866]), .Q(\modmult_1/xin[866] ) );
  DFF \modmult_1/xreg_reg[865]  ( .D(\modmult_1/xin[864] ), .CLK(clk), .RST(
        start_in[0]), .I(c[865]), .Q(\modmult_1/xin[865] ) );
  DFF \modmult_1/xreg_reg[864]  ( .D(\modmult_1/xin[863] ), .CLK(clk), .RST(
        start_in[0]), .I(c[864]), .Q(\modmult_1/xin[864] ) );
  DFF \modmult_1/xreg_reg[863]  ( .D(\modmult_1/xin[862] ), .CLK(clk), .RST(
        start_in[0]), .I(c[863]), .Q(\modmult_1/xin[863] ) );
  DFF \modmult_1/xreg_reg[862]  ( .D(\modmult_1/xin[861] ), .CLK(clk), .RST(
        start_in[0]), .I(c[862]), .Q(\modmult_1/xin[862] ) );
  DFF \modmult_1/xreg_reg[861]  ( .D(\modmult_1/xin[860] ), .CLK(clk), .RST(
        start_in[0]), .I(c[861]), .Q(\modmult_1/xin[861] ) );
  DFF \modmult_1/xreg_reg[860]  ( .D(\modmult_1/xin[859] ), .CLK(clk), .RST(
        start_in[0]), .I(c[860]), .Q(\modmult_1/xin[860] ) );
  DFF \modmult_1/xreg_reg[859]  ( .D(\modmult_1/xin[858] ), .CLK(clk), .RST(
        start_in[0]), .I(c[859]), .Q(\modmult_1/xin[859] ) );
  DFF \modmult_1/xreg_reg[858]  ( .D(\modmult_1/xin[857] ), .CLK(clk), .RST(
        start_in[0]), .I(c[858]), .Q(\modmult_1/xin[858] ) );
  DFF \modmult_1/xreg_reg[857]  ( .D(\modmult_1/xin[856] ), .CLK(clk), .RST(
        start_in[0]), .I(c[857]), .Q(\modmult_1/xin[857] ) );
  DFF \modmult_1/xreg_reg[856]  ( .D(\modmult_1/xin[855] ), .CLK(clk), .RST(
        start_in[0]), .I(c[856]), .Q(\modmult_1/xin[856] ) );
  DFF \modmult_1/xreg_reg[855]  ( .D(\modmult_1/xin[854] ), .CLK(clk), .RST(
        start_in[0]), .I(c[855]), .Q(\modmult_1/xin[855] ) );
  DFF \modmult_1/xreg_reg[854]  ( .D(\modmult_1/xin[853] ), .CLK(clk), .RST(
        start_in[0]), .I(c[854]), .Q(\modmult_1/xin[854] ) );
  DFF \modmult_1/xreg_reg[853]  ( .D(\modmult_1/xin[852] ), .CLK(clk), .RST(
        start_in[0]), .I(c[853]), .Q(\modmult_1/xin[853] ) );
  DFF \modmult_1/xreg_reg[852]  ( .D(\modmult_1/xin[851] ), .CLK(clk), .RST(
        start_in[0]), .I(c[852]), .Q(\modmult_1/xin[852] ) );
  DFF \modmult_1/xreg_reg[851]  ( .D(\modmult_1/xin[850] ), .CLK(clk), .RST(
        start_in[0]), .I(c[851]), .Q(\modmult_1/xin[851] ) );
  DFF \modmult_1/xreg_reg[850]  ( .D(\modmult_1/xin[849] ), .CLK(clk), .RST(
        start_in[0]), .I(c[850]), .Q(\modmult_1/xin[850] ) );
  DFF \modmult_1/xreg_reg[849]  ( .D(\modmult_1/xin[848] ), .CLK(clk), .RST(
        start_in[0]), .I(c[849]), .Q(\modmult_1/xin[849] ) );
  DFF \modmult_1/xreg_reg[848]  ( .D(\modmult_1/xin[847] ), .CLK(clk), .RST(
        start_in[0]), .I(c[848]), .Q(\modmult_1/xin[848] ) );
  DFF \modmult_1/xreg_reg[847]  ( .D(\modmult_1/xin[846] ), .CLK(clk), .RST(
        start_in[0]), .I(c[847]), .Q(\modmult_1/xin[847] ) );
  DFF \modmult_1/xreg_reg[846]  ( .D(\modmult_1/xin[845] ), .CLK(clk), .RST(
        start_in[0]), .I(c[846]), .Q(\modmult_1/xin[846] ) );
  DFF \modmult_1/xreg_reg[845]  ( .D(\modmult_1/xin[844] ), .CLK(clk), .RST(
        start_in[0]), .I(c[845]), .Q(\modmult_1/xin[845] ) );
  DFF \modmult_1/xreg_reg[844]  ( .D(\modmult_1/xin[843] ), .CLK(clk), .RST(
        start_in[0]), .I(c[844]), .Q(\modmult_1/xin[844] ) );
  DFF \modmult_1/xreg_reg[843]  ( .D(\modmult_1/xin[842] ), .CLK(clk), .RST(
        start_in[0]), .I(c[843]), .Q(\modmult_1/xin[843] ) );
  DFF \modmult_1/xreg_reg[842]  ( .D(\modmult_1/xin[841] ), .CLK(clk), .RST(
        start_in[0]), .I(c[842]), .Q(\modmult_1/xin[842] ) );
  DFF \modmult_1/xreg_reg[841]  ( .D(\modmult_1/xin[840] ), .CLK(clk), .RST(
        start_in[0]), .I(c[841]), .Q(\modmult_1/xin[841] ) );
  DFF \modmult_1/xreg_reg[840]  ( .D(\modmult_1/xin[839] ), .CLK(clk), .RST(
        start_in[0]), .I(c[840]), .Q(\modmult_1/xin[840] ) );
  DFF \modmult_1/xreg_reg[839]  ( .D(\modmult_1/xin[838] ), .CLK(clk), .RST(
        start_in[0]), .I(c[839]), .Q(\modmult_1/xin[839] ) );
  DFF \modmult_1/xreg_reg[838]  ( .D(\modmult_1/xin[837] ), .CLK(clk), .RST(
        start_in[0]), .I(c[838]), .Q(\modmult_1/xin[838] ) );
  DFF \modmult_1/xreg_reg[837]  ( .D(\modmult_1/xin[836] ), .CLK(clk), .RST(
        start_in[0]), .I(c[837]), .Q(\modmult_1/xin[837] ) );
  DFF \modmult_1/xreg_reg[836]  ( .D(\modmult_1/xin[835] ), .CLK(clk), .RST(
        start_in[0]), .I(c[836]), .Q(\modmult_1/xin[836] ) );
  DFF \modmult_1/xreg_reg[835]  ( .D(\modmult_1/xin[834] ), .CLK(clk), .RST(
        start_in[0]), .I(c[835]), .Q(\modmult_1/xin[835] ) );
  DFF \modmult_1/xreg_reg[834]  ( .D(\modmult_1/xin[833] ), .CLK(clk), .RST(
        start_in[0]), .I(c[834]), .Q(\modmult_1/xin[834] ) );
  DFF \modmult_1/xreg_reg[833]  ( .D(\modmult_1/xin[832] ), .CLK(clk), .RST(
        start_in[0]), .I(c[833]), .Q(\modmult_1/xin[833] ) );
  DFF \modmult_1/xreg_reg[832]  ( .D(\modmult_1/xin[831] ), .CLK(clk), .RST(
        start_in[0]), .I(c[832]), .Q(\modmult_1/xin[832] ) );
  DFF \modmult_1/xreg_reg[831]  ( .D(\modmult_1/xin[830] ), .CLK(clk), .RST(
        start_in[0]), .I(c[831]), .Q(\modmult_1/xin[831] ) );
  DFF \modmult_1/xreg_reg[830]  ( .D(\modmult_1/xin[829] ), .CLK(clk), .RST(
        start_in[0]), .I(c[830]), .Q(\modmult_1/xin[830] ) );
  DFF \modmult_1/xreg_reg[829]  ( .D(\modmult_1/xin[828] ), .CLK(clk), .RST(
        start_in[0]), .I(c[829]), .Q(\modmult_1/xin[829] ) );
  DFF \modmult_1/xreg_reg[828]  ( .D(\modmult_1/xin[827] ), .CLK(clk), .RST(
        start_in[0]), .I(c[828]), .Q(\modmult_1/xin[828] ) );
  DFF \modmult_1/xreg_reg[827]  ( .D(\modmult_1/xin[826] ), .CLK(clk), .RST(
        start_in[0]), .I(c[827]), .Q(\modmult_1/xin[827] ) );
  DFF \modmult_1/xreg_reg[826]  ( .D(\modmult_1/xin[825] ), .CLK(clk), .RST(
        start_in[0]), .I(c[826]), .Q(\modmult_1/xin[826] ) );
  DFF \modmult_1/xreg_reg[825]  ( .D(\modmult_1/xin[824] ), .CLK(clk), .RST(
        start_in[0]), .I(c[825]), .Q(\modmult_1/xin[825] ) );
  DFF \modmult_1/xreg_reg[824]  ( .D(\modmult_1/xin[823] ), .CLK(clk), .RST(
        start_in[0]), .I(c[824]), .Q(\modmult_1/xin[824] ) );
  DFF \modmult_1/xreg_reg[823]  ( .D(\modmult_1/xin[822] ), .CLK(clk), .RST(
        start_in[0]), .I(c[823]), .Q(\modmult_1/xin[823] ) );
  DFF \modmult_1/xreg_reg[822]  ( .D(\modmult_1/xin[821] ), .CLK(clk), .RST(
        start_in[0]), .I(c[822]), .Q(\modmult_1/xin[822] ) );
  DFF \modmult_1/xreg_reg[821]  ( .D(\modmult_1/xin[820] ), .CLK(clk), .RST(
        start_in[0]), .I(c[821]), .Q(\modmult_1/xin[821] ) );
  DFF \modmult_1/xreg_reg[820]  ( .D(\modmult_1/xin[819] ), .CLK(clk), .RST(
        start_in[0]), .I(c[820]), .Q(\modmult_1/xin[820] ) );
  DFF \modmult_1/xreg_reg[819]  ( .D(\modmult_1/xin[818] ), .CLK(clk), .RST(
        start_in[0]), .I(c[819]), .Q(\modmult_1/xin[819] ) );
  DFF \modmult_1/xreg_reg[818]  ( .D(\modmult_1/xin[817] ), .CLK(clk), .RST(
        start_in[0]), .I(c[818]), .Q(\modmult_1/xin[818] ) );
  DFF \modmult_1/xreg_reg[817]  ( .D(\modmult_1/xin[816] ), .CLK(clk), .RST(
        start_in[0]), .I(c[817]), .Q(\modmult_1/xin[817] ) );
  DFF \modmult_1/xreg_reg[816]  ( .D(\modmult_1/xin[815] ), .CLK(clk), .RST(
        start_in[0]), .I(c[816]), .Q(\modmult_1/xin[816] ) );
  DFF \modmult_1/xreg_reg[815]  ( .D(\modmult_1/xin[814] ), .CLK(clk), .RST(
        start_in[0]), .I(c[815]), .Q(\modmult_1/xin[815] ) );
  DFF \modmult_1/xreg_reg[814]  ( .D(\modmult_1/xin[813] ), .CLK(clk), .RST(
        start_in[0]), .I(c[814]), .Q(\modmult_1/xin[814] ) );
  DFF \modmult_1/xreg_reg[813]  ( .D(\modmult_1/xin[812] ), .CLK(clk), .RST(
        start_in[0]), .I(c[813]), .Q(\modmult_1/xin[813] ) );
  DFF \modmult_1/xreg_reg[812]  ( .D(\modmult_1/xin[811] ), .CLK(clk), .RST(
        start_in[0]), .I(c[812]), .Q(\modmult_1/xin[812] ) );
  DFF \modmult_1/xreg_reg[811]  ( .D(\modmult_1/xin[810] ), .CLK(clk), .RST(
        start_in[0]), .I(c[811]), .Q(\modmult_1/xin[811] ) );
  DFF \modmult_1/xreg_reg[810]  ( .D(\modmult_1/xin[809] ), .CLK(clk), .RST(
        start_in[0]), .I(c[810]), .Q(\modmult_1/xin[810] ) );
  DFF \modmult_1/xreg_reg[809]  ( .D(\modmult_1/xin[808] ), .CLK(clk), .RST(
        start_in[0]), .I(c[809]), .Q(\modmult_1/xin[809] ) );
  DFF \modmult_1/xreg_reg[808]  ( .D(\modmult_1/xin[807] ), .CLK(clk), .RST(
        start_in[0]), .I(c[808]), .Q(\modmult_1/xin[808] ) );
  DFF \modmult_1/xreg_reg[807]  ( .D(\modmult_1/xin[806] ), .CLK(clk), .RST(
        start_in[0]), .I(c[807]), .Q(\modmult_1/xin[807] ) );
  DFF \modmult_1/xreg_reg[806]  ( .D(\modmult_1/xin[805] ), .CLK(clk), .RST(
        start_in[0]), .I(c[806]), .Q(\modmult_1/xin[806] ) );
  DFF \modmult_1/xreg_reg[805]  ( .D(\modmult_1/xin[804] ), .CLK(clk), .RST(
        start_in[0]), .I(c[805]), .Q(\modmult_1/xin[805] ) );
  DFF \modmult_1/xreg_reg[804]  ( .D(\modmult_1/xin[803] ), .CLK(clk), .RST(
        start_in[0]), .I(c[804]), .Q(\modmult_1/xin[804] ) );
  DFF \modmult_1/xreg_reg[803]  ( .D(\modmult_1/xin[802] ), .CLK(clk), .RST(
        start_in[0]), .I(c[803]), .Q(\modmult_1/xin[803] ) );
  DFF \modmult_1/xreg_reg[802]  ( .D(\modmult_1/xin[801] ), .CLK(clk), .RST(
        start_in[0]), .I(c[802]), .Q(\modmult_1/xin[802] ) );
  DFF \modmult_1/xreg_reg[801]  ( .D(\modmult_1/xin[800] ), .CLK(clk), .RST(
        start_in[0]), .I(c[801]), .Q(\modmult_1/xin[801] ) );
  DFF \modmult_1/xreg_reg[800]  ( .D(\modmult_1/xin[799] ), .CLK(clk), .RST(
        start_in[0]), .I(c[800]), .Q(\modmult_1/xin[800] ) );
  DFF \modmult_1/xreg_reg[799]  ( .D(\modmult_1/xin[798] ), .CLK(clk), .RST(
        start_in[0]), .I(c[799]), .Q(\modmult_1/xin[799] ) );
  DFF \modmult_1/xreg_reg[798]  ( .D(\modmult_1/xin[797] ), .CLK(clk), .RST(
        start_in[0]), .I(c[798]), .Q(\modmult_1/xin[798] ) );
  DFF \modmult_1/xreg_reg[797]  ( .D(\modmult_1/xin[796] ), .CLK(clk), .RST(
        start_in[0]), .I(c[797]), .Q(\modmult_1/xin[797] ) );
  DFF \modmult_1/xreg_reg[796]  ( .D(\modmult_1/xin[795] ), .CLK(clk), .RST(
        start_in[0]), .I(c[796]), .Q(\modmult_1/xin[796] ) );
  DFF \modmult_1/xreg_reg[795]  ( .D(\modmult_1/xin[794] ), .CLK(clk), .RST(
        start_in[0]), .I(c[795]), .Q(\modmult_1/xin[795] ) );
  DFF \modmult_1/xreg_reg[794]  ( .D(\modmult_1/xin[793] ), .CLK(clk), .RST(
        start_in[0]), .I(c[794]), .Q(\modmult_1/xin[794] ) );
  DFF \modmult_1/xreg_reg[793]  ( .D(\modmult_1/xin[792] ), .CLK(clk), .RST(
        start_in[0]), .I(c[793]), .Q(\modmult_1/xin[793] ) );
  DFF \modmult_1/xreg_reg[792]  ( .D(\modmult_1/xin[791] ), .CLK(clk), .RST(
        start_in[0]), .I(c[792]), .Q(\modmult_1/xin[792] ) );
  DFF \modmult_1/xreg_reg[791]  ( .D(\modmult_1/xin[790] ), .CLK(clk), .RST(
        start_in[0]), .I(c[791]), .Q(\modmult_1/xin[791] ) );
  DFF \modmult_1/xreg_reg[790]  ( .D(\modmult_1/xin[789] ), .CLK(clk), .RST(
        start_in[0]), .I(c[790]), .Q(\modmult_1/xin[790] ) );
  DFF \modmult_1/xreg_reg[789]  ( .D(\modmult_1/xin[788] ), .CLK(clk), .RST(
        start_in[0]), .I(c[789]), .Q(\modmult_1/xin[789] ) );
  DFF \modmult_1/xreg_reg[788]  ( .D(\modmult_1/xin[787] ), .CLK(clk), .RST(
        start_in[0]), .I(c[788]), .Q(\modmult_1/xin[788] ) );
  DFF \modmult_1/xreg_reg[787]  ( .D(\modmult_1/xin[786] ), .CLK(clk), .RST(
        start_in[0]), .I(c[787]), .Q(\modmult_1/xin[787] ) );
  DFF \modmult_1/xreg_reg[786]  ( .D(\modmult_1/xin[785] ), .CLK(clk), .RST(
        start_in[0]), .I(c[786]), .Q(\modmult_1/xin[786] ) );
  DFF \modmult_1/xreg_reg[785]  ( .D(\modmult_1/xin[784] ), .CLK(clk), .RST(
        start_in[0]), .I(c[785]), .Q(\modmult_1/xin[785] ) );
  DFF \modmult_1/xreg_reg[784]  ( .D(\modmult_1/xin[783] ), .CLK(clk), .RST(
        start_in[0]), .I(c[784]), .Q(\modmult_1/xin[784] ) );
  DFF \modmult_1/xreg_reg[783]  ( .D(\modmult_1/xin[782] ), .CLK(clk), .RST(
        start_in[0]), .I(c[783]), .Q(\modmult_1/xin[783] ) );
  DFF \modmult_1/xreg_reg[782]  ( .D(\modmult_1/xin[781] ), .CLK(clk), .RST(
        start_in[0]), .I(c[782]), .Q(\modmult_1/xin[782] ) );
  DFF \modmult_1/xreg_reg[781]  ( .D(\modmult_1/xin[780] ), .CLK(clk), .RST(
        start_in[0]), .I(c[781]), .Q(\modmult_1/xin[781] ) );
  DFF \modmult_1/xreg_reg[780]  ( .D(\modmult_1/xin[779] ), .CLK(clk), .RST(
        start_in[0]), .I(c[780]), .Q(\modmult_1/xin[780] ) );
  DFF \modmult_1/xreg_reg[779]  ( .D(\modmult_1/xin[778] ), .CLK(clk), .RST(
        start_in[0]), .I(c[779]), .Q(\modmult_1/xin[779] ) );
  DFF \modmult_1/xreg_reg[778]  ( .D(\modmult_1/xin[777] ), .CLK(clk), .RST(
        start_in[0]), .I(c[778]), .Q(\modmult_1/xin[778] ) );
  DFF \modmult_1/xreg_reg[777]  ( .D(\modmult_1/xin[776] ), .CLK(clk), .RST(
        start_in[0]), .I(c[777]), .Q(\modmult_1/xin[777] ) );
  DFF \modmult_1/xreg_reg[776]  ( .D(\modmult_1/xin[775] ), .CLK(clk), .RST(
        start_in[0]), .I(c[776]), .Q(\modmult_1/xin[776] ) );
  DFF \modmult_1/xreg_reg[775]  ( .D(\modmult_1/xin[774] ), .CLK(clk), .RST(
        start_in[0]), .I(c[775]), .Q(\modmult_1/xin[775] ) );
  DFF \modmult_1/xreg_reg[774]  ( .D(\modmult_1/xin[773] ), .CLK(clk), .RST(
        start_in[0]), .I(c[774]), .Q(\modmult_1/xin[774] ) );
  DFF \modmult_1/xreg_reg[773]  ( .D(\modmult_1/xin[772] ), .CLK(clk), .RST(
        start_in[0]), .I(c[773]), .Q(\modmult_1/xin[773] ) );
  DFF \modmult_1/xreg_reg[772]  ( .D(\modmult_1/xin[771] ), .CLK(clk), .RST(
        start_in[0]), .I(c[772]), .Q(\modmult_1/xin[772] ) );
  DFF \modmult_1/xreg_reg[771]  ( .D(\modmult_1/xin[770] ), .CLK(clk), .RST(
        start_in[0]), .I(c[771]), .Q(\modmult_1/xin[771] ) );
  DFF \modmult_1/xreg_reg[770]  ( .D(\modmult_1/xin[769] ), .CLK(clk), .RST(
        start_in[0]), .I(c[770]), .Q(\modmult_1/xin[770] ) );
  DFF \modmult_1/xreg_reg[769]  ( .D(\modmult_1/xin[768] ), .CLK(clk), .RST(
        start_in[0]), .I(c[769]), .Q(\modmult_1/xin[769] ) );
  DFF \modmult_1/xreg_reg[768]  ( .D(\modmult_1/xin[767] ), .CLK(clk), .RST(
        start_in[0]), .I(c[768]), .Q(\modmult_1/xin[768] ) );
  DFF \modmult_1/xreg_reg[767]  ( .D(\modmult_1/xin[766] ), .CLK(clk), .RST(
        start_in[0]), .I(c[767]), .Q(\modmult_1/xin[767] ) );
  DFF \modmult_1/xreg_reg[766]  ( .D(\modmult_1/xin[765] ), .CLK(clk), .RST(
        start_in[0]), .I(c[766]), .Q(\modmult_1/xin[766] ) );
  DFF \modmult_1/xreg_reg[765]  ( .D(\modmult_1/xin[764] ), .CLK(clk), .RST(
        start_in[0]), .I(c[765]), .Q(\modmult_1/xin[765] ) );
  DFF \modmult_1/xreg_reg[764]  ( .D(\modmult_1/xin[763] ), .CLK(clk), .RST(
        start_in[0]), .I(c[764]), .Q(\modmult_1/xin[764] ) );
  DFF \modmult_1/xreg_reg[763]  ( .D(\modmult_1/xin[762] ), .CLK(clk), .RST(
        start_in[0]), .I(c[763]), .Q(\modmult_1/xin[763] ) );
  DFF \modmult_1/xreg_reg[762]  ( .D(\modmult_1/xin[761] ), .CLK(clk), .RST(
        start_in[0]), .I(c[762]), .Q(\modmult_1/xin[762] ) );
  DFF \modmult_1/xreg_reg[761]  ( .D(\modmult_1/xin[760] ), .CLK(clk), .RST(
        start_in[0]), .I(c[761]), .Q(\modmult_1/xin[761] ) );
  DFF \modmult_1/xreg_reg[760]  ( .D(\modmult_1/xin[759] ), .CLK(clk), .RST(
        start_in[0]), .I(c[760]), .Q(\modmult_1/xin[760] ) );
  DFF \modmult_1/xreg_reg[759]  ( .D(\modmult_1/xin[758] ), .CLK(clk), .RST(
        start_in[0]), .I(c[759]), .Q(\modmult_1/xin[759] ) );
  DFF \modmult_1/xreg_reg[758]  ( .D(\modmult_1/xin[757] ), .CLK(clk), .RST(
        start_in[0]), .I(c[758]), .Q(\modmult_1/xin[758] ) );
  DFF \modmult_1/xreg_reg[757]  ( .D(\modmult_1/xin[756] ), .CLK(clk), .RST(
        start_in[0]), .I(c[757]), .Q(\modmult_1/xin[757] ) );
  DFF \modmult_1/xreg_reg[756]  ( .D(\modmult_1/xin[755] ), .CLK(clk), .RST(
        start_in[0]), .I(c[756]), .Q(\modmult_1/xin[756] ) );
  DFF \modmult_1/xreg_reg[755]  ( .D(\modmult_1/xin[754] ), .CLK(clk), .RST(
        start_in[0]), .I(c[755]), .Q(\modmult_1/xin[755] ) );
  DFF \modmult_1/xreg_reg[754]  ( .D(\modmult_1/xin[753] ), .CLK(clk), .RST(
        start_in[0]), .I(c[754]), .Q(\modmult_1/xin[754] ) );
  DFF \modmult_1/xreg_reg[753]  ( .D(\modmult_1/xin[752] ), .CLK(clk), .RST(
        start_in[0]), .I(c[753]), .Q(\modmult_1/xin[753] ) );
  DFF \modmult_1/xreg_reg[752]  ( .D(\modmult_1/xin[751] ), .CLK(clk), .RST(
        start_in[0]), .I(c[752]), .Q(\modmult_1/xin[752] ) );
  DFF \modmult_1/xreg_reg[751]  ( .D(\modmult_1/xin[750] ), .CLK(clk), .RST(
        start_in[0]), .I(c[751]), .Q(\modmult_1/xin[751] ) );
  DFF \modmult_1/xreg_reg[750]  ( .D(\modmult_1/xin[749] ), .CLK(clk), .RST(
        start_in[0]), .I(c[750]), .Q(\modmult_1/xin[750] ) );
  DFF \modmult_1/xreg_reg[749]  ( .D(\modmult_1/xin[748] ), .CLK(clk), .RST(
        start_in[0]), .I(c[749]), .Q(\modmult_1/xin[749] ) );
  DFF \modmult_1/xreg_reg[748]  ( .D(\modmult_1/xin[747] ), .CLK(clk), .RST(
        start_in[0]), .I(c[748]), .Q(\modmult_1/xin[748] ) );
  DFF \modmult_1/xreg_reg[747]  ( .D(\modmult_1/xin[746] ), .CLK(clk), .RST(
        start_in[0]), .I(c[747]), .Q(\modmult_1/xin[747] ) );
  DFF \modmult_1/xreg_reg[746]  ( .D(\modmult_1/xin[745] ), .CLK(clk), .RST(
        start_in[0]), .I(c[746]), .Q(\modmult_1/xin[746] ) );
  DFF \modmult_1/xreg_reg[745]  ( .D(\modmult_1/xin[744] ), .CLK(clk), .RST(
        start_in[0]), .I(c[745]), .Q(\modmult_1/xin[745] ) );
  DFF \modmult_1/xreg_reg[744]  ( .D(\modmult_1/xin[743] ), .CLK(clk), .RST(
        start_in[0]), .I(c[744]), .Q(\modmult_1/xin[744] ) );
  DFF \modmult_1/xreg_reg[743]  ( .D(\modmult_1/xin[742] ), .CLK(clk), .RST(
        start_in[0]), .I(c[743]), .Q(\modmult_1/xin[743] ) );
  DFF \modmult_1/xreg_reg[742]  ( .D(\modmult_1/xin[741] ), .CLK(clk), .RST(
        start_in[0]), .I(c[742]), .Q(\modmult_1/xin[742] ) );
  DFF \modmult_1/xreg_reg[741]  ( .D(\modmult_1/xin[740] ), .CLK(clk), .RST(
        start_in[0]), .I(c[741]), .Q(\modmult_1/xin[741] ) );
  DFF \modmult_1/xreg_reg[740]  ( .D(\modmult_1/xin[739] ), .CLK(clk), .RST(
        start_in[0]), .I(c[740]), .Q(\modmult_1/xin[740] ) );
  DFF \modmult_1/xreg_reg[739]  ( .D(\modmult_1/xin[738] ), .CLK(clk), .RST(
        start_in[0]), .I(c[739]), .Q(\modmult_1/xin[739] ) );
  DFF \modmult_1/xreg_reg[738]  ( .D(\modmult_1/xin[737] ), .CLK(clk), .RST(
        start_in[0]), .I(c[738]), .Q(\modmult_1/xin[738] ) );
  DFF \modmult_1/xreg_reg[737]  ( .D(\modmult_1/xin[736] ), .CLK(clk), .RST(
        start_in[0]), .I(c[737]), .Q(\modmult_1/xin[737] ) );
  DFF \modmult_1/xreg_reg[736]  ( .D(\modmult_1/xin[735] ), .CLK(clk), .RST(
        start_in[0]), .I(c[736]), .Q(\modmult_1/xin[736] ) );
  DFF \modmult_1/xreg_reg[735]  ( .D(\modmult_1/xin[734] ), .CLK(clk), .RST(
        start_in[0]), .I(c[735]), .Q(\modmult_1/xin[735] ) );
  DFF \modmult_1/xreg_reg[734]  ( .D(\modmult_1/xin[733] ), .CLK(clk), .RST(
        start_in[0]), .I(c[734]), .Q(\modmult_1/xin[734] ) );
  DFF \modmult_1/xreg_reg[733]  ( .D(\modmult_1/xin[732] ), .CLK(clk), .RST(
        start_in[0]), .I(c[733]), .Q(\modmult_1/xin[733] ) );
  DFF \modmult_1/xreg_reg[732]  ( .D(\modmult_1/xin[731] ), .CLK(clk), .RST(
        start_in[0]), .I(c[732]), .Q(\modmult_1/xin[732] ) );
  DFF \modmult_1/xreg_reg[731]  ( .D(\modmult_1/xin[730] ), .CLK(clk), .RST(
        start_in[0]), .I(c[731]), .Q(\modmult_1/xin[731] ) );
  DFF \modmult_1/xreg_reg[730]  ( .D(\modmult_1/xin[729] ), .CLK(clk), .RST(
        start_in[0]), .I(c[730]), .Q(\modmult_1/xin[730] ) );
  DFF \modmult_1/xreg_reg[729]  ( .D(\modmult_1/xin[728] ), .CLK(clk), .RST(
        start_in[0]), .I(c[729]), .Q(\modmult_1/xin[729] ) );
  DFF \modmult_1/xreg_reg[728]  ( .D(\modmult_1/xin[727] ), .CLK(clk), .RST(
        start_in[0]), .I(c[728]), .Q(\modmult_1/xin[728] ) );
  DFF \modmult_1/xreg_reg[727]  ( .D(\modmult_1/xin[726] ), .CLK(clk), .RST(
        start_in[0]), .I(c[727]), .Q(\modmult_1/xin[727] ) );
  DFF \modmult_1/xreg_reg[726]  ( .D(\modmult_1/xin[725] ), .CLK(clk), .RST(
        start_in[0]), .I(c[726]), .Q(\modmult_1/xin[726] ) );
  DFF \modmult_1/xreg_reg[725]  ( .D(\modmult_1/xin[724] ), .CLK(clk), .RST(
        start_in[0]), .I(c[725]), .Q(\modmult_1/xin[725] ) );
  DFF \modmult_1/xreg_reg[724]  ( .D(\modmult_1/xin[723] ), .CLK(clk), .RST(
        start_in[0]), .I(c[724]), .Q(\modmult_1/xin[724] ) );
  DFF \modmult_1/xreg_reg[723]  ( .D(\modmult_1/xin[722] ), .CLK(clk), .RST(
        start_in[0]), .I(c[723]), .Q(\modmult_1/xin[723] ) );
  DFF \modmult_1/xreg_reg[722]  ( .D(\modmult_1/xin[721] ), .CLK(clk), .RST(
        start_in[0]), .I(c[722]), .Q(\modmult_1/xin[722] ) );
  DFF \modmult_1/xreg_reg[721]  ( .D(\modmult_1/xin[720] ), .CLK(clk), .RST(
        start_in[0]), .I(c[721]), .Q(\modmult_1/xin[721] ) );
  DFF \modmult_1/xreg_reg[720]  ( .D(\modmult_1/xin[719] ), .CLK(clk), .RST(
        start_in[0]), .I(c[720]), .Q(\modmult_1/xin[720] ) );
  DFF \modmult_1/xreg_reg[719]  ( .D(\modmult_1/xin[718] ), .CLK(clk), .RST(
        start_in[0]), .I(c[719]), .Q(\modmult_1/xin[719] ) );
  DFF \modmult_1/xreg_reg[718]  ( .D(\modmult_1/xin[717] ), .CLK(clk), .RST(
        start_in[0]), .I(c[718]), .Q(\modmult_1/xin[718] ) );
  DFF \modmult_1/xreg_reg[717]  ( .D(\modmult_1/xin[716] ), .CLK(clk), .RST(
        start_in[0]), .I(c[717]), .Q(\modmult_1/xin[717] ) );
  DFF \modmult_1/xreg_reg[716]  ( .D(\modmult_1/xin[715] ), .CLK(clk), .RST(
        start_in[0]), .I(c[716]), .Q(\modmult_1/xin[716] ) );
  DFF \modmult_1/xreg_reg[715]  ( .D(\modmult_1/xin[714] ), .CLK(clk), .RST(
        start_in[0]), .I(c[715]), .Q(\modmult_1/xin[715] ) );
  DFF \modmult_1/xreg_reg[714]  ( .D(\modmult_1/xin[713] ), .CLK(clk), .RST(
        start_in[0]), .I(c[714]), .Q(\modmult_1/xin[714] ) );
  DFF \modmult_1/xreg_reg[713]  ( .D(\modmult_1/xin[712] ), .CLK(clk), .RST(
        start_in[0]), .I(c[713]), .Q(\modmult_1/xin[713] ) );
  DFF \modmult_1/xreg_reg[712]  ( .D(\modmult_1/xin[711] ), .CLK(clk), .RST(
        start_in[0]), .I(c[712]), .Q(\modmult_1/xin[712] ) );
  DFF \modmult_1/xreg_reg[711]  ( .D(\modmult_1/xin[710] ), .CLK(clk), .RST(
        start_in[0]), .I(c[711]), .Q(\modmult_1/xin[711] ) );
  DFF \modmult_1/xreg_reg[710]  ( .D(\modmult_1/xin[709] ), .CLK(clk), .RST(
        start_in[0]), .I(c[710]), .Q(\modmult_1/xin[710] ) );
  DFF \modmult_1/xreg_reg[709]  ( .D(\modmult_1/xin[708] ), .CLK(clk), .RST(
        start_in[0]), .I(c[709]), .Q(\modmult_1/xin[709] ) );
  DFF \modmult_1/xreg_reg[708]  ( .D(\modmult_1/xin[707] ), .CLK(clk), .RST(
        start_in[0]), .I(c[708]), .Q(\modmult_1/xin[708] ) );
  DFF \modmult_1/xreg_reg[707]  ( .D(\modmult_1/xin[706] ), .CLK(clk), .RST(
        start_in[0]), .I(c[707]), .Q(\modmult_1/xin[707] ) );
  DFF \modmult_1/xreg_reg[706]  ( .D(\modmult_1/xin[705] ), .CLK(clk), .RST(
        start_in[0]), .I(c[706]), .Q(\modmult_1/xin[706] ) );
  DFF \modmult_1/xreg_reg[705]  ( .D(\modmult_1/xin[704] ), .CLK(clk), .RST(
        start_in[0]), .I(c[705]), .Q(\modmult_1/xin[705] ) );
  DFF \modmult_1/xreg_reg[704]  ( .D(\modmult_1/xin[703] ), .CLK(clk), .RST(
        start_in[0]), .I(c[704]), .Q(\modmult_1/xin[704] ) );
  DFF \modmult_1/xreg_reg[703]  ( .D(\modmult_1/xin[702] ), .CLK(clk), .RST(
        start_in[0]), .I(c[703]), .Q(\modmult_1/xin[703] ) );
  DFF \modmult_1/xreg_reg[702]  ( .D(\modmult_1/xin[701] ), .CLK(clk), .RST(
        start_in[0]), .I(c[702]), .Q(\modmult_1/xin[702] ) );
  DFF \modmult_1/xreg_reg[701]  ( .D(\modmult_1/xin[700] ), .CLK(clk), .RST(
        start_in[0]), .I(c[701]), .Q(\modmult_1/xin[701] ) );
  DFF \modmult_1/xreg_reg[700]  ( .D(\modmult_1/xin[699] ), .CLK(clk), .RST(
        start_in[0]), .I(c[700]), .Q(\modmult_1/xin[700] ) );
  DFF \modmult_1/xreg_reg[699]  ( .D(\modmult_1/xin[698] ), .CLK(clk), .RST(
        start_in[0]), .I(c[699]), .Q(\modmult_1/xin[699] ) );
  DFF \modmult_1/xreg_reg[698]  ( .D(\modmult_1/xin[697] ), .CLK(clk), .RST(
        start_in[0]), .I(c[698]), .Q(\modmult_1/xin[698] ) );
  DFF \modmult_1/xreg_reg[697]  ( .D(\modmult_1/xin[696] ), .CLK(clk), .RST(
        start_in[0]), .I(c[697]), .Q(\modmult_1/xin[697] ) );
  DFF \modmult_1/xreg_reg[696]  ( .D(\modmult_1/xin[695] ), .CLK(clk), .RST(
        start_in[0]), .I(c[696]), .Q(\modmult_1/xin[696] ) );
  DFF \modmult_1/xreg_reg[695]  ( .D(\modmult_1/xin[694] ), .CLK(clk), .RST(
        start_in[0]), .I(c[695]), .Q(\modmult_1/xin[695] ) );
  DFF \modmult_1/xreg_reg[694]  ( .D(\modmult_1/xin[693] ), .CLK(clk), .RST(
        start_in[0]), .I(c[694]), .Q(\modmult_1/xin[694] ) );
  DFF \modmult_1/xreg_reg[693]  ( .D(\modmult_1/xin[692] ), .CLK(clk), .RST(
        start_in[0]), .I(c[693]), .Q(\modmult_1/xin[693] ) );
  DFF \modmult_1/xreg_reg[692]  ( .D(\modmult_1/xin[691] ), .CLK(clk), .RST(
        start_in[0]), .I(c[692]), .Q(\modmult_1/xin[692] ) );
  DFF \modmult_1/xreg_reg[691]  ( .D(\modmult_1/xin[690] ), .CLK(clk), .RST(
        start_in[0]), .I(c[691]), .Q(\modmult_1/xin[691] ) );
  DFF \modmult_1/xreg_reg[690]  ( .D(\modmult_1/xin[689] ), .CLK(clk), .RST(
        start_in[0]), .I(c[690]), .Q(\modmult_1/xin[690] ) );
  DFF \modmult_1/xreg_reg[689]  ( .D(\modmult_1/xin[688] ), .CLK(clk), .RST(
        start_in[0]), .I(c[689]), .Q(\modmult_1/xin[689] ) );
  DFF \modmult_1/xreg_reg[688]  ( .D(\modmult_1/xin[687] ), .CLK(clk), .RST(
        start_in[0]), .I(c[688]), .Q(\modmult_1/xin[688] ) );
  DFF \modmult_1/xreg_reg[687]  ( .D(\modmult_1/xin[686] ), .CLK(clk), .RST(
        start_in[0]), .I(c[687]), .Q(\modmult_1/xin[687] ) );
  DFF \modmult_1/xreg_reg[686]  ( .D(\modmult_1/xin[685] ), .CLK(clk), .RST(
        start_in[0]), .I(c[686]), .Q(\modmult_1/xin[686] ) );
  DFF \modmult_1/xreg_reg[685]  ( .D(\modmult_1/xin[684] ), .CLK(clk), .RST(
        start_in[0]), .I(c[685]), .Q(\modmult_1/xin[685] ) );
  DFF \modmult_1/xreg_reg[684]  ( .D(\modmult_1/xin[683] ), .CLK(clk), .RST(
        start_in[0]), .I(c[684]), .Q(\modmult_1/xin[684] ) );
  DFF \modmult_1/xreg_reg[683]  ( .D(\modmult_1/xin[682] ), .CLK(clk), .RST(
        start_in[0]), .I(c[683]), .Q(\modmult_1/xin[683] ) );
  DFF \modmult_1/xreg_reg[682]  ( .D(\modmult_1/xin[681] ), .CLK(clk), .RST(
        start_in[0]), .I(c[682]), .Q(\modmult_1/xin[682] ) );
  DFF \modmult_1/xreg_reg[681]  ( .D(\modmult_1/xin[680] ), .CLK(clk), .RST(
        start_in[0]), .I(c[681]), .Q(\modmult_1/xin[681] ) );
  DFF \modmult_1/xreg_reg[680]  ( .D(\modmult_1/xin[679] ), .CLK(clk), .RST(
        start_in[0]), .I(c[680]), .Q(\modmult_1/xin[680] ) );
  DFF \modmult_1/xreg_reg[679]  ( .D(\modmult_1/xin[678] ), .CLK(clk), .RST(
        start_in[0]), .I(c[679]), .Q(\modmult_1/xin[679] ) );
  DFF \modmult_1/xreg_reg[678]  ( .D(\modmult_1/xin[677] ), .CLK(clk), .RST(
        start_in[0]), .I(c[678]), .Q(\modmult_1/xin[678] ) );
  DFF \modmult_1/xreg_reg[677]  ( .D(\modmult_1/xin[676] ), .CLK(clk), .RST(
        start_in[0]), .I(c[677]), .Q(\modmult_1/xin[677] ) );
  DFF \modmult_1/xreg_reg[676]  ( .D(\modmult_1/xin[675] ), .CLK(clk), .RST(
        start_in[0]), .I(c[676]), .Q(\modmult_1/xin[676] ) );
  DFF \modmult_1/xreg_reg[675]  ( .D(\modmult_1/xin[674] ), .CLK(clk), .RST(
        start_in[0]), .I(c[675]), .Q(\modmult_1/xin[675] ) );
  DFF \modmult_1/xreg_reg[674]  ( .D(\modmult_1/xin[673] ), .CLK(clk), .RST(
        start_in[0]), .I(c[674]), .Q(\modmult_1/xin[674] ) );
  DFF \modmult_1/xreg_reg[673]  ( .D(\modmult_1/xin[672] ), .CLK(clk), .RST(
        start_in[0]), .I(c[673]), .Q(\modmult_1/xin[673] ) );
  DFF \modmult_1/xreg_reg[672]  ( .D(\modmult_1/xin[671] ), .CLK(clk), .RST(
        start_in[0]), .I(c[672]), .Q(\modmult_1/xin[672] ) );
  DFF \modmult_1/xreg_reg[671]  ( .D(\modmult_1/xin[670] ), .CLK(clk), .RST(
        start_in[0]), .I(c[671]), .Q(\modmult_1/xin[671] ) );
  DFF \modmult_1/xreg_reg[670]  ( .D(\modmult_1/xin[669] ), .CLK(clk), .RST(
        start_in[0]), .I(c[670]), .Q(\modmult_1/xin[670] ) );
  DFF \modmult_1/xreg_reg[669]  ( .D(\modmult_1/xin[668] ), .CLK(clk), .RST(
        start_in[0]), .I(c[669]), .Q(\modmult_1/xin[669] ) );
  DFF \modmult_1/xreg_reg[668]  ( .D(\modmult_1/xin[667] ), .CLK(clk), .RST(
        start_in[0]), .I(c[668]), .Q(\modmult_1/xin[668] ) );
  DFF \modmult_1/xreg_reg[667]  ( .D(\modmult_1/xin[666] ), .CLK(clk), .RST(
        start_in[0]), .I(c[667]), .Q(\modmult_1/xin[667] ) );
  DFF \modmult_1/xreg_reg[666]  ( .D(\modmult_1/xin[665] ), .CLK(clk), .RST(
        start_in[0]), .I(c[666]), .Q(\modmult_1/xin[666] ) );
  DFF \modmult_1/xreg_reg[665]  ( .D(\modmult_1/xin[664] ), .CLK(clk), .RST(
        start_in[0]), .I(c[665]), .Q(\modmult_1/xin[665] ) );
  DFF \modmult_1/xreg_reg[664]  ( .D(\modmult_1/xin[663] ), .CLK(clk), .RST(
        start_in[0]), .I(c[664]), .Q(\modmult_1/xin[664] ) );
  DFF \modmult_1/xreg_reg[663]  ( .D(\modmult_1/xin[662] ), .CLK(clk), .RST(
        start_in[0]), .I(c[663]), .Q(\modmult_1/xin[663] ) );
  DFF \modmult_1/xreg_reg[662]  ( .D(\modmult_1/xin[661] ), .CLK(clk), .RST(
        start_in[0]), .I(c[662]), .Q(\modmult_1/xin[662] ) );
  DFF \modmult_1/xreg_reg[661]  ( .D(\modmult_1/xin[660] ), .CLK(clk), .RST(
        start_in[0]), .I(c[661]), .Q(\modmult_1/xin[661] ) );
  DFF \modmult_1/xreg_reg[660]  ( .D(\modmult_1/xin[659] ), .CLK(clk), .RST(
        start_in[0]), .I(c[660]), .Q(\modmult_1/xin[660] ) );
  DFF \modmult_1/xreg_reg[659]  ( .D(\modmult_1/xin[658] ), .CLK(clk), .RST(
        start_in[0]), .I(c[659]), .Q(\modmult_1/xin[659] ) );
  DFF \modmult_1/xreg_reg[658]  ( .D(\modmult_1/xin[657] ), .CLK(clk), .RST(
        start_in[0]), .I(c[658]), .Q(\modmult_1/xin[658] ) );
  DFF \modmult_1/xreg_reg[657]  ( .D(\modmult_1/xin[656] ), .CLK(clk), .RST(
        start_in[0]), .I(c[657]), .Q(\modmult_1/xin[657] ) );
  DFF \modmult_1/xreg_reg[656]  ( .D(\modmult_1/xin[655] ), .CLK(clk), .RST(
        start_in[0]), .I(c[656]), .Q(\modmult_1/xin[656] ) );
  DFF \modmult_1/xreg_reg[655]  ( .D(\modmult_1/xin[654] ), .CLK(clk), .RST(
        start_in[0]), .I(c[655]), .Q(\modmult_1/xin[655] ) );
  DFF \modmult_1/xreg_reg[654]  ( .D(\modmult_1/xin[653] ), .CLK(clk), .RST(
        start_in[0]), .I(c[654]), .Q(\modmult_1/xin[654] ) );
  DFF \modmult_1/xreg_reg[653]  ( .D(\modmult_1/xin[652] ), .CLK(clk), .RST(
        start_in[0]), .I(c[653]), .Q(\modmult_1/xin[653] ) );
  DFF \modmult_1/xreg_reg[652]  ( .D(\modmult_1/xin[651] ), .CLK(clk), .RST(
        start_in[0]), .I(c[652]), .Q(\modmult_1/xin[652] ) );
  DFF \modmult_1/xreg_reg[651]  ( .D(\modmult_1/xin[650] ), .CLK(clk), .RST(
        start_in[0]), .I(c[651]), .Q(\modmult_1/xin[651] ) );
  DFF \modmult_1/xreg_reg[650]  ( .D(\modmult_1/xin[649] ), .CLK(clk), .RST(
        start_in[0]), .I(c[650]), .Q(\modmult_1/xin[650] ) );
  DFF \modmult_1/xreg_reg[649]  ( .D(\modmult_1/xin[648] ), .CLK(clk), .RST(
        start_in[0]), .I(c[649]), .Q(\modmult_1/xin[649] ) );
  DFF \modmult_1/xreg_reg[648]  ( .D(\modmult_1/xin[647] ), .CLK(clk), .RST(
        start_in[0]), .I(c[648]), .Q(\modmult_1/xin[648] ) );
  DFF \modmult_1/xreg_reg[647]  ( .D(\modmult_1/xin[646] ), .CLK(clk), .RST(
        start_in[0]), .I(c[647]), .Q(\modmult_1/xin[647] ) );
  DFF \modmult_1/xreg_reg[646]  ( .D(\modmult_1/xin[645] ), .CLK(clk), .RST(
        start_in[0]), .I(c[646]), .Q(\modmult_1/xin[646] ) );
  DFF \modmult_1/xreg_reg[645]  ( .D(\modmult_1/xin[644] ), .CLK(clk), .RST(
        start_in[0]), .I(c[645]), .Q(\modmult_1/xin[645] ) );
  DFF \modmult_1/xreg_reg[644]  ( .D(\modmult_1/xin[643] ), .CLK(clk), .RST(
        start_in[0]), .I(c[644]), .Q(\modmult_1/xin[644] ) );
  DFF \modmult_1/xreg_reg[643]  ( .D(\modmult_1/xin[642] ), .CLK(clk), .RST(
        start_in[0]), .I(c[643]), .Q(\modmult_1/xin[643] ) );
  DFF \modmult_1/xreg_reg[642]  ( .D(\modmult_1/xin[641] ), .CLK(clk), .RST(
        start_in[0]), .I(c[642]), .Q(\modmult_1/xin[642] ) );
  DFF \modmult_1/xreg_reg[641]  ( .D(\modmult_1/xin[640] ), .CLK(clk), .RST(
        start_in[0]), .I(c[641]), .Q(\modmult_1/xin[641] ) );
  DFF \modmult_1/xreg_reg[640]  ( .D(\modmult_1/xin[639] ), .CLK(clk), .RST(
        start_in[0]), .I(c[640]), .Q(\modmult_1/xin[640] ) );
  DFF \modmult_1/xreg_reg[639]  ( .D(\modmult_1/xin[638] ), .CLK(clk), .RST(
        start_in[0]), .I(c[639]), .Q(\modmult_1/xin[639] ) );
  DFF \modmult_1/xreg_reg[638]  ( .D(\modmult_1/xin[637] ), .CLK(clk), .RST(
        start_in[0]), .I(c[638]), .Q(\modmult_1/xin[638] ) );
  DFF \modmult_1/xreg_reg[637]  ( .D(\modmult_1/xin[636] ), .CLK(clk), .RST(
        start_in[0]), .I(c[637]), .Q(\modmult_1/xin[637] ) );
  DFF \modmult_1/xreg_reg[636]  ( .D(\modmult_1/xin[635] ), .CLK(clk), .RST(
        start_in[0]), .I(c[636]), .Q(\modmult_1/xin[636] ) );
  DFF \modmult_1/xreg_reg[635]  ( .D(\modmult_1/xin[634] ), .CLK(clk), .RST(
        start_in[0]), .I(c[635]), .Q(\modmult_1/xin[635] ) );
  DFF \modmult_1/xreg_reg[634]  ( .D(\modmult_1/xin[633] ), .CLK(clk), .RST(
        start_in[0]), .I(c[634]), .Q(\modmult_1/xin[634] ) );
  DFF \modmult_1/xreg_reg[633]  ( .D(\modmult_1/xin[632] ), .CLK(clk), .RST(
        start_in[0]), .I(c[633]), .Q(\modmult_1/xin[633] ) );
  DFF \modmult_1/xreg_reg[632]  ( .D(\modmult_1/xin[631] ), .CLK(clk), .RST(
        start_in[0]), .I(c[632]), .Q(\modmult_1/xin[632] ) );
  DFF \modmult_1/xreg_reg[631]  ( .D(\modmult_1/xin[630] ), .CLK(clk), .RST(
        start_in[0]), .I(c[631]), .Q(\modmult_1/xin[631] ) );
  DFF \modmult_1/xreg_reg[630]  ( .D(\modmult_1/xin[629] ), .CLK(clk), .RST(
        start_in[0]), .I(c[630]), .Q(\modmult_1/xin[630] ) );
  DFF \modmult_1/xreg_reg[629]  ( .D(\modmult_1/xin[628] ), .CLK(clk), .RST(
        start_in[0]), .I(c[629]), .Q(\modmult_1/xin[629] ) );
  DFF \modmult_1/xreg_reg[628]  ( .D(\modmult_1/xin[627] ), .CLK(clk), .RST(
        start_in[0]), .I(c[628]), .Q(\modmult_1/xin[628] ) );
  DFF \modmult_1/xreg_reg[627]  ( .D(\modmult_1/xin[626] ), .CLK(clk), .RST(
        start_in[0]), .I(c[627]), .Q(\modmult_1/xin[627] ) );
  DFF \modmult_1/xreg_reg[626]  ( .D(\modmult_1/xin[625] ), .CLK(clk), .RST(
        start_in[0]), .I(c[626]), .Q(\modmult_1/xin[626] ) );
  DFF \modmult_1/xreg_reg[625]  ( .D(\modmult_1/xin[624] ), .CLK(clk), .RST(
        start_in[0]), .I(c[625]), .Q(\modmult_1/xin[625] ) );
  DFF \modmult_1/xreg_reg[624]  ( .D(\modmult_1/xin[623] ), .CLK(clk), .RST(
        start_in[0]), .I(c[624]), .Q(\modmult_1/xin[624] ) );
  DFF \modmult_1/xreg_reg[623]  ( .D(\modmult_1/xin[622] ), .CLK(clk), .RST(
        start_in[0]), .I(c[623]), .Q(\modmult_1/xin[623] ) );
  DFF \modmult_1/xreg_reg[622]  ( .D(\modmult_1/xin[621] ), .CLK(clk), .RST(
        start_in[0]), .I(c[622]), .Q(\modmult_1/xin[622] ) );
  DFF \modmult_1/xreg_reg[621]  ( .D(\modmult_1/xin[620] ), .CLK(clk), .RST(
        start_in[0]), .I(c[621]), .Q(\modmult_1/xin[621] ) );
  DFF \modmult_1/xreg_reg[620]  ( .D(\modmult_1/xin[619] ), .CLK(clk), .RST(
        start_in[0]), .I(c[620]), .Q(\modmult_1/xin[620] ) );
  DFF \modmult_1/xreg_reg[619]  ( .D(\modmult_1/xin[618] ), .CLK(clk), .RST(
        start_in[0]), .I(c[619]), .Q(\modmult_1/xin[619] ) );
  DFF \modmult_1/xreg_reg[618]  ( .D(\modmult_1/xin[617] ), .CLK(clk), .RST(
        start_in[0]), .I(c[618]), .Q(\modmult_1/xin[618] ) );
  DFF \modmult_1/xreg_reg[617]  ( .D(\modmult_1/xin[616] ), .CLK(clk), .RST(
        start_in[0]), .I(c[617]), .Q(\modmult_1/xin[617] ) );
  DFF \modmult_1/xreg_reg[616]  ( .D(\modmult_1/xin[615] ), .CLK(clk), .RST(
        start_in[0]), .I(c[616]), .Q(\modmult_1/xin[616] ) );
  DFF \modmult_1/xreg_reg[615]  ( .D(\modmult_1/xin[614] ), .CLK(clk), .RST(
        start_in[0]), .I(c[615]), .Q(\modmult_1/xin[615] ) );
  DFF \modmult_1/xreg_reg[614]  ( .D(\modmult_1/xin[613] ), .CLK(clk), .RST(
        start_in[0]), .I(c[614]), .Q(\modmult_1/xin[614] ) );
  DFF \modmult_1/xreg_reg[613]  ( .D(\modmult_1/xin[612] ), .CLK(clk), .RST(
        start_in[0]), .I(c[613]), .Q(\modmult_1/xin[613] ) );
  DFF \modmult_1/xreg_reg[612]  ( .D(\modmult_1/xin[611] ), .CLK(clk), .RST(
        start_in[0]), .I(c[612]), .Q(\modmult_1/xin[612] ) );
  DFF \modmult_1/xreg_reg[611]  ( .D(\modmult_1/xin[610] ), .CLK(clk), .RST(
        start_in[0]), .I(c[611]), .Q(\modmult_1/xin[611] ) );
  DFF \modmult_1/xreg_reg[610]  ( .D(\modmult_1/xin[609] ), .CLK(clk), .RST(
        start_in[0]), .I(c[610]), .Q(\modmult_1/xin[610] ) );
  DFF \modmult_1/xreg_reg[609]  ( .D(\modmult_1/xin[608] ), .CLK(clk), .RST(
        start_in[0]), .I(c[609]), .Q(\modmult_1/xin[609] ) );
  DFF \modmult_1/xreg_reg[608]  ( .D(\modmult_1/xin[607] ), .CLK(clk), .RST(
        start_in[0]), .I(c[608]), .Q(\modmult_1/xin[608] ) );
  DFF \modmult_1/xreg_reg[607]  ( .D(\modmult_1/xin[606] ), .CLK(clk), .RST(
        start_in[0]), .I(c[607]), .Q(\modmult_1/xin[607] ) );
  DFF \modmult_1/xreg_reg[606]  ( .D(\modmult_1/xin[605] ), .CLK(clk), .RST(
        start_in[0]), .I(c[606]), .Q(\modmult_1/xin[606] ) );
  DFF \modmult_1/xreg_reg[605]  ( .D(\modmult_1/xin[604] ), .CLK(clk), .RST(
        start_in[0]), .I(c[605]), .Q(\modmult_1/xin[605] ) );
  DFF \modmult_1/xreg_reg[604]  ( .D(\modmult_1/xin[603] ), .CLK(clk), .RST(
        start_in[0]), .I(c[604]), .Q(\modmult_1/xin[604] ) );
  DFF \modmult_1/xreg_reg[603]  ( .D(\modmult_1/xin[602] ), .CLK(clk), .RST(
        start_in[0]), .I(c[603]), .Q(\modmult_1/xin[603] ) );
  DFF \modmult_1/xreg_reg[602]  ( .D(\modmult_1/xin[601] ), .CLK(clk), .RST(
        start_in[0]), .I(c[602]), .Q(\modmult_1/xin[602] ) );
  DFF \modmult_1/xreg_reg[601]  ( .D(\modmult_1/xin[600] ), .CLK(clk), .RST(
        start_in[0]), .I(c[601]), .Q(\modmult_1/xin[601] ) );
  DFF \modmult_1/xreg_reg[600]  ( .D(\modmult_1/xin[599] ), .CLK(clk), .RST(
        start_in[0]), .I(c[600]), .Q(\modmult_1/xin[600] ) );
  DFF \modmult_1/xreg_reg[599]  ( .D(\modmult_1/xin[598] ), .CLK(clk), .RST(
        start_in[0]), .I(c[599]), .Q(\modmult_1/xin[599] ) );
  DFF \modmult_1/xreg_reg[598]  ( .D(\modmult_1/xin[597] ), .CLK(clk), .RST(
        start_in[0]), .I(c[598]), .Q(\modmult_1/xin[598] ) );
  DFF \modmult_1/xreg_reg[597]  ( .D(\modmult_1/xin[596] ), .CLK(clk), .RST(
        start_in[0]), .I(c[597]), .Q(\modmult_1/xin[597] ) );
  DFF \modmult_1/xreg_reg[596]  ( .D(\modmult_1/xin[595] ), .CLK(clk), .RST(
        start_in[0]), .I(c[596]), .Q(\modmult_1/xin[596] ) );
  DFF \modmult_1/xreg_reg[595]  ( .D(\modmult_1/xin[594] ), .CLK(clk), .RST(
        start_in[0]), .I(c[595]), .Q(\modmult_1/xin[595] ) );
  DFF \modmult_1/xreg_reg[594]  ( .D(\modmult_1/xin[593] ), .CLK(clk), .RST(
        start_in[0]), .I(c[594]), .Q(\modmult_1/xin[594] ) );
  DFF \modmult_1/xreg_reg[593]  ( .D(\modmult_1/xin[592] ), .CLK(clk), .RST(
        start_in[0]), .I(c[593]), .Q(\modmult_1/xin[593] ) );
  DFF \modmult_1/xreg_reg[592]  ( .D(\modmult_1/xin[591] ), .CLK(clk), .RST(
        start_in[0]), .I(c[592]), .Q(\modmult_1/xin[592] ) );
  DFF \modmult_1/xreg_reg[591]  ( .D(\modmult_1/xin[590] ), .CLK(clk), .RST(
        start_in[0]), .I(c[591]), .Q(\modmult_1/xin[591] ) );
  DFF \modmult_1/xreg_reg[590]  ( .D(\modmult_1/xin[589] ), .CLK(clk), .RST(
        start_in[0]), .I(c[590]), .Q(\modmult_1/xin[590] ) );
  DFF \modmult_1/xreg_reg[589]  ( .D(\modmult_1/xin[588] ), .CLK(clk), .RST(
        start_in[0]), .I(c[589]), .Q(\modmult_1/xin[589] ) );
  DFF \modmult_1/xreg_reg[588]  ( .D(\modmult_1/xin[587] ), .CLK(clk), .RST(
        start_in[0]), .I(c[588]), .Q(\modmult_1/xin[588] ) );
  DFF \modmult_1/xreg_reg[587]  ( .D(\modmult_1/xin[586] ), .CLK(clk), .RST(
        start_in[0]), .I(c[587]), .Q(\modmult_1/xin[587] ) );
  DFF \modmult_1/xreg_reg[586]  ( .D(\modmult_1/xin[585] ), .CLK(clk), .RST(
        start_in[0]), .I(c[586]), .Q(\modmult_1/xin[586] ) );
  DFF \modmult_1/xreg_reg[585]  ( .D(\modmult_1/xin[584] ), .CLK(clk), .RST(
        start_in[0]), .I(c[585]), .Q(\modmult_1/xin[585] ) );
  DFF \modmult_1/xreg_reg[584]  ( .D(\modmult_1/xin[583] ), .CLK(clk), .RST(
        start_in[0]), .I(c[584]), .Q(\modmult_1/xin[584] ) );
  DFF \modmult_1/xreg_reg[583]  ( .D(\modmult_1/xin[582] ), .CLK(clk), .RST(
        start_in[0]), .I(c[583]), .Q(\modmult_1/xin[583] ) );
  DFF \modmult_1/xreg_reg[582]  ( .D(\modmult_1/xin[581] ), .CLK(clk), .RST(
        start_in[0]), .I(c[582]), .Q(\modmult_1/xin[582] ) );
  DFF \modmult_1/xreg_reg[581]  ( .D(\modmult_1/xin[580] ), .CLK(clk), .RST(
        start_in[0]), .I(c[581]), .Q(\modmult_1/xin[581] ) );
  DFF \modmult_1/xreg_reg[580]  ( .D(\modmult_1/xin[579] ), .CLK(clk), .RST(
        start_in[0]), .I(c[580]), .Q(\modmult_1/xin[580] ) );
  DFF \modmult_1/xreg_reg[579]  ( .D(\modmult_1/xin[578] ), .CLK(clk), .RST(
        start_in[0]), .I(c[579]), .Q(\modmult_1/xin[579] ) );
  DFF \modmult_1/xreg_reg[578]  ( .D(\modmult_1/xin[577] ), .CLK(clk), .RST(
        start_in[0]), .I(c[578]), .Q(\modmult_1/xin[578] ) );
  DFF \modmult_1/xreg_reg[577]  ( .D(\modmult_1/xin[576] ), .CLK(clk), .RST(
        start_in[0]), .I(c[577]), .Q(\modmult_1/xin[577] ) );
  DFF \modmult_1/xreg_reg[576]  ( .D(\modmult_1/xin[575] ), .CLK(clk), .RST(
        start_in[0]), .I(c[576]), .Q(\modmult_1/xin[576] ) );
  DFF \modmult_1/xreg_reg[575]  ( .D(\modmult_1/xin[574] ), .CLK(clk), .RST(
        start_in[0]), .I(c[575]), .Q(\modmult_1/xin[575] ) );
  DFF \modmult_1/xreg_reg[574]  ( .D(\modmult_1/xin[573] ), .CLK(clk), .RST(
        start_in[0]), .I(c[574]), .Q(\modmult_1/xin[574] ) );
  DFF \modmult_1/xreg_reg[573]  ( .D(\modmult_1/xin[572] ), .CLK(clk), .RST(
        start_in[0]), .I(c[573]), .Q(\modmult_1/xin[573] ) );
  DFF \modmult_1/xreg_reg[572]  ( .D(\modmult_1/xin[571] ), .CLK(clk), .RST(
        start_in[0]), .I(c[572]), .Q(\modmult_1/xin[572] ) );
  DFF \modmult_1/xreg_reg[571]  ( .D(\modmult_1/xin[570] ), .CLK(clk), .RST(
        start_in[0]), .I(c[571]), .Q(\modmult_1/xin[571] ) );
  DFF \modmult_1/xreg_reg[570]  ( .D(\modmult_1/xin[569] ), .CLK(clk), .RST(
        start_in[0]), .I(c[570]), .Q(\modmult_1/xin[570] ) );
  DFF \modmult_1/xreg_reg[569]  ( .D(\modmult_1/xin[568] ), .CLK(clk), .RST(
        start_in[0]), .I(c[569]), .Q(\modmult_1/xin[569] ) );
  DFF \modmult_1/xreg_reg[568]  ( .D(\modmult_1/xin[567] ), .CLK(clk), .RST(
        start_in[0]), .I(c[568]), .Q(\modmult_1/xin[568] ) );
  DFF \modmult_1/xreg_reg[567]  ( .D(\modmult_1/xin[566] ), .CLK(clk), .RST(
        start_in[0]), .I(c[567]), .Q(\modmult_1/xin[567] ) );
  DFF \modmult_1/xreg_reg[566]  ( .D(\modmult_1/xin[565] ), .CLK(clk), .RST(
        start_in[0]), .I(c[566]), .Q(\modmult_1/xin[566] ) );
  DFF \modmult_1/xreg_reg[565]  ( .D(\modmult_1/xin[564] ), .CLK(clk), .RST(
        start_in[0]), .I(c[565]), .Q(\modmult_1/xin[565] ) );
  DFF \modmult_1/xreg_reg[564]  ( .D(\modmult_1/xin[563] ), .CLK(clk), .RST(
        start_in[0]), .I(c[564]), .Q(\modmult_1/xin[564] ) );
  DFF \modmult_1/xreg_reg[563]  ( .D(\modmult_1/xin[562] ), .CLK(clk), .RST(
        start_in[0]), .I(c[563]), .Q(\modmult_1/xin[563] ) );
  DFF \modmult_1/xreg_reg[562]  ( .D(\modmult_1/xin[561] ), .CLK(clk), .RST(
        start_in[0]), .I(c[562]), .Q(\modmult_1/xin[562] ) );
  DFF \modmult_1/xreg_reg[561]  ( .D(\modmult_1/xin[560] ), .CLK(clk), .RST(
        start_in[0]), .I(c[561]), .Q(\modmult_1/xin[561] ) );
  DFF \modmult_1/xreg_reg[560]  ( .D(\modmult_1/xin[559] ), .CLK(clk), .RST(
        start_in[0]), .I(c[560]), .Q(\modmult_1/xin[560] ) );
  DFF \modmult_1/xreg_reg[559]  ( .D(\modmult_1/xin[558] ), .CLK(clk), .RST(
        start_in[0]), .I(c[559]), .Q(\modmult_1/xin[559] ) );
  DFF \modmult_1/xreg_reg[558]  ( .D(\modmult_1/xin[557] ), .CLK(clk), .RST(
        start_in[0]), .I(c[558]), .Q(\modmult_1/xin[558] ) );
  DFF \modmult_1/xreg_reg[557]  ( .D(\modmult_1/xin[556] ), .CLK(clk), .RST(
        start_in[0]), .I(c[557]), .Q(\modmult_1/xin[557] ) );
  DFF \modmult_1/xreg_reg[556]  ( .D(\modmult_1/xin[555] ), .CLK(clk), .RST(
        start_in[0]), .I(c[556]), .Q(\modmult_1/xin[556] ) );
  DFF \modmult_1/xreg_reg[555]  ( .D(\modmult_1/xin[554] ), .CLK(clk), .RST(
        start_in[0]), .I(c[555]), .Q(\modmult_1/xin[555] ) );
  DFF \modmult_1/xreg_reg[554]  ( .D(\modmult_1/xin[553] ), .CLK(clk), .RST(
        start_in[0]), .I(c[554]), .Q(\modmult_1/xin[554] ) );
  DFF \modmult_1/xreg_reg[553]  ( .D(\modmult_1/xin[552] ), .CLK(clk), .RST(
        start_in[0]), .I(c[553]), .Q(\modmult_1/xin[553] ) );
  DFF \modmult_1/xreg_reg[552]  ( .D(\modmult_1/xin[551] ), .CLK(clk), .RST(
        start_in[0]), .I(c[552]), .Q(\modmult_1/xin[552] ) );
  DFF \modmult_1/xreg_reg[551]  ( .D(\modmult_1/xin[550] ), .CLK(clk), .RST(
        start_in[0]), .I(c[551]), .Q(\modmult_1/xin[551] ) );
  DFF \modmult_1/xreg_reg[550]  ( .D(\modmult_1/xin[549] ), .CLK(clk), .RST(
        start_in[0]), .I(c[550]), .Q(\modmult_1/xin[550] ) );
  DFF \modmult_1/xreg_reg[549]  ( .D(\modmult_1/xin[548] ), .CLK(clk), .RST(
        start_in[0]), .I(c[549]), .Q(\modmult_1/xin[549] ) );
  DFF \modmult_1/xreg_reg[548]  ( .D(\modmult_1/xin[547] ), .CLK(clk), .RST(
        start_in[0]), .I(c[548]), .Q(\modmult_1/xin[548] ) );
  DFF \modmult_1/xreg_reg[547]  ( .D(\modmult_1/xin[546] ), .CLK(clk), .RST(
        start_in[0]), .I(c[547]), .Q(\modmult_1/xin[547] ) );
  DFF \modmult_1/xreg_reg[546]  ( .D(\modmult_1/xin[545] ), .CLK(clk), .RST(
        start_in[0]), .I(c[546]), .Q(\modmult_1/xin[546] ) );
  DFF \modmult_1/xreg_reg[545]  ( .D(\modmult_1/xin[544] ), .CLK(clk), .RST(
        start_in[0]), .I(c[545]), .Q(\modmult_1/xin[545] ) );
  DFF \modmult_1/xreg_reg[544]  ( .D(\modmult_1/xin[543] ), .CLK(clk), .RST(
        start_in[0]), .I(c[544]), .Q(\modmult_1/xin[544] ) );
  DFF \modmult_1/xreg_reg[543]  ( .D(\modmult_1/xin[542] ), .CLK(clk), .RST(
        start_in[0]), .I(c[543]), .Q(\modmult_1/xin[543] ) );
  DFF \modmult_1/xreg_reg[542]  ( .D(\modmult_1/xin[541] ), .CLK(clk), .RST(
        start_in[0]), .I(c[542]), .Q(\modmult_1/xin[542] ) );
  DFF \modmult_1/xreg_reg[541]  ( .D(\modmult_1/xin[540] ), .CLK(clk), .RST(
        start_in[0]), .I(c[541]), .Q(\modmult_1/xin[541] ) );
  DFF \modmult_1/xreg_reg[540]  ( .D(\modmult_1/xin[539] ), .CLK(clk), .RST(
        start_in[0]), .I(c[540]), .Q(\modmult_1/xin[540] ) );
  DFF \modmult_1/xreg_reg[539]  ( .D(\modmult_1/xin[538] ), .CLK(clk), .RST(
        start_in[0]), .I(c[539]), .Q(\modmult_1/xin[539] ) );
  DFF \modmult_1/xreg_reg[538]  ( .D(\modmult_1/xin[537] ), .CLK(clk), .RST(
        start_in[0]), .I(c[538]), .Q(\modmult_1/xin[538] ) );
  DFF \modmult_1/xreg_reg[537]  ( .D(\modmult_1/xin[536] ), .CLK(clk), .RST(
        start_in[0]), .I(c[537]), .Q(\modmult_1/xin[537] ) );
  DFF \modmult_1/xreg_reg[536]  ( .D(\modmult_1/xin[535] ), .CLK(clk), .RST(
        start_in[0]), .I(c[536]), .Q(\modmult_1/xin[536] ) );
  DFF \modmult_1/xreg_reg[535]  ( .D(\modmult_1/xin[534] ), .CLK(clk), .RST(
        start_in[0]), .I(c[535]), .Q(\modmult_1/xin[535] ) );
  DFF \modmult_1/xreg_reg[534]  ( .D(\modmult_1/xin[533] ), .CLK(clk), .RST(
        start_in[0]), .I(c[534]), .Q(\modmult_1/xin[534] ) );
  DFF \modmult_1/xreg_reg[533]  ( .D(\modmult_1/xin[532] ), .CLK(clk), .RST(
        start_in[0]), .I(c[533]), .Q(\modmult_1/xin[533] ) );
  DFF \modmult_1/xreg_reg[532]  ( .D(\modmult_1/xin[531] ), .CLK(clk), .RST(
        start_in[0]), .I(c[532]), .Q(\modmult_1/xin[532] ) );
  DFF \modmult_1/xreg_reg[531]  ( .D(\modmult_1/xin[530] ), .CLK(clk), .RST(
        start_in[0]), .I(c[531]), .Q(\modmult_1/xin[531] ) );
  DFF \modmult_1/xreg_reg[530]  ( .D(\modmult_1/xin[529] ), .CLK(clk), .RST(
        start_in[0]), .I(c[530]), .Q(\modmult_1/xin[530] ) );
  DFF \modmult_1/xreg_reg[529]  ( .D(\modmult_1/xin[528] ), .CLK(clk), .RST(
        start_in[0]), .I(c[529]), .Q(\modmult_1/xin[529] ) );
  DFF \modmult_1/xreg_reg[528]  ( .D(\modmult_1/xin[527] ), .CLK(clk), .RST(
        start_in[0]), .I(c[528]), .Q(\modmult_1/xin[528] ) );
  DFF \modmult_1/xreg_reg[527]  ( .D(\modmult_1/xin[526] ), .CLK(clk), .RST(
        start_in[0]), .I(c[527]), .Q(\modmult_1/xin[527] ) );
  DFF \modmult_1/xreg_reg[526]  ( .D(\modmult_1/xin[525] ), .CLK(clk), .RST(
        start_in[0]), .I(c[526]), .Q(\modmult_1/xin[526] ) );
  DFF \modmult_1/xreg_reg[525]  ( .D(\modmult_1/xin[524] ), .CLK(clk), .RST(
        start_in[0]), .I(c[525]), .Q(\modmult_1/xin[525] ) );
  DFF \modmult_1/xreg_reg[524]  ( .D(\modmult_1/xin[523] ), .CLK(clk), .RST(
        start_in[0]), .I(c[524]), .Q(\modmult_1/xin[524] ) );
  DFF \modmult_1/xreg_reg[523]  ( .D(\modmult_1/xin[522] ), .CLK(clk), .RST(
        start_in[0]), .I(c[523]), .Q(\modmult_1/xin[523] ) );
  DFF \modmult_1/xreg_reg[522]  ( .D(\modmult_1/xin[521] ), .CLK(clk), .RST(
        start_in[0]), .I(c[522]), .Q(\modmult_1/xin[522] ) );
  DFF \modmult_1/xreg_reg[521]  ( .D(\modmult_1/xin[520] ), .CLK(clk), .RST(
        start_in[0]), .I(c[521]), .Q(\modmult_1/xin[521] ) );
  DFF \modmult_1/xreg_reg[520]  ( .D(\modmult_1/xin[519] ), .CLK(clk), .RST(
        start_in[0]), .I(c[520]), .Q(\modmult_1/xin[520] ) );
  DFF \modmult_1/xreg_reg[519]  ( .D(\modmult_1/xin[518] ), .CLK(clk), .RST(
        start_in[0]), .I(c[519]), .Q(\modmult_1/xin[519] ) );
  DFF \modmult_1/xreg_reg[518]  ( .D(\modmult_1/xin[517] ), .CLK(clk), .RST(
        start_in[0]), .I(c[518]), .Q(\modmult_1/xin[518] ) );
  DFF \modmult_1/xreg_reg[517]  ( .D(\modmult_1/xin[516] ), .CLK(clk), .RST(
        start_in[0]), .I(c[517]), .Q(\modmult_1/xin[517] ) );
  DFF \modmult_1/xreg_reg[516]  ( .D(\modmult_1/xin[515] ), .CLK(clk), .RST(
        start_in[0]), .I(c[516]), .Q(\modmult_1/xin[516] ) );
  DFF \modmult_1/xreg_reg[515]  ( .D(\modmult_1/xin[514] ), .CLK(clk), .RST(
        start_in[0]), .I(c[515]), .Q(\modmult_1/xin[515] ) );
  DFF \modmult_1/xreg_reg[514]  ( .D(\modmult_1/xin[513] ), .CLK(clk), .RST(
        start_in[0]), .I(c[514]), .Q(\modmult_1/xin[514] ) );
  DFF \modmult_1/xreg_reg[513]  ( .D(\modmult_1/xin[512] ), .CLK(clk), .RST(
        start_in[0]), .I(c[513]), .Q(\modmult_1/xin[513] ) );
  DFF \modmult_1/xreg_reg[512]  ( .D(\modmult_1/xin[511] ), .CLK(clk), .RST(
        start_in[0]), .I(c[512]), .Q(\modmult_1/xin[512] ) );
  DFF \modmult_1/xreg_reg[511]  ( .D(\modmult_1/xin[510] ), .CLK(clk), .RST(
        start_in[0]), .I(c[511]), .Q(\modmult_1/xin[511] ) );
  DFF \modmult_1/xreg_reg[510]  ( .D(\modmult_1/xin[509] ), .CLK(clk), .RST(
        start_in[0]), .I(c[510]), .Q(\modmult_1/xin[510] ) );
  DFF \modmult_1/xreg_reg[509]  ( .D(\modmult_1/xin[508] ), .CLK(clk), .RST(
        start_in[0]), .I(c[509]), .Q(\modmult_1/xin[509] ) );
  DFF \modmult_1/xreg_reg[508]  ( .D(\modmult_1/xin[507] ), .CLK(clk), .RST(
        start_in[0]), .I(c[508]), .Q(\modmult_1/xin[508] ) );
  DFF \modmult_1/xreg_reg[507]  ( .D(\modmult_1/xin[506] ), .CLK(clk), .RST(
        start_in[0]), .I(c[507]), .Q(\modmult_1/xin[507] ) );
  DFF \modmult_1/xreg_reg[506]  ( .D(\modmult_1/xin[505] ), .CLK(clk), .RST(
        start_in[0]), .I(c[506]), .Q(\modmult_1/xin[506] ) );
  DFF \modmult_1/xreg_reg[505]  ( .D(\modmult_1/xin[504] ), .CLK(clk), .RST(
        start_in[0]), .I(c[505]), .Q(\modmult_1/xin[505] ) );
  DFF \modmult_1/xreg_reg[504]  ( .D(\modmult_1/xin[503] ), .CLK(clk), .RST(
        start_in[0]), .I(c[504]), .Q(\modmult_1/xin[504] ) );
  DFF \modmult_1/xreg_reg[503]  ( .D(\modmult_1/xin[502] ), .CLK(clk), .RST(
        start_in[0]), .I(c[503]), .Q(\modmult_1/xin[503] ) );
  DFF \modmult_1/xreg_reg[502]  ( .D(\modmult_1/xin[501] ), .CLK(clk), .RST(
        start_in[0]), .I(c[502]), .Q(\modmult_1/xin[502] ) );
  DFF \modmult_1/xreg_reg[501]  ( .D(\modmult_1/xin[500] ), .CLK(clk), .RST(
        start_in[0]), .I(c[501]), .Q(\modmult_1/xin[501] ) );
  DFF \modmult_1/xreg_reg[500]  ( .D(\modmult_1/xin[499] ), .CLK(clk), .RST(
        start_in[0]), .I(c[500]), .Q(\modmult_1/xin[500] ) );
  DFF \modmult_1/xreg_reg[499]  ( .D(\modmult_1/xin[498] ), .CLK(clk), .RST(
        start_in[0]), .I(c[499]), .Q(\modmult_1/xin[499] ) );
  DFF \modmult_1/xreg_reg[498]  ( .D(\modmult_1/xin[497] ), .CLK(clk), .RST(
        start_in[0]), .I(c[498]), .Q(\modmult_1/xin[498] ) );
  DFF \modmult_1/xreg_reg[497]  ( .D(\modmult_1/xin[496] ), .CLK(clk), .RST(
        start_in[0]), .I(c[497]), .Q(\modmult_1/xin[497] ) );
  DFF \modmult_1/xreg_reg[496]  ( .D(\modmult_1/xin[495] ), .CLK(clk), .RST(
        start_in[0]), .I(c[496]), .Q(\modmult_1/xin[496] ) );
  DFF \modmult_1/xreg_reg[495]  ( .D(\modmult_1/xin[494] ), .CLK(clk), .RST(
        start_in[0]), .I(c[495]), .Q(\modmult_1/xin[495] ) );
  DFF \modmult_1/xreg_reg[494]  ( .D(\modmult_1/xin[493] ), .CLK(clk), .RST(
        start_in[0]), .I(c[494]), .Q(\modmult_1/xin[494] ) );
  DFF \modmult_1/xreg_reg[493]  ( .D(\modmult_1/xin[492] ), .CLK(clk), .RST(
        start_in[0]), .I(c[493]), .Q(\modmult_1/xin[493] ) );
  DFF \modmult_1/xreg_reg[492]  ( .D(\modmult_1/xin[491] ), .CLK(clk), .RST(
        start_in[0]), .I(c[492]), .Q(\modmult_1/xin[492] ) );
  DFF \modmult_1/xreg_reg[491]  ( .D(\modmult_1/xin[490] ), .CLK(clk), .RST(
        start_in[0]), .I(c[491]), .Q(\modmult_1/xin[491] ) );
  DFF \modmult_1/xreg_reg[490]  ( .D(\modmult_1/xin[489] ), .CLK(clk), .RST(
        start_in[0]), .I(c[490]), .Q(\modmult_1/xin[490] ) );
  DFF \modmult_1/xreg_reg[489]  ( .D(\modmult_1/xin[488] ), .CLK(clk), .RST(
        start_in[0]), .I(c[489]), .Q(\modmult_1/xin[489] ) );
  DFF \modmult_1/xreg_reg[488]  ( .D(\modmult_1/xin[487] ), .CLK(clk), .RST(
        start_in[0]), .I(c[488]), .Q(\modmult_1/xin[488] ) );
  DFF \modmult_1/xreg_reg[487]  ( .D(\modmult_1/xin[486] ), .CLK(clk), .RST(
        start_in[0]), .I(c[487]), .Q(\modmult_1/xin[487] ) );
  DFF \modmult_1/xreg_reg[486]  ( .D(\modmult_1/xin[485] ), .CLK(clk), .RST(
        start_in[0]), .I(c[486]), .Q(\modmult_1/xin[486] ) );
  DFF \modmult_1/xreg_reg[485]  ( .D(\modmult_1/xin[484] ), .CLK(clk), .RST(
        start_in[0]), .I(c[485]), .Q(\modmult_1/xin[485] ) );
  DFF \modmult_1/xreg_reg[484]  ( .D(\modmult_1/xin[483] ), .CLK(clk), .RST(
        start_in[0]), .I(c[484]), .Q(\modmult_1/xin[484] ) );
  DFF \modmult_1/xreg_reg[483]  ( .D(\modmult_1/xin[482] ), .CLK(clk), .RST(
        start_in[0]), .I(c[483]), .Q(\modmult_1/xin[483] ) );
  DFF \modmult_1/xreg_reg[482]  ( .D(\modmult_1/xin[481] ), .CLK(clk), .RST(
        start_in[0]), .I(c[482]), .Q(\modmult_1/xin[482] ) );
  DFF \modmult_1/xreg_reg[481]  ( .D(\modmult_1/xin[480] ), .CLK(clk), .RST(
        start_in[0]), .I(c[481]), .Q(\modmult_1/xin[481] ) );
  DFF \modmult_1/xreg_reg[480]  ( .D(\modmult_1/xin[479] ), .CLK(clk), .RST(
        start_in[0]), .I(c[480]), .Q(\modmult_1/xin[480] ) );
  DFF \modmult_1/xreg_reg[479]  ( .D(\modmult_1/xin[478] ), .CLK(clk), .RST(
        start_in[0]), .I(c[479]), .Q(\modmult_1/xin[479] ) );
  DFF \modmult_1/xreg_reg[478]  ( .D(\modmult_1/xin[477] ), .CLK(clk), .RST(
        start_in[0]), .I(c[478]), .Q(\modmult_1/xin[478] ) );
  DFF \modmult_1/xreg_reg[477]  ( .D(\modmult_1/xin[476] ), .CLK(clk), .RST(
        start_in[0]), .I(c[477]), .Q(\modmult_1/xin[477] ) );
  DFF \modmult_1/xreg_reg[476]  ( .D(\modmult_1/xin[475] ), .CLK(clk), .RST(
        start_in[0]), .I(c[476]), .Q(\modmult_1/xin[476] ) );
  DFF \modmult_1/xreg_reg[475]  ( .D(\modmult_1/xin[474] ), .CLK(clk), .RST(
        start_in[0]), .I(c[475]), .Q(\modmult_1/xin[475] ) );
  DFF \modmult_1/xreg_reg[474]  ( .D(\modmult_1/xin[473] ), .CLK(clk), .RST(
        start_in[0]), .I(c[474]), .Q(\modmult_1/xin[474] ) );
  DFF \modmult_1/xreg_reg[473]  ( .D(\modmult_1/xin[472] ), .CLK(clk), .RST(
        start_in[0]), .I(c[473]), .Q(\modmult_1/xin[473] ) );
  DFF \modmult_1/xreg_reg[472]  ( .D(\modmult_1/xin[471] ), .CLK(clk), .RST(
        start_in[0]), .I(c[472]), .Q(\modmult_1/xin[472] ) );
  DFF \modmult_1/xreg_reg[471]  ( .D(\modmult_1/xin[470] ), .CLK(clk), .RST(
        start_in[0]), .I(c[471]), .Q(\modmult_1/xin[471] ) );
  DFF \modmult_1/xreg_reg[470]  ( .D(\modmult_1/xin[469] ), .CLK(clk), .RST(
        start_in[0]), .I(c[470]), .Q(\modmult_1/xin[470] ) );
  DFF \modmult_1/xreg_reg[469]  ( .D(\modmult_1/xin[468] ), .CLK(clk), .RST(
        start_in[0]), .I(c[469]), .Q(\modmult_1/xin[469] ) );
  DFF \modmult_1/xreg_reg[468]  ( .D(\modmult_1/xin[467] ), .CLK(clk), .RST(
        start_in[0]), .I(c[468]), .Q(\modmult_1/xin[468] ) );
  DFF \modmult_1/xreg_reg[467]  ( .D(\modmult_1/xin[466] ), .CLK(clk), .RST(
        start_in[0]), .I(c[467]), .Q(\modmult_1/xin[467] ) );
  DFF \modmult_1/xreg_reg[466]  ( .D(\modmult_1/xin[465] ), .CLK(clk), .RST(
        start_in[0]), .I(c[466]), .Q(\modmult_1/xin[466] ) );
  DFF \modmult_1/xreg_reg[465]  ( .D(\modmult_1/xin[464] ), .CLK(clk), .RST(
        start_in[0]), .I(c[465]), .Q(\modmult_1/xin[465] ) );
  DFF \modmult_1/xreg_reg[464]  ( .D(\modmult_1/xin[463] ), .CLK(clk), .RST(
        start_in[0]), .I(c[464]), .Q(\modmult_1/xin[464] ) );
  DFF \modmult_1/xreg_reg[463]  ( .D(\modmult_1/xin[462] ), .CLK(clk), .RST(
        start_in[0]), .I(c[463]), .Q(\modmult_1/xin[463] ) );
  DFF \modmult_1/xreg_reg[462]  ( .D(\modmult_1/xin[461] ), .CLK(clk), .RST(
        start_in[0]), .I(c[462]), .Q(\modmult_1/xin[462] ) );
  DFF \modmult_1/xreg_reg[461]  ( .D(\modmult_1/xin[460] ), .CLK(clk), .RST(
        start_in[0]), .I(c[461]), .Q(\modmult_1/xin[461] ) );
  DFF \modmult_1/xreg_reg[460]  ( .D(\modmult_1/xin[459] ), .CLK(clk), .RST(
        start_in[0]), .I(c[460]), .Q(\modmult_1/xin[460] ) );
  DFF \modmult_1/xreg_reg[459]  ( .D(\modmult_1/xin[458] ), .CLK(clk), .RST(
        start_in[0]), .I(c[459]), .Q(\modmult_1/xin[459] ) );
  DFF \modmult_1/xreg_reg[458]  ( .D(\modmult_1/xin[457] ), .CLK(clk), .RST(
        start_in[0]), .I(c[458]), .Q(\modmult_1/xin[458] ) );
  DFF \modmult_1/xreg_reg[457]  ( .D(\modmult_1/xin[456] ), .CLK(clk), .RST(
        start_in[0]), .I(c[457]), .Q(\modmult_1/xin[457] ) );
  DFF \modmult_1/xreg_reg[456]  ( .D(\modmult_1/xin[455] ), .CLK(clk), .RST(
        start_in[0]), .I(c[456]), .Q(\modmult_1/xin[456] ) );
  DFF \modmult_1/xreg_reg[455]  ( .D(\modmult_1/xin[454] ), .CLK(clk), .RST(
        start_in[0]), .I(c[455]), .Q(\modmult_1/xin[455] ) );
  DFF \modmult_1/xreg_reg[454]  ( .D(\modmult_1/xin[453] ), .CLK(clk), .RST(
        start_in[0]), .I(c[454]), .Q(\modmult_1/xin[454] ) );
  DFF \modmult_1/xreg_reg[453]  ( .D(\modmult_1/xin[452] ), .CLK(clk), .RST(
        start_in[0]), .I(c[453]), .Q(\modmult_1/xin[453] ) );
  DFF \modmult_1/xreg_reg[452]  ( .D(\modmult_1/xin[451] ), .CLK(clk), .RST(
        start_in[0]), .I(c[452]), .Q(\modmult_1/xin[452] ) );
  DFF \modmult_1/xreg_reg[451]  ( .D(\modmult_1/xin[450] ), .CLK(clk), .RST(
        start_in[0]), .I(c[451]), .Q(\modmult_1/xin[451] ) );
  DFF \modmult_1/xreg_reg[450]  ( .D(\modmult_1/xin[449] ), .CLK(clk), .RST(
        start_in[0]), .I(c[450]), .Q(\modmult_1/xin[450] ) );
  DFF \modmult_1/xreg_reg[449]  ( .D(\modmult_1/xin[448] ), .CLK(clk), .RST(
        start_in[0]), .I(c[449]), .Q(\modmult_1/xin[449] ) );
  DFF \modmult_1/xreg_reg[448]  ( .D(\modmult_1/xin[447] ), .CLK(clk), .RST(
        start_in[0]), .I(c[448]), .Q(\modmult_1/xin[448] ) );
  DFF \modmult_1/xreg_reg[447]  ( .D(\modmult_1/xin[446] ), .CLK(clk), .RST(
        start_in[0]), .I(c[447]), .Q(\modmult_1/xin[447] ) );
  DFF \modmult_1/xreg_reg[446]  ( .D(\modmult_1/xin[445] ), .CLK(clk), .RST(
        start_in[0]), .I(c[446]), .Q(\modmult_1/xin[446] ) );
  DFF \modmult_1/xreg_reg[445]  ( .D(\modmult_1/xin[444] ), .CLK(clk), .RST(
        start_in[0]), .I(c[445]), .Q(\modmult_1/xin[445] ) );
  DFF \modmult_1/xreg_reg[444]  ( .D(\modmult_1/xin[443] ), .CLK(clk), .RST(
        start_in[0]), .I(c[444]), .Q(\modmult_1/xin[444] ) );
  DFF \modmult_1/xreg_reg[443]  ( .D(\modmult_1/xin[442] ), .CLK(clk), .RST(
        start_in[0]), .I(c[443]), .Q(\modmult_1/xin[443] ) );
  DFF \modmult_1/xreg_reg[442]  ( .D(\modmult_1/xin[441] ), .CLK(clk), .RST(
        start_in[0]), .I(c[442]), .Q(\modmult_1/xin[442] ) );
  DFF \modmult_1/xreg_reg[441]  ( .D(\modmult_1/xin[440] ), .CLK(clk), .RST(
        start_in[0]), .I(c[441]), .Q(\modmult_1/xin[441] ) );
  DFF \modmult_1/xreg_reg[440]  ( .D(\modmult_1/xin[439] ), .CLK(clk), .RST(
        start_in[0]), .I(c[440]), .Q(\modmult_1/xin[440] ) );
  DFF \modmult_1/xreg_reg[439]  ( .D(\modmult_1/xin[438] ), .CLK(clk), .RST(
        start_in[0]), .I(c[439]), .Q(\modmult_1/xin[439] ) );
  DFF \modmult_1/xreg_reg[438]  ( .D(\modmult_1/xin[437] ), .CLK(clk), .RST(
        start_in[0]), .I(c[438]), .Q(\modmult_1/xin[438] ) );
  DFF \modmult_1/xreg_reg[437]  ( .D(\modmult_1/xin[436] ), .CLK(clk), .RST(
        start_in[0]), .I(c[437]), .Q(\modmult_1/xin[437] ) );
  DFF \modmult_1/xreg_reg[436]  ( .D(\modmult_1/xin[435] ), .CLK(clk), .RST(
        start_in[0]), .I(c[436]), .Q(\modmult_1/xin[436] ) );
  DFF \modmult_1/xreg_reg[435]  ( .D(\modmult_1/xin[434] ), .CLK(clk), .RST(
        start_in[0]), .I(c[435]), .Q(\modmult_1/xin[435] ) );
  DFF \modmult_1/xreg_reg[434]  ( .D(\modmult_1/xin[433] ), .CLK(clk), .RST(
        start_in[0]), .I(c[434]), .Q(\modmult_1/xin[434] ) );
  DFF \modmult_1/xreg_reg[433]  ( .D(\modmult_1/xin[432] ), .CLK(clk), .RST(
        start_in[0]), .I(c[433]), .Q(\modmult_1/xin[433] ) );
  DFF \modmult_1/xreg_reg[432]  ( .D(\modmult_1/xin[431] ), .CLK(clk), .RST(
        start_in[0]), .I(c[432]), .Q(\modmult_1/xin[432] ) );
  DFF \modmult_1/xreg_reg[431]  ( .D(\modmult_1/xin[430] ), .CLK(clk), .RST(
        start_in[0]), .I(c[431]), .Q(\modmult_1/xin[431] ) );
  DFF \modmult_1/xreg_reg[430]  ( .D(\modmult_1/xin[429] ), .CLK(clk), .RST(
        start_in[0]), .I(c[430]), .Q(\modmult_1/xin[430] ) );
  DFF \modmult_1/xreg_reg[429]  ( .D(\modmult_1/xin[428] ), .CLK(clk), .RST(
        start_in[0]), .I(c[429]), .Q(\modmult_1/xin[429] ) );
  DFF \modmult_1/xreg_reg[428]  ( .D(\modmult_1/xin[427] ), .CLK(clk), .RST(
        start_in[0]), .I(c[428]), .Q(\modmult_1/xin[428] ) );
  DFF \modmult_1/xreg_reg[427]  ( .D(\modmult_1/xin[426] ), .CLK(clk), .RST(
        start_in[0]), .I(c[427]), .Q(\modmult_1/xin[427] ) );
  DFF \modmult_1/xreg_reg[426]  ( .D(\modmult_1/xin[425] ), .CLK(clk), .RST(
        start_in[0]), .I(c[426]), .Q(\modmult_1/xin[426] ) );
  DFF \modmult_1/xreg_reg[425]  ( .D(\modmult_1/xin[424] ), .CLK(clk), .RST(
        start_in[0]), .I(c[425]), .Q(\modmult_1/xin[425] ) );
  DFF \modmult_1/xreg_reg[424]  ( .D(\modmult_1/xin[423] ), .CLK(clk), .RST(
        start_in[0]), .I(c[424]), .Q(\modmult_1/xin[424] ) );
  DFF \modmult_1/xreg_reg[423]  ( .D(\modmult_1/xin[422] ), .CLK(clk), .RST(
        start_in[0]), .I(c[423]), .Q(\modmult_1/xin[423] ) );
  DFF \modmult_1/xreg_reg[422]  ( .D(\modmult_1/xin[421] ), .CLK(clk), .RST(
        start_in[0]), .I(c[422]), .Q(\modmult_1/xin[422] ) );
  DFF \modmult_1/xreg_reg[421]  ( .D(\modmult_1/xin[420] ), .CLK(clk), .RST(
        start_in[0]), .I(c[421]), .Q(\modmult_1/xin[421] ) );
  DFF \modmult_1/xreg_reg[420]  ( .D(\modmult_1/xin[419] ), .CLK(clk), .RST(
        start_in[0]), .I(c[420]), .Q(\modmult_1/xin[420] ) );
  DFF \modmult_1/xreg_reg[419]  ( .D(\modmult_1/xin[418] ), .CLK(clk), .RST(
        start_in[0]), .I(c[419]), .Q(\modmult_1/xin[419] ) );
  DFF \modmult_1/xreg_reg[418]  ( .D(\modmult_1/xin[417] ), .CLK(clk), .RST(
        start_in[0]), .I(c[418]), .Q(\modmult_1/xin[418] ) );
  DFF \modmult_1/xreg_reg[417]  ( .D(\modmult_1/xin[416] ), .CLK(clk), .RST(
        start_in[0]), .I(c[417]), .Q(\modmult_1/xin[417] ) );
  DFF \modmult_1/xreg_reg[416]  ( .D(\modmult_1/xin[415] ), .CLK(clk), .RST(
        start_in[0]), .I(c[416]), .Q(\modmult_1/xin[416] ) );
  DFF \modmult_1/xreg_reg[415]  ( .D(\modmult_1/xin[414] ), .CLK(clk), .RST(
        start_in[0]), .I(c[415]), .Q(\modmult_1/xin[415] ) );
  DFF \modmult_1/xreg_reg[414]  ( .D(\modmult_1/xin[413] ), .CLK(clk), .RST(
        start_in[0]), .I(c[414]), .Q(\modmult_1/xin[414] ) );
  DFF \modmult_1/xreg_reg[413]  ( .D(\modmult_1/xin[412] ), .CLK(clk), .RST(
        start_in[0]), .I(c[413]), .Q(\modmult_1/xin[413] ) );
  DFF \modmult_1/xreg_reg[412]  ( .D(\modmult_1/xin[411] ), .CLK(clk), .RST(
        start_in[0]), .I(c[412]), .Q(\modmult_1/xin[412] ) );
  DFF \modmult_1/xreg_reg[411]  ( .D(\modmult_1/xin[410] ), .CLK(clk), .RST(
        start_in[0]), .I(c[411]), .Q(\modmult_1/xin[411] ) );
  DFF \modmult_1/xreg_reg[410]  ( .D(\modmult_1/xin[409] ), .CLK(clk), .RST(
        start_in[0]), .I(c[410]), .Q(\modmult_1/xin[410] ) );
  DFF \modmult_1/xreg_reg[409]  ( .D(\modmult_1/xin[408] ), .CLK(clk), .RST(
        start_in[0]), .I(c[409]), .Q(\modmult_1/xin[409] ) );
  DFF \modmult_1/xreg_reg[408]  ( .D(\modmult_1/xin[407] ), .CLK(clk), .RST(
        start_in[0]), .I(c[408]), .Q(\modmult_1/xin[408] ) );
  DFF \modmult_1/xreg_reg[407]  ( .D(\modmult_1/xin[406] ), .CLK(clk), .RST(
        start_in[0]), .I(c[407]), .Q(\modmult_1/xin[407] ) );
  DFF \modmult_1/xreg_reg[406]  ( .D(\modmult_1/xin[405] ), .CLK(clk), .RST(
        start_in[0]), .I(c[406]), .Q(\modmult_1/xin[406] ) );
  DFF \modmult_1/xreg_reg[405]  ( .D(\modmult_1/xin[404] ), .CLK(clk), .RST(
        start_in[0]), .I(c[405]), .Q(\modmult_1/xin[405] ) );
  DFF \modmult_1/xreg_reg[404]  ( .D(\modmult_1/xin[403] ), .CLK(clk), .RST(
        start_in[0]), .I(c[404]), .Q(\modmult_1/xin[404] ) );
  DFF \modmult_1/xreg_reg[403]  ( .D(\modmult_1/xin[402] ), .CLK(clk), .RST(
        start_in[0]), .I(c[403]), .Q(\modmult_1/xin[403] ) );
  DFF \modmult_1/xreg_reg[402]  ( .D(\modmult_1/xin[401] ), .CLK(clk), .RST(
        start_in[0]), .I(c[402]), .Q(\modmult_1/xin[402] ) );
  DFF \modmult_1/xreg_reg[401]  ( .D(\modmult_1/xin[400] ), .CLK(clk), .RST(
        start_in[0]), .I(c[401]), .Q(\modmult_1/xin[401] ) );
  DFF \modmult_1/xreg_reg[400]  ( .D(\modmult_1/xin[399] ), .CLK(clk), .RST(
        start_in[0]), .I(c[400]), .Q(\modmult_1/xin[400] ) );
  DFF \modmult_1/xreg_reg[399]  ( .D(\modmult_1/xin[398] ), .CLK(clk), .RST(
        start_in[0]), .I(c[399]), .Q(\modmult_1/xin[399] ) );
  DFF \modmult_1/xreg_reg[398]  ( .D(\modmult_1/xin[397] ), .CLK(clk), .RST(
        start_in[0]), .I(c[398]), .Q(\modmult_1/xin[398] ) );
  DFF \modmult_1/xreg_reg[397]  ( .D(\modmult_1/xin[396] ), .CLK(clk), .RST(
        start_in[0]), .I(c[397]), .Q(\modmult_1/xin[397] ) );
  DFF \modmult_1/xreg_reg[396]  ( .D(\modmult_1/xin[395] ), .CLK(clk), .RST(
        start_in[0]), .I(c[396]), .Q(\modmult_1/xin[396] ) );
  DFF \modmult_1/xreg_reg[395]  ( .D(\modmult_1/xin[394] ), .CLK(clk), .RST(
        start_in[0]), .I(c[395]), .Q(\modmult_1/xin[395] ) );
  DFF \modmult_1/xreg_reg[394]  ( .D(\modmult_1/xin[393] ), .CLK(clk), .RST(
        start_in[0]), .I(c[394]), .Q(\modmult_1/xin[394] ) );
  DFF \modmult_1/xreg_reg[393]  ( .D(\modmult_1/xin[392] ), .CLK(clk), .RST(
        start_in[0]), .I(c[393]), .Q(\modmult_1/xin[393] ) );
  DFF \modmult_1/xreg_reg[392]  ( .D(\modmult_1/xin[391] ), .CLK(clk), .RST(
        start_in[0]), .I(c[392]), .Q(\modmult_1/xin[392] ) );
  DFF \modmult_1/xreg_reg[391]  ( .D(\modmult_1/xin[390] ), .CLK(clk), .RST(
        start_in[0]), .I(c[391]), .Q(\modmult_1/xin[391] ) );
  DFF \modmult_1/xreg_reg[390]  ( .D(\modmult_1/xin[389] ), .CLK(clk), .RST(
        start_in[0]), .I(c[390]), .Q(\modmult_1/xin[390] ) );
  DFF \modmult_1/xreg_reg[389]  ( .D(\modmult_1/xin[388] ), .CLK(clk), .RST(
        start_in[0]), .I(c[389]), .Q(\modmult_1/xin[389] ) );
  DFF \modmult_1/xreg_reg[388]  ( .D(\modmult_1/xin[387] ), .CLK(clk), .RST(
        start_in[0]), .I(c[388]), .Q(\modmult_1/xin[388] ) );
  DFF \modmult_1/xreg_reg[387]  ( .D(\modmult_1/xin[386] ), .CLK(clk), .RST(
        start_in[0]), .I(c[387]), .Q(\modmult_1/xin[387] ) );
  DFF \modmult_1/xreg_reg[386]  ( .D(\modmult_1/xin[385] ), .CLK(clk), .RST(
        start_in[0]), .I(c[386]), .Q(\modmult_1/xin[386] ) );
  DFF \modmult_1/xreg_reg[385]  ( .D(\modmult_1/xin[384] ), .CLK(clk), .RST(
        start_in[0]), .I(c[385]), .Q(\modmult_1/xin[385] ) );
  DFF \modmult_1/xreg_reg[384]  ( .D(\modmult_1/xin[383] ), .CLK(clk), .RST(
        start_in[0]), .I(c[384]), .Q(\modmult_1/xin[384] ) );
  DFF \modmult_1/xreg_reg[383]  ( .D(\modmult_1/xin[382] ), .CLK(clk), .RST(
        start_in[0]), .I(c[383]), .Q(\modmult_1/xin[383] ) );
  DFF \modmult_1/xreg_reg[382]  ( .D(\modmult_1/xin[381] ), .CLK(clk), .RST(
        start_in[0]), .I(c[382]), .Q(\modmult_1/xin[382] ) );
  DFF \modmult_1/xreg_reg[381]  ( .D(\modmult_1/xin[380] ), .CLK(clk), .RST(
        start_in[0]), .I(c[381]), .Q(\modmult_1/xin[381] ) );
  DFF \modmult_1/xreg_reg[380]  ( .D(\modmult_1/xin[379] ), .CLK(clk), .RST(
        start_in[0]), .I(c[380]), .Q(\modmult_1/xin[380] ) );
  DFF \modmult_1/xreg_reg[379]  ( .D(\modmult_1/xin[378] ), .CLK(clk), .RST(
        start_in[0]), .I(c[379]), .Q(\modmult_1/xin[379] ) );
  DFF \modmult_1/xreg_reg[378]  ( .D(\modmult_1/xin[377] ), .CLK(clk), .RST(
        start_in[0]), .I(c[378]), .Q(\modmult_1/xin[378] ) );
  DFF \modmult_1/xreg_reg[377]  ( .D(\modmult_1/xin[376] ), .CLK(clk), .RST(
        start_in[0]), .I(c[377]), .Q(\modmult_1/xin[377] ) );
  DFF \modmult_1/xreg_reg[376]  ( .D(\modmult_1/xin[375] ), .CLK(clk), .RST(
        start_in[0]), .I(c[376]), .Q(\modmult_1/xin[376] ) );
  DFF \modmult_1/xreg_reg[375]  ( .D(\modmult_1/xin[374] ), .CLK(clk), .RST(
        start_in[0]), .I(c[375]), .Q(\modmult_1/xin[375] ) );
  DFF \modmult_1/xreg_reg[374]  ( .D(\modmult_1/xin[373] ), .CLK(clk), .RST(
        start_in[0]), .I(c[374]), .Q(\modmult_1/xin[374] ) );
  DFF \modmult_1/xreg_reg[373]  ( .D(\modmult_1/xin[372] ), .CLK(clk), .RST(
        start_in[0]), .I(c[373]), .Q(\modmult_1/xin[373] ) );
  DFF \modmult_1/xreg_reg[372]  ( .D(\modmult_1/xin[371] ), .CLK(clk), .RST(
        start_in[0]), .I(c[372]), .Q(\modmult_1/xin[372] ) );
  DFF \modmult_1/xreg_reg[371]  ( .D(\modmult_1/xin[370] ), .CLK(clk), .RST(
        start_in[0]), .I(c[371]), .Q(\modmult_1/xin[371] ) );
  DFF \modmult_1/xreg_reg[370]  ( .D(\modmult_1/xin[369] ), .CLK(clk), .RST(
        start_in[0]), .I(c[370]), .Q(\modmult_1/xin[370] ) );
  DFF \modmult_1/xreg_reg[369]  ( .D(\modmult_1/xin[368] ), .CLK(clk), .RST(
        start_in[0]), .I(c[369]), .Q(\modmult_1/xin[369] ) );
  DFF \modmult_1/xreg_reg[368]  ( .D(\modmult_1/xin[367] ), .CLK(clk), .RST(
        start_in[0]), .I(c[368]), .Q(\modmult_1/xin[368] ) );
  DFF \modmult_1/xreg_reg[367]  ( .D(\modmult_1/xin[366] ), .CLK(clk), .RST(
        start_in[0]), .I(c[367]), .Q(\modmult_1/xin[367] ) );
  DFF \modmult_1/xreg_reg[366]  ( .D(\modmult_1/xin[365] ), .CLK(clk), .RST(
        start_in[0]), .I(c[366]), .Q(\modmult_1/xin[366] ) );
  DFF \modmult_1/xreg_reg[365]  ( .D(\modmult_1/xin[364] ), .CLK(clk), .RST(
        start_in[0]), .I(c[365]), .Q(\modmult_1/xin[365] ) );
  DFF \modmult_1/xreg_reg[364]  ( .D(\modmult_1/xin[363] ), .CLK(clk), .RST(
        start_in[0]), .I(c[364]), .Q(\modmult_1/xin[364] ) );
  DFF \modmult_1/xreg_reg[363]  ( .D(\modmult_1/xin[362] ), .CLK(clk), .RST(
        start_in[0]), .I(c[363]), .Q(\modmult_1/xin[363] ) );
  DFF \modmult_1/xreg_reg[362]  ( .D(\modmult_1/xin[361] ), .CLK(clk), .RST(
        start_in[0]), .I(c[362]), .Q(\modmult_1/xin[362] ) );
  DFF \modmult_1/xreg_reg[361]  ( .D(\modmult_1/xin[360] ), .CLK(clk), .RST(
        start_in[0]), .I(c[361]), .Q(\modmult_1/xin[361] ) );
  DFF \modmult_1/xreg_reg[360]  ( .D(\modmult_1/xin[359] ), .CLK(clk), .RST(
        start_in[0]), .I(c[360]), .Q(\modmult_1/xin[360] ) );
  DFF \modmult_1/xreg_reg[359]  ( .D(\modmult_1/xin[358] ), .CLK(clk), .RST(
        start_in[0]), .I(c[359]), .Q(\modmult_1/xin[359] ) );
  DFF \modmult_1/xreg_reg[358]  ( .D(\modmult_1/xin[357] ), .CLK(clk), .RST(
        start_in[0]), .I(c[358]), .Q(\modmult_1/xin[358] ) );
  DFF \modmult_1/xreg_reg[357]  ( .D(\modmult_1/xin[356] ), .CLK(clk), .RST(
        start_in[0]), .I(c[357]), .Q(\modmult_1/xin[357] ) );
  DFF \modmult_1/xreg_reg[356]  ( .D(\modmult_1/xin[355] ), .CLK(clk), .RST(
        start_in[0]), .I(c[356]), .Q(\modmult_1/xin[356] ) );
  DFF \modmult_1/xreg_reg[355]  ( .D(\modmult_1/xin[354] ), .CLK(clk), .RST(
        start_in[0]), .I(c[355]), .Q(\modmult_1/xin[355] ) );
  DFF \modmult_1/xreg_reg[354]  ( .D(\modmult_1/xin[353] ), .CLK(clk), .RST(
        start_in[0]), .I(c[354]), .Q(\modmult_1/xin[354] ) );
  DFF \modmult_1/xreg_reg[353]  ( .D(\modmult_1/xin[352] ), .CLK(clk), .RST(
        start_in[0]), .I(c[353]), .Q(\modmult_1/xin[353] ) );
  DFF \modmult_1/xreg_reg[352]  ( .D(\modmult_1/xin[351] ), .CLK(clk), .RST(
        start_in[0]), .I(c[352]), .Q(\modmult_1/xin[352] ) );
  DFF \modmult_1/xreg_reg[351]  ( .D(\modmult_1/xin[350] ), .CLK(clk), .RST(
        start_in[0]), .I(c[351]), .Q(\modmult_1/xin[351] ) );
  DFF \modmult_1/xreg_reg[350]  ( .D(\modmult_1/xin[349] ), .CLK(clk), .RST(
        start_in[0]), .I(c[350]), .Q(\modmult_1/xin[350] ) );
  DFF \modmult_1/xreg_reg[349]  ( .D(\modmult_1/xin[348] ), .CLK(clk), .RST(
        start_in[0]), .I(c[349]), .Q(\modmult_1/xin[349] ) );
  DFF \modmult_1/xreg_reg[348]  ( .D(\modmult_1/xin[347] ), .CLK(clk), .RST(
        start_in[0]), .I(c[348]), .Q(\modmult_1/xin[348] ) );
  DFF \modmult_1/xreg_reg[347]  ( .D(\modmult_1/xin[346] ), .CLK(clk), .RST(
        start_in[0]), .I(c[347]), .Q(\modmult_1/xin[347] ) );
  DFF \modmult_1/xreg_reg[346]  ( .D(\modmult_1/xin[345] ), .CLK(clk), .RST(
        start_in[0]), .I(c[346]), .Q(\modmult_1/xin[346] ) );
  DFF \modmult_1/xreg_reg[345]  ( .D(\modmult_1/xin[344] ), .CLK(clk), .RST(
        start_in[0]), .I(c[345]), .Q(\modmult_1/xin[345] ) );
  DFF \modmult_1/xreg_reg[344]  ( .D(\modmult_1/xin[343] ), .CLK(clk), .RST(
        start_in[0]), .I(c[344]), .Q(\modmult_1/xin[344] ) );
  DFF \modmult_1/xreg_reg[343]  ( .D(\modmult_1/xin[342] ), .CLK(clk), .RST(
        start_in[0]), .I(c[343]), .Q(\modmult_1/xin[343] ) );
  DFF \modmult_1/xreg_reg[342]  ( .D(\modmult_1/xin[341] ), .CLK(clk), .RST(
        start_in[0]), .I(c[342]), .Q(\modmult_1/xin[342] ) );
  DFF \modmult_1/xreg_reg[341]  ( .D(\modmult_1/xin[340] ), .CLK(clk), .RST(
        start_in[0]), .I(c[341]), .Q(\modmult_1/xin[341] ) );
  DFF \modmult_1/xreg_reg[340]  ( .D(\modmult_1/xin[339] ), .CLK(clk), .RST(
        start_in[0]), .I(c[340]), .Q(\modmult_1/xin[340] ) );
  DFF \modmult_1/xreg_reg[339]  ( .D(\modmult_1/xin[338] ), .CLK(clk), .RST(
        start_in[0]), .I(c[339]), .Q(\modmult_1/xin[339] ) );
  DFF \modmult_1/xreg_reg[338]  ( .D(\modmult_1/xin[337] ), .CLK(clk), .RST(
        start_in[0]), .I(c[338]), .Q(\modmult_1/xin[338] ) );
  DFF \modmult_1/xreg_reg[337]  ( .D(\modmult_1/xin[336] ), .CLK(clk), .RST(
        start_in[0]), .I(c[337]), .Q(\modmult_1/xin[337] ) );
  DFF \modmult_1/xreg_reg[336]  ( .D(\modmult_1/xin[335] ), .CLK(clk), .RST(
        start_in[0]), .I(c[336]), .Q(\modmult_1/xin[336] ) );
  DFF \modmult_1/xreg_reg[335]  ( .D(\modmult_1/xin[334] ), .CLK(clk), .RST(
        start_in[0]), .I(c[335]), .Q(\modmult_1/xin[335] ) );
  DFF \modmult_1/xreg_reg[334]  ( .D(\modmult_1/xin[333] ), .CLK(clk), .RST(
        start_in[0]), .I(c[334]), .Q(\modmult_1/xin[334] ) );
  DFF \modmult_1/xreg_reg[333]  ( .D(\modmult_1/xin[332] ), .CLK(clk), .RST(
        start_in[0]), .I(c[333]), .Q(\modmult_1/xin[333] ) );
  DFF \modmult_1/xreg_reg[332]  ( .D(\modmult_1/xin[331] ), .CLK(clk), .RST(
        start_in[0]), .I(c[332]), .Q(\modmult_1/xin[332] ) );
  DFF \modmult_1/xreg_reg[331]  ( .D(\modmult_1/xin[330] ), .CLK(clk), .RST(
        start_in[0]), .I(c[331]), .Q(\modmult_1/xin[331] ) );
  DFF \modmult_1/xreg_reg[330]  ( .D(\modmult_1/xin[329] ), .CLK(clk), .RST(
        start_in[0]), .I(c[330]), .Q(\modmult_1/xin[330] ) );
  DFF \modmult_1/xreg_reg[329]  ( .D(\modmult_1/xin[328] ), .CLK(clk), .RST(
        start_in[0]), .I(c[329]), .Q(\modmult_1/xin[329] ) );
  DFF \modmult_1/xreg_reg[328]  ( .D(\modmult_1/xin[327] ), .CLK(clk), .RST(
        start_in[0]), .I(c[328]), .Q(\modmult_1/xin[328] ) );
  DFF \modmult_1/xreg_reg[327]  ( .D(\modmult_1/xin[326] ), .CLK(clk), .RST(
        start_in[0]), .I(c[327]), .Q(\modmult_1/xin[327] ) );
  DFF \modmult_1/xreg_reg[326]  ( .D(\modmult_1/xin[325] ), .CLK(clk), .RST(
        start_in[0]), .I(c[326]), .Q(\modmult_1/xin[326] ) );
  DFF \modmult_1/xreg_reg[325]  ( .D(\modmult_1/xin[324] ), .CLK(clk), .RST(
        start_in[0]), .I(c[325]), .Q(\modmult_1/xin[325] ) );
  DFF \modmult_1/xreg_reg[324]  ( .D(\modmult_1/xin[323] ), .CLK(clk), .RST(
        start_in[0]), .I(c[324]), .Q(\modmult_1/xin[324] ) );
  DFF \modmult_1/xreg_reg[323]  ( .D(\modmult_1/xin[322] ), .CLK(clk), .RST(
        start_in[0]), .I(c[323]), .Q(\modmult_1/xin[323] ) );
  DFF \modmult_1/xreg_reg[322]  ( .D(\modmult_1/xin[321] ), .CLK(clk), .RST(
        start_in[0]), .I(c[322]), .Q(\modmult_1/xin[322] ) );
  DFF \modmult_1/xreg_reg[321]  ( .D(\modmult_1/xin[320] ), .CLK(clk), .RST(
        start_in[0]), .I(c[321]), .Q(\modmult_1/xin[321] ) );
  DFF \modmult_1/xreg_reg[320]  ( .D(\modmult_1/xin[319] ), .CLK(clk), .RST(
        start_in[0]), .I(c[320]), .Q(\modmult_1/xin[320] ) );
  DFF \modmult_1/xreg_reg[319]  ( .D(\modmult_1/xin[318] ), .CLK(clk), .RST(
        start_in[0]), .I(c[319]), .Q(\modmult_1/xin[319] ) );
  DFF \modmult_1/xreg_reg[318]  ( .D(\modmult_1/xin[317] ), .CLK(clk), .RST(
        start_in[0]), .I(c[318]), .Q(\modmult_1/xin[318] ) );
  DFF \modmult_1/xreg_reg[317]  ( .D(\modmult_1/xin[316] ), .CLK(clk), .RST(
        start_in[0]), .I(c[317]), .Q(\modmult_1/xin[317] ) );
  DFF \modmult_1/xreg_reg[316]  ( .D(\modmult_1/xin[315] ), .CLK(clk), .RST(
        start_in[0]), .I(c[316]), .Q(\modmult_1/xin[316] ) );
  DFF \modmult_1/xreg_reg[315]  ( .D(\modmult_1/xin[314] ), .CLK(clk), .RST(
        start_in[0]), .I(c[315]), .Q(\modmult_1/xin[315] ) );
  DFF \modmult_1/xreg_reg[314]  ( .D(\modmult_1/xin[313] ), .CLK(clk), .RST(
        start_in[0]), .I(c[314]), .Q(\modmult_1/xin[314] ) );
  DFF \modmult_1/xreg_reg[313]  ( .D(\modmult_1/xin[312] ), .CLK(clk), .RST(
        start_in[0]), .I(c[313]), .Q(\modmult_1/xin[313] ) );
  DFF \modmult_1/xreg_reg[312]  ( .D(\modmult_1/xin[311] ), .CLK(clk), .RST(
        start_in[0]), .I(c[312]), .Q(\modmult_1/xin[312] ) );
  DFF \modmult_1/xreg_reg[311]  ( .D(\modmult_1/xin[310] ), .CLK(clk), .RST(
        start_in[0]), .I(c[311]), .Q(\modmult_1/xin[311] ) );
  DFF \modmult_1/xreg_reg[310]  ( .D(\modmult_1/xin[309] ), .CLK(clk), .RST(
        start_in[0]), .I(c[310]), .Q(\modmult_1/xin[310] ) );
  DFF \modmult_1/xreg_reg[309]  ( .D(\modmult_1/xin[308] ), .CLK(clk), .RST(
        start_in[0]), .I(c[309]), .Q(\modmult_1/xin[309] ) );
  DFF \modmult_1/xreg_reg[308]  ( .D(\modmult_1/xin[307] ), .CLK(clk), .RST(
        start_in[0]), .I(c[308]), .Q(\modmult_1/xin[308] ) );
  DFF \modmult_1/xreg_reg[307]  ( .D(\modmult_1/xin[306] ), .CLK(clk), .RST(
        start_in[0]), .I(c[307]), .Q(\modmult_1/xin[307] ) );
  DFF \modmult_1/xreg_reg[306]  ( .D(\modmult_1/xin[305] ), .CLK(clk), .RST(
        start_in[0]), .I(c[306]), .Q(\modmult_1/xin[306] ) );
  DFF \modmult_1/xreg_reg[305]  ( .D(\modmult_1/xin[304] ), .CLK(clk), .RST(
        start_in[0]), .I(c[305]), .Q(\modmult_1/xin[305] ) );
  DFF \modmult_1/xreg_reg[304]  ( .D(\modmult_1/xin[303] ), .CLK(clk), .RST(
        start_in[0]), .I(c[304]), .Q(\modmult_1/xin[304] ) );
  DFF \modmult_1/xreg_reg[303]  ( .D(\modmult_1/xin[302] ), .CLK(clk), .RST(
        start_in[0]), .I(c[303]), .Q(\modmult_1/xin[303] ) );
  DFF \modmult_1/xreg_reg[302]  ( .D(\modmult_1/xin[301] ), .CLK(clk), .RST(
        start_in[0]), .I(c[302]), .Q(\modmult_1/xin[302] ) );
  DFF \modmult_1/xreg_reg[301]  ( .D(\modmult_1/xin[300] ), .CLK(clk), .RST(
        start_in[0]), .I(c[301]), .Q(\modmult_1/xin[301] ) );
  DFF \modmult_1/xreg_reg[300]  ( .D(\modmult_1/xin[299] ), .CLK(clk), .RST(
        start_in[0]), .I(c[300]), .Q(\modmult_1/xin[300] ) );
  DFF \modmult_1/xreg_reg[299]  ( .D(\modmult_1/xin[298] ), .CLK(clk), .RST(
        start_in[0]), .I(c[299]), .Q(\modmult_1/xin[299] ) );
  DFF \modmult_1/xreg_reg[298]  ( .D(\modmult_1/xin[297] ), .CLK(clk), .RST(
        start_in[0]), .I(c[298]), .Q(\modmult_1/xin[298] ) );
  DFF \modmult_1/xreg_reg[297]  ( .D(\modmult_1/xin[296] ), .CLK(clk), .RST(
        start_in[0]), .I(c[297]), .Q(\modmult_1/xin[297] ) );
  DFF \modmult_1/xreg_reg[296]  ( .D(\modmult_1/xin[295] ), .CLK(clk), .RST(
        start_in[0]), .I(c[296]), .Q(\modmult_1/xin[296] ) );
  DFF \modmult_1/xreg_reg[295]  ( .D(\modmult_1/xin[294] ), .CLK(clk), .RST(
        start_in[0]), .I(c[295]), .Q(\modmult_1/xin[295] ) );
  DFF \modmult_1/xreg_reg[294]  ( .D(\modmult_1/xin[293] ), .CLK(clk), .RST(
        start_in[0]), .I(c[294]), .Q(\modmult_1/xin[294] ) );
  DFF \modmult_1/xreg_reg[293]  ( .D(\modmult_1/xin[292] ), .CLK(clk), .RST(
        start_in[0]), .I(c[293]), .Q(\modmult_1/xin[293] ) );
  DFF \modmult_1/xreg_reg[292]  ( .D(\modmult_1/xin[291] ), .CLK(clk), .RST(
        start_in[0]), .I(c[292]), .Q(\modmult_1/xin[292] ) );
  DFF \modmult_1/xreg_reg[291]  ( .D(\modmult_1/xin[290] ), .CLK(clk), .RST(
        start_in[0]), .I(c[291]), .Q(\modmult_1/xin[291] ) );
  DFF \modmult_1/xreg_reg[290]  ( .D(\modmult_1/xin[289] ), .CLK(clk), .RST(
        start_in[0]), .I(c[290]), .Q(\modmult_1/xin[290] ) );
  DFF \modmult_1/xreg_reg[289]  ( .D(\modmult_1/xin[288] ), .CLK(clk), .RST(
        start_in[0]), .I(c[289]), .Q(\modmult_1/xin[289] ) );
  DFF \modmult_1/xreg_reg[288]  ( .D(\modmult_1/xin[287] ), .CLK(clk), .RST(
        start_in[0]), .I(c[288]), .Q(\modmult_1/xin[288] ) );
  DFF \modmult_1/xreg_reg[287]  ( .D(\modmult_1/xin[286] ), .CLK(clk), .RST(
        start_in[0]), .I(c[287]), .Q(\modmult_1/xin[287] ) );
  DFF \modmult_1/xreg_reg[286]  ( .D(\modmult_1/xin[285] ), .CLK(clk), .RST(
        start_in[0]), .I(c[286]), .Q(\modmult_1/xin[286] ) );
  DFF \modmult_1/xreg_reg[285]  ( .D(\modmult_1/xin[284] ), .CLK(clk), .RST(
        start_in[0]), .I(c[285]), .Q(\modmult_1/xin[285] ) );
  DFF \modmult_1/xreg_reg[284]  ( .D(\modmult_1/xin[283] ), .CLK(clk), .RST(
        start_in[0]), .I(c[284]), .Q(\modmult_1/xin[284] ) );
  DFF \modmult_1/xreg_reg[283]  ( .D(\modmult_1/xin[282] ), .CLK(clk), .RST(
        start_in[0]), .I(c[283]), .Q(\modmult_1/xin[283] ) );
  DFF \modmult_1/xreg_reg[282]  ( .D(\modmult_1/xin[281] ), .CLK(clk), .RST(
        start_in[0]), .I(c[282]), .Q(\modmult_1/xin[282] ) );
  DFF \modmult_1/xreg_reg[281]  ( .D(\modmult_1/xin[280] ), .CLK(clk), .RST(
        start_in[0]), .I(c[281]), .Q(\modmult_1/xin[281] ) );
  DFF \modmult_1/xreg_reg[280]  ( .D(\modmult_1/xin[279] ), .CLK(clk), .RST(
        start_in[0]), .I(c[280]), .Q(\modmult_1/xin[280] ) );
  DFF \modmult_1/xreg_reg[279]  ( .D(\modmult_1/xin[278] ), .CLK(clk), .RST(
        start_in[0]), .I(c[279]), .Q(\modmult_1/xin[279] ) );
  DFF \modmult_1/xreg_reg[278]  ( .D(\modmult_1/xin[277] ), .CLK(clk), .RST(
        start_in[0]), .I(c[278]), .Q(\modmult_1/xin[278] ) );
  DFF \modmult_1/xreg_reg[277]  ( .D(\modmult_1/xin[276] ), .CLK(clk), .RST(
        start_in[0]), .I(c[277]), .Q(\modmult_1/xin[277] ) );
  DFF \modmult_1/xreg_reg[276]  ( .D(\modmult_1/xin[275] ), .CLK(clk), .RST(
        start_in[0]), .I(c[276]), .Q(\modmult_1/xin[276] ) );
  DFF \modmult_1/xreg_reg[275]  ( .D(\modmult_1/xin[274] ), .CLK(clk), .RST(
        start_in[0]), .I(c[275]), .Q(\modmult_1/xin[275] ) );
  DFF \modmult_1/xreg_reg[274]  ( .D(\modmult_1/xin[273] ), .CLK(clk), .RST(
        start_in[0]), .I(c[274]), .Q(\modmult_1/xin[274] ) );
  DFF \modmult_1/xreg_reg[273]  ( .D(\modmult_1/xin[272] ), .CLK(clk), .RST(
        start_in[0]), .I(c[273]), .Q(\modmult_1/xin[273] ) );
  DFF \modmult_1/xreg_reg[272]  ( .D(\modmult_1/xin[271] ), .CLK(clk), .RST(
        start_in[0]), .I(c[272]), .Q(\modmult_1/xin[272] ) );
  DFF \modmult_1/xreg_reg[271]  ( .D(\modmult_1/xin[270] ), .CLK(clk), .RST(
        start_in[0]), .I(c[271]), .Q(\modmult_1/xin[271] ) );
  DFF \modmult_1/xreg_reg[270]  ( .D(\modmult_1/xin[269] ), .CLK(clk), .RST(
        start_in[0]), .I(c[270]), .Q(\modmult_1/xin[270] ) );
  DFF \modmult_1/xreg_reg[269]  ( .D(\modmult_1/xin[268] ), .CLK(clk), .RST(
        start_in[0]), .I(c[269]), .Q(\modmult_1/xin[269] ) );
  DFF \modmult_1/xreg_reg[268]  ( .D(\modmult_1/xin[267] ), .CLK(clk), .RST(
        start_in[0]), .I(c[268]), .Q(\modmult_1/xin[268] ) );
  DFF \modmult_1/xreg_reg[267]  ( .D(\modmult_1/xin[266] ), .CLK(clk), .RST(
        start_in[0]), .I(c[267]), .Q(\modmult_1/xin[267] ) );
  DFF \modmult_1/xreg_reg[266]  ( .D(\modmult_1/xin[265] ), .CLK(clk), .RST(
        start_in[0]), .I(c[266]), .Q(\modmult_1/xin[266] ) );
  DFF \modmult_1/xreg_reg[265]  ( .D(\modmult_1/xin[264] ), .CLK(clk), .RST(
        start_in[0]), .I(c[265]), .Q(\modmult_1/xin[265] ) );
  DFF \modmult_1/xreg_reg[264]  ( .D(\modmult_1/xin[263] ), .CLK(clk), .RST(
        start_in[0]), .I(c[264]), .Q(\modmult_1/xin[264] ) );
  DFF \modmult_1/xreg_reg[263]  ( .D(\modmult_1/xin[262] ), .CLK(clk), .RST(
        start_in[0]), .I(c[263]), .Q(\modmult_1/xin[263] ) );
  DFF \modmult_1/xreg_reg[262]  ( .D(\modmult_1/xin[261] ), .CLK(clk), .RST(
        start_in[0]), .I(c[262]), .Q(\modmult_1/xin[262] ) );
  DFF \modmult_1/xreg_reg[261]  ( .D(\modmult_1/xin[260] ), .CLK(clk), .RST(
        start_in[0]), .I(c[261]), .Q(\modmult_1/xin[261] ) );
  DFF \modmult_1/xreg_reg[260]  ( .D(\modmult_1/xin[259] ), .CLK(clk), .RST(
        start_in[0]), .I(c[260]), .Q(\modmult_1/xin[260] ) );
  DFF \modmult_1/xreg_reg[259]  ( .D(\modmult_1/xin[258] ), .CLK(clk), .RST(
        start_in[0]), .I(c[259]), .Q(\modmult_1/xin[259] ) );
  DFF \modmult_1/xreg_reg[258]  ( .D(\modmult_1/xin[257] ), .CLK(clk), .RST(
        start_in[0]), .I(c[258]), .Q(\modmult_1/xin[258] ) );
  DFF \modmult_1/xreg_reg[257]  ( .D(\modmult_1/xin[256] ), .CLK(clk), .RST(
        start_in[0]), .I(c[257]), .Q(\modmult_1/xin[257] ) );
  DFF \modmult_1/xreg_reg[256]  ( .D(\modmult_1/xin[255] ), .CLK(clk), .RST(
        start_in[0]), .I(c[256]), .Q(\modmult_1/xin[256] ) );
  DFF \modmult_1/xreg_reg[255]  ( .D(\modmult_1/xin[254] ), .CLK(clk), .RST(
        start_in[0]), .I(c[255]), .Q(\modmult_1/xin[255] ) );
  DFF \modmult_1/xreg_reg[254]  ( .D(\modmult_1/xin[253] ), .CLK(clk), .RST(
        start_in[0]), .I(c[254]), .Q(\modmult_1/xin[254] ) );
  DFF \modmult_1/xreg_reg[253]  ( .D(\modmult_1/xin[252] ), .CLK(clk), .RST(
        start_in[0]), .I(c[253]), .Q(\modmult_1/xin[253] ) );
  DFF \modmult_1/xreg_reg[252]  ( .D(\modmult_1/xin[251] ), .CLK(clk), .RST(
        start_in[0]), .I(c[252]), .Q(\modmult_1/xin[252] ) );
  DFF \modmult_1/xreg_reg[251]  ( .D(\modmult_1/xin[250] ), .CLK(clk), .RST(
        start_in[0]), .I(c[251]), .Q(\modmult_1/xin[251] ) );
  DFF \modmult_1/xreg_reg[250]  ( .D(\modmult_1/xin[249] ), .CLK(clk), .RST(
        start_in[0]), .I(c[250]), .Q(\modmult_1/xin[250] ) );
  DFF \modmult_1/xreg_reg[249]  ( .D(\modmult_1/xin[248] ), .CLK(clk), .RST(
        start_in[0]), .I(c[249]), .Q(\modmult_1/xin[249] ) );
  DFF \modmult_1/xreg_reg[248]  ( .D(\modmult_1/xin[247] ), .CLK(clk), .RST(
        start_in[0]), .I(c[248]), .Q(\modmult_1/xin[248] ) );
  DFF \modmult_1/xreg_reg[247]  ( .D(\modmult_1/xin[246] ), .CLK(clk), .RST(
        start_in[0]), .I(c[247]), .Q(\modmult_1/xin[247] ) );
  DFF \modmult_1/xreg_reg[246]  ( .D(\modmult_1/xin[245] ), .CLK(clk), .RST(
        start_in[0]), .I(c[246]), .Q(\modmult_1/xin[246] ) );
  DFF \modmult_1/xreg_reg[245]  ( .D(\modmult_1/xin[244] ), .CLK(clk), .RST(
        start_in[0]), .I(c[245]), .Q(\modmult_1/xin[245] ) );
  DFF \modmult_1/xreg_reg[244]  ( .D(\modmult_1/xin[243] ), .CLK(clk), .RST(
        start_in[0]), .I(c[244]), .Q(\modmult_1/xin[244] ) );
  DFF \modmult_1/xreg_reg[243]  ( .D(\modmult_1/xin[242] ), .CLK(clk), .RST(
        start_in[0]), .I(c[243]), .Q(\modmult_1/xin[243] ) );
  DFF \modmult_1/xreg_reg[242]  ( .D(\modmult_1/xin[241] ), .CLK(clk), .RST(
        start_in[0]), .I(c[242]), .Q(\modmult_1/xin[242] ) );
  DFF \modmult_1/xreg_reg[241]  ( .D(\modmult_1/xin[240] ), .CLK(clk), .RST(
        start_in[0]), .I(c[241]), .Q(\modmult_1/xin[241] ) );
  DFF \modmult_1/xreg_reg[240]  ( .D(\modmult_1/xin[239] ), .CLK(clk), .RST(
        start_in[0]), .I(c[240]), .Q(\modmult_1/xin[240] ) );
  DFF \modmult_1/xreg_reg[239]  ( .D(\modmult_1/xin[238] ), .CLK(clk), .RST(
        start_in[0]), .I(c[239]), .Q(\modmult_1/xin[239] ) );
  DFF \modmult_1/xreg_reg[238]  ( .D(\modmult_1/xin[237] ), .CLK(clk), .RST(
        start_in[0]), .I(c[238]), .Q(\modmult_1/xin[238] ) );
  DFF \modmult_1/xreg_reg[237]  ( .D(\modmult_1/xin[236] ), .CLK(clk), .RST(
        start_in[0]), .I(c[237]), .Q(\modmult_1/xin[237] ) );
  DFF \modmult_1/xreg_reg[236]  ( .D(\modmult_1/xin[235] ), .CLK(clk), .RST(
        start_in[0]), .I(c[236]), .Q(\modmult_1/xin[236] ) );
  DFF \modmult_1/xreg_reg[235]  ( .D(\modmult_1/xin[234] ), .CLK(clk), .RST(
        start_in[0]), .I(c[235]), .Q(\modmult_1/xin[235] ) );
  DFF \modmult_1/xreg_reg[234]  ( .D(\modmult_1/xin[233] ), .CLK(clk), .RST(
        start_in[0]), .I(c[234]), .Q(\modmult_1/xin[234] ) );
  DFF \modmult_1/xreg_reg[233]  ( .D(\modmult_1/xin[232] ), .CLK(clk), .RST(
        start_in[0]), .I(c[233]), .Q(\modmult_1/xin[233] ) );
  DFF \modmult_1/xreg_reg[232]  ( .D(\modmult_1/xin[231] ), .CLK(clk), .RST(
        start_in[0]), .I(c[232]), .Q(\modmult_1/xin[232] ) );
  DFF \modmult_1/xreg_reg[231]  ( .D(\modmult_1/xin[230] ), .CLK(clk), .RST(
        start_in[0]), .I(c[231]), .Q(\modmult_1/xin[231] ) );
  DFF \modmult_1/xreg_reg[230]  ( .D(\modmult_1/xin[229] ), .CLK(clk), .RST(
        start_in[0]), .I(c[230]), .Q(\modmult_1/xin[230] ) );
  DFF \modmult_1/xreg_reg[229]  ( .D(\modmult_1/xin[228] ), .CLK(clk), .RST(
        start_in[0]), .I(c[229]), .Q(\modmult_1/xin[229] ) );
  DFF \modmult_1/xreg_reg[228]  ( .D(\modmult_1/xin[227] ), .CLK(clk), .RST(
        start_in[0]), .I(c[228]), .Q(\modmult_1/xin[228] ) );
  DFF \modmult_1/xreg_reg[227]  ( .D(\modmult_1/xin[226] ), .CLK(clk), .RST(
        start_in[0]), .I(c[227]), .Q(\modmult_1/xin[227] ) );
  DFF \modmult_1/xreg_reg[226]  ( .D(\modmult_1/xin[225] ), .CLK(clk), .RST(
        start_in[0]), .I(c[226]), .Q(\modmult_1/xin[226] ) );
  DFF \modmult_1/xreg_reg[225]  ( .D(\modmult_1/xin[224] ), .CLK(clk), .RST(
        start_in[0]), .I(c[225]), .Q(\modmult_1/xin[225] ) );
  DFF \modmult_1/xreg_reg[224]  ( .D(\modmult_1/xin[223] ), .CLK(clk), .RST(
        start_in[0]), .I(c[224]), .Q(\modmult_1/xin[224] ) );
  DFF \modmult_1/xreg_reg[223]  ( .D(\modmult_1/xin[222] ), .CLK(clk), .RST(
        start_in[0]), .I(c[223]), .Q(\modmult_1/xin[223] ) );
  DFF \modmult_1/xreg_reg[222]  ( .D(\modmult_1/xin[221] ), .CLK(clk), .RST(
        start_in[0]), .I(c[222]), .Q(\modmult_1/xin[222] ) );
  DFF \modmult_1/xreg_reg[221]  ( .D(\modmult_1/xin[220] ), .CLK(clk), .RST(
        start_in[0]), .I(c[221]), .Q(\modmult_1/xin[221] ) );
  DFF \modmult_1/xreg_reg[220]  ( .D(\modmult_1/xin[219] ), .CLK(clk), .RST(
        start_in[0]), .I(c[220]), .Q(\modmult_1/xin[220] ) );
  DFF \modmult_1/xreg_reg[219]  ( .D(\modmult_1/xin[218] ), .CLK(clk), .RST(
        start_in[0]), .I(c[219]), .Q(\modmult_1/xin[219] ) );
  DFF \modmult_1/xreg_reg[218]  ( .D(\modmult_1/xin[217] ), .CLK(clk), .RST(
        start_in[0]), .I(c[218]), .Q(\modmult_1/xin[218] ) );
  DFF \modmult_1/xreg_reg[217]  ( .D(\modmult_1/xin[216] ), .CLK(clk), .RST(
        start_in[0]), .I(c[217]), .Q(\modmult_1/xin[217] ) );
  DFF \modmult_1/xreg_reg[216]  ( .D(\modmult_1/xin[215] ), .CLK(clk), .RST(
        start_in[0]), .I(c[216]), .Q(\modmult_1/xin[216] ) );
  DFF \modmult_1/xreg_reg[215]  ( .D(\modmult_1/xin[214] ), .CLK(clk), .RST(
        start_in[0]), .I(c[215]), .Q(\modmult_1/xin[215] ) );
  DFF \modmult_1/xreg_reg[214]  ( .D(\modmult_1/xin[213] ), .CLK(clk), .RST(
        start_in[0]), .I(c[214]), .Q(\modmult_1/xin[214] ) );
  DFF \modmult_1/xreg_reg[213]  ( .D(\modmult_1/xin[212] ), .CLK(clk), .RST(
        start_in[0]), .I(c[213]), .Q(\modmult_1/xin[213] ) );
  DFF \modmult_1/xreg_reg[212]  ( .D(\modmult_1/xin[211] ), .CLK(clk), .RST(
        start_in[0]), .I(c[212]), .Q(\modmult_1/xin[212] ) );
  DFF \modmult_1/xreg_reg[211]  ( .D(\modmult_1/xin[210] ), .CLK(clk), .RST(
        start_in[0]), .I(c[211]), .Q(\modmult_1/xin[211] ) );
  DFF \modmult_1/xreg_reg[210]  ( .D(\modmult_1/xin[209] ), .CLK(clk), .RST(
        start_in[0]), .I(c[210]), .Q(\modmult_1/xin[210] ) );
  DFF \modmult_1/xreg_reg[209]  ( .D(\modmult_1/xin[208] ), .CLK(clk), .RST(
        start_in[0]), .I(c[209]), .Q(\modmult_1/xin[209] ) );
  DFF \modmult_1/xreg_reg[208]  ( .D(\modmult_1/xin[207] ), .CLK(clk), .RST(
        start_in[0]), .I(c[208]), .Q(\modmult_1/xin[208] ) );
  DFF \modmult_1/xreg_reg[207]  ( .D(\modmult_1/xin[206] ), .CLK(clk), .RST(
        start_in[0]), .I(c[207]), .Q(\modmult_1/xin[207] ) );
  DFF \modmult_1/xreg_reg[206]  ( .D(\modmult_1/xin[205] ), .CLK(clk), .RST(
        start_in[0]), .I(c[206]), .Q(\modmult_1/xin[206] ) );
  DFF \modmult_1/xreg_reg[205]  ( .D(\modmult_1/xin[204] ), .CLK(clk), .RST(
        start_in[0]), .I(c[205]), .Q(\modmult_1/xin[205] ) );
  DFF \modmult_1/xreg_reg[204]  ( .D(\modmult_1/xin[203] ), .CLK(clk), .RST(
        start_in[0]), .I(c[204]), .Q(\modmult_1/xin[204] ) );
  DFF \modmult_1/xreg_reg[203]  ( .D(\modmult_1/xin[202] ), .CLK(clk), .RST(
        start_in[0]), .I(c[203]), .Q(\modmult_1/xin[203] ) );
  DFF \modmult_1/xreg_reg[202]  ( .D(\modmult_1/xin[201] ), .CLK(clk), .RST(
        start_in[0]), .I(c[202]), .Q(\modmult_1/xin[202] ) );
  DFF \modmult_1/xreg_reg[201]  ( .D(\modmult_1/xin[200] ), .CLK(clk), .RST(
        start_in[0]), .I(c[201]), .Q(\modmult_1/xin[201] ) );
  DFF \modmult_1/xreg_reg[200]  ( .D(\modmult_1/xin[199] ), .CLK(clk), .RST(
        start_in[0]), .I(c[200]), .Q(\modmult_1/xin[200] ) );
  DFF \modmult_1/xreg_reg[199]  ( .D(\modmult_1/xin[198] ), .CLK(clk), .RST(
        start_in[0]), .I(c[199]), .Q(\modmult_1/xin[199] ) );
  DFF \modmult_1/xreg_reg[198]  ( .D(\modmult_1/xin[197] ), .CLK(clk), .RST(
        start_in[0]), .I(c[198]), .Q(\modmult_1/xin[198] ) );
  DFF \modmult_1/xreg_reg[197]  ( .D(\modmult_1/xin[196] ), .CLK(clk), .RST(
        start_in[0]), .I(c[197]), .Q(\modmult_1/xin[197] ) );
  DFF \modmult_1/xreg_reg[196]  ( .D(\modmult_1/xin[195] ), .CLK(clk), .RST(
        start_in[0]), .I(c[196]), .Q(\modmult_1/xin[196] ) );
  DFF \modmult_1/xreg_reg[195]  ( .D(\modmult_1/xin[194] ), .CLK(clk), .RST(
        start_in[0]), .I(c[195]), .Q(\modmult_1/xin[195] ) );
  DFF \modmult_1/xreg_reg[194]  ( .D(\modmult_1/xin[193] ), .CLK(clk), .RST(
        start_in[0]), .I(c[194]), .Q(\modmult_1/xin[194] ) );
  DFF \modmult_1/xreg_reg[193]  ( .D(\modmult_1/xin[192] ), .CLK(clk), .RST(
        start_in[0]), .I(c[193]), .Q(\modmult_1/xin[193] ) );
  DFF \modmult_1/xreg_reg[192]  ( .D(\modmult_1/xin[191] ), .CLK(clk), .RST(
        start_in[0]), .I(c[192]), .Q(\modmult_1/xin[192] ) );
  DFF \modmult_1/xreg_reg[191]  ( .D(\modmult_1/xin[190] ), .CLK(clk), .RST(
        start_in[0]), .I(c[191]), .Q(\modmult_1/xin[191] ) );
  DFF \modmult_1/xreg_reg[190]  ( .D(\modmult_1/xin[189] ), .CLK(clk), .RST(
        start_in[0]), .I(c[190]), .Q(\modmult_1/xin[190] ) );
  DFF \modmult_1/xreg_reg[189]  ( .D(\modmult_1/xin[188] ), .CLK(clk), .RST(
        start_in[0]), .I(c[189]), .Q(\modmult_1/xin[189] ) );
  DFF \modmult_1/xreg_reg[188]  ( .D(\modmult_1/xin[187] ), .CLK(clk), .RST(
        start_in[0]), .I(c[188]), .Q(\modmult_1/xin[188] ) );
  DFF \modmult_1/xreg_reg[187]  ( .D(\modmult_1/xin[186] ), .CLK(clk), .RST(
        start_in[0]), .I(c[187]), .Q(\modmult_1/xin[187] ) );
  DFF \modmult_1/xreg_reg[186]  ( .D(\modmult_1/xin[185] ), .CLK(clk), .RST(
        start_in[0]), .I(c[186]), .Q(\modmult_1/xin[186] ) );
  DFF \modmult_1/xreg_reg[185]  ( .D(\modmult_1/xin[184] ), .CLK(clk), .RST(
        start_in[0]), .I(c[185]), .Q(\modmult_1/xin[185] ) );
  DFF \modmult_1/xreg_reg[184]  ( .D(\modmult_1/xin[183] ), .CLK(clk), .RST(
        start_in[0]), .I(c[184]), .Q(\modmult_1/xin[184] ) );
  DFF \modmult_1/xreg_reg[183]  ( .D(\modmult_1/xin[182] ), .CLK(clk), .RST(
        start_in[0]), .I(c[183]), .Q(\modmult_1/xin[183] ) );
  DFF \modmult_1/xreg_reg[182]  ( .D(\modmult_1/xin[181] ), .CLK(clk), .RST(
        start_in[0]), .I(c[182]), .Q(\modmult_1/xin[182] ) );
  DFF \modmult_1/xreg_reg[181]  ( .D(\modmult_1/xin[180] ), .CLK(clk), .RST(
        start_in[0]), .I(c[181]), .Q(\modmult_1/xin[181] ) );
  DFF \modmult_1/xreg_reg[180]  ( .D(\modmult_1/xin[179] ), .CLK(clk), .RST(
        start_in[0]), .I(c[180]), .Q(\modmult_1/xin[180] ) );
  DFF \modmult_1/xreg_reg[179]  ( .D(\modmult_1/xin[178] ), .CLK(clk), .RST(
        start_in[0]), .I(c[179]), .Q(\modmult_1/xin[179] ) );
  DFF \modmult_1/xreg_reg[178]  ( .D(\modmult_1/xin[177] ), .CLK(clk), .RST(
        start_in[0]), .I(c[178]), .Q(\modmult_1/xin[178] ) );
  DFF \modmult_1/xreg_reg[177]  ( .D(\modmult_1/xin[176] ), .CLK(clk), .RST(
        start_in[0]), .I(c[177]), .Q(\modmult_1/xin[177] ) );
  DFF \modmult_1/xreg_reg[176]  ( .D(\modmult_1/xin[175] ), .CLK(clk), .RST(
        start_in[0]), .I(c[176]), .Q(\modmult_1/xin[176] ) );
  DFF \modmult_1/xreg_reg[175]  ( .D(\modmult_1/xin[174] ), .CLK(clk), .RST(
        start_in[0]), .I(c[175]), .Q(\modmult_1/xin[175] ) );
  DFF \modmult_1/xreg_reg[174]  ( .D(\modmult_1/xin[173] ), .CLK(clk), .RST(
        start_in[0]), .I(c[174]), .Q(\modmult_1/xin[174] ) );
  DFF \modmult_1/xreg_reg[173]  ( .D(\modmult_1/xin[172] ), .CLK(clk), .RST(
        start_in[0]), .I(c[173]), .Q(\modmult_1/xin[173] ) );
  DFF \modmult_1/xreg_reg[172]  ( .D(\modmult_1/xin[171] ), .CLK(clk), .RST(
        start_in[0]), .I(c[172]), .Q(\modmult_1/xin[172] ) );
  DFF \modmult_1/xreg_reg[171]  ( .D(\modmult_1/xin[170] ), .CLK(clk), .RST(
        start_in[0]), .I(c[171]), .Q(\modmult_1/xin[171] ) );
  DFF \modmult_1/xreg_reg[170]  ( .D(\modmult_1/xin[169] ), .CLK(clk), .RST(
        start_in[0]), .I(c[170]), .Q(\modmult_1/xin[170] ) );
  DFF \modmult_1/xreg_reg[169]  ( .D(\modmult_1/xin[168] ), .CLK(clk), .RST(
        start_in[0]), .I(c[169]), .Q(\modmult_1/xin[169] ) );
  DFF \modmult_1/xreg_reg[168]  ( .D(\modmult_1/xin[167] ), .CLK(clk), .RST(
        start_in[0]), .I(c[168]), .Q(\modmult_1/xin[168] ) );
  DFF \modmult_1/xreg_reg[167]  ( .D(\modmult_1/xin[166] ), .CLK(clk), .RST(
        start_in[0]), .I(c[167]), .Q(\modmult_1/xin[167] ) );
  DFF \modmult_1/xreg_reg[166]  ( .D(\modmult_1/xin[165] ), .CLK(clk), .RST(
        start_in[0]), .I(c[166]), .Q(\modmult_1/xin[166] ) );
  DFF \modmult_1/xreg_reg[165]  ( .D(\modmult_1/xin[164] ), .CLK(clk), .RST(
        start_in[0]), .I(c[165]), .Q(\modmult_1/xin[165] ) );
  DFF \modmult_1/xreg_reg[164]  ( .D(\modmult_1/xin[163] ), .CLK(clk), .RST(
        start_in[0]), .I(c[164]), .Q(\modmult_1/xin[164] ) );
  DFF \modmult_1/xreg_reg[163]  ( .D(\modmult_1/xin[162] ), .CLK(clk), .RST(
        start_in[0]), .I(c[163]), .Q(\modmult_1/xin[163] ) );
  DFF \modmult_1/xreg_reg[162]  ( .D(\modmult_1/xin[161] ), .CLK(clk), .RST(
        start_in[0]), .I(c[162]), .Q(\modmult_1/xin[162] ) );
  DFF \modmult_1/xreg_reg[161]  ( .D(\modmult_1/xin[160] ), .CLK(clk), .RST(
        start_in[0]), .I(c[161]), .Q(\modmult_1/xin[161] ) );
  DFF \modmult_1/xreg_reg[160]  ( .D(\modmult_1/xin[159] ), .CLK(clk), .RST(
        start_in[0]), .I(c[160]), .Q(\modmult_1/xin[160] ) );
  DFF \modmult_1/xreg_reg[159]  ( .D(\modmult_1/xin[158] ), .CLK(clk), .RST(
        start_in[0]), .I(c[159]), .Q(\modmult_1/xin[159] ) );
  DFF \modmult_1/xreg_reg[158]  ( .D(\modmult_1/xin[157] ), .CLK(clk), .RST(
        start_in[0]), .I(c[158]), .Q(\modmult_1/xin[158] ) );
  DFF \modmult_1/xreg_reg[157]  ( .D(\modmult_1/xin[156] ), .CLK(clk), .RST(
        start_in[0]), .I(c[157]), .Q(\modmult_1/xin[157] ) );
  DFF \modmult_1/xreg_reg[156]  ( .D(\modmult_1/xin[155] ), .CLK(clk), .RST(
        start_in[0]), .I(c[156]), .Q(\modmult_1/xin[156] ) );
  DFF \modmult_1/xreg_reg[155]  ( .D(\modmult_1/xin[154] ), .CLK(clk), .RST(
        start_in[0]), .I(c[155]), .Q(\modmult_1/xin[155] ) );
  DFF \modmult_1/xreg_reg[154]  ( .D(\modmult_1/xin[153] ), .CLK(clk), .RST(
        start_in[0]), .I(c[154]), .Q(\modmult_1/xin[154] ) );
  DFF \modmult_1/xreg_reg[153]  ( .D(\modmult_1/xin[152] ), .CLK(clk), .RST(
        start_in[0]), .I(c[153]), .Q(\modmult_1/xin[153] ) );
  DFF \modmult_1/xreg_reg[152]  ( .D(\modmult_1/xin[151] ), .CLK(clk), .RST(
        start_in[0]), .I(c[152]), .Q(\modmult_1/xin[152] ) );
  DFF \modmult_1/xreg_reg[151]  ( .D(\modmult_1/xin[150] ), .CLK(clk), .RST(
        start_in[0]), .I(c[151]), .Q(\modmult_1/xin[151] ) );
  DFF \modmult_1/xreg_reg[150]  ( .D(\modmult_1/xin[149] ), .CLK(clk), .RST(
        start_in[0]), .I(c[150]), .Q(\modmult_1/xin[150] ) );
  DFF \modmult_1/xreg_reg[149]  ( .D(\modmult_1/xin[148] ), .CLK(clk), .RST(
        start_in[0]), .I(c[149]), .Q(\modmult_1/xin[149] ) );
  DFF \modmult_1/xreg_reg[148]  ( .D(\modmult_1/xin[147] ), .CLK(clk), .RST(
        start_in[0]), .I(c[148]), .Q(\modmult_1/xin[148] ) );
  DFF \modmult_1/xreg_reg[147]  ( .D(\modmult_1/xin[146] ), .CLK(clk), .RST(
        start_in[0]), .I(c[147]), .Q(\modmult_1/xin[147] ) );
  DFF \modmult_1/xreg_reg[146]  ( .D(\modmult_1/xin[145] ), .CLK(clk), .RST(
        start_in[0]), .I(c[146]), .Q(\modmult_1/xin[146] ) );
  DFF \modmult_1/xreg_reg[145]  ( .D(\modmult_1/xin[144] ), .CLK(clk), .RST(
        start_in[0]), .I(c[145]), .Q(\modmult_1/xin[145] ) );
  DFF \modmult_1/xreg_reg[144]  ( .D(\modmult_1/xin[143] ), .CLK(clk), .RST(
        start_in[0]), .I(c[144]), .Q(\modmult_1/xin[144] ) );
  DFF \modmult_1/xreg_reg[143]  ( .D(\modmult_1/xin[142] ), .CLK(clk), .RST(
        start_in[0]), .I(c[143]), .Q(\modmult_1/xin[143] ) );
  DFF \modmult_1/xreg_reg[142]  ( .D(\modmult_1/xin[141] ), .CLK(clk), .RST(
        start_in[0]), .I(c[142]), .Q(\modmult_1/xin[142] ) );
  DFF \modmult_1/xreg_reg[141]  ( .D(\modmult_1/xin[140] ), .CLK(clk), .RST(
        start_in[0]), .I(c[141]), .Q(\modmult_1/xin[141] ) );
  DFF \modmult_1/xreg_reg[140]  ( .D(\modmult_1/xin[139] ), .CLK(clk), .RST(
        start_in[0]), .I(c[140]), .Q(\modmult_1/xin[140] ) );
  DFF \modmult_1/xreg_reg[139]  ( .D(\modmult_1/xin[138] ), .CLK(clk), .RST(
        start_in[0]), .I(c[139]), .Q(\modmult_1/xin[139] ) );
  DFF \modmult_1/xreg_reg[138]  ( .D(\modmult_1/xin[137] ), .CLK(clk), .RST(
        start_in[0]), .I(c[138]), .Q(\modmult_1/xin[138] ) );
  DFF \modmult_1/xreg_reg[137]  ( .D(\modmult_1/xin[136] ), .CLK(clk), .RST(
        start_in[0]), .I(c[137]), .Q(\modmult_1/xin[137] ) );
  DFF \modmult_1/xreg_reg[136]  ( .D(\modmult_1/xin[135] ), .CLK(clk), .RST(
        start_in[0]), .I(c[136]), .Q(\modmult_1/xin[136] ) );
  DFF \modmult_1/xreg_reg[135]  ( .D(\modmult_1/xin[134] ), .CLK(clk), .RST(
        start_in[0]), .I(c[135]), .Q(\modmult_1/xin[135] ) );
  DFF \modmult_1/xreg_reg[134]  ( .D(\modmult_1/xin[133] ), .CLK(clk), .RST(
        start_in[0]), .I(c[134]), .Q(\modmult_1/xin[134] ) );
  DFF \modmult_1/xreg_reg[133]  ( .D(\modmult_1/xin[132] ), .CLK(clk), .RST(
        start_in[0]), .I(c[133]), .Q(\modmult_1/xin[133] ) );
  DFF \modmult_1/xreg_reg[132]  ( .D(\modmult_1/xin[131] ), .CLK(clk), .RST(
        start_in[0]), .I(c[132]), .Q(\modmult_1/xin[132] ) );
  DFF \modmult_1/xreg_reg[131]  ( .D(\modmult_1/xin[130] ), .CLK(clk), .RST(
        start_in[0]), .I(c[131]), .Q(\modmult_1/xin[131] ) );
  DFF \modmult_1/xreg_reg[130]  ( .D(\modmult_1/xin[129] ), .CLK(clk), .RST(
        start_in[0]), .I(c[130]), .Q(\modmult_1/xin[130] ) );
  DFF \modmult_1/xreg_reg[129]  ( .D(\modmult_1/xin[128] ), .CLK(clk), .RST(
        start_in[0]), .I(c[129]), .Q(\modmult_1/xin[129] ) );
  DFF \modmult_1/xreg_reg[128]  ( .D(\modmult_1/xin[127] ), .CLK(clk), .RST(
        start_in[0]), .I(c[128]), .Q(\modmult_1/xin[128] ) );
  DFF \modmult_1/xreg_reg[127]  ( .D(\modmult_1/xin[126] ), .CLK(clk), .RST(
        start_in[0]), .I(c[127]), .Q(\modmult_1/xin[127] ) );
  DFF \modmult_1/xreg_reg[126]  ( .D(\modmult_1/xin[125] ), .CLK(clk), .RST(
        start_in[0]), .I(c[126]), .Q(\modmult_1/xin[126] ) );
  DFF \modmult_1/xreg_reg[125]  ( .D(\modmult_1/xin[124] ), .CLK(clk), .RST(
        start_in[0]), .I(c[125]), .Q(\modmult_1/xin[125] ) );
  DFF \modmult_1/xreg_reg[124]  ( .D(\modmult_1/xin[123] ), .CLK(clk), .RST(
        start_in[0]), .I(c[124]), .Q(\modmult_1/xin[124] ) );
  DFF \modmult_1/xreg_reg[123]  ( .D(\modmult_1/xin[122] ), .CLK(clk), .RST(
        start_in[0]), .I(c[123]), .Q(\modmult_1/xin[123] ) );
  DFF \modmult_1/xreg_reg[122]  ( .D(\modmult_1/xin[121] ), .CLK(clk), .RST(
        start_in[0]), .I(c[122]), .Q(\modmult_1/xin[122] ) );
  DFF \modmult_1/xreg_reg[121]  ( .D(\modmult_1/xin[120] ), .CLK(clk), .RST(
        start_in[0]), .I(c[121]), .Q(\modmult_1/xin[121] ) );
  DFF \modmult_1/xreg_reg[120]  ( .D(\modmult_1/xin[119] ), .CLK(clk), .RST(
        start_in[0]), .I(c[120]), .Q(\modmult_1/xin[120] ) );
  DFF \modmult_1/xreg_reg[119]  ( .D(\modmult_1/xin[118] ), .CLK(clk), .RST(
        start_in[0]), .I(c[119]), .Q(\modmult_1/xin[119] ) );
  DFF \modmult_1/xreg_reg[118]  ( .D(\modmult_1/xin[117] ), .CLK(clk), .RST(
        start_in[0]), .I(c[118]), .Q(\modmult_1/xin[118] ) );
  DFF \modmult_1/xreg_reg[117]  ( .D(\modmult_1/xin[116] ), .CLK(clk), .RST(
        start_in[0]), .I(c[117]), .Q(\modmult_1/xin[117] ) );
  DFF \modmult_1/xreg_reg[116]  ( .D(\modmult_1/xin[115] ), .CLK(clk), .RST(
        start_in[0]), .I(c[116]), .Q(\modmult_1/xin[116] ) );
  DFF \modmult_1/xreg_reg[115]  ( .D(\modmult_1/xin[114] ), .CLK(clk), .RST(
        start_in[0]), .I(c[115]), .Q(\modmult_1/xin[115] ) );
  DFF \modmult_1/xreg_reg[114]  ( .D(\modmult_1/xin[113] ), .CLK(clk), .RST(
        start_in[0]), .I(c[114]), .Q(\modmult_1/xin[114] ) );
  DFF \modmult_1/xreg_reg[113]  ( .D(\modmult_1/xin[112] ), .CLK(clk), .RST(
        start_in[0]), .I(c[113]), .Q(\modmult_1/xin[113] ) );
  DFF \modmult_1/xreg_reg[112]  ( .D(\modmult_1/xin[111] ), .CLK(clk), .RST(
        start_in[0]), .I(c[112]), .Q(\modmult_1/xin[112] ) );
  DFF \modmult_1/xreg_reg[111]  ( .D(\modmult_1/xin[110] ), .CLK(clk), .RST(
        start_in[0]), .I(c[111]), .Q(\modmult_1/xin[111] ) );
  DFF \modmult_1/xreg_reg[110]  ( .D(\modmult_1/xin[109] ), .CLK(clk), .RST(
        start_in[0]), .I(c[110]), .Q(\modmult_1/xin[110] ) );
  DFF \modmult_1/xreg_reg[109]  ( .D(\modmult_1/xin[108] ), .CLK(clk), .RST(
        start_in[0]), .I(c[109]), .Q(\modmult_1/xin[109] ) );
  DFF \modmult_1/xreg_reg[108]  ( .D(\modmult_1/xin[107] ), .CLK(clk), .RST(
        start_in[0]), .I(c[108]), .Q(\modmult_1/xin[108] ) );
  DFF \modmult_1/xreg_reg[107]  ( .D(\modmult_1/xin[106] ), .CLK(clk), .RST(
        start_in[0]), .I(c[107]), .Q(\modmult_1/xin[107] ) );
  DFF \modmult_1/xreg_reg[106]  ( .D(\modmult_1/xin[105] ), .CLK(clk), .RST(
        start_in[0]), .I(c[106]), .Q(\modmult_1/xin[106] ) );
  DFF \modmult_1/xreg_reg[105]  ( .D(\modmult_1/xin[104] ), .CLK(clk), .RST(
        start_in[0]), .I(c[105]), .Q(\modmult_1/xin[105] ) );
  DFF \modmult_1/xreg_reg[104]  ( .D(\modmult_1/xin[103] ), .CLK(clk), .RST(
        start_in[0]), .I(c[104]), .Q(\modmult_1/xin[104] ) );
  DFF \modmult_1/xreg_reg[103]  ( .D(\modmult_1/xin[102] ), .CLK(clk), .RST(
        start_in[0]), .I(c[103]), .Q(\modmult_1/xin[103] ) );
  DFF \modmult_1/xreg_reg[102]  ( .D(\modmult_1/xin[101] ), .CLK(clk), .RST(
        start_in[0]), .I(c[102]), .Q(\modmult_1/xin[102] ) );
  DFF \modmult_1/xreg_reg[101]  ( .D(\modmult_1/xin[100] ), .CLK(clk), .RST(
        start_in[0]), .I(c[101]), .Q(\modmult_1/xin[101] ) );
  DFF \modmult_1/xreg_reg[100]  ( .D(\modmult_1/xin[99] ), .CLK(clk), .RST(
        start_in[0]), .I(c[100]), .Q(\modmult_1/xin[100] ) );
  DFF \modmult_1/xreg_reg[99]  ( .D(\modmult_1/xin[98] ), .CLK(clk), .RST(
        start_in[0]), .I(c[99]), .Q(\modmult_1/xin[99] ) );
  DFF \modmult_1/xreg_reg[98]  ( .D(\modmult_1/xin[97] ), .CLK(clk), .RST(
        start_in[0]), .I(c[98]), .Q(\modmult_1/xin[98] ) );
  DFF \modmult_1/xreg_reg[97]  ( .D(\modmult_1/xin[96] ), .CLK(clk), .RST(
        start_in[0]), .I(c[97]), .Q(\modmult_1/xin[97] ) );
  DFF \modmult_1/xreg_reg[96]  ( .D(\modmult_1/xin[95] ), .CLK(clk), .RST(
        start_in[0]), .I(c[96]), .Q(\modmult_1/xin[96] ) );
  DFF \modmult_1/xreg_reg[95]  ( .D(\modmult_1/xin[94] ), .CLK(clk), .RST(
        start_in[0]), .I(c[95]), .Q(\modmult_1/xin[95] ) );
  DFF \modmult_1/xreg_reg[94]  ( .D(\modmult_1/xin[93] ), .CLK(clk), .RST(
        start_in[0]), .I(c[94]), .Q(\modmult_1/xin[94] ) );
  DFF \modmult_1/xreg_reg[93]  ( .D(\modmult_1/xin[92] ), .CLK(clk), .RST(
        start_in[0]), .I(c[93]), .Q(\modmult_1/xin[93] ) );
  DFF \modmult_1/xreg_reg[92]  ( .D(\modmult_1/xin[91] ), .CLK(clk), .RST(
        start_in[0]), .I(c[92]), .Q(\modmult_1/xin[92] ) );
  DFF \modmult_1/xreg_reg[91]  ( .D(\modmult_1/xin[90] ), .CLK(clk), .RST(
        start_in[0]), .I(c[91]), .Q(\modmult_1/xin[91] ) );
  DFF \modmult_1/xreg_reg[90]  ( .D(\modmult_1/xin[89] ), .CLK(clk), .RST(
        start_in[0]), .I(c[90]), .Q(\modmult_1/xin[90] ) );
  DFF \modmult_1/xreg_reg[89]  ( .D(\modmult_1/xin[88] ), .CLK(clk), .RST(
        start_in[0]), .I(c[89]), .Q(\modmult_1/xin[89] ) );
  DFF \modmult_1/xreg_reg[88]  ( .D(\modmult_1/xin[87] ), .CLK(clk), .RST(
        start_in[0]), .I(c[88]), .Q(\modmult_1/xin[88] ) );
  DFF \modmult_1/xreg_reg[87]  ( .D(\modmult_1/xin[86] ), .CLK(clk), .RST(
        start_in[0]), .I(c[87]), .Q(\modmult_1/xin[87] ) );
  DFF \modmult_1/xreg_reg[86]  ( .D(\modmult_1/xin[85] ), .CLK(clk), .RST(
        start_in[0]), .I(c[86]), .Q(\modmult_1/xin[86] ) );
  DFF \modmult_1/xreg_reg[85]  ( .D(\modmult_1/xin[84] ), .CLK(clk), .RST(
        start_in[0]), .I(c[85]), .Q(\modmult_1/xin[85] ) );
  DFF \modmult_1/xreg_reg[84]  ( .D(\modmult_1/xin[83] ), .CLK(clk), .RST(
        start_in[0]), .I(c[84]), .Q(\modmult_1/xin[84] ) );
  DFF \modmult_1/xreg_reg[83]  ( .D(\modmult_1/xin[82] ), .CLK(clk), .RST(
        start_in[0]), .I(c[83]), .Q(\modmult_1/xin[83] ) );
  DFF \modmult_1/xreg_reg[82]  ( .D(\modmult_1/xin[81] ), .CLK(clk), .RST(
        start_in[0]), .I(c[82]), .Q(\modmult_1/xin[82] ) );
  DFF \modmult_1/xreg_reg[81]  ( .D(\modmult_1/xin[80] ), .CLK(clk), .RST(
        start_in[0]), .I(c[81]), .Q(\modmult_1/xin[81] ) );
  DFF \modmult_1/xreg_reg[80]  ( .D(\modmult_1/xin[79] ), .CLK(clk), .RST(
        start_in[0]), .I(c[80]), .Q(\modmult_1/xin[80] ) );
  DFF \modmult_1/xreg_reg[79]  ( .D(\modmult_1/xin[78] ), .CLK(clk), .RST(
        start_in[0]), .I(c[79]), .Q(\modmult_1/xin[79] ) );
  DFF \modmult_1/xreg_reg[78]  ( .D(\modmult_1/xin[77] ), .CLK(clk), .RST(
        start_in[0]), .I(c[78]), .Q(\modmult_1/xin[78] ) );
  DFF \modmult_1/xreg_reg[77]  ( .D(\modmult_1/xin[76] ), .CLK(clk), .RST(
        start_in[0]), .I(c[77]), .Q(\modmult_1/xin[77] ) );
  DFF \modmult_1/xreg_reg[76]  ( .D(\modmult_1/xin[75] ), .CLK(clk), .RST(
        start_in[0]), .I(c[76]), .Q(\modmult_1/xin[76] ) );
  DFF \modmult_1/xreg_reg[75]  ( .D(\modmult_1/xin[74] ), .CLK(clk), .RST(
        start_in[0]), .I(c[75]), .Q(\modmult_1/xin[75] ) );
  DFF \modmult_1/xreg_reg[74]  ( .D(\modmult_1/xin[73] ), .CLK(clk), .RST(
        start_in[0]), .I(c[74]), .Q(\modmult_1/xin[74] ) );
  DFF \modmult_1/xreg_reg[73]  ( .D(\modmult_1/xin[72] ), .CLK(clk), .RST(
        start_in[0]), .I(c[73]), .Q(\modmult_1/xin[73] ) );
  DFF \modmult_1/xreg_reg[72]  ( .D(\modmult_1/xin[71] ), .CLK(clk), .RST(
        start_in[0]), .I(c[72]), .Q(\modmult_1/xin[72] ) );
  DFF \modmult_1/xreg_reg[71]  ( .D(\modmult_1/xin[70] ), .CLK(clk), .RST(
        start_in[0]), .I(c[71]), .Q(\modmult_1/xin[71] ) );
  DFF \modmult_1/xreg_reg[70]  ( .D(\modmult_1/xin[69] ), .CLK(clk), .RST(
        start_in[0]), .I(c[70]), .Q(\modmult_1/xin[70] ) );
  DFF \modmult_1/xreg_reg[69]  ( .D(\modmult_1/xin[68] ), .CLK(clk), .RST(
        start_in[0]), .I(c[69]), .Q(\modmult_1/xin[69] ) );
  DFF \modmult_1/xreg_reg[68]  ( .D(\modmult_1/xin[67] ), .CLK(clk), .RST(
        start_in[0]), .I(c[68]), .Q(\modmult_1/xin[68] ) );
  DFF \modmult_1/xreg_reg[67]  ( .D(\modmult_1/xin[66] ), .CLK(clk), .RST(
        start_in[0]), .I(c[67]), .Q(\modmult_1/xin[67] ) );
  DFF \modmult_1/xreg_reg[66]  ( .D(\modmult_1/xin[65] ), .CLK(clk), .RST(
        start_in[0]), .I(c[66]), .Q(\modmult_1/xin[66] ) );
  DFF \modmult_1/xreg_reg[65]  ( .D(\modmult_1/xin[64] ), .CLK(clk), .RST(
        start_in[0]), .I(c[65]), .Q(\modmult_1/xin[65] ) );
  DFF \modmult_1/xreg_reg[64]  ( .D(\modmult_1/xin[63] ), .CLK(clk), .RST(
        start_in[0]), .I(c[64]), .Q(\modmult_1/xin[64] ) );
  DFF \modmult_1/xreg_reg[63]  ( .D(\modmult_1/xin[62] ), .CLK(clk), .RST(
        start_in[0]), .I(c[63]), .Q(\modmult_1/xin[63] ) );
  DFF \modmult_1/xreg_reg[62]  ( .D(\modmult_1/xin[61] ), .CLK(clk), .RST(
        start_in[0]), .I(c[62]), .Q(\modmult_1/xin[62] ) );
  DFF \modmult_1/xreg_reg[61]  ( .D(\modmult_1/xin[60] ), .CLK(clk), .RST(
        start_in[0]), .I(c[61]), .Q(\modmult_1/xin[61] ) );
  DFF \modmult_1/xreg_reg[60]  ( .D(\modmult_1/xin[59] ), .CLK(clk), .RST(
        start_in[0]), .I(c[60]), .Q(\modmult_1/xin[60] ) );
  DFF \modmult_1/xreg_reg[59]  ( .D(\modmult_1/xin[58] ), .CLK(clk), .RST(
        start_in[0]), .I(c[59]), .Q(\modmult_1/xin[59] ) );
  DFF \modmult_1/xreg_reg[58]  ( .D(\modmult_1/xin[57] ), .CLK(clk), .RST(
        start_in[0]), .I(c[58]), .Q(\modmult_1/xin[58] ) );
  DFF \modmult_1/xreg_reg[57]  ( .D(\modmult_1/xin[56] ), .CLK(clk), .RST(
        start_in[0]), .I(c[57]), .Q(\modmult_1/xin[57] ) );
  DFF \modmult_1/xreg_reg[56]  ( .D(\modmult_1/xin[55] ), .CLK(clk), .RST(
        start_in[0]), .I(c[56]), .Q(\modmult_1/xin[56] ) );
  DFF \modmult_1/xreg_reg[55]  ( .D(\modmult_1/xin[54] ), .CLK(clk), .RST(
        start_in[0]), .I(c[55]), .Q(\modmult_1/xin[55] ) );
  DFF \modmult_1/xreg_reg[54]  ( .D(\modmult_1/xin[53] ), .CLK(clk), .RST(
        start_in[0]), .I(c[54]), .Q(\modmult_1/xin[54] ) );
  DFF \modmult_1/xreg_reg[53]  ( .D(\modmult_1/xin[52] ), .CLK(clk), .RST(
        start_in[0]), .I(c[53]), .Q(\modmult_1/xin[53] ) );
  DFF \modmult_1/xreg_reg[52]  ( .D(\modmult_1/xin[51] ), .CLK(clk), .RST(
        start_in[0]), .I(c[52]), .Q(\modmult_1/xin[52] ) );
  DFF \modmult_1/xreg_reg[51]  ( .D(\modmult_1/xin[50] ), .CLK(clk), .RST(
        start_in[0]), .I(c[51]), .Q(\modmult_1/xin[51] ) );
  DFF \modmult_1/xreg_reg[50]  ( .D(\modmult_1/xin[49] ), .CLK(clk), .RST(
        start_in[0]), .I(c[50]), .Q(\modmult_1/xin[50] ) );
  DFF \modmult_1/xreg_reg[49]  ( .D(\modmult_1/xin[48] ), .CLK(clk), .RST(
        start_in[0]), .I(c[49]), .Q(\modmult_1/xin[49] ) );
  DFF \modmult_1/xreg_reg[48]  ( .D(\modmult_1/xin[47] ), .CLK(clk), .RST(
        start_in[0]), .I(c[48]), .Q(\modmult_1/xin[48] ) );
  DFF \modmult_1/xreg_reg[47]  ( .D(\modmult_1/xin[46] ), .CLK(clk), .RST(
        start_in[0]), .I(c[47]), .Q(\modmult_1/xin[47] ) );
  DFF \modmult_1/xreg_reg[46]  ( .D(\modmult_1/xin[45] ), .CLK(clk), .RST(
        start_in[0]), .I(c[46]), .Q(\modmult_1/xin[46] ) );
  DFF \modmult_1/xreg_reg[45]  ( .D(\modmult_1/xin[44] ), .CLK(clk), .RST(
        start_in[0]), .I(c[45]), .Q(\modmult_1/xin[45] ) );
  DFF \modmult_1/xreg_reg[44]  ( .D(\modmult_1/xin[43] ), .CLK(clk), .RST(
        start_in[0]), .I(c[44]), .Q(\modmult_1/xin[44] ) );
  DFF \modmult_1/xreg_reg[43]  ( .D(\modmult_1/xin[42] ), .CLK(clk), .RST(
        start_in[0]), .I(c[43]), .Q(\modmult_1/xin[43] ) );
  DFF \modmult_1/xreg_reg[42]  ( .D(\modmult_1/xin[41] ), .CLK(clk), .RST(
        start_in[0]), .I(c[42]), .Q(\modmult_1/xin[42] ) );
  DFF \modmult_1/xreg_reg[41]  ( .D(\modmult_1/xin[40] ), .CLK(clk), .RST(
        start_in[0]), .I(c[41]), .Q(\modmult_1/xin[41] ) );
  DFF \modmult_1/xreg_reg[40]  ( .D(\modmult_1/xin[39] ), .CLK(clk), .RST(
        start_in[0]), .I(c[40]), .Q(\modmult_1/xin[40] ) );
  DFF \modmult_1/xreg_reg[39]  ( .D(\modmult_1/xin[38] ), .CLK(clk), .RST(
        start_in[0]), .I(c[39]), .Q(\modmult_1/xin[39] ) );
  DFF \modmult_1/xreg_reg[38]  ( .D(\modmult_1/xin[37] ), .CLK(clk), .RST(
        start_in[0]), .I(c[38]), .Q(\modmult_1/xin[38] ) );
  DFF \modmult_1/xreg_reg[37]  ( .D(\modmult_1/xin[36] ), .CLK(clk), .RST(
        start_in[0]), .I(c[37]), .Q(\modmult_1/xin[37] ) );
  DFF \modmult_1/xreg_reg[36]  ( .D(\modmult_1/xin[35] ), .CLK(clk), .RST(
        start_in[0]), .I(c[36]), .Q(\modmult_1/xin[36] ) );
  DFF \modmult_1/xreg_reg[35]  ( .D(\modmult_1/xin[34] ), .CLK(clk), .RST(
        start_in[0]), .I(c[35]), .Q(\modmult_1/xin[35] ) );
  DFF \modmult_1/xreg_reg[34]  ( .D(\modmult_1/xin[33] ), .CLK(clk), .RST(
        start_in[0]), .I(c[34]), .Q(\modmult_1/xin[34] ) );
  DFF \modmult_1/xreg_reg[33]  ( .D(\modmult_1/xin[32] ), .CLK(clk), .RST(
        start_in[0]), .I(c[33]), .Q(\modmult_1/xin[33] ) );
  DFF \modmult_1/xreg_reg[32]  ( .D(\modmult_1/xin[31] ), .CLK(clk), .RST(
        start_in[0]), .I(c[32]), .Q(\modmult_1/xin[32] ) );
  DFF \modmult_1/xreg_reg[31]  ( .D(\modmult_1/xin[30] ), .CLK(clk), .RST(
        start_in[0]), .I(c[31]), .Q(\modmult_1/xin[31] ) );
  DFF \modmult_1/xreg_reg[30]  ( .D(\modmult_1/xin[29] ), .CLK(clk), .RST(
        start_in[0]), .I(c[30]), .Q(\modmult_1/xin[30] ) );
  DFF \modmult_1/xreg_reg[29]  ( .D(\modmult_1/xin[28] ), .CLK(clk), .RST(
        start_in[0]), .I(c[29]), .Q(\modmult_1/xin[29] ) );
  DFF \modmult_1/xreg_reg[28]  ( .D(\modmult_1/xin[27] ), .CLK(clk), .RST(
        start_in[0]), .I(c[28]), .Q(\modmult_1/xin[28] ) );
  DFF \modmult_1/xreg_reg[27]  ( .D(\modmult_1/xin[26] ), .CLK(clk), .RST(
        start_in[0]), .I(c[27]), .Q(\modmult_1/xin[27] ) );
  DFF \modmult_1/xreg_reg[26]  ( .D(\modmult_1/xin[25] ), .CLK(clk), .RST(
        start_in[0]), .I(c[26]), .Q(\modmult_1/xin[26] ) );
  DFF \modmult_1/xreg_reg[25]  ( .D(\modmult_1/xin[24] ), .CLK(clk), .RST(
        start_in[0]), .I(c[25]), .Q(\modmult_1/xin[25] ) );
  DFF \modmult_1/xreg_reg[24]  ( .D(\modmult_1/xin[23] ), .CLK(clk), .RST(
        start_in[0]), .I(c[24]), .Q(\modmult_1/xin[24] ) );
  DFF \modmult_1/xreg_reg[23]  ( .D(\modmult_1/xin[22] ), .CLK(clk), .RST(
        start_in[0]), .I(c[23]), .Q(\modmult_1/xin[23] ) );
  DFF \modmult_1/xreg_reg[22]  ( .D(\modmult_1/xin[21] ), .CLK(clk), .RST(
        start_in[0]), .I(c[22]), .Q(\modmult_1/xin[22] ) );
  DFF \modmult_1/xreg_reg[21]  ( .D(\modmult_1/xin[20] ), .CLK(clk), .RST(
        start_in[0]), .I(c[21]), .Q(\modmult_1/xin[21] ) );
  DFF \modmult_1/xreg_reg[20]  ( .D(\modmult_1/xin[19] ), .CLK(clk), .RST(
        start_in[0]), .I(c[20]), .Q(\modmult_1/xin[20] ) );
  DFF \modmult_1/xreg_reg[19]  ( .D(\modmult_1/xin[18] ), .CLK(clk), .RST(
        start_in[0]), .I(c[19]), .Q(\modmult_1/xin[19] ) );
  DFF \modmult_1/xreg_reg[18]  ( .D(\modmult_1/xin[17] ), .CLK(clk), .RST(
        start_in[0]), .I(c[18]), .Q(\modmult_1/xin[18] ) );
  DFF \modmult_1/xreg_reg[17]  ( .D(\modmult_1/xin[16] ), .CLK(clk), .RST(
        start_in[0]), .I(c[17]), .Q(\modmult_1/xin[17] ) );
  DFF \modmult_1/xreg_reg[16]  ( .D(\modmult_1/xin[15] ), .CLK(clk), .RST(
        start_in[0]), .I(c[16]), .Q(\modmult_1/xin[16] ) );
  DFF \modmult_1/xreg_reg[15]  ( .D(\modmult_1/xin[14] ), .CLK(clk), .RST(
        start_in[0]), .I(c[15]), .Q(\modmult_1/xin[15] ) );
  DFF \modmult_1/xreg_reg[14]  ( .D(\modmult_1/xin[13] ), .CLK(clk), .RST(
        start_in[0]), .I(c[14]), .Q(\modmult_1/xin[14] ) );
  DFF \modmult_1/xreg_reg[13]  ( .D(\modmult_1/xin[12] ), .CLK(clk), .RST(
        start_in[0]), .I(c[13]), .Q(\modmult_1/xin[13] ) );
  DFF \modmult_1/xreg_reg[12]  ( .D(\modmult_1/xin[11] ), .CLK(clk), .RST(
        start_in[0]), .I(c[12]), .Q(\modmult_1/xin[12] ) );
  DFF \modmult_1/xreg_reg[11]  ( .D(\modmult_1/xin[10] ), .CLK(clk), .RST(
        start_in[0]), .I(c[11]), .Q(\modmult_1/xin[11] ) );
  DFF \modmult_1/xreg_reg[10]  ( .D(\modmult_1/xin[9] ), .CLK(clk), .RST(
        start_in[0]), .I(c[10]), .Q(\modmult_1/xin[10] ) );
  DFF \modmult_1/xreg_reg[9]  ( .D(\modmult_1/xin[8] ), .CLK(clk), .RST(
        start_in[0]), .I(c[9]), .Q(\modmult_1/xin[9] ) );
  DFF \modmult_1/xreg_reg[8]  ( .D(\modmult_1/xin[7] ), .CLK(clk), .RST(
        start_in[0]), .I(c[8]), .Q(\modmult_1/xin[8] ) );
  DFF \modmult_1/xreg_reg[7]  ( .D(\modmult_1/xin[6] ), .CLK(clk), .RST(
        start_in[0]), .I(c[7]), .Q(\modmult_1/xin[7] ) );
  DFF \modmult_1/xreg_reg[6]  ( .D(\modmult_1/xin[5] ), .CLK(clk), .RST(
        start_in[0]), .I(c[6]), .Q(\modmult_1/xin[6] ) );
  DFF \modmult_1/xreg_reg[5]  ( .D(\modmult_1/xin[4] ), .CLK(clk), .RST(
        start_in[0]), .I(c[5]), .Q(\modmult_1/xin[5] ) );
  DFF \modmult_1/xreg_reg[4]  ( .D(\modmult_1/xin[3] ), .CLK(clk), .RST(
        start_in[0]), .I(c[4]), .Q(\modmult_1/xin[4] ) );
  DFF \modmult_1/xreg_reg[3]  ( .D(\modmult_1/xin[2] ), .CLK(clk), .RST(
        start_in[0]), .I(c[3]), .Q(\modmult_1/xin[3] ) );
  DFF \modmult_1/xreg_reg[2]  ( .D(\modmult_1/xin[1] ), .CLK(clk), .RST(
        start_in[0]), .I(c[2]), .Q(\modmult_1/xin[2] ) );
  DFF \modmult_1/xreg_reg[1]  ( .D(\modmult_1/xin[0] ), .CLK(clk), .RST(
        start_in[0]), .I(c[1]), .Q(\modmult_1/xin[1] ) );
  DFF \modmult_1/xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start_in[0]), .I(
        c[0]), .Q(\modmult_1/xin[0] ) );
  XOR U1036 ( .A(start_in[1023]), .B(mul_pow), .Z(n8) );
  NANDN U1037 ( .A(first_one), .B(n1033), .Z(n6) );
  NAND U1038 ( .A(n1034), .B(ein[1023]), .Z(n1033) );
  AND U1039 ( .A(start_in[1023]), .B(mul_pow), .Z(n1034) );
  XOR U1040 ( .A(n1035), .B(n1036), .Z(\modmult_1/zout[0][1024] ) );
  XOR U1041 ( .A(n1037), .B(n1038), .Z(n1036) );
  ANDN U1042 ( .B(n1039), .A(n1040), .Z(n1037) );
  XOR U1043 ( .A(n1041), .B(n1042), .Z(n1039) );
  XOR U1044 ( .A(ein[8]), .B(n1043), .Z(ereg_next[9]) );
  AND U1045 ( .A(mul_pow), .B(n1044), .Z(n1043) );
  XOR U1046 ( .A(ein[9]), .B(ein[8]), .Z(n1044) );
  XOR U1047 ( .A(ein[98]), .B(n1045), .Z(ereg_next[99]) );
  AND U1048 ( .A(mul_pow), .B(n1046), .Z(n1045) );
  XOR U1049 ( .A(ein[99]), .B(ein[98]), .Z(n1046) );
  XOR U1050 ( .A(ein[998]), .B(n1047), .Z(ereg_next[999]) );
  AND U1051 ( .A(mul_pow), .B(n1048), .Z(n1047) );
  XOR U1052 ( .A(ein[999]), .B(ein[998]), .Z(n1048) );
  XOR U1053 ( .A(ein[997]), .B(n1049), .Z(ereg_next[998]) );
  AND U1054 ( .A(mul_pow), .B(n1050), .Z(n1049) );
  XOR U1055 ( .A(ein[998]), .B(ein[997]), .Z(n1050) );
  XOR U1056 ( .A(ein[996]), .B(n1051), .Z(ereg_next[997]) );
  AND U1057 ( .A(mul_pow), .B(n1052), .Z(n1051) );
  XOR U1058 ( .A(ein[997]), .B(ein[996]), .Z(n1052) );
  XOR U1059 ( .A(ein[995]), .B(n1053), .Z(ereg_next[996]) );
  AND U1060 ( .A(mul_pow), .B(n1054), .Z(n1053) );
  XOR U1061 ( .A(ein[996]), .B(ein[995]), .Z(n1054) );
  XOR U1062 ( .A(ein[994]), .B(n1055), .Z(ereg_next[995]) );
  AND U1063 ( .A(mul_pow), .B(n1056), .Z(n1055) );
  XOR U1064 ( .A(ein[995]), .B(ein[994]), .Z(n1056) );
  XOR U1065 ( .A(ein[993]), .B(n1057), .Z(ereg_next[994]) );
  AND U1066 ( .A(mul_pow), .B(n1058), .Z(n1057) );
  XOR U1067 ( .A(ein[994]), .B(ein[993]), .Z(n1058) );
  XOR U1068 ( .A(ein[992]), .B(n1059), .Z(ereg_next[993]) );
  AND U1069 ( .A(mul_pow), .B(n1060), .Z(n1059) );
  XOR U1070 ( .A(ein[993]), .B(ein[992]), .Z(n1060) );
  XOR U1071 ( .A(ein[991]), .B(n1061), .Z(ereg_next[992]) );
  AND U1072 ( .A(mul_pow), .B(n1062), .Z(n1061) );
  XOR U1073 ( .A(ein[992]), .B(ein[991]), .Z(n1062) );
  XOR U1074 ( .A(ein[990]), .B(n1063), .Z(ereg_next[991]) );
  AND U1075 ( .A(mul_pow), .B(n1064), .Z(n1063) );
  XOR U1076 ( .A(ein[991]), .B(ein[990]), .Z(n1064) );
  XOR U1077 ( .A(ein[989]), .B(n1065), .Z(ereg_next[990]) );
  AND U1078 ( .A(mul_pow), .B(n1066), .Z(n1065) );
  XOR U1079 ( .A(ein[990]), .B(ein[989]), .Z(n1066) );
  XOR U1080 ( .A(ein[97]), .B(n1067), .Z(ereg_next[98]) );
  AND U1081 ( .A(mul_pow), .B(n1068), .Z(n1067) );
  XOR U1082 ( .A(ein[98]), .B(ein[97]), .Z(n1068) );
  XOR U1083 ( .A(ein[988]), .B(n1069), .Z(ereg_next[989]) );
  AND U1084 ( .A(mul_pow), .B(n1070), .Z(n1069) );
  XOR U1085 ( .A(ein[989]), .B(ein[988]), .Z(n1070) );
  XOR U1086 ( .A(ein[987]), .B(n1071), .Z(ereg_next[988]) );
  AND U1087 ( .A(mul_pow), .B(n1072), .Z(n1071) );
  XOR U1088 ( .A(ein[988]), .B(ein[987]), .Z(n1072) );
  XOR U1089 ( .A(ein[986]), .B(n1073), .Z(ereg_next[987]) );
  AND U1090 ( .A(mul_pow), .B(n1074), .Z(n1073) );
  XOR U1091 ( .A(ein[987]), .B(ein[986]), .Z(n1074) );
  XOR U1092 ( .A(ein[985]), .B(n1075), .Z(ereg_next[986]) );
  AND U1093 ( .A(mul_pow), .B(n1076), .Z(n1075) );
  XOR U1094 ( .A(ein[986]), .B(ein[985]), .Z(n1076) );
  XOR U1095 ( .A(ein[984]), .B(n1077), .Z(ereg_next[985]) );
  AND U1096 ( .A(mul_pow), .B(n1078), .Z(n1077) );
  XOR U1097 ( .A(ein[985]), .B(ein[984]), .Z(n1078) );
  XOR U1098 ( .A(ein[983]), .B(n1079), .Z(ereg_next[984]) );
  AND U1099 ( .A(mul_pow), .B(n1080), .Z(n1079) );
  XOR U1100 ( .A(ein[984]), .B(ein[983]), .Z(n1080) );
  XOR U1101 ( .A(ein[982]), .B(n1081), .Z(ereg_next[983]) );
  AND U1102 ( .A(mul_pow), .B(n1082), .Z(n1081) );
  XOR U1103 ( .A(ein[983]), .B(ein[982]), .Z(n1082) );
  XOR U1104 ( .A(ein[981]), .B(n1083), .Z(ereg_next[982]) );
  AND U1105 ( .A(mul_pow), .B(n1084), .Z(n1083) );
  XOR U1106 ( .A(ein[982]), .B(ein[981]), .Z(n1084) );
  XOR U1107 ( .A(ein[980]), .B(n1085), .Z(ereg_next[981]) );
  AND U1108 ( .A(mul_pow), .B(n1086), .Z(n1085) );
  XOR U1109 ( .A(ein[981]), .B(ein[980]), .Z(n1086) );
  XOR U1110 ( .A(ein[979]), .B(n1087), .Z(ereg_next[980]) );
  AND U1111 ( .A(mul_pow), .B(n1088), .Z(n1087) );
  XOR U1112 ( .A(ein[980]), .B(ein[979]), .Z(n1088) );
  XOR U1113 ( .A(ein[96]), .B(n1089), .Z(ereg_next[97]) );
  AND U1114 ( .A(mul_pow), .B(n1090), .Z(n1089) );
  XOR U1115 ( .A(ein[97]), .B(ein[96]), .Z(n1090) );
  XOR U1116 ( .A(ein[978]), .B(n1091), .Z(ereg_next[979]) );
  AND U1117 ( .A(mul_pow), .B(n1092), .Z(n1091) );
  XOR U1118 ( .A(ein[979]), .B(ein[978]), .Z(n1092) );
  XOR U1119 ( .A(ein[977]), .B(n1093), .Z(ereg_next[978]) );
  AND U1120 ( .A(mul_pow), .B(n1094), .Z(n1093) );
  XOR U1121 ( .A(ein[978]), .B(ein[977]), .Z(n1094) );
  XOR U1122 ( .A(ein[976]), .B(n1095), .Z(ereg_next[977]) );
  AND U1123 ( .A(mul_pow), .B(n1096), .Z(n1095) );
  XOR U1124 ( .A(ein[977]), .B(ein[976]), .Z(n1096) );
  XOR U1125 ( .A(ein[975]), .B(n1097), .Z(ereg_next[976]) );
  AND U1126 ( .A(mul_pow), .B(n1098), .Z(n1097) );
  XOR U1127 ( .A(ein[976]), .B(ein[975]), .Z(n1098) );
  XOR U1128 ( .A(ein[974]), .B(n1099), .Z(ereg_next[975]) );
  AND U1129 ( .A(mul_pow), .B(n1100), .Z(n1099) );
  XOR U1130 ( .A(ein[975]), .B(ein[974]), .Z(n1100) );
  XOR U1131 ( .A(ein[973]), .B(n1101), .Z(ereg_next[974]) );
  AND U1132 ( .A(mul_pow), .B(n1102), .Z(n1101) );
  XOR U1133 ( .A(ein[974]), .B(ein[973]), .Z(n1102) );
  XOR U1134 ( .A(ein[972]), .B(n1103), .Z(ereg_next[973]) );
  AND U1135 ( .A(mul_pow), .B(n1104), .Z(n1103) );
  XOR U1136 ( .A(ein[973]), .B(ein[972]), .Z(n1104) );
  XOR U1137 ( .A(ein[971]), .B(n1105), .Z(ereg_next[972]) );
  AND U1138 ( .A(mul_pow), .B(n1106), .Z(n1105) );
  XOR U1139 ( .A(ein[972]), .B(ein[971]), .Z(n1106) );
  XOR U1140 ( .A(ein[970]), .B(n1107), .Z(ereg_next[971]) );
  AND U1141 ( .A(mul_pow), .B(n1108), .Z(n1107) );
  XOR U1142 ( .A(ein[971]), .B(ein[970]), .Z(n1108) );
  XOR U1143 ( .A(ein[969]), .B(n1109), .Z(ereg_next[970]) );
  AND U1144 ( .A(mul_pow), .B(n1110), .Z(n1109) );
  XOR U1145 ( .A(ein[970]), .B(ein[969]), .Z(n1110) );
  XOR U1146 ( .A(ein[95]), .B(n1111), .Z(ereg_next[96]) );
  AND U1147 ( .A(mul_pow), .B(n1112), .Z(n1111) );
  XOR U1148 ( .A(ein[96]), .B(ein[95]), .Z(n1112) );
  XOR U1149 ( .A(ein[968]), .B(n1113), .Z(ereg_next[969]) );
  AND U1150 ( .A(mul_pow), .B(n1114), .Z(n1113) );
  XOR U1151 ( .A(ein[969]), .B(ein[968]), .Z(n1114) );
  XOR U1152 ( .A(ein[967]), .B(n1115), .Z(ereg_next[968]) );
  AND U1153 ( .A(mul_pow), .B(n1116), .Z(n1115) );
  XOR U1154 ( .A(ein[968]), .B(ein[967]), .Z(n1116) );
  XOR U1155 ( .A(ein[966]), .B(n1117), .Z(ereg_next[967]) );
  AND U1156 ( .A(mul_pow), .B(n1118), .Z(n1117) );
  XOR U1157 ( .A(ein[967]), .B(ein[966]), .Z(n1118) );
  XOR U1158 ( .A(ein[965]), .B(n1119), .Z(ereg_next[966]) );
  AND U1159 ( .A(mul_pow), .B(n1120), .Z(n1119) );
  XOR U1160 ( .A(ein[966]), .B(ein[965]), .Z(n1120) );
  XOR U1161 ( .A(ein[964]), .B(n1121), .Z(ereg_next[965]) );
  AND U1162 ( .A(mul_pow), .B(n1122), .Z(n1121) );
  XOR U1163 ( .A(ein[965]), .B(ein[964]), .Z(n1122) );
  XOR U1164 ( .A(ein[963]), .B(n1123), .Z(ereg_next[964]) );
  AND U1165 ( .A(mul_pow), .B(n1124), .Z(n1123) );
  XOR U1166 ( .A(ein[964]), .B(ein[963]), .Z(n1124) );
  XOR U1167 ( .A(ein[962]), .B(n1125), .Z(ereg_next[963]) );
  AND U1168 ( .A(mul_pow), .B(n1126), .Z(n1125) );
  XOR U1169 ( .A(ein[963]), .B(ein[962]), .Z(n1126) );
  XOR U1170 ( .A(ein[961]), .B(n1127), .Z(ereg_next[962]) );
  AND U1171 ( .A(mul_pow), .B(n1128), .Z(n1127) );
  XOR U1172 ( .A(ein[962]), .B(ein[961]), .Z(n1128) );
  XOR U1173 ( .A(ein[960]), .B(n1129), .Z(ereg_next[961]) );
  AND U1174 ( .A(mul_pow), .B(n1130), .Z(n1129) );
  XOR U1175 ( .A(ein[961]), .B(ein[960]), .Z(n1130) );
  XOR U1176 ( .A(ein[959]), .B(n1131), .Z(ereg_next[960]) );
  AND U1177 ( .A(mul_pow), .B(n1132), .Z(n1131) );
  XOR U1178 ( .A(ein[960]), .B(ein[959]), .Z(n1132) );
  XOR U1179 ( .A(ein[94]), .B(n1133), .Z(ereg_next[95]) );
  AND U1180 ( .A(mul_pow), .B(n1134), .Z(n1133) );
  XOR U1181 ( .A(ein[95]), .B(ein[94]), .Z(n1134) );
  XOR U1182 ( .A(ein[958]), .B(n1135), .Z(ereg_next[959]) );
  AND U1183 ( .A(mul_pow), .B(n1136), .Z(n1135) );
  XOR U1184 ( .A(ein[959]), .B(ein[958]), .Z(n1136) );
  XOR U1185 ( .A(ein[957]), .B(n1137), .Z(ereg_next[958]) );
  AND U1186 ( .A(mul_pow), .B(n1138), .Z(n1137) );
  XOR U1187 ( .A(ein[958]), .B(ein[957]), .Z(n1138) );
  XOR U1188 ( .A(ein[956]), .B(n1139), .Z(ereg_next[957]) );
  AND U1189 ( .A(mul_pow), .B(n1140), .Z(n1139) );
  XOR U1190 ( .A(ein[957]), .B(ein[956]), .Z(n1140) );
  XOR U1191 ( .A(ein[955]), .B(n1141), .Z(ereg_next[956]) );
  AND U1192 ( .A(mul_pow), .B(n1142), .Z(n1141) );
  XOR U1193 ( .A(ein[956]), .B(ein[955]), .Z(n1142) );
  XOR U1194 ( .A(ein[954]), .B(n1143), .Z(ereg_next[955]) );
  AND U1195 ( .A(mul_pow), .B(n1144), .Z(n1143) );
  XOR U1196 ( .A(ein[955]), .B(ein[954]), .Z(n1144) );
  XOR U1197 ( .A(ein[953]), .B(n1145), .Z(ereg_next[954]) );
  AND U1198 ( .A(mul_pow), .B(n1146), .Z(n1145) );
  XOR U1199 ( .A(ein[954]), .B(ein[953]), .Z(n1146) );
  XOR U1200 ( .A(ein[952]), .B(n1147), .Z(ereg_next[953]) );
  AND U1201 ( .A(mul_pow), .B(n1148), .Z(n1147) );
  XOR U1202 ( .A(ein[953]), .B(ein[952]), .Z(n1148) );
  XOR U1203 ( .A(ein[951]), .B(n1149), .Z(ereg_next[952]) );
  AND U1204 ( .A(mul_pow), .B(n1150), .Z(n1149) );
  XOR U1205 ( .A(ein[952]), .B(ein[951]), .Z(n1150) );
  XOR U1206 ( .A(ein[950]), .B(n1151), .Z(ereg_next[951]) );
  AND U1207 ( .A(mul_pow), .B(n1152), .Z(n1151) );
  XOR U1208 ( .A(ein[951]), .B(ein[950]), .Z(n1152) );
  XOR U1209 ( .A(ein[949]), .B(n1153), .Z(ereg_next[950]) );
  AND U1210 ( .A(mul_pow), .B(n1154), .Z(n1153) );
  XOR U1211 ( .A(ein[950]), .B(ein[949]), .Z(n1154) );
  XOR U1212 ( .A(ein[93]), .B(n1155), .Z(ereg_next[94]) );
  AND U1213 ( .A(mul_pow), .B(n1156), .Z(n1155) );
  XOR U1214 ( .A(ein[94]), .B(ein[93]), .Z(n1156) );
  XOR U1215 ( .A(ein[948]), .B(n1157), .Z(ereg_next[949]) );
  AND U1216 ( .A(mul_pow), .B(n1158), .Z(n1157) );
  XOR U1217 ( .A(ein[949]), .B(ein[948]), .Z(n1158) );
  XOR U1218 ( .A(ein[947]), .B(n1159), .Z(ereg_next[948]) );
  AND U1219 ( .A(mul_pow), .B(n1160), .Z(n1159) );
  XOR U1220 ( .A(ein[948]), .B(ein[947]), .Z(n1160) );
  XOR U1221 ( .A(ein[946]), .B(n1161), .Z(ereg_next[947]) );
  AND U1222 ( .A(mul_pow), .B(n1162), .Z(n1161) );
  XOR U1223 ( .A(ein[947]), .B(ein[946]), .Z(n1162) );
  XOR U1224 ( .A(ein[945]), .B(n1163), .Z(ereg_next[946]) );
  AND U1225 ( .A(mul_pow), .B(n1164), .Z(n1163) );
  XOR U1226 ( .A(ein[946]), .B(ein[945]), .Z(n1164) );
  XOR U1227 ( .A(ein[944]), .B(n1165), .Z(ereg_next[945]) );
  AND U1228 ( .A(mul_pow), .B(n1166), .Z(n1165) );
  XOR U1229 ( .A(ein[945]), .B(ein[944]), .Z(n1166) );
  XOR U1230 ( .A(ein[943]), .B(n1167), .Z(ereg_next[944]) );
  AND U1231 ( .A(mul_pow), .B(n1168), .Z(n1167) );
  XOR U1232 ( .A(ein[944]), .B(ein[943]), .Z(n1168) );
  XOR U1233 ( .A(ein[942]), .B(n1169), .Z(ereg_next[943]) );
  AND U1234 ( .A(mul_pow), .B(n1170), .Z(n1169) );
  XOR U1235 ( .A(ein[943]), .B(ein[942]), .Z(n1170) );
  XOR U1236 ( .A(ein[941]), .B(n1171), .Z(ereg_next[942]) );
  AND U1237 ( .A(mul_pow), .B(n1172), .Z(n1171) );
  XOR U1238 ( .A(ein[942]), .B(ein[941]), .Z(n1172) );
  XOR U1239 ( .A(ein[940]), .B(n1173), .Z(ereg_next[941]) );
  AND U1240 ( .A(mul_pow), .B(n1174), .Z(n1173) );
  XOR U1241 ( .A(ein[941]), .B(ein[940]), .Z(n1174) );
  XOR U1242 ( .A(ein[939]), .B(n1175), .Z(ereg_next[940]) );
  AND U1243 ( .A(mul_pow), .B(n1176), .Z(n1175) );
  XOR U1244 ( .A(ein[940]), .B(ein[939]), .Z(n1176) );
  XOR U1245 ( .A(ein[92]), .B(n1177), .Z(ereg_next[93]) );
  AND U1246 ( .A(mul_pow), .B(n1178), .Z(n1177) );
  XOR U1247 ( .A(ein[93]), .B(ein[92]), .Z(n1178) );
  XOR U1248 ( .A(ein[938]), .B(n1179), .Z(ereg_next[939]) );
  AND U1249 ( .A(mul_pow), .B(n1180), .Z(n1179) );
  XOR U1250 ( .A(ein[939]), .B(ein[938]), .Z(n1180) );
  XOR U1251 ( .A(ein[937]), .B(n1181), .Z(ereg_next[938]) );
  AND U1252 ( .A(mul_pow), .B(n1182), .Z(n1181) );
  XOR U1253 ( .A(ein[938]), .B(ein[937]), .Z(n1182) );
  XOR U1254 ( .A(ein[936]), .B(n1183), .Z(ereg_next[937]) );
  AND U1255 ( .A(mul_pow), .B(n1184), .Z(n1183) );
  XOR U1256 ( .A(ein[937]), .B(ein[936]), .Z(n1184) );
  XOR U1257 ( .A(ein[935]), .B(n1185), .Z(ereg_next[936]) );
  AND U1258 ( .A(mul_pow), .B(n1186), .Z(n1185) );
  XOR U1259 ( .A(ein[936]), .B(ein[935]), .Z(n1186) );
  XOR U1260 ( .A(ein[934]), .B(n1187), .Z(ereg_next[935]) );
  AND U1261 ( .A(mul_pow), .B(n1188), .Z(n1187) );
  XOR U1262 ( .A(ein[935]), .B(ein[934]), .Z(n1188) );
  XOR U1263 ( .A(ein[933]), .B(n1189), .Z(ereg_next[934]) );
  AND U1264 ( .A(mul_pow), .B(n1190), .Z(n1189) );
  XOR U1265 ( .A(ein[934]), .B(ein[933]), .Z(n1190) );
  XOR U1266 ( .A(ein[932]), .B(n1191), .Z(ereg_next[933]) );
  AND U1267 ( .A(mul_pow), .B(n1192), .Z(n1191) );
  XOR U1268 ( .A(ein[933]), .B(ein[932]), .Z(n1192) );
  XOR U1269 ( .A(ein[931]), .B(n1193), .Z(ereg_next[932]) );
  AND U1270 ( .A(mul_pow), .B(n1194), .Z(n1193) );
  XOR U1271 ( .A(ein[932]), .B(ein[931]), .Z(n1194) );
  XOR U1272 ( .A(ein[930]), .B(n1195), .Z(ereg_next[931]) );
  AND U1273 ( .A(mul_pow), .B(n1196), .Z(n1195) );
  XOR U1274 ( .A(ein[931]), .B(ein[930]), .Z(n1196) );
  XOR U1275 ( .A(ein[929]), .B(n1197), .Z(ereg_next[930]) );
  AND U1276 ( .A(mul_pow), .B(n1198), .Z(n1197) );
  XOR U1277 ( .A(ein[930]), .B(ein[929]), .Z(n1198) );
  XOR U1278 ( .A(ein[91]), .B(n1199), .Z(ereg_next[92]) );
  AND U1279 ( .A(mul_pow), .B(n1200), .Z(n1199) );
  XOR U1280 ( .A(ein[92]), .B(ein[91]), .Z(n1200) );
  XOR U1281 ( .A(ein[928]), .B(n1201), .Z(ereg_next[929]) );
  AND U1282 ( .A(mul_pow), .B(n1202), .Z(n1201) );
  XOR U1283 ( .A(ein[929]), .B(ein[928]), .Z(n1202) );
  XOR U1284 ( .A(ein[927]), .B(n1203), .Z(ereg_next[928]) );
  AND U1285 ( .A(mul_pow), .B(n1204), .Z(n1203) );
  XOR U1286 ( .A(ein[928]), .B(ein[927]), .Z(n1204) );
  XOR U1287 ( .A(ein[926]), .B(n1205), .Z(ereg_next[927]) );
  AND U1288 ( .A(mul_pow), .B(n1206), .Z(n1205) );
  XOR U1289 ( .A(ein[927]), .B(ein[926]), .Z(n1206) );
  XOR U1290 ( .A(ein[925]), .B(n1207), .Z(ereg_next[926]) );
  AND U1291 ( .A(mul_pow), .B(n1208), .Z(n1207) );
  XOR U1292 ( .A(ein[926]), .B(ein[925]), .Z(n1208) );
  XOR U1293 ( .A(ein[924]), .B(n1209), .Z(ereg_next[925]) );
  AND U1294 ( .A(mul_pow), .B(n1210), .Z(n1209) );
  XOR U1295 ( .A(ein[925]), .B(ein[924]), .Z(n1210) );
  XOR U1296 ( .A(ein[923]), .B(n1211), .Z(ereg_next[924]) );
  AND U1297 ( .A(mul_pow), .B(n1212), .Z(n1211) );
  XOR U1298 ( .A(ein[924]), .B(ein[923]), .Z(n1212) );
  XOR U1299 ( .A(ein[922]), .B(n1213), .Z(ereg_next[923]) );
  AND U1300 ( .A(mul_pow), .B(n1214), .Z(n1213) );
  XOR U1301 ( .A(ein[923]), .B(ein[922]), .Z(n1214) );
  XOR U1302 ( .A(ein[921]), .B(n1215), .Z(ereg_next[922]) );
  AND U1303 ( .A(mul_pow), .B(n1216), .Z(n1215) );
  XOR U1304 ( .A(ein[922]), .B(ein[921]), .Z(n1216) );
  XOR U1305 ( .A(ein[920]), .B(n1217), .Z(ereg_next[921]) );
  AND U1306 ( .A(mul_pow), .B(n1218), .Z(n1217) );
  XOR U1307 ( .A(ein[921]), .B(ein[920]), .Z(n1218) );
  XOR U1308 ( .A(ein[919]), .B(n1219), .Z(ereg_next[920]) );
  AND U1309 ( .A(mul_pow), .B(n1220), .Z(n1219) );
  XOR U1310 ( .A(ein[920]), .B(ein[919]), .Z(n1220) );
  XOR U1311 ( .A(ein[90]), .B(n1221), .Z(ereg_next[91]) );
  AND U1312 ( .A(mul_pow), .B(n1222), .Z(n1221) );
  XOR U1313 ( .A(ein[91]), .B(ein[90]), .Z(n1222) );
  XOR U1314 ( .A(ein[918]), .B(n1223), .Z(ereg_next[919]) );
  AND U1315 ( .A(mul_pow), .B(n1224), .Z(n1223) );
  XOR U1316 ( .A(ein[919]), .B(ein[918]), .Z(n1224) );
  XOR U1317 ( .A(ein[917]), .B(n1225), .Z(ereg_next[918]) );
  AND U1318 ( .A(mul_pow), .B(n1226), .Z(n1225) );
  XOR U1319 ( .A(ein[918]), .B(ein[917]), .Z(n1226) );
  XOR U1320 ( .A(ein[916]), .B(n1227), .Z(ereg_next[917]) );
  AND U1321 ( .A(mul_pow), .B(n1228), .Z(n1227) );
  XOR U1322 ( .A(ein[917]), .B(ein[916]), .Z(n1228) );
  XOR U1323 ( .A(ein[915]), .B(n1229), .Z(ereg_next[916]) );
  AND U1324 ( .A(mul_pow), .B(n1230), .Z(n1229) );
  XOR U1325 ( .A(ein[916]), .B(ein[915]), .Z(n1230) );
  XOR U1326 ( .A(ein[914]), .B(n1231), .Z(ereg_next[915]) );
  AND U1327 ( .A(mul_pow), .B(n1232), .Z(n1231) );
  XOR U1328 ( .A(ein[915]), .B(ein[914]), .Z(n1232) );
  XOR U1329 ( .A(ein[913]), .B(n1233), .Z(ereg_next[914]) );
  AND U1330 ( .A(mul_pow), .B(n1234), .Z(n1233) );
  XOR U1331 ( .A(ein[914]), .B(ein[913]), .Z(n1234) );
  XOR U1332 ( .A(ein[912]), .B(n1235), .Z(ereg_next[913]) );
  AND U1333 ( .A(mul_pow), .B(n1236), .Z(n1235) );
  XOR U1334 ( .A(ein[913]), .B(ein[912]), .Z(n1236) );
  XOR U1335 ( .A(ein[911]), .B(n1237), .Z(ereg_next[912]) );
  AND U1336 ( .A(mul_pow), .B(n1238), .Z(n1237) );
  XOR U1337 ( .A(ein[912]), .B(ein[911]), .Z(n1238) );
  XOR U1338 ( .A(ein[910]), .B(n1239), .Z(ereg_next[911]) );
  AND U1339 ( .A(mul_pow), .B(n1240), .Z(n1239) );
  XOR U1340 ( .A(ein[911]), .B(ein[910]), .Z(n1240) );
  XOR U1341 ( .A(ein[909]), .B(n1241), .Z(ereg_next[910]) );
  AND U1342 ( .A(mul_pow), .B(n1242), .Z(n1241) );
  XOR U1343 ( .A(ein[910]), .B(ein[909]), .Z(n1242) );
  XOR U1344 ( .A(ein[89]), .B(n1243), .Z(ereg_next[90]) );
  AND U1345 ( .A(mul_pow), .B(n1244), .Z(n1243) );
  XOR U1346 ( .A(ein[90]), .B(ein[89]), .Z(n1244) );
  XOR U1347 ( .A(ein[908]), .B(n1245), .Z(ereg_next[909]) );
  AND U1348 ( .A(mul_pow), .B(n1246), .Z(n1245) );
  XOR U1349 ( .A(ein[909]), .B(ein[908]), .Z(n1246) );
  XOR U1350 ( .A(ein[907]), .B(n1247), .Z(ereg_next[908]) );
  AND U1351 ( .A(mul_pow), .B(n1248), .Z(n1247) );
  XOR U1352 ( .A(ein[908]), .B(ein[907]), .Z(n1248) );
  XOR U1353 ( .A(ein[906]), .B(n1249), .Z(ereg_next[907]) );
  AND U1354 ( .A(mul_pow), .B(n1250), .Z(n1249) );
  XOR U1355 ( .A(ein[907]), .B(ein[906]), .Z(n1250) );
  XOR U1356 ( .A(ein[905]), .B(n1251), .Z(ereg_next[906]) );
  AND U1357 ( .A(mul_pow), .B(n1252), .Z(n1251) );
  XOR U1358 ( .A(ein[906]), .B(ein[905]), .Z(n1252) );
  XOR U1359 ( .A(ein[904]), .B(n1253), .Z(ereg_next[905]) );
  AND U1360 ( .A(mul_pow), .B(n1254), .Z(n1253) );
  XOR U1361 ( .A(ein[905]), .B(ein[904]), .Z(n1254) );
  XOR U1362 ( .A(ein[903]), .B(n1255), .Z(ereg_next[904]) );
  AND U1363 ( .A(mul_pow), .B(n1256), .Z(n1255) );
  XOR U1364 ( .A(ein[904]), .B(ein[903]), .Z(n1256) );
  XOR U1365 ( .A(ein[902]), .B(n1257), .Z(ereg_next[903]) );
  AND U1366 ( .A(mul_pow), .B(n1258), .Z(n1257) );
  XOR U1367 ( .A(ein[903]), .B(ein[902]), .Z(n1258) );
  XOR U1368 ( .A(ein[901]), .B(n1259), .Z(ereg_next[902]) );
  AND U1369 ( .A(mul_pow), .B(n1260), .Z(n1259) );
  XOR U1370 ( .A(ein[902]), .B(ein[901]), .Z(n1260) );
  XOR U1371 ( .A(ein[900]), .B(n1261), .Z(ereg_next[901]) );
  AND U1372 ( .A(mul_pow), .B(n1262), .Z(n1261) );
  XOR U1373 ( .A(ein[901]), .B(ein[900]), .Z(n1262) );
  XOR U1374 ( .A(ein[899]), .B(n1263), .Z(ereg_next[900]) );
  AND U1375 ( .A(mul_pow), .B(n1264), .Z(n1263) );
  XOR U1376 ( .A(ein[900]), .B(ein[899]), .Z(n1264) );
  XOR U1377 ( .A(ein[7]), .B(n1265), .Z(ereg_next[8]) );
  AND U1378 ( .A(mul_pow), .B(n1266), .Z(n1265) );
  XOR U1379 ( .A(ein[8]), .B(ein[7]), .Z(n1266) );
  XOR U1380 ( .A(ein[88]), .B(n1267), .Z(ereg_next[89]) );
  AND U1381 ( .A(mul_pow), .B(n1268), .Z(n1267) );
  XOR U1382 ( .A(ein[89]), .B(ein[88]), .Z(n1268) );
  XOR U1383 ( .A(ein[898]), .B(n1269), .Z(ereg_next[899]) );
  AND U1384 ( .A(mul_pow), .B(n1270), .Z(n1269) );
  XOR U1385 ( .A(ein[899]), .B(ein[898]), .Z(n1270) );
  XOR U1386 ( .A(ein[897]), .B(n1271), .Z(ereg_next[898]) );
  AND U1387 ( .A(mul_pow), .B(n1272), .Z(n1271) );
  XOR U1388 ( .A(ein[898]), .B(ein[897]), .Z(n1272) );
  XOR U1389 ( .A(ein[896]), .B(n1273), .Z(ereg_next[897]) );
  AND U1390 ( .A(mul_pow), .B(n1274), .Z(n1273) );
  XOR U1391 ( .A(ein[897]), .B(ein[896]), .Z(n1274) );
  XOR U1392 ( .A(ein[895]), .B(n1275), .Z(ereg_next[896]) );
  AND U1393 ( .A(mul_pow), .B(n1276), .Z(n1275) );
  XOR U1394 ( .A(ein[896]), .B(ein[895]), .Z(n1276) );
  XOR U1395 ( .A(ein[894]), .B(n1277), .Z(ereg_next[895]) );
  AND U1396 ( .A(mul_pow), .B(n1278), .Z(n1277) );
  XOR U1397 ( .A(ein[895]), .B(ein[894]), .Z(n1278) );
  XOR U1398 ( .A(ein[893]), .B(n1279), .Z(ereg_next[894]) );
  AND U1399 ( .A(mul_pow), .B(n1280), .Z(n1279) );
  XOR U1400 ( .A(ein[894]), .B(ein[893]), .Z(n1280) );
  XOR U1401 ( .A(ein[892]), .B(n1281), .Z(ereg_next[893]) );
  AND U1402 ( .A(mul_pow), .B(n1282), .Z(n1281) );
  XOR U1403 ( .A(ein[893]), .B(ein[892]), .Z(n1282) );
  XOR U1404 ( .A(ein[891]), .B(n1283), .Z(ereg_next[892]) );
  AND U1405 ( .A(mul_pow), .B(n1284), .Z(n1283) );
  XOR U1406 ( .A(ein[892]), .B(ein[891]), .Z(n1284) );
  XOR U1407 ( .A(ein[890]), .B(n1285), .Z(ereg_next[891]) );
  AND U1408 ( .A(mul_pow), .B(n1286), .Z(n1285) );
  XOR U1409 ( .A(ein[891]), .B(ein[890]), .Z(n1286) );
  XOR U1410 ( .A(ein[889]), .B(n1287), .Z(ereg_next[890]) );
  AND U1411 ( .A(mul_pow), .B(n1288), .Z(n1287) );
  XOR U1412 ( .A(ein[890]), .B(ein[889]), .Z(n1288) );
  XOR U1413 ( .A(ein[87]), .B(n1289), .Z(ereg_next[88]) );
  AND U1414 ( .A(mul_pow), .B(n1290), .Z(n1289) );
  XOR U1415 ( .A(ein[88]), .B(ein[87]), .Z(n1290) );
  XOR U1416 ( .A(ein[888]), .B(n1291), .Z(ereg_next[889]) );
  AND U1417 ( .A(mul_pow), .B(n1292), .Z(n1291) );
  XOR U1418 ( .A(ein[889]), .B(ein[888]), .Z(n1292) );
  XOR U1419 ( .A(ein[887]), .B(n1293), .Z(ereg_next[888]) );
  AND U1420 ( .A(mul_pow), .B(n1294), .Z(n1293) );
  XOR U1421 ( .A(ein[888]), .B(ein[887]), .Z(n1294) );
  XOR U1422 ( .A(ein[886]), .B(n1295), .Z(ereg_next[887]) );
  AND U1423 ( .A(mul_pow), .B(n1296), .Z(n1295) );
  XOR U1424 ( .A(ein[887]), .B(ein[886]), .Z(n1296) );
  XOR U1425 ( .A(ein[885]), .B(n1297), .Z(ereg_next[886]) );
  AND U1426 ( .A(mul_pow), .B(n1298), .Z(n1297) );
  XOR U1427 ( .A(ein[886]), .B(ein[885]), .Z(n1298) );
  XOR U1428 ( .A(ein[884]), .B(n1299), .Z(ereg_next[885]) );
  AND U1429 ( .A(mul_pow), .B(n1300), .Z(n1299) );
  XOR U1430 ( .A(ein[885]), .B(ein[884]), .Z(n1300) );
  XOR U1431 ( .A(ein[883]), .B(n1301), .Z(ereg_next[884]) );
  AND U1432 ( .A(mul_pow), .B(n1302), .Z(n1301) );
  XOR U1433 ( .A(ein[884]), .B(ein[883]), .Z(n1302) );
  XOR U1434 ( .A(ein[882]), .B(n1303), .Z(ereg_next[883]) );
  AND U1435 ( .A(mul_pow), .B(n1304), .Z(n1303) );
  XOR U1436 ( .A(ein[883]), .B(ein[882]), .Z(n1304) );
  XOR U1437 ( .A(ein[881]), .B(n1305), .Z(ereg_next[882]) );
  AND U1438 ( .A(mul_pow), .B(n1306), .Z(n1305) );
  XOR U1439 ( .A(ein[882]), .B(ein[881]), .Z(n1306) );
  XOR U1440 ( .A(ein[880]), .B(n1307), .Z(ereg_next[881]) );
  AND U1441 ( .A(mul_pow), .B(n1308), .Z(n1307) );
  XOR U1442 ( .A(ein[881]), .B(ein[880]), .Z(n1308) );
  XOR U1443 ( .A(ein[879]), .B(n1309), .Z(ereg_next[880]) );
  AND U1444 ( .A(mul_pow), .B(n1310), .Z(n1309) );
  XOR U1445 ( .A(ein[880]), .B(ein[879]), .Z(n1310) );
  XOR U1446 ( .A(ein[86]), .B(n1311), .Z(ereg_next[87]) );
  AND U1447 ( .A(mul_pow), .B(n1312), .Z(n1311) );
  XOR U1448 ( .A(ein[87]), .B(ein[86]), .Z(n1312) );
  XOR U1449 ( .A(ein[878]), .B(n1313), .Z(ereg_next[879]) );
  AND U1450 ( .A(mul_pow), .B(n1314), .Z(n1313) );
  XOR U1451 ( .A(ein[879]), .B(ein[878]), .Z(n1314) );
  XOR U1452 ( .A(ein[877]), .B(n1315), .Z(ereg_next[878]) );
  AND U1453 ( .A(mul_pow), .B(n1316), .Z(n1315) );
  XOR U1454 ( .A(ein[878]), .B(ein[877]), .Z(n1316) );
  XOR U1455 ( .A(ein[876]), .B(n1317), .Z(ereg_next[877]) );
  AND U1456 ( .A(mul_pow), .B(n1318), .Z(n1317) );
  XOR U1457 ( .A(ein[877]), .B(ein[876]), .Z(n1318) );
  XOR U1458 ( .A(ein[875]), .B(n1319), .Z(ereg_next[876]) );
  AND U1459 ( .A(mul_pow), .B(n1320), .Z(n1319) );
  XOR U1460 ( .A(ein[876]), .B(ein[875]), .Z(n1320) );
  XOR U1461 ( .A(ein[874]), .B(n1321), .Z(ereg_next[875]) );
  AND U1462 ( .A(mul_pow), .B(n1322), .Z(n1321) );
  XOR U1463 ( .A(ein[875]), .B(ein[874]), .Z(n1322) );
  XOR U1464 ( .A(ein[873]), .B(n1323), .Z(ereg_next[874]) );
  AND U1465 ( .A(mul_pow), .B(n1324), .Z(n1323) );
  XOR U1466 ( .A(ein[874]), .B(ein[873]), .Z(n1324) );
  XOR U1467 ( .A(ein[872]), .B(n1325), .Z(ereg_next[873]) );
  AND U1468 ( .A(mul_pow), .B(n1326), .Z(n1325) );
  XOR U1469 ( .A(ein[873]), .B(ein[872]), .Z(n1326) );
  XOR U1470 ( .A(ein[871]), .B(n1327), .Z(ereg_next[872]) );
  AND U1471 ( .A(mul_pow), .B(n1328), .Z(n1327) );
  XOR U1472 ( .A(ein[872]), .B(ein[871]), .Z(n1328) );
  XOR U1473 ( .A(ein[870]), .B(n1329), .Z(ereg_next[871]) );
  AND U1474 ( .A(mul_pow), .B(n1330), .Z(n1329) );
  XOR U1475 ( .A(ein[871]), .B(ein[870]), .Z(n1330) );
  XOR U1476 ( .A(ein[869]), .B(n1331), .Z(ereg_next[870]) );
  AND U1477 ( .A(mul_pow), .B(n1332), .Z(n1331) );
  XOR U1478 ( .A(ein[870]), .B(ein[869]), .Z(n1332) );
  XOR U1479 ( .A(ein[85]), .B(n1333), .Z(ereg_next[86]) );
  AND U1480 ( .A(mul_pow), .B(n1334), .Z(n1333) );
  XOR U1481 ( .A(ein[86]), .B(ein[85]), .Z(n1334) );
  XOR U1482 ( .A(ein[868]), .B(n1335), .Z(ereg_next[869]) );
  AND U1483 ( .A(mul_pow), .B(n1336), .Z(n1335) );
  XOR U1484 ( .A(ein[869]), .B(ein[868]), .Z(n1336) );
  XOR U1485 ( .A(ein[867]), .B(n1337), .Z(ereg_next[868]) );
  AND U1486 ( .A(mul_pow), .B(n1338), .Z(n1337) );
  XOR U1487 ( .A(ein[868]), .B(ein[867]), .Z(n1338) );
  XOR U1488 ( .A(ein[866]), .B(n1339), .Z(ereg_next[867]) );
  AND U1489 ( .A(mul_pow), .B(n1340), .Z(n1339) );
  XOR U1490 ( .A(ein[867]), .B(ein[866]), .Z(n1340) );
  XOR U1491 ( .A(ein[865]), .B(n1341), .Z(ereg_next[866]) );
  AND U1492 ( .A(mul_pow), .B(n1342), .Z(n1341) );
  XOR U1493 ( .A(ein[866]), .B(ein[865]), .Z(n1342) );
  XOR U1494 ( .A(ein[864]), .B(n1343), .Z(ereg_next[865]) );
  AND U1495 ( .A(mul_pow), .B(n1344), .Z(n1343) );
  XOR U1496 ( .A(ein[865]), .B(ein[864]), .Z(n1344) );
  XOR U1497 ( .A(ein[863]), .B(n1345), .Z(ereg_next[864]) );
  AND U1498 ( .A(mul_pow), .B(n1346), .Z(n1345) );
  XOR U1499 ( .A(ein[864]), .B(ein[863]), .Z(n1346) );
  XOR U1500 ( .A(ein[862]), .B(n1347), .Z(ereg_next[863]) );
  AND U1501 ( .A(mul_pow), .B(n1348), .Z(n1347) );
  XOR U1502 ( .A(ein[863]), .B(ein[862]), .Z(n1348) );
  XOR U1503 ( .A(ein[861]), .B(n1349), .Z(ereg_next[862]) );
  AND U1504 ( .A(mul_pow), .B(n1350), .Z(n1349) );
  XOR U1505 ( .A(ein[862]), .B(ein[861]), .Z(n1350) );
  XOR U1506 ( .A(ein[860]), .B(n1351), .Z(ereg_next[861]) );
  AND U1507 ( .A(mul_pow), .B(n1352), .Z(n1351) );
  XOR U1508 ( .A(ein[861]), .B(ein[860]), .Z(n1352) );
  XOR U1509 ( .A(ein[859]), .B(n1353), .Z(ereg_next[860]) );
  AND U1510 ( .A(mul_pow), .B(n1354), .Z(n1353) );
  XOR U1511 ( .A(ein[860]), .B(ein[859]), .Z(n1354) );
  XOR U1512 ( .A(ein[84]), .B(n1355), .Z(ereg_next[85]) );
  AND U1513 ( .A(mul_pow), .B(n1356), .Z(n1355) );
  XOR U1514 ( .A(ein[85]), .B(ein[84]), .Z(n1356) );
  XOR U1515 ( .A(ein[858]), .B(n1357), .Z(ereg_next[859]) );
  AND U1516 ( .A(mul_pow), .B(n1358), .Z(n1357) );
  XOR U1517 ( .A(ein[859]), .B(ein[858]), .Z(n1358) );
  XOR U1518 ( .A(ein[857]), .B(n1359), .Z(ereg_next[858]) );
  AND U1519 ( .A(mul_pow), .B(n1360), .Z(n1359) );
  XOR U1520 ( .A(ein[858]), .B(ein[857]), .Z(n1360) );
  XOR U1521 ( .A(ein[856]), .B(n1361), .Z(ereg_next[857]) );
  AND U1522 ( .A(mul_pow), .B(n1362), .Z(n1361) );
  XOR U1523 ( .A(ein[857]), .B(ein[856]), .Z(n1362) );
  XOR U1524 ( .A(ein[855]), .B(n1363), .Z(ereg_next[856]) );
  AND U1525 ( .A(mul_pow), .B(n1364), .Z(n1363) );
  XOR U1526 ( .A(ein[856]), .B(ein[855]), .Z(n1364) );
  XOR U1527 ( .A(ein[854]), .B(n1365), .Z(ereg_next[855]) );
  AND U1528 ( .A(mul_pow), .B(n1366), .Z(n1365) );
  XOR U1529 ( .A(ein[855]), .B(ein[854]), .Z(n1366) );
  XOR U1530 ( .A(ein[853]), .B(n1367), .Z(ereg_next[854]) );
  AND U1531 ( .A(mul_pow), .B(n1368), .Z(n1367) );
  XOR U1532 ( .A(ein[854]), .B(ein[853]), .Z(n1368) );
  XOR U1533 ( .A(ein[852]), .B(n1369), .Z(ereg_next[853]) );
  AND U1534 ( .A(mul_pow), .B(n1370), .Z(n1369) );
  XOR U1535 ( .A(ein[853]), .B(ein[852]), .Z(n1370) );
  XOR U1536 ( .A(ein[851]), .B(n1371), .Z(ereg_next[852]) );
  AND U1537 ( .A(mul_pow), .B(n1372), .Z(n1371) );
  XOR U1538 ( .A(ein[852]), .B(ein[851]), .Z(n1372) );
  XOR U1539 ( .A(ein[850]), .B(n1373), .Z(ereg_next[851]) );
  AND U1540 ( .A(mul_pow), .B(n1374), .Z(n1373) );
  XOR U1541 ( .A(ein[851]), .B(ein[850]), .Z(n1374) );
  XOR U1542 ( .A(ein[849]), .B(n1375), .Z(ereg_next[850]) );
  AND U1543 ( .A(mul_pow), .B(n1376), .Z(n1375) );
  XOR U1544 ( .A(ein[850]), .B(ein[849]), .Z(n1376) );
  XOR U1545 ( .A(ein[83]), .B(n1377), .Z(ereg_next[84]) );
  AND U1546 ( .A(mul_pow), .B(n1378), .Z(n1377) );
  XOR U1547 ( .A(ein[84]), .B(ein[83]), .Z(n1378) );
  XOR U1548 ( .A(ein[848]), .B(n1379), .Z(ereg_next[849]) );
  AND U1549 ( .A(mul_pow), .B(n1380), .Z(n1379) );
  XOR U1550 ( .A(ein[849]), .B(ein[848]), .Z(n1380) );
  XOR U1551 ( .A(ein[847]), .B(n1381), .Z(ereg_next[848]) );
  AND U1552 ( .A(mul_pow), .B(n1382), .Z(n1381) );
  XOR U1553 ( .A(ein[848]), .B(ein[847]), .Z(n1382) );
  XOR U1554 ( .A(ein[846]), .B(n1383), .Z(ereg_next[847]) );
  AND U1555 ( .A(mul_pow), .B(n1384), .Z(n1383) );
  XOR U1556 ( .A(ein[847]), .B(ein[846]), .Z(n1384) );
  XOR U1557 ( .A(ein[845]), .B(n1385), .Z(ereg_next[846]) );
  AND U1558 ( .A(mul_pow), .B(n1386), .Z(n1385) );
  XOR U1559 ( .A(ein[846]), .B(ein[845]), .Z(n1386) );
  XOR U1560 ( .A(ein[844]), .B(n1387), .Z(ereg_next[845]) );
  AND U1561 ( .A(mul_pow), .B(n1388), .Z(n1387) );
  XOR U1562 ( .A(ein[845]), .B(ein[844]), .Z(n1388) );
  XOR U1563 ( .A(ein[843]), .B(n1389), .Z(ereg_next[844]) );
  AND U1564 ( .A(mul_pow), .B(n1390), .Z(n1389) );
  XOR U1565 ( .A(ein[844]), .B(ein[843]), .Z(n1390) );
  XOR U1566 ( .A(ein[842]), .B(n1391), .Z(ereg_next[843]) );
  AND U1567 ( .A(mul_pow), .B(n1392), .Z(n1391) );
  XOR U1568 ( .A(ein[843]), .B(ein[842]), .Z(n1392) );
  XOR U1569 ( .A(ein[841]), .B(n1393), .Z(ereg_next[842]) );
  AND U1570 ( .A(mul_pow), .B(n1394), .Z(n1393) );
  XOR U1571 ( .A(ein[842]), .B(ein[841]), .Z(n1394) );
  XOR U1572 ( .A(ein[840]), .B(n1395), .Z(ereg_next[841]) );
  AND U1573 ( .A(mul_pow), .B(n1396), .Z(n1395) );
  XOR U1574 ( .A(ein[841]), .B(ein[840]), .Z(n1396) );
  XOR U1575 ( .A(ein[839]), .B(n1397), .Z(ereg_next[840]) );
  AND U1576 ( .A(mul_pow), .B(n1398), .Z(n1397) );
  XOR U1577 ( .A(ein[840]), .B(ein[839]), .Z(n1398) );
  XOR U1578 ( .A(ein[82]), .B(n1399), .Z(ereg_next[83]) );
  AND U1579 ( .A(mul_pow), .B(n1400), .Z(n1399) );
  XOR U1580 ( .A(ein[83]), .B(ein[82]), .Z(n1400) );
  XOR U1581 ( .A(ein[838]), .B(n1401), .Z(ereg_next[839]) );
  AND U1582 ( .A(mul_pow), .B(n1402), .Z(n1401) );
  XOR U1583 ( .A(ein[839]), .B(ein[838]), .Z(n1402) );
  XOR U1584 ( .A(ein[837]), .B(n1403), .Z(ereg_next[838]) );
  AND U1585 ( .A(mul_pow), .B(n1404), .Z(n1403) );
  XOR U1586 ( .A(ein[838]), .B(ein[837]), .Z(n1404) );
  XOR U1587 ( .A(ein[836]), .B(n1405), .Z(ereg_next[837]) );
  AND U1588 ( .A(mul_pow), .B(n1406), .Z(n1405) );
  XOR U1589 ( .A(ein[837]), .B(ein[836]), .Z(n1406) );
  XOR U1590 ( .A(ein[835]), .B(n1407), .Z(ereg_next[836]) );
  AND U1591 ( .A(mul_pow), .B(n1408), .Z(n1407) );
  XOR U1592 ( .A(ein[836]), .B(ein[835]), .Z(n1408) );
  XOR U1593 ( .A(ein[834]), .B(n1409), .Z(ereg_next[835]) );
  AND U1594 ( .A(mul_pow), .B(n1410), .Z(n1409) );
  XOR U1595 ( .A(ein[835]), .B(ein[834]), .Z(n1410) );
  XOR U1596 ( .A(ein[833]), .B(n1411), .Z(ereg_next[834]) );
  AND U1597 ( .A(mul_pow), .B(n1412), .Z(n1411) );
  XOR U1598 ( .A(ein[834]), .B(ein[833]), .Z(n1412) );
  XOR U1599 ( .A(ein[832]), .B(n1413), .Z(ereg_next[833]) );
  AND U1600 ( .A(mul_pow), .B(n1414), .Z(n1413) );
  XOR U1601 ( .A(ein[833]), .B(ein[832]), .Z(n1414) );
  XOR U1602 ( .A(ein[831]), .B(n1415), .Z(ereg_next[832]) );
  AND U1603 ( .A(mul_pow), .B(n1416), .Z(n1415) );
  XOR U1604 ( .A(ein[832]), .B(ein[831]), .Z(n1416) );
  XOR U1605 ( .A(ein[830]), .B(n1417), .Z(ereg_next[831]) );
  AND U1606 ( .A(mul_pow), .B(n1418), .Z(n1417) );
  XOR U1607 ( .A(ein[831]), .B(ein[830]), .Z(n1418) );
  XOR U1608 ( .A(ein[829]), .B(n1419), .Z(ereg_next[830]) );
  AND U1609 ( .A(mul_pow), .B(n1420), .Z(n1419) );
  XOR U1610 ( .A(ein[830]), .B(ein[829]), .Z(n1420) );
  XOR U1611 ( .A(ein[81]), .B(n1421), .Z(ereg_next[82]) );
  AND U1612 ( .A(mul_pow), .B(n1422), .Z(n1421) );
  XOR U1613 ( .A(ein[82]), .B(ein[81]), .Z(n1422) );
  XOR U1614 ( .A(ein[828]), .B(n1423), .Z(ereg_next[829]) );
  AND U1615 ( .A(mul_pow), .B(n1424), .Z(n1423) );
  XOR U1616 ( .A(ein[829]), .B(ein[828]), .Z(n1424) );
  XOR U1617 ( .A(ein[827]), .B(n1425), .Z(ereg_next[828]) );
  AND U1618 ( .A(mul_pow), .B(n1426), .Z(n1425) );
  XOR U1619 ( .A(ein[828]), .B(ein[827]), .Z(n1426) );
  XOR U1620 ( .A(ein[826]), .B(n1427), .Z(ereg_next[827]) );
  AND U1621 ( .A(mul_pow), .B(n1428), .Z(n1427) );
  XOR U1622 ( .A(ein[827]), .B(ein[826]), .Z(n1428) );
  XOR U1623 ( .A(ein[825]), .B(n1429), .Z(ereg_next[826]) );
  AND U1624 ( .A(mul_pow), .B(n1430), .Z(n1429) );
  XOR U1625 ( .A(ein[826]), .B(ein[825]), .Z(n1430) );
  XOR U1626 ( .A(ein[824]), .B(n1431), .Z(ereg_next[825]) );
  AND U1627 ( .A(mul_pow), .B(n1432), .Z(n1431) );
  XOR U1628 ( .A(ein[825]), .B(ein[824]), .Z(n1432) );
  XOR U1629 ( .A(ein[823]), .B(n1433), .Z(ereg_next[824]) );
  AND U1630 ( .A(mul_pow), .B(n1434), .Z(n1433) );
  XOR U1631 ( .A(ein[824]), .B(ein[823]), .Z(n1434) );
  XOR U1632 ( .A(ein[822]), .B(n1435), .Z(ereg_next[823]) );
  AND U1633 ( .A(mul_pow), .B(n1436), .Z(n1435) );
  XOR U1634 ( .A(ein[823]), .B(ein[822]), .Z(n1436) );
  XOR U1635 ( .A(ein[821]), .B(n1437), .Z(ereg_next[822]) );
  AND U1636 ( .A(mul_pow), .B(n1438), .Z(n1437) );
  XOR U1637 ( .A(ein[822]), .B(ein[821]), .Z(n1438) );
  XOR U1638 ( .A(ein[820]), .B(n1439), .Z(ereg_next[821]) );
  AND U1639 ( .A(mul_pow), .B(n1440), .Z(n1439) );
  XOR U1640 ( .A(ein[821]), .B(ein[820]), .Z(n1440) );
  XOR U1641 ( .A(ein[819]), .B(n1441), .Z(ereg_next[820]) );
  AND U1642 ( .A(mul_pow), .B(n1442), .Z(n1441) );
  XOR U1643 ( .A(ein[820]), .B(ein[819]), .Z(n1442) );
  XOR U1644 ( .A(ein[80]), .B(n1443), .Z(ereg_next[81]) );
  AND U1645 ( .A(mul_pow), .B(n1444), .Z(n1443) );
  XOR U1646 ( .A(ein[81]), .B(ein[80]), .Z(n1444) );
  XOR U1647 ( .A(ein[818]), .B(n1445), .Z(ereg_next[819]) );
  AND U1648 ( .A(mul_pow), .B(n1446), .Z(n1445) );
  XOR U1649 ( .A(ein[819]), .B(ein[818]), .Z(n1446) );
  XOR U1650 ( .A(ein[817]), .B(n1447), .Z(ereg_next[818]) );
  AND U1651 ( .A(mul_pow), .B(n1448), .Z(n1447) );
  XOR U1652 ( .A(ein[818]), .B(ein[817]), .Z(n1448) );
  XOR U1653 ( .A(ein[816]), .B(n1449), .Z(ereg_next[817]) );
  AND U1654 ( .A(mul_pow), .B(n1450), .Z(n1449) );
  XOR U1655 ( .A(ein[817]), .B(ein[816]), .Z(n1450) );
  XOR U1656 ( .A(ein[815]), .B(n1451), .Z(ereg_next[816]) );
  AND U1657 ( .A(mul_pow), .B(n1452), .Z(n1451) );
  XOR U1658 ( .A(ein[816]), .B(ein[815]), .Z(n1452) );
  XOR U1659 ( .A(ein[814]), .B(n1453), .Z(ereg_next[815]) );
  AND U1660 ( .A(mul_pow), .B(n1454), .Z(n1453) );
  XOR U1661 ( .A(ein[815]), .B(ein[814]), .Z(n1454) );
  XOR U1662 ( .A(ein[813]), .B(n1455), .Z(ereg_next[814]) );
  AND U1663 ( .A(mul_pow), .B(n1456), .Z(n1455) );
  XOR U1664 ( .A(ein[814]), .B(ein[813]), .Z(n1456) );
  XOR U1665 ( .A(ein[812]), .B(n1457), .Z(ereg_next[813]) );
  AND U1666 ( .A(mul_pow), .B(n1458), .Z(n1457) );
  XOR U1667 ( .A(ein[813]), .B(ein[812]), .Z(n1458) );
  XOR U1668 ( .A(ein[811]), .B(n1459), .Z(ereg_next[812]) );
  AND U1669 ( .A(mul_pow), .B(n1460), .Z(n1459) );
  XOR U1670 ( .A(ein[812]), .B(ein[811]), .Z(n1460) );
  XOR U1671 ( .A(ein[810]), .B(n1461), .Z(ereg_next[811]) );
  AND U1672 ( .A(mul_pow), .B(n1462), .Z(n1461) );
  XOR U1673 ( .A(ein[811]), .B(ein[810]), .Z(n1462) );
  XOR U1674 ( .A(ein[809]), .B(n1463), .Z(ereg_next[810]) );
  AND U1675 ( .A(mul_pow), .B(n1464), .Z(n1463) );
  XOR U1676 ( .A(ein[810]), .B(ein[809]), .Z(n1464) );
  XOR U1677 ( .A(ein[79]), .B(n1465), .Z(ereg_next[80]) );
  AND U1678 ( .A(mul_pow), .B(n1466), .Z(n1465) );
  XOR U1679 ( .A(ein[80]), .B(ein[79]), .Z(n1466) );
  XOR U1680 ( .A(ein[808]), .B(n1467), .Z(ereg_next[809]) );
  AND U1681 ( .A(mul_pow), .B(n1468), .Z(n1467) );
  XOR U1682 ( .A(ein[809]), .B(ein[808]), .Z(n1468) );
  XOR U1683 ( .A(ein[807]), .B(n1469), .Z(ereg_next[808]) );
  AND U1684 ( .A(mul_pow), .B(n1470), .Z(n1469) );
  XOR U1685 ( .A(ein[808]), .B(ein[807]), .Z(n1470) );
  XOR U1686 ( .A(ein[806]), .B(n1471), .Z(ereg_next[807]) );
  AND U1687 ( .A(mul_pow), .B(n1472), .Z(n1471) );
  XOR U1688 ( .A(ein[807]), .B(ein[806]), .Z(n1472) );
  XOR U1689 ( .A(ein[805]), .B(n1473), .Z(ereg_next[806]) );
  AND U1690 ( .A(mul_pow), .B(n1474), .Z(n1473) );
  XOR U1691 ( .A(ein[806]), .B(ein[805]), .Z(n1474) );
  XOR U1692 ( .A(ein[804]), .B(n1475), .Z(ereg_next[805]) );
  AND U1693 ( .A(mul_pow), .B(n1476), .Z(n1475) );
  XOR U1694 ( .A(ein[805]), .B(ein[804]), .Z(n1476) );
  XOR U1695 ( .A(ein[803]), .B(n1477), .Z(ereg_next[804]) );
  AND U1696 ( .A(mul_pow), .B(n1478), .Z(n1477) );
  XOR U1697 ( .A(ein[804]), .B(ein[803]), .Z(n1478) );
  XOR U1698 ( .A(ein[802]), .B(n1479), .Z(ereg_next[803]) );
  AND U1699 ( .A(mul_pow), .B(n1480), .Z(n1479) );
  XOR U1700 ( .A(ein[803]), .B(ein[802]), .Z(n1480) );
  XOR U1701 ( .A(ein[801]), .B(n1481), .Z(ereg_next[802]) );
  AND U1702 ( .A(mul_pow), .B(n1482), .Z(n1481) );
  XOR U1703 ( .A(ein[802]), .B(ein[801]), .Z(n1482) );
  XOR U1704 ( .A(ein[800]), .B(n1483), .Z(ereg_next[801]) );
  AND U1705 ( .A(mul_pow), .B(n1484), .Z(n1483) );
  XOR U1706 ( .A(ein[801]), .B(ein[800]), .Z(n1484) );
  XOR U1707 ( .A(ein[799]), .B(n1485), .Z(ereg_next[800]) );
  AND U1708 ( .A(mul_pow), .B(n1486), .Z(n1485) );
  XOR U1709 ( .A(ein[800]), .B(ein[799]), .Z(n1486) );
  XOR U1710 ( .A(ein[6]), .B(n1487), .Z(ereg_next[7]) );
  AND U1711 ( .A(mul_pow), .B(n1488), .Z(n1487) );
  XOR U1712 ( .A(ein[7]), .B(ein[6]), .Z(n1488) );
  XOR U1713 ( .A(ein[78]), .B(n1489), .Z(ereg_next[79]) );
  AND U1714 ( .A(mul_pow), .B(n1490), .Z(n1489) );
  XOR U1715 ( .A(ein[79]), .B(ein[78]), .Z(n1490) );
  XOR U1716 ( .A(ein[798]), .B(n1491), .Z(ereg_next[799]) );
  AND U1717 ( .A(mul_pow), .B(n1492), .Z(n1491) );
  XOR U1718 ( .A(ein[799]), .B(ein[798]), .Z(n1492) );
  XOR U1719 ( .A(ein[797]), .B(n1493), .Z(ereg_next[798]) );
  AND U1720 ( .A(mul_pow), .B(n1494), .Z(n1493) );
  XOR U1721 ( .A(ein[798]), .B(ein[797]), .Z(n1494) );
  XOR U1722 ( .A(ein[796]), .B(n1495), .Z(ereg_next[797]) );
  AND U1723 ( .A(mul_pow), .B(n1496), .Z(n1495) );
  XOR U1724 ( .A(ein[797]), .B(ein[796]), .Z(n1496) );
  XOR U1725 ( .A(ein[795]), .B(n1497), .Z(ereg_next[796]) );
  AND U1726 ( .A(mul_pow), .B(n1498), .Z(n1497) );
  XOR U1727 ( .A(ein[796]), .B(ein[795]), .Z(n1498) );
  XOR U1728 ( .A(ein[794]), .B(n1499), .Z(ereg_next[795]) );
  AND U1729 ( .A(mul_pow), .B(n1500), .Z(n1499) );
  XOR U1730 ( .A(ein[795]), .B(ein[794]), .Z(n1500) );
  XOR U1731 ( .A(ein[793]), .B(n1501), .Z(ereg_next[794]) );
  AND U1732 ( .A(mul_pow), .B(n1502), .Z(n1501) );
  XOR U1733 ( .A(ein[794]), .B(ein[793]), .Z(n1502) );
  XOR U1734 ( .A(ein[792]), .B(n1503), .Z(ereg_next[793]) );
  AND U1735 ( .A(mul_pow), .B(n1504), .Z(n1503) );
  XOR U1736 ( .A(ein[793]), .B(ein[792]), .Z(n1504) );
  XOR U1737 ( .A(ein[791]), .B(n1505), .Z(ereg_next[792]) );
  AND U1738 ( .A(mul_pow), .B(n1506), .Z(n1505) );
  XOR U1739 ( .A(ein[792]), .B(ein[791]), .Z(n1506) );
  XOR U1740 ( .A(ein[790]), .B(n1507), .Z(ereg_next[791]) );
  AND U1741 ( .A(mul_pow), .B(n1508), .Z(n1507) );
  XOR U1742 ( .A(ein[791]), .B(ein[790]), .Z(n1508) );
  XOR U1743 ( .A(ein[789]), .B(n1509), .Z(ereg_next[790]) );
  AND U1744 ( .A(mul_pow), .B(n1510), .Z(n1509) );
  XOR U1745 ( .A(ein[790]), .B(ein[789]), .Z(n1510) );
  XOR U1746 ( .A(ein[77]), .B(n1511), .Z(ereg_next[78]) );
  AND U1747 ( .A(mul_pow), .B(n1512), .Z(n1511) );
  XOR U1748 ( .A(ein[78]), .B(ein[77]), .Z(n1512) );
  XOR U1749 ( .A(ein[788]), .B(n1513), .Z(ereg_next[789]) );
  AND U1750 ( .A(mul_pow), .B(n1514), .Z(n1513) );
  XOR U1751 ( .A(ein[789]), .B(ein[788]), .Z(n1514) );
  XOR U1752 ( .A(ein[787]), .B(n1515), .Z(ereg_next[788]) );
  AND U1753 ( .A(mul_pow), .B(n1516), .Z(n1515) );
  XOR U1754 ( .A(ein[788]), .B(ein[787]), .Z(n1516) );
  XOR U1755 ( .A(ein[786]), .B(n1517), .Z(ereg_next[787]) );
  AND U1756 ( .A(mul_pow), .B(n1518), .Z(n1517) );
  XOR U1757 ( .A(ein[787]), .B(ein[786]), .Z(n1518) );
  XOR U1758 ( .A(ein[785]), .B(n1519), .Z(ereg_next[786]) );
  AND U1759 ( .A(mul_pow), .B(n1520), .Z(n1519) );
  XOR U1760 ( .A(ein[786]), .B(ein[785]), .Z(n1520) );
  XOR U1761 ( .A(ein[784]), .B(n1521), .Z(ereg_next[785]) );
  AND U1762 ( .A(mul_pow), .B(n1522), .Z(n1521) );
  XOR U1763 ( .A(ein[785]), .B(ein[784]), .Z(n1522) );
  XOR U1764 ( .A(ein[783]), .B(n1523), .Z(ereg_next[784]) );
  AND U1765 ( .A(mul_pow), .B(n1524), .Z(n1523) );
  XOR U1766 ( .A(ein[784]), .B(ein[783]), .Z(n1524) );
  XOR U1767 ( .A(ein[782]), .B(n1525), .Z(ereg_next[783]) );
  AND U1768 ( .A(mul_pow), .B(n1526), .Z(n1525) );
  XOR U1769 ( .A(ein[783]), .B(ein[782]), .Z(n1526) );
  XOR U1770 ( .A(ein[781]), .B(n1527), .Z(ereg_next[782]) );
  AND U1771 ( .A(mul_pow), .B(n1528), .Z(n1527) );
  XOR U1772 ( .A(ein[782]), .B(ein[781]), .Z(n1528) );
  XOR U1773 ( .A(ein[780]), .B(n1529), .Z(ereg_next[781]) );
  AND U1774 ( .A(mul_pow), .B(n1530), .Z(n1529) );
  XOR U1775 ( .A(ein[781]), .B(ein[780]), .Z(n1530) );
  XOR U1776 ( .A(ein[779]), .B(n1531), .Z(ereg_next[780]) );
  AND U1777 ( .A(mul_pow), .B(n1532), .Z(n1531) );
  XOR U1778 ( .A(ein[780]), .B(ein[779]), .Z(n1532) );
  XOR U1779 ( .A(ein[76]), .B(n1533), .Z(ereg_next[77]) );
  AND U1780 ( .A(mul_pow), .B(n1534), .Z(n1533) );
  XOR U1781 ( .A(ein[77]), .B(ein[76]), .Z(n1534) );
  XOR U1782 ( .A(ein[778]), .B(n1535), .Z(ereg_next[779]) );
  AND U1783 ( .A(mul_pow), .B(n1536), .Z(n1535) );
  XOR U1784 ( .A(ein[779]), .B(ein[778]), .Z(n1536) );
  XOR U1785 ( .A(ein[777]), .B(n1537), .Z(ereg_next[778]) );
  AND U1786 ( .A(mul_pow), .B(n1538), .Z(n1537) );
  XOR U1787 ( .A(ein[778]), .B(ein[777]), .Z(n1538) );
  XOR U1788 ( .A(ein[776]), .B(n1539), .Z(ereg_next[777]) );
  AND U1789 ( .A(mul_pow), .B(n1540), .Z(n1539) );
  XOR U1790 ( .A(ein[777]), .B(ein[776]), .Z(n1540) );
  XOR U1791 ( .A(ein[775]), .B(n1541), .Z(ereg_next[776]) );
  AND U1792 ( .A(mul_pow), .B(n1542), .Z(n1541) );
  XOR U1793 ( .A(ein[776]), .B(ein[775]), .Z(n1542) );
  XOR U1794 ( .A(ein[774]), .B(n1543), .Z(ereg_next[775]) );
  AND U1795 ( .A(mul_pow), .B(n1544), .Z(n1543) );
  XOR U1796 ( .A(ein[775]), .B(ein[774]), .Z(n1544) );
  XOR U1797 ( .A(ein[773]), .B(n1545), .Z(ereg_next[774]) );
  AND U1798 ( .A(mul_pow), .B(n1546), .Z(n1545) );
  XOR U1799 ( .A(ein[774]), .B(ein[773]), .Z(n1546) );
  XOR U1800 ( .A(ein[772]), .B(n1547), .Z(ereg_next[773]) );
  AND U1801 ( .A(mul_pow), .B(n1548), .Z(n1547) );
  XOR U1802 ( .A(ein[773]), .B(ein[772]), .Z(n1548) );
  XOR U1803 ( .A(ein[771]), .B(n1549), .Z(ereg_next[772]) );
  AND U1804 ( .A(mul_pow), .B(n1550), .Z(n1549) );
  XOR U1805 ( .A(ein[772]), .B(ein[771]), .Z(n1550) );
  XOR U1806 ( .A(ein[770]), .B(n1551), .Z(ereg_next[771]) );
  AND U1807 ( .A(mul_pow), .B(n1552), .Z(n1551) );
  XOR U1808 ( .A(ein[771]), .B(ein[770]), .Z(n1552) );
  XOR U1809 ( .A(ein[769]), .B(n1553), .Z(ereg_next[770]) );
  AND U1810 ( .A(mul_pow), .B(n1554), .Z(n1553) );
  XOR U1811 ( .A(ein[770]), .B(ein[769]), .Z(n1554) );
  XOR U1812 ( .A(ein[75]), .B(n1555), .Z(ereg_next[76]) );
  AND U1813 ( .A(mul_pow), .B(n1556), .Z(n1555) );
  XOR U1814 ( .A(ein[76]), .B(ein[75]), .Z(n1556) );
  XOR U1815 ( .A(ein[768]), .B(n1557), .Z(ereg_next[769]) );
  AND U1816 ( .A(mul_pow), .B(n1558), .Z(n1557) );
  XOR U1817 ( .A(ein[769]), .B(ein[768]), .Z(n1558) );
  XOR U1818 ( .A(ein[767]), .B(n1559), .Z(ereg_next[768]) );
  AND U1819 ( .A(mul_pow), .B(n1560), .Z(n1559) );
  XOR U1820 ( .A(ein[768]), .B(ein[767]), .Z(n1560) );
  XOR U1821 ( .A(ein[766]), .B(n1561), .Z(ereg_next[767]) );
  AND U1822 ( .A(mul_pow), .B(n1562), .Z(n1561) );
  XOR U1823 ( .A(ein[767]), .B(ein[766]), .Z(n1562) );
  XOR U1824 ( .A(ein[765]), .B(n1563), .Z(ereg_next[766]) );
  AND U1825 ( .A(mul_pow), .B(n1564), .Z(n1563) );
  XOR U1826 ( .A(ein[766]), .B(ein[765]), .Z(n1564) );
  XOR U1827 ( .A(ein[764]), .B(n1565), .Z(ereg_next[765]) );
  AND U1828 ( .A(mul_pow), .B(n1566), .Z(n1565) );
  XOR U1829 ( .A(ein[765]), .B(ein[764]), .Z(n1566) );
  XOR U1830 ( .A(ein[763]), .B(n1567), .Z(ereg_next[764]) );
  AND U1831 ( .A(mul_pow), .B(n1568), .Z(n1567) );
  XOR U1832 ( .A(ein[764]), .B(ein[763]), .Z(n1568) );
  XOR U1833 ( .A(ein[762]), .B(n1569), .Z(ereg_next[763]) );
  AND U1834 ( .A(mul_pow), .B(n1570), .Z(n1569) );
  XOR U1835 ( .A(ein[763]), .B(ein[762]), .Z(n1570) );
  XOR U1836 ( .A(ein[761]), .B(n1571), .Z(ereg_next[762]) );
  AND U1837 ( .A(mul_pow), .B(n1572), .Z(n1571) );
  XOR U1838 ( .A(ein[762]), .B(ein[761]), .Z(n1572) );
  XOR U1839 ( .A(ein[760]), .B(n1573), .Z(ereg_next[761]) );
  AND U1840 ( .A(mul_pow), .B(n1574), .Z(n1573) );
  XOR U1841 ( .A(ein[761]), .B(ein[760]), .Z(n1574) );
  XOR U1842 ( .A(ein[759]), .B(n1575), .Z(ereg_next[760]) );
  AND U1843 ( .A(mul_pow), .B(n1576), .Z(n1575) );
  XOR U1844 ( .A(ein[760]), .B(ein[759]), .Z(n1576) );
  XOR U1845 ( .A(ein[74]), .B(n1577), .Z(ereg_next[75]) );
  AND U1846 ( .A(mul_pow), .B(n1578), .Z(n1577) );
  XOR U1847 ( .A(ein[75]), .B(ein[74]), .Z(n1578) );
  XOR U1848 ( .A(ein[758]), .B(n1579), .Z(ereg_next[759]) );
  AND U1849 ( .A(mul_pow), .B(n1580), .Z(n1579) );
  XOR U1850 ( .A(ein[759]), .B(ein[758]), .Z(n1580) );
  XOR U1851 ( .A(ein[757]), .B(n1581), .Z(ereg_next[758]) );
  AND U1852 ( .A(mul_pow), .B(n1582), .Z(n1581) );
  XOR U1853 ( .A(ein[758]), .B(ein[757]), .Z(n1582) );
  XOR U1854 ( .A(ein[756]), .B(n1583), .Z(ereg_next[757]) );
  AND U1855 ( .A(mul_pow), .B(n1584), .Z(n1583) );
  XOR U1856 ( .A(ein[757]), .B(ein[756]), .Z(n1584) );
  XOR U1857 ( .A(ein[755]), .B(n1585), .Z(ereg_next[756]) );
  AND U1858 ( .A(mul_pow), .B(n1586), .Z(n1585) );
  XOR U1859 ( .A(ein[756]), .B(ein[755]), .Z(n1586) );
  XOR U1860 ( .A(ein[754]), .B(n1587), .Z(ereg_next[755]) );
  AND U1861 ( .A(mul_pow), .B(n1588), .Z(n1587) );
  XOR U1862 ( .A(ein[755]), .B(ein[754]), .Z(n1588) );
  XOR U1863 ( .A(ein[753]), .B(n1589), .Z(ereg_next[754]) );
  AND U1864 ( .A(mul_pow), .B(n1590), .Z(n1589) );
  XOR U1865 ( .A(ein[754]), .B(ein[753]), .Z(n1590) );
  XOR U1866 ( .A(ein[752]), .B(n1591), .Z(ereg_next[753]) );
  AND U1867 ( .A(mul_pow), .B(n1592), .Z(n1591) );
  XOR U1868 ( .A(ein[753]), .B(ein[752]), .Z(n1592) );
  XOR U1869 ( .A(ein[751]), .B(n1593), .Z(ereg_next[752]) );
  AND U1870 ( .A(mul_pow), .B(n1594), .Z(n1593) );
  XOR U1871 ( .A(ein[752]), .B(ein[751]), .Z(n1594) );
  XOR U1872 ( .A(ein[750]), .B(n1595), .Z(ereg_next[751]) );
  AND U1873 ( .A(mul_pow), .B(n1596), .Z(n1595) );
  XOR U1874 ( .A(ein[751]), .B(ein[750]), .Z(n1596) );
  XOR U1875 ( .A(ein[749]), .B(n1597), .Z(ereg_next[750]) );
  AND U1876 ( .A(mul_pow), .B(n1598), .Z(n1597) );
  XOR U1877 ( .A(ein[750]), .B(ein[749]), .Z(n1598) );
  XOR U1878 ( .A(ein[73]), .B(n1599), .Z(ereg_next[74]) );
  AND U1879 ( .A(mul_pow), .B(n1600), .Z(n1599) );
  XOR U1880 ( .A(ein[74]), .B(ein[73]), .Z(n1600) );
  XOR U1881 ( .A(ein[748]), .B(n1601), .Z(ereg_next[749]) );
  AND U1882 ( .A(mul_pow), .B(n1602), .Z(n1601) );
  XOR U1883 ( .A(ein[749]), .B(ein[748]), .Z(n1602) );
  XOR U1884 ( .A(ein[747]), .B(n1603), .Z(ereg_next[748]) );
  AND U1885 ( .A(mul_pow), .B(n1604), .Z(n1603) );
  XOR U1886 ( .A(ein[748]), .B(ein[747]), .Z(n1604) );
  XOR U1887 ( .A(ein[746]), .B(n1605), .Z(ereg_next[747]) );
  AND U1888 ( .A(mul_pow), .B(n1606), .Z(n1605) );
  XOR U1889 ( .A(ein[747]), .B(ein[746]), .Z(n1606) );
  XOR U1890 ( .A(ein[745]), .B(n1607), .Z(ereg_next[746]) );
  AND U1891 ( .A(mul_pow), .B(n1608), .Z(n1607) );
  XOR U1892 ( .A(ein[746]), .B(ein[745]), .Z(n1608) );
  XOR U1893 ( .A(ein[744]), .B(n1609), .Z(ereg_next[745]) );
  AND U1894 ( .A(mul_pow), .B(n1610), .Z(n1609) );
  XOR U1895 ( .A(ein[745]), .B(ein[744]), .Z(n1610) );
  XOR U1896 ( .A(ein[743]), .B(n1611), .Z(ereg_next[744]) );
  AND U1897 ( .A(mul_pow), .B(n1612), .Z(n1611) );
  XOR U1898 ( .A(ein[744]), .B(ein[743]), .Z(n1612) );
  XOR U1899 ( .A(ein[742]), .B(n1613), .Z(ereg_next[743]) );
  AND U1900 ( .A(mul_pow), .B(n1614), .Z(n1613) );
  XOR U1901 ( .A(ein[743]), .B(ein[742]), .Z(n1614) );
  XOR U1902 ( .A(ein[741]), .B(n1615), .Z(ereg_next[742]) );
  AND U1903 ( .A(mul_pow), .B(n1616), .Z(n1615) );
  XOR U1904 ( .A(ein[742]), .B(ein[741]), .Z(n1616) );
  XOR U1905 ( .A(ein[740]), .B(n1617), .Z(ereg_next[741]) );
  AND U1906 ( .A(mul_pow), .B(n1618), .Z(n1617) );
  XOR U1907 ( .A(ein[741]), .B(ein[740]), .Z(n1618) );
  XOR U1908 ( .A(ein[739]), .B(n1619), .Z(ereg_next[740]) );
  AND U1909 ( .A(mul_pow), .B(n1620), .Z(n1619) );
  XOR U1910 ( .A(ein[740]), .B(ein[739]), .Z(n1620) );
  XOR U1911 ( .A(ein[72]), .B(n1621), .Z(ereg_next[73]) );
  AND U1912 ( .A(mul_pow), .B(n1622), .Z(n1621) );
  XOR U1913 ( .A(ein[73]), .B(ein[72]), .Z(n1622) );
  XOR U1914 ( .A(ein[738]), .B(n1623), .Z(ereg_next[739]) );
  AND U1915 ( .A(mul_pow), .B(n1624), .Z(n1623) );
  XOR U1916 ( .A(ein[739]), .B(ein[738]), .Z(n1624) );
  XOR U1917 ( .A(ein[737]), .B(n1625), .Z(ereg_next[738]) );
  AND U1918 ( .A(mul_pow), .B(n1626), .Z(n1625) );
  XOR U1919 ( .A(ein[738]), .B(ein[737]), .Z(n1626) );
  XOR U1920 ( .A(ein[736]), .B(n1627), .Z(ereg_next[737]) );
  AND U1921 ( .A(mul_pow), .B(n1628), .Z(n1627) );
  XOR U1922 ( .A(ein[737]), .B(ein[736]), .Z(n1628) );
  XOR U1923 ( .A(ein[735]), .B(n1629), .Z(ereg_next[736]) );
  AND U1924 ( .A(mul_pow), .B(n1630), .Z(n1629) );
  XOR U1925 ( .A(ein[736]), .B(ein[735]), .Z(n1630) );
  XOR U1926 ( .A(ein[734]), .B(n1631), .Z(ereg_next[735]) );
  AND U1927 ( .A(mul_pow), .B(n1632), .Z(n1631) );
  XOR U1928 ( .A(ein[735]), .B(ein[734]), .Z(n1632) );
  XOR U1929 ( .A(ein[733]), .B(n1633), .Z(ereg_next[734]) );
  AND U1930 ( .A(mul_pow), .B(n1634), .Z(n1633) );
  XOR U1931 ( .A(ein[734]), .B(ein[733]), .Z(n1634) );
  XOR U1932 ( .A(ein[732]), .B(n1635), .Z(ereg_next[733]) );
  AND U1933 ( .A(mul_pow), .B(n1636), .Z(n1635) );
  XOR U1934 ( .A(ein[733]), .B(ein[732]), .Z(n1636) );
  XOR U1935 ( .A(ein[731]), .B(n1637), .Z(ereg_next[732]) );
  AND U1936 ( .A(mul_pow), .B(n1638), .Z(n1637) );
  XOR U1937 ( .A(ein[732]), .B(ein[731]), .Z(n1638) );
  XOR U1938 ( .A(ein[730]), .B(n1639), .Z(ereg_next[731]) );
  AND U1939 ( .A(mul_pow), .B(n1640), .Z(n1639) );
  XOR U1940 ( .A(ein[731]), .B(ein[730]), .Z(n1640) );
  XOR U1941 ( .A(ein[729]), .B(n1641), .Z(ereg_next[730]) );
  AND U1942 ( .A(mul_pow), .B(n1642), .Z(n1641) );
  XOR U1943 ( .A(ein[730]), .B(ein[729]), .Z(n1642) );
  XOR U1944 ( .A(ein[71]), .B(n1643), .Z(ereg_next[72]) );
  AND U1945 ( .A(mul_pow), .B(n1644), .Z(n1643) );
  XOR U1946 ( .A(ein[72]), .B(ein[71]), .Z(n1644) );
  XOR U1947 ( .A(ein[728]), .B(n1645), .Z(ereg_next[729]) );
  AND U1948 ( .A(mul_pow), .B(n1646), .Z(n1645) );
  XOR U1949 ( .A(ein[729]), .B(ein[728]), .Z(n1646) );
  XOR U1950 ( .A(ein[727]), .B(n1647), .Z(ereg_next[728]) );
  AND U1951 ( .A(mul_pow), .B(n1648), .Z(n1647) );
  XOR U1952 ( .A(ein[728]), .B(ein[727]), .Z(n1648) );
  XOR U1953 ( .A(ein[726]), .B(n1649), .Z(ereg_next[727]) );
  AND U1954 ( .A(mul_pow), .B(n1650), .Z(n1649) );
  XOR U1955 ( .A(ein[727]), .B(ein[726]), .Z(n1650) );
  XOR U1956 ( .A(ein[725]), .B(n1651), .Z(ereg_next[726]) );
  AND U1957 ( .A(mul_pow), .B(n1652), .Z(n1651) );
  XOR U1958 ( .A(ein[726]), .B(ein[725]), .Z(n1652) );
  XOR U1959 ( .A(ein[724]), .B(n1653), .Z(ereg_next[725]) );
  AND U1960 ( .A(mul_pow), .B(n1654), .Z(n1653) );
  XOR U1961 ( .A(ein[725]), .B(ein[724]), .Z(n1654) );
  XOR U1962 ( .A(ein[723]), .B(n1655), .Z(ereg_next[724]) );
  AND U1963 ( .A(mul_pow), .B(n1656), .Z(n1655) );
  XOR U1964 ( .A(ein[724]), .B(ein[723]), .Z(n1656) );
  XOR U1965 ( .A(ein[722]), .B(n1657), .Z(ereg_next[723]) );
  AND U1966 ( .A(mul_pow), .B(n1658), .Z(n1657) );
  XOR U1967 ( .A(ein[723]), .B(ein[722]), .Z(n1658) );
  XOR U1968 ( .A(ein[721]), .B(n1659), .Z(ereg_next[722]) );
  AND U1969 ( .A(mul_pow), .B(n1660), .Z(n1659) );
  XOR U1970 ( .A(ein[722]), .B(ein[721]), .Z(n1660) );
  XOR U1971 ( .A(ein[720]), .B(n1661), .Z(ereg_next[721]) );
  AND U1972 ( .A(mul_pow), .B(n1662), .Z(n1661) );
  XOR U1973 ( .A(ein[721]), .B(ein[720]), .Z(n1662) );
  XOR U1974 ( .A(ein[719]), .B(n1663), .Z(ereg_next[720]) );
  AND U1975 ( .A(mul_pow), .B(n1664), .Z(n1663) );
  XOR U1976 ( .A(ein[720]), .B(ein[719]), .Z(n1664) );
  XOR U1977 ( .A(ein[70]), .B(n1665), .Z(ereg_next[71]) );
  AND U1978 ( .A(mul_pow), .B(n1666), .Z(n1665) );
  XOR U1979 ( .A(ein[71]), .B(ein[70]), .Z(n1666) );
  XOR U1980 ( .A(ein[718]), .B(n1667), .Z(ereg_next[719]) );
  AND U1981 ( .A(mul_pow), .B(n1668), .Z(n1667) );
  XOR U1982 ( .A(ein[719]), .B(ein[718]), .Z(n1668) );
  XOR U1983 ( .A(ein[717]), .B(n1669), .Z(ereg_next[718]) );
  AND U1984 ( .A(mul_pow), .B(n1670), .Z(n1669) );
  XOR U1985 ( .A(ein[718]), .B(ein[717]), .Z(n1670) );
  XOR U1986 ( .A(ein[716]), .B(n1671), .Z(ereg_next[717]) );
  AND U1987 ( .A(mul_pow), .B(n1672), .Z(n1671) );
  XOR U1988 ( .A(ein[717]), .B(ein[716]), .Z(n1672) );
  XOR U1989 ( .A(ein[715]), .B(n1673), .Z(ereg_next[716]) );
  AND U1990 ( .A(mul_pow), .B(n1674), .Z(n1673) );
  XOR U1991 ( .A(ein[716]), .B(ein[715]), .Z(n1674) );
  XOR U1992 ( .A(ein[714]), .B(n1675), .Z(ereg_next[715]) );
  AND U1993 ( .A(mul_pow), .B(n1676), .Z(n1675) );
  XOR U1994 ( .A(ein[715]), .B(ein[714]), .Z(n1676) );
  XOR U1995 ( .A(ein[713]), .B(n1677), .Z(ereg_next[714]) );
  AND U1996 ( .A(mul_pow), .B(n1678), .Z(n1677) );
  XOR U1997 ( .A(ein[714]), .B(ein[713]), .Z(n1678) );
  XOR U1998 ( .A(ein[712]), .B(n1679), .Z(ereg_next[713]) );
  AND U1999 ( .A(mul_pow), .B(n1680), .Z(n1679) );
  XOR U2000 ( .A(ein[713]), .B(ein[712]), .Z(n1680) );
  XOR U2001 ( .A(ein[711]), .B(n1681), .Z(ereg_next[712]) );
  AND U2002 ( .A(mul_pow), .B(n1682), .Z(n1681) );
  XOR U2003 ( .A(ein[712]), .B(ein[711]), .Z(n1682) );
  XOR U2004 ( .A(ein[710]), .B(n1683), .Z(ereg_next[711]) );
  AND U2005 ( .A(mul_pow), .B(n1684), .Z(n1683) );
  XOR U2006 ( .A(ein[711]), .B(ein[710]), .Z(n1684) );
  XOR U2007 ( .A(ein[709]), .B(n1685), .Z(ereg_next[710]) );
  AND U2008 ( .A(mul_pow), .B(n1686), .Z(n1685) );
  XOR U2009 ( .A(ein[710]), .B(ein[709]), .Z(n1686) );
  XOR U2010 ( .A(ein[69]), .B(n1687), .Z(ereg_next[70]) );
  AND U2011 ( .A(mul_pow), .B(n1688), .Z(n1687) );
  XOR U2012 ( .A(ein[70]), .B(ein[69]), .Z(n1688) );
  XOR U2013 ( .A(ein[708]), .B(n1689), .Z(ereg_next[709]) );
  AND U2014 ( .A(mul_pow), .B(n1690), .Z(n1689) );
  XOR U2015 ( .A(ein[709]), .B(ein[708]), .Z(n1690) );
  XOR U2016 ( .A(ein[707]), .B(n1691), .Z(ereg_next[708]) );
  AND U2017 ( .A(mul_pow), .B(n1692), .Z(n1691) );
  XOR U2018 ( .A(ein[708]), .B(ein[707]), .Z(n1692) );
  XOR U2019 ( .A(ein[706]), .B(n1693), .Z(ereg_next[707]) );
  AND U2020 ( .A(mul_pow), .B(n1694), .Z(n1693) );
  XOR U2021 ( .A(ein[707]), .B(ein[706]), .Z(n1694) );
  XOR U2022 ( .A(ein[705]), .B(n1695), .Z(ereg_next[706]) );
  AND U2023 ( .A(mul_pow), .B(n1696), .Z(n1695) );
  XOR U2024 ( .A(ein[706]), .B(ein[705]), .Z(n1696) );
  XOR U2025 ( .A(ein[704]), .B(n1697), .Z(ereg_next[705]) );
  AND U2026 ( .A(mul_pow), .B(n1698), .Z(n1697) );
  XOR U2027 ( .A(ein[705]), .B(ein[704]), .Z(n1698) );
  XOR U2028 ( .A(ein[703]), .B(n1699), .Z(ereg_next[704]) );
  AND U2029 ( .A(mul_pow), .B(n1700), .Z(n1699) );
  XOR U2030 ( .A(ein[704]), .B(ein[703]), .Z(n1700) );
  XOR U2031 ( .A(ein[702]), .B(n1701), .Z(ereg_next[703]) );
  AND U2032 ( .A(mul_pow), .B(n1702), .Z(n1701) );
  XOR U2033 ( .A(ein[703]), .B(ein[702]), .Z(n1702) );
  XOR U2034 ( .A(ein[701]), .B(n1703), .Z(ereg_next[702]) );
  AND U2035 ( .A(mul_pow), .B(n1704), .Z(n1703) );
  XOR U2036 ( .A(ein[702]), .B(ein[701]), .Z(n1704) );
  XOR U2037 ( .A(ein[700]), .B(n1705), .Z(ereg_next[701]) );
  AND U2038 ( .A(mul_pow), .B(n1706), .Z(n1705) );
  XOR U2039 ( .A(ein[701]), .B(ein[700]), .Z(n1706) );
  XOR U2040 ( .A(ein[699]), .B(n1707), .Z(ereg_next[700]) );
  AND U2041 ( .A(mul_pow), .B(n1708), .Z(n1707) );
  XOR U2042 ( .A(ein[700]), .B(ein[699]), .Z(n1708) );
  XOR U2043 ( .A(ein[5]), .B(n1709), .Z(ereg_next[6]) );
  AND U2044 ( .A(mul_pow), .B(n1710), .Z(n1709) );
  XOR U2045 ( .A(ein[6]), .B(ein[5]), .Z(n1710) );
  XOR U2046 ( .A(ein[68]), .B(n1711), .Z(ereg_next[69]) );
  AND U2047 ( .A(mul_pow), .B(n1712), .Z(n1711) );
  XOR U2048 ( .A(ein[69]), .B(ein[68]), .Z(n1712) );
  XOR U2049 ( .A(ein[698]), .B(n1713), .Z(ereg_next[699]) );
  AND U2050 ( .A(mul_pow), .B(n1714), .Z(n1713) );
  XOR U2051 ( .A(ein[699]), .B(ein[698]), .Z(n1714) );
  XOR U2052 ( .A(ein[697]), .B(n1715), .Z(ereg_next[698]) );
  AND U2053 ( .A(mul_pow), .B(n1716), .Z(n1715) );
  XOR U2054 ( .A(ein[698]), .B(ein[697]), .Z(n1716) );
  XOR U2055 ( .A(ein[696]), .B(n1717), .Z(ereg_next[697]) );
  AND U2056 ( .A(mul_pow), .B(n1718), .Z(n1717) );
  XOR U2057 ( .A(ein[697]), .B(ein[696]), .Z(n1718) );
  XOR U2058 ( .A(ein[695]), .B(n1719), .Z(ereg_next[696]) );
  AND U2059 ( .A(mul_pow), .B(n1720), .Z(n1719) );
  XOR U2060 ( .A(ein[696]), .B(ein[695]), .Z(n1720) );
  XOR U2061 ( .A(ein[694]), .B(n1721), .Z(ereg_next[695]) );
  AND U2062 ( .A(mul_pow), .B(n1722), .Z(n1721) );
  XOR U2063 ( .A(ein[695]), .B(ein[694]), .Z(n1722) );
  XOR U2064 ( .A(ein[693]), .B(n1723), .Z(ereg_next[694]) );
  AND U2065 ( .A(mul_pow), .B(n1724), .Z(n1723) );
  XOR U2066 ( .A(ein[694]), .B(ein[693]), .Z(n1724) );
  XOR U2067 ( .A(ein[692]), .B(n1725), .Z(ereg_next[693]) );
  AND U2068 ( .A(mul_pow), .B(n1726), .Z(n1725) );
  XOR U2069 ( .A(ein[693]), .B(ein[692]), .Z(n1726) );
  XOR U2070 ( .A(ein[691]), .B(n1727), .Z(ereg_next[692]) );
  AND U2071 ( .A(mul_pow), .B(n1728), .Z(n1727) );
  XOR U2072 ( .A(ein[692]), .B(ein[691]), .Z(n1728) );
  XOR U2073 ( .A(ein[690]), .B(n1729), .Z(ereg_next[691]) );
  AND U2074 ( .A(mul_pow), .B(n1730), .Z(n1729) );
  XOR U2075 ( .A(ein[691]), .B(ein[690]), .Z(n1730) );
  XOR U2076 ( .A(ein[689]), .B(n1731), .Z(ereg_next[690]) );
  AND U2077 ( .A(mul_pow), .B(n1732), .Z(n1731) );
  XOR U2078 ( .A(ein[690]), .B(ein[689]), .Z(n1732) );
  XOR U2079 ( .A(ein[67]), .B(n1733), .Z(ereg_next[68]) );
  AND U2080 ( .A(mul_pow), .B(n1734), .Z(n1733) );
  XOR U2081 ( .A(ein[68]), .B(ein[67]), .Z(n1734) );
  XOR U2082 ( .A(ein[688]), .B(n1735), .Z(ereg_next[689]) );
  AND U2083 ( .A(mul_pow), .B(n1736), .Z(n1735) );
  XOR U2084 ( .A(ein[689]), .B(ein[688]), .Z(n1736) );
  XOR U2085 ( .A(ein[687]), .B(n1737), .Z(ereg_next[688]) );
  AND U2086 ( .A(mul_pow), .B(n1738), .Z(n1737) );
  XOR U2087 ( .A(ein[688]), .B(ein[687]), .Z(n1738) );
  XOR U2088 ( .A(ein[686]), .B(n1739), .Z(ereg_next[687]) );
  AND U2089 ( .A(mul_pow), .B(n1740), .Z(n1739) );
  XOR U2090 ( .A(ein[687]), .B(ein[686]), .Z(n1740) );
  XOR U2091 ( .A(ein[685]), .B(n1741), .Z(ereg_next[686]) );
  AND U2092 ( .A(mul_pow), .B(n1742), .Z(n1741) );
  XOR U2093 ( .A(ein[686]), .B(ein[685]), .Z(n1742) );
  XOR U2094 ( .A(ein[684]), .B(n1743), .Z(ereg_next[685]) );
  AND U2095 ( .A(mul_pow), .B(n1744), .Z(n1743) );
  XOR U2096 ( .A(ein[685]), .B(ein[684]), .Z(n1744) );
  XOR U2097 ( .A(ein[683]), .B(n1745), .Z(ereg_next[684]) );
  AND U2098 ( .A(mul_pow), .B(n1746), .Z(n1745) );
  XOR U2099 ( .A(ein[684]), .B(ein[683]), .Z(n1746) );
  XOR U2100 ( .A(ein[682]), .B(n1747), .Z(ereg_next[683]) );
  AND U2101 ( .A(mul_pow), .B(n1748), .Z(n1747) );
  XOR U2102 ( .A(ein[683]), .B(ein[682]), .Z(n1748) );
  XOR U2103 ( .A(ein[681]), .B(n1749), .Z(ereg_next[682]) );
  AND U2104 ( .A(mul_pow), .B(n1750), .Z(n1749) );
  XOR U2105 ( .A(ein[682]), .B(ein[681]), .Z(n1750) );
  XOR U2106 ( .A(ein[680]), .B(n1751), .Z(ereg_next[681]) );
  AND U2107 ( .A(mul_pow), .B(n1752), .Z(n1751) );
  XOR U2108 ( .A(ein[681]), .B(ein[680]), .Z(n1752) );
  XOR U2109 ( .A(ein[679]), .B(n1753), .Z(ereg_next[680]) );
  AND U2110 ( .A(mul_pow), .B(n1754), .Z(n1753) );
  XOR U2111 ( .A(ein[680]), .B(ein[679]), .Z(n1754) );
  XOR U2112 ( .A(ein[66]), .B(n1755), .Z(ereg_next[67]) );
  AND U2113 ( .A(mul_pow), .B(n1756), .Z(n1755) );
  XOR U2114 ( .A(ein[67]), .B(ein[66]), .Z(n1756) );
  XOR U2115 ( .A(ein[678]), .B(n1757), .Z(ereg_next[679]) );
  AND U2116 ( .A(mul_pow), .B(n1758), .Z(n1757) );
  XOR U2117 ( .A(ein[679]), .B(ein[678]), .Z(n1758) );
  XOR U2118 ( .A(ein[677]), .B(n1759), .Z(ereg_next[678]) );
  AND U2119 ( .A(mul_pow), .B(n1760), .Z(n1759) );
  XOR U2120 ( .A(ein[678]), .B(ein[677]), .Z(n1760) );
  XOR U2121 ( .A(ein[676]), .B(n1761), .Z(ereg_next[677]) );
  AND U2122 ( .A(mul_pow), .B(n1762), .Z(n1761) );
  XOR U2123 ( .A(ein[677]), .B(ein[676]), .Z(n1762) );
  XOR U2124 ( .A(ein[675]), .B(n1763), .Z(ereg_next[676]) );
  AND U2125 ( .A(mul_pow), .B(n1764), .Z(n1763) );
  XOR U2126 ( .A(ein[676]), .B(ein[675]), .Z(n1764) );
  XOR U2127 ( .A(ein[674]), .B(n1765), .Z(ereg_next[675]) );
  AND U2128 ( .A(mul_pow), .B(n1766), .Z(n1765) );
  XOR U2129 ( .A(ein[675]), .B(ein[674]), .Z(n1766) );
  XOR U2130 ( .A(ein[673]), .B(n1767), .Z(ereg_next[674]) );
  AND U2131 ( .A(mul_pow), .B(n1768), .Z(n1767) );
  XOR U2132 ( .A(ein[674]), .B(ein[673]), .Z(n1768) );
  XOR U2133 ( .A(ein[672]), .B(n1769), .Z(ereg_next[673]) );
  AND U2134 ( .A(mul_pow), .B(n1770), .Z(n1769) );
  XOR U2135 ( .A(ein[673]), .B(ein[672]), .Z(n1770) );
  XOR U2136 ( .A(ein[671]), .B(n1771), .Z(ereg_next[672]) );
  AND U2137 ( .A(mul_pow), .B(n1772), .Z(n1771) );
  XOR U2138 ( .A(ein[672]), .B(ein[671]), .Z(n1772) );
  XOR U2139 ( .A(ein[670]), .B(n1773), .Z(ereg_next[671]) );
  AND U2140 ( .A(mul_pow), .B(n1774), .Z(n1773) );
  XOR U2141 ( .A(ein[671]), .B(ein[670]), .Z(n1774) );
  XOR U2142 ( .A(ein[669]), .B(n1775), .Z(ereg_next[670]) );
  AND U2143 ( .A(mul_pow), .B(n1776), .Z(n1775) );
  XOR U2144 ( .A(ein[670]), .B(ein[669]), .Z(n1776) );
  XOR U2145 ( .A(ein[65]), .B(n1777), .Z(ereg_next[66]) );
  AND U2146 ( .A(mul_pow), .B(n1778), .Z(n1777) );
  XOR U2147 ( .A(ein[66]), .B(ein[65]), .Z(n1778) );
  XOR U2148 ( .A(ein[668]), .B(n1779), .Z(ereg_next[669]) );
  AND U2149 ( .A(mul_pow), .B(n1780), .Z(n1779) );
  XOR U2150 ( .A(ein[669]), .B(ein[668]), .Z(n1780) );
  XOR U2151 ( .A(ein[667]), .B(n1781), .Z(ereg_next[668]) );
  AND U2152 ( .A(mul_pow), .B(n1782), .Z(n1781) );
  XOR U2153 ( .A(ein[668]), .B(ein[667]), .Z(n1782) );
  XOR U2154 ( .A(ein[666]), .B(n1783), .Z(ereg_next[667]) );
  AND U2155 ( .A(mul_pow), .B(n1784), .Z(n1783) );
  XOR U2156 ( .A(ein[667]), .B(ein[666]), .Z(n1784) );
  XOR U2157 ( .A(ein[665]), .B(n1785), .Z(ereg_next[666]) );
  AND U2158 ( .A(mul_pow), .B(n1786), .Z(n1785) );
  XOR U2159 ( .A(ein[666]), .B(ein[665]), .Z(n1786) );
  XOR U2160 ( .A(ein[664]), .B(n1787), .Z(ereg_next[665]) );
  AND U2161 ( .A(mul_pow), .B(n1788), .Z(n1787) );
  XOR U2162 ( .A(ein[665]), .B(ein[664]), .Z(n1788) );
  XOR U2163 ( .A(ein[663]), .B(n1789), .Z(ereg_next[664]) );
  AND U2164 ( .A(mul_pow), .B(n1790), .Z(n1789) );
  XOR U2165 ( .A(ein[664]), .B(ein[663]), .Z(n1790) );
  XOR U2166 ( .A(ein[662]), .B(n1791), .Z(ereg_next[663]) );
  AND U2167 ( .A(mul_pow), .B(n1792), .Z(n1791) );
  XOR U2168 ( .A(ein[663]), .B(ein[662]), .Z(n1792) );
  XOR U2169 ( .A(ein[661]), .B(n1793), .Z(ereg_next[662]) );
  AND U2170 ( .A(mul_pow), .B(n1794), .Z(n1793) );
  XOR U2171 ( .A(ein[662]), .B(ein[661]), .Z(n1794) );
  XOR U2172 ( .A(ein[660]), .B(n1795), .Z(ereg_next[661]) );
  AND U2173 ( .A(mul_pow), .B(n1796), .Z(n1795) );
  XOR U2174 ( .A(ein[661]), .B(ein[660]), .Z(n1796) );
  XOR U2175 ( .A(ein[659]), .B(n1797), .Z(ereg_next[660]) );
  AND U2176 ( .A(mul_pow), .B(n1798), .Z(n1797) );
  XOR U2177 ( .A(ein[660]), .B(ein[659]), .Z(n1798) );
  XOR U2178 ( .A(ein[64]), .B(n1799), .Z(ereg_next[65]) );
  AND U2179 ( .A(mul_pow), .B(n1800), .Z(n1799) );
  XOR U2180 ( .A(ein[65]), .B(ein[64]), .Z(n1800) );
  XOR U2181 ( .A(ein[658]), .B(n1801), .Z(ereg_next[659]) );
  AND U2182 ( .A(mul_pow), .B(n1802), .Z(n1801) );
  XOR U2183 ( .A(ein[659]), .B(ein[658]), .Z(n1802) );
  XOR U2184 ( .A(ein[657]), .B(n1803), .Z(ereg_next[658]) );
  AND U2185 ( .A(mul_pow), .B(n1804), .Z(n1803) );
  XOR U2186 ( .A(ein[658]), .B(ein[657]), .Z(n1804) );
  XOR U2187 ( .A(ein[656]), .B(n1805), .Z(ereg_next[657]) );
  AND U2188 ( .A(mul_pow), .B(n1806), .Z(n1805) );
  XOR U2189 ( .A(ein[657]), .B(ein[656]), .Z(n1806) );
  XOR U2190 ( .A(ein[655]), .B(n1807), .Z(ereg_next[656]) );
  AND U2191 ( .A(mul_pow), .B(n1808), .Z(n1807) );
  XOR U2192 ( .A(ein[656]), .B(ein[655]), .Z(n1808) );
  XOR U2193 ( .A(ein[654]), .B(n1809), .Z(ereg_next[655]) );
  AND U2194 ( .A(mul_pow), .B(n1810), .Z(n1809) );
  XOR U2195 ( .A(ein[655]), .B(ein[654]), .Z(n1810) );
  XOR U2196 ( .A(ein[653]), .B(n1811), .Z(ereg_next[654]) );
  AND U2197 ( .A(mul_pow), .B(n1812), .Z(n1811) );
  XOR U2198 ( .A(ein[654]), .B(ein[653]), .Z(n1812) );
  XOR U2199 ( .A(ein[652]), .B(n1813), .Z(ereg_next[653]) );
  AND U2200 ( .A(mul_pow), .B(n1814), .Z(n1813) );
  XOR U2201 ( .A(ein[653]), .B(ein[652]), .Z(n1814) );
  XOR U2202 ( .A(ein[651]), .B(n1815), .Z(ereg_next[652]) );
  AND U2203 ( .A(mul_pow), .B(n1816), .Z(n1815) );
  XOR U2204 ( .A(ein[652]), .B(ein[651]), .Z(n1816) );
  XOR U2205 ( .A(ein[650]), .B(n1817), .Z(ereg_next[651]) );
  AND U2206 ( .A(mul_pow), .B(n1818), .Z(n1817) );
  XOR U2207 ( .A(ein[651]), .B(ein[650]), .Z(n1818) );
  XOR U2208 ( .A(ein[649]), .B(n1819), .Z(ereg_next[650]) );
  AND U2209 ( .A(mul_pow), .B(n1820), .Z(n1819) );
  XOR U2210 ( .A(ein[650]), .B(ein[649]), .Z(n1820) );
  XOR U2211 ( .A(ein[63]), .B(n1821), .Z(ereg_next[64]) );
  AND U2212 ( .A(mul_pow), .B(n1822), .Z(n1821) );
  XOR U2213 ( .A(ein[64]), .B(ein[63]), .Z(n1822) );
  XOR U2214 ( .A(ein[648]), .B(n1823), .Z(ereg_next[649]) );
  AND U2215 ( .A(mul_pow), .B(n1824), .Z(n1823) );
  XOR U2216 ( .A(ein[649]), .B(ein[648]), .Z(n1824) );
  XOR U2217 ( .A(ein[647]), .B(n1825), .Z(ereg_next[648]) );
  AND U2218 ( .A(mul_pow), .B(n1826), .Z(n1825) );
  XOR U2219 ( .A(ein[648]), .B(ein[647]), .Z(n1826) );
  XOR U2220 ( .A(ein[646]), .B(n1827), .Z(ereg_next[647]) );
  AND U2221 ( .A(mul_pow), .B(n1828), .Z(n1827) );
  XOR U2222 ( .A(ein[647]), .B(ein[646]), .Z(n1828) );
  XOR U2223 ( .A(ein[645]), .B(n1829), .Z(ereg_next[646]) );
  AND U2224 ( .A(mul_pow), .B(n1830), .Z(n1829) );
  XOR U2225 ( .A(ein[646]), .B(ein[645]), .Z(n1830) );
  XOR U2226 ( .A(ein[644]), .B(n1831), .Z(ereg_next[645]) );
  AND U2227 ( .A(mul_pow), .B(n1832), .Z(n1831) );
  XOR U2228 ( .A(ein[645]), .B(ein[644]), .Z(n1832) );
  XOR U2229 ( .A(ein[643]), .B(n1833), .Z(ereg_next[644]) );
  AND U2230 ( .A(mul_pow), .B(n1834), .Z(n1833) );
  XOR U2231 ( .A(ein[644]), .B(ein[643]), .Z(n1834) );
  XOR U2232 ( .A(ein[642]), .B(n1835), .Z(ereg_next[643]) );
  AND U2233 ( .A(mul_pow), .B(n1836), .Z(n1835) );
  XOR U2234 ( .A(ein[643]), .B(ein[642]), .Z(n1836) );
  XOR U2235 ( .A(ein[641]), .B(n1837), .Z(ereg_next[642]) );
  AND U2236 ( .A(mul_pow), .B(n1838), .Z(n1837) );
  XOR U2237 ( .A(ein[642]), .B(ein[641]), .Z(n1838) );
  XOR U2238 ( .A(ein[640]), .B(n1839), .Z(ereg_next[641]) );
  AND U2239 ( .A(mul_pow), .B(n1840), .Z(n1839) );
  XOR U2240 ( .A(ein[641]), .B(ein[640]), .Z(n1840) );
  XOR U2241 ( .A(ein[639]), .B(n1841), .Z(ereg_next[640]) );
  AND U2242 ( .A(mul_pow), .B(n1842), .Z(n1841) );
  XOR U2243 ( .A(ein[640]), .B(ein[639]), .Z(n1842) );
  XOR U2244 ( .A(ein[62]), .B(n1843), .Z(ereg_next[63]) );
  AND U2245 ( .A(mul_pow), .B(n1844), .Z(n1843) );
  XOR U2246 ( .A(ein[63]), .B(ein[62]), .Z(n1844) );
  XOR U2247 ( .A(ein[638]), .B(n1845), .Z(ereg_next[639]) );
  AND U2248 ( .A(mul_pow), .B(n1846), .Z(n1845) );
  XOR U2249 ( .A(ein[639]), .B(ein[638]), .Z(n1846) );
  XOR U2250 ( .A(ein[637]), .B(n1847), .Z(ereg_next[638]) );
  AND U2251 ( .A(mul_pow), .B(n1848), .Z(n1847) );
  XOR U2252 ( .A(ein[638]), .B(ein[637]), .Z(n1848) );
  XOR U2253 ( .A(ein[636]), .B(n1849), .Z(ereg_next[637]) );
  AND U2254 ( .A(mul_pow), .B(n1850), .Z(n1849) );
  XOR U2255 ( .A(ein[637]), .B(ein[636]), .Z(n1850) );
  XOR U2256 ( .A(ein[635]), .B(n1851), .Z(ereg_next[636]) );
  AND U2257 ( .A(mul_pow), .B(n1852), .Z(n1851) );
  XOR U2258 ( .A(ein[636]), .B(ein[635]), .Z(n1852) );
  XOR U2259 ( .A(ein[634]), .B(n1853), .Z(ereg_next[635]) );
  AND U2260 ( .A(mul_pow), .B(n1854), .Z(n1853) );
  XOR U2261 ( .A(ein[635]), .B(ein[634]), .Z(n1854) );
  XOR U2262 ( .A(ein[633]), .B(n1855), .Z(ereg_next[634]) );
  AND U2263 ( .A(mul_pow), .B(n1856), .Z(n1855) );
  XOR U2264 ( .A(ein[634]), .B(ein[633]), .Z(n1856) );
  XOR U2265 ( .A(ein[632]), .B(n1857), .Z(ereg_next[633]) );
  AND U2266 ( .A(mul_pow), .B(n1858), .Z(n1857) );
  XOR U2267 ( .A(ein[633]), .B(ein[632]), .Z(n1858) );
  XOR U2268 ( .A(ein[631]), .B(n1859), .Z(ereg_next[632]) );
  AND U2269 ( .A(mul_pow), .B(n1860), .Z(n1859) );
  XOR U2270 ( .A(ein[632]), .B(ein[631]), .Z(n1860) );
  XOR U2271 ( .A(ein[630]), .B(n1861), .Z(ereg_next[631]) );
  AND U2272 ( .A(mul_pow), .B(n1862), .Z(n1861) );
  XOR U2273 ( .A(ein[631]), .B(ein[630]), .Z(n1862) );
  XOR U2274 ( .A(ein[629]), .B(n1863), .Z(ereg_next[630]) );
  AND U2275 ( .A(mul_pow), .B(n1864), .Z(n1863) );
  XOR U2276 ( .A(ein[630]), .B(ein[629]), .Z(n1864) );
  XOR U2277 ( .A(ein[61]), .B(n1865), .Z(ereg_next[62]) );
  AND U2278 ( .A(mul_pow), .B(n1866), .Z(n1865) );
  XOR U2279 ( .A(ein[62]), .B(ein[61]), .Z(n1866) );
  XOR U2280 ( .A(ein[628]), .B(n1867), .Z(ereg_next[629]) );
  AND U2281 ( .A(mul_pow), .B(n1868), .Z(n1867) );
  XOR U2282 ( .A(ein[629]), .B(ein[628]), .Z(n1868) );
  XOR U2283 ( .A(ein[627]), .B(n1869), .Z(ereg_next[628]) );
  AND U2284 ( .A(mul_pow), .B(n1870), .Z(n1869) );
  XOR U2285 ( .A(ein[628]), .B(ein[627]), .Z(n1870) );
  XOR U2286 ( .A(ein[626]), .B(n1871), .Z(ereg_next[627]) );
  AND U2287 ( .A(mul_pow), .B(n1872), .Z(n1871) );
  XOR U2288 ( .A(ein[627]), .B(ein[626]), .Z(n1872) );
  XOR U2289 ( .A(ein[625]), .B(n1873), .Z(ereg_next[626]) );
  AND U2290 ( .A(mul_pow), .B(n1874), .Z(n1873) );
  XOR U2291 ( .A(ein[626]), .B(ein[625]), .Z(n1874) );
  XOR U2292 ( .A(ein[624]), .B(n1875), .Z(ereg_next[625]) );
  AND U2293 ( .A(mul_pow), .B(n1876), .Z(n1875) );
  XOR U2294 ( .A(ein[625]), .B(ein[624]), .Z(n1876) );
  XOR U2295 ( .A(ein[623]), .B(n1877), .Z(ereg_next[624]) );
  AND U2296 ( .A(mul_pow), .B(n1878), .Z(n1877) );
  XOR U2297 ( .A(ein[624]), .B(ein[623]), .Z(n1878) );
  XOR U2298 ( .A(ein[622]), .B(n1879), .Z(ereg_next[623]) );
  AND U2299 ( .A(mul_pow), .B(n1880), .Z(n1879) );
  XOR U2300 ( .A(ein[623]), .B(ein[622]), .Z(n1880) );
  XOR U2301 ( .A(ein[621]), .B(n1881), .Z(ereg_next[622]) );
  AND U2302 ( .A(mul_pow), .B(n1882), .Z(n1881) );
  XOR U2303 ( .A(ein[622]), .B(ein[621]), .Z(n1882) );
  XOR U2304 ( .A(ein[620]), .B(n1883), .Z(ereg_next[621]) );
  AND U2305 ( .A(mul_pow), .B(n1884), .Z(n1883) );
  XOR U2306 ( .A(ein[621]), .B(ein[620]), .Z(n1884) );
  XOR U2307 ( .A(ein[619]), .B(n1885), .Z(ereg_next[620]) );
  AND U2308 ( .A(mul_pow), .B(n1886), .Z(n1885) );
  XOR U2309 ( .A(ein[620]), .B(ein[619]), .Z(n1886) );
  XOR U2310 ( .A(ein[60]), .B(n1887), .Z(ereg_next[61]) );
  AND U2311 ( .A(mul_pow), .B(n1888), .Z(n1887) );
  XOR U2312 ( .A(ein[61]), .B(ein[60]), .Z(n1888) );
  XOR U2313 ( .A(ein[618]), .B(n1889), .Z(ereg_next[619]) );
  AND U2314 ( .A(mul_pow), .B(n1890), .Z(n1889) );
  XOR U2315 ( .A(ein[619]), .B(ein[618]), .Z(n1890) );
  XOR U2316 ( .A(ein[617]), .B(n1891), .Z(ereg_next[618]) );
  AND U2317 ( .A(mul_pow), .B(n1892), .Z(n1891) );
  XOR U2318 ( .A(ein[618]), .B(ein[617]), .Z(n1892) );
  XOR U2319 ( .A(ein[616]), .B(n1893), .Z(ereg_next[617]) );
  AND U2320 ( .A(mul_pow), .B(n1894), .Z(n1893) );
  XOR U2321 ( .A(ein[617]), .B(ein[616]), .Z(n1894) );
  XOR U2322 ( .A(ein[615]), .B(n1895), .Z(ereg_next[616]) );
  AND U2323 ( .A(mul_pow), .B(n1896), .Z(n1895) );
  XOR U2324 ( .A(ein[616]), .B(ein[615]), .Z(n1896) );
  XOR U2325 ( .A(ein[614]), .B(n1897), .Z(ereg_next[615]) );
  AND U2326 ( .A(mul_pow), .B(n1898), .Z(n1897) );
  XOR U2327 ( .A(ein[615]), .B(ein[614]), .Z(n1898) );
  XOR U2328 ( .A(ein[613]), .B(n1899), .Z(ereg_next[614]) );
  AND U2329 ( .A(mul_pow), .B(n1900), .Z(n1899) );
  XOR U2330 ( .A(ein[614]), .B(ein[613]), .Z(n1900) );
  XOR U2331 ( .A(ein[612]), .B(n1901), .Z(ereg_next[613]) );
  AND U2332 ( .A(mul_pow), .B(n1902), .Z(n1901) );
  XOR U2333 ( .A(ein[613]), .B(ein[612]), .Z(n1902) );
  XOR U2334 ( .A(ein[611]), .B(n1903), .Z(ereg_next[612]) );
  AND U2335 ( .A(mul_pow), .B(n1904), .Z(n1903) );
  XOR U2336 ( .A(ein[612]), .B(ein[611]), .Z(n1904) );
  XOR U2337 ( .A(ein[610]), .B(n1905), .Z(ereg_next[611]) );
  AND U2338 ( .A(mul_pow), .B(n1906), .Z(n1905) );
  XOR U2339 ( .A(ein[611]), .B(ein[610]), .Z(n1906) );
  XOR U2340 ( .A(ein[609]), .B(n1907), .Z(ereg_next[610]) );
  AND U2341 ( .A(mul_pow), .B(n1908), .Z(n1907) );
  XOR U2342 ( .A(ein[610]), .B(ein[609]), .Z(n1908) );
  XOR U2343 ( .A(ein[59]), .B(n1909), .Z(ereg_next[60]) );
  AND U2344 ( .A(mul_pow), .B(n1910), .Z(n1909) );
  XOR U2345 ( .A(ein[60]), .B(ein[59]), .Z(n1910) );
  XOR U2346 ( .A(ein[608]), .B(n1911), .Z(ereg_next[609]) );
  AND U2347 ( .A(mul_pow), .B(n1912), .Z(n1911) );
  XOR U2348 ( .A(ein[609]), .B(ein[608]), .Z(n1912) );
  XOR U2349 ( .A(ein[607]), .B(n1913), .Z(ereg_next[608]) );
  AND U2350 ( .A(mul_pow), .B(n1914), .Z(n1913) );
  XOR U2351 ( .A(ein[608]), .B(ein[607]), .Z(n1914) );
  XOR U2352 ( .A(ein[606]), .B(n1915), .Z(ereg_next[607]) );
  AND U2353 ( .A(mul_pow), .B(n1916), .Z(n1915) );
  XOR U2354 ( .A(ein[607]), .B(ein[606]), .Z(n1916) );
  XOR U2355 ( .A(ein[605]), .B(n1917), .Z(ereg_next[606]) );
  AND U2356 ( .A(mul_pow), .B(n1918), .Z(n1917) );
  XOR U2357 ( .A(ein[606]), .B(ein[605]), .Z(n1918) );
  XOR U2358 ( .A(ein[604]), .B(n1919), .Z(ereg_next[605]) );
  AND U2359 ( .A(mul_pow), .B(n1920), .Z(n1919) );
  XOR U2360 ( .A(ein[605]), .B(ein[604]), .Z(n1920) );
  XOR U2361 ( .A(ein[603]), .B(n1921), .Z(ereg_next[604]) );
  AND U2362 ( .A(mul_pow), .B(n1922), .Z(n1921) );
  XOR U2363 ( .A(ein[604]), .B(ein[603]), .Z(n1922) );
  XOR U2364 ( .A(ein[602]), .B(n1923), .Z(ereg_next[603]) );
  AND U2365 ( .A(mul_pow), .B(n1924), .Z(n1923) );
  XOR U2366 ( .A(ein[603]), .B(ein[602]), .Z(n1924) );
  XOR U2367 ( .A(ein[601]), .B(n1925), .Z(ereg_next[602]) );
  AND U2368 ( .A(mul_pow), .B(n1926), .Z(n1925) );
  XOR U2369 ( .A(ein[602]), .B(ein[601]), .Z(n1926) );
  XOR U2370 ( .A(ein[600]), .B(n1927), .Z(ereg_next[601]) );
  AND U2371 ( .A(mul_pow), .B(n1928), .Z(n1927) );
  XOR U2372 ( .A(ein[601]), .B(ein[600]), .Z(n1928) );
  XOR U2373 ( .A(ein[599]), .B(n1929), .Z(ereg_next[600]) );
  AND U2374 ( .A(mul_pow), .B(n1930), .Z(n1929) );
  XOR U2375 ( .A(ein[600]), .B(ein[599]), .Z(n1930) );
  XOR U2376 ( .A(ein[4]), .B(n1931), .Z(ereg_next[5]) );
  AND U2377 ( .A(mul_pow), .B(n1932), .Z(n1931) );
  XOR U2378 ( .A(ein[5]), .B(ein[4]), .Z(n1932) );
  XOR U2379 ( .A(ein[58]), .B(n1933), .Z(ereg_next[59]) );
  AND U2380 ( .A(mul_pow), .B(n1934), .Z(n1933) );
  XOR U2381 ( .A(ein[59]), .B(ein[58]), .Z(n1934) );
  XOR U2382 ( .A(ein[598]), .B(n1935), .Z(ereg_next[599]) );
  AND U2383 ( .A(mul_pow), .B(n1936), .Z(n1935) );
  XOR U2384 ( .A(ein[599]), .B(ein[598]), .Z(n1936) );
  XOR U2385 ( .A(ein[597]), .B(n1937), .Z(ereg_next[598]) );
  AND U2386 ( .A(mul_pow), .B(n1938), .Z(n1937) );
  XOR U2387 ( .A(ein[598]), .B(ein[597]), .Z(n1938) );
  XOR U2388 ( .A(ein[596]), .B(n1939), .Z(ereg_next[597]) );
  AND U2389 ( .A(mul_pow), .B(n1940), .Z(n1939) );
  XOR U2390 ( .A(ein[597]), .B(ein[596]), .Z(n1940) );
  XOR U2391 ( .A(ein[595]), .B(n1941), .Z(ereg_next[596]) );
  AND U2392 ( .A(mul_pow), .B(n1942), .Z(n1941) );
  XOR U2393 ( .A(ein[596]), .B(ein[595]), .Z(n1942) );
  XOR U2394 ( .A(ein[594]), .B(n1943), .Z(ereg_next[595]) );
  AND U2395 ( .A(mul_pow), .B(n1944), .Z(n1943) );
  XOR U2396 ( .A(ein[595]), .B(ein[594]), .Z(n1944) );
  XOR U2397 ( .A(ein[593]), .B(n1945), .Z(ereg_next[594]) );
  AND U2398 ( .A(mul_pow), .B(n1946), .Z(n1945) );
  XOR U2399 ( .A(ein[594]), .B(ein[593]), .Z(n1946) );
  XOR U2400 ( .A(ein[592]), .B(n1947), .Z(ereg_next[593]) );
  AND U2401 ( .A(mul_pow), .B(n1948), .Z(n1947) );
  XOR U2402 ( .A(ein[593]), .B(ein[592]), .Z(n1948) );
  XOR U2403 ( .A(ein[591]), .B(n1949), .Z(ereg_next[592]) );
  AND U2404 ( .A(mul_pow), .B(n1950), .Z(n1949) );
  XOR U2405 ( .A(ein[592]), .B(ein[591]), .Z(n1950) );
  XOR U2406 ( .A(ein[590]), .B(n1951), .Z(ereg_next[591]) );
  AND U2407 ( .A(mul_pow), .B(n1952), .Z(n1951) );
  XOR U2408 ( .A(ein[591]), .B(ein[590]), .Z(n1952) );
  XOR U2409 ( .A(ein[589]), .B(n1953), .Z(ereg_next[590]) );
  AND U2410 ( .A(mul_pow), .B(n1954), .Z(n1953) );
  XOR U2411 ( .A(ein[590]), .B(ein[589]), .Z(n1954) );
  XOR U2412 ( .A(ein[57]), .B(n1955), .Z(ereg_next[58]) );
  AND U2413 ( .A(mul_pow), .B(n1956), .Z(n1955) );
  XOR U2414 ( .A(ein[58]), .B(ein[57]), .Z(n1956) );
  XOR U2415 ( .A(ein[588]), .B(n1957), .Z(ereg_next[589]) );
  AND U2416 ( .A(mul_pow), .B(n1958), .Z(n1957) );
  XOR U2417 ( .A(ein[589]), .B(ein[588]), .Z(n1958) );
  XOR U2418 ( .A(ein[587]), .B(n1959), .Z(ereg_next[588]) );
  AND U2419 ( .A(mul_pow), .B(n1960), .Z(n1959) );
  XOR U2420 ( .A(ein[588]), .B(ein[587]), .Z(n1960) );
  XOR U2421 ( .A(ein[586]), .B(n1961), .Z(ereg_next[587]) );
  AND U2422 ( .A(mul_pow), .B(n1962), .Z(n1961) );
  XOR U2423 ( .A(ein[587]), .B(ein[586]), .Z(n1962) );
  XOR U2424 ( .A(ein[585]), .B(n1963), .Z(ereg_next[586]) );
  AND U2425 ( .A(mul_pow), .B(n1964), .Z(n1963) );
  XOR U2426 ( .A(ein[586]), .B(ein[585]), .Z(n1964) );
  XOR U2427 ( .A(ein[584]), .B(n1965), .Z(ereg_next[585]) );
  AND U2428 ( .A(mul_pow), .B(n1966), .Z(n1965) );
  XOR U2429 ( .A(ein[585]), .B(ein[584]), .Z(n1966) );
  XOR U2430 ( .A(ein[583]), .B(n1967), .Z(ereg_next[584]) );
  AND U2431 ( .A(mul_pow), .B(n1968), .Z(n1967) );
  XOR U2432 ( .A(ein[584]), .B(ein[583]), .Z(n1968) );
  XOR U2433 ( .A(ein[582]), .B(n1969), .Z(ereg_next[583]) );
  AND U2434 ( .A(mul_pow), .B(n1970), .Z(n1969) );
  XOR U2435 ( .A(ein[583]), .B(ein[582]), .Z(n1970) );
  XOR U2436 ( .A(ein[581]), .B(n1971), .Z(ereg_next[582]) );
  AND U2437 ( .A(mul_pow), .B(n1972), .Z(n1971) );
  XOR U2438 ( .A(ein[582]), .B(ein[581]), .Z(n1972) );
  XOR U2439 ( .A(ein[580]), .B(n1973), .Z(ereg_next[581]) );
  AND U2440 ( .A(mul_pow), .B(n1974), .Z(n1973) );
  XOR U2441 ( .A(ein[581]), .B(ein[580]), .Z(n1974) );
  XOR U2442 ( .A(ein[579]), .B(n1975), .Z(ereg_next[580]) );
  AND U2443 ( .A(mul_pow), .B(n1976), .Z(n1975) );
  XOR U2444 ( .A(ein[580]), .B(ein[579]), .Z(n1976) );
  XOR U2445 ( .A(ein[56]), .B(n1977), .Z(ereg_next[57]) );
  AND U2446 ( .A(mul_pow), .B(n1978), .Z(n1977) );
  XOR U2447 ( .A(ein[57]), .B(ein[56]), .Z(n1978) );
  XOR U2448 ( .A(ein[578]), .B(n1979), .Z(ereg_next[579]) );
  AND U2449 ( .A(mul_pow), .B(n1980), .Z(n1979) );
  XOR U2450 ( .A(ein[579]), .B(ein[578]), .Z(n1980) );
  XOR U2451 ( .A(ein[577]), .B(n1981), .Z(ereg_next[578]) );
  AND U2452 ( .A(mul_pow), .B(n1982), .Z(n1981) );
  XOR U2453 ( .A(ein[578]), .B(ein[577]), .Z(n1982) );
  XOR U2454 ( .A(ein[576]), .B(n1983), .Z(ereg_next[577]) );
  AND U2455 ( .A(mul_pow), .B(n1984), .Z(n1983) );
  XOR U2456 ( .A(ein[577]), .B(ein[576]), .Z(n1984) );
  XOR U2457 ( .A(ein[575]), .B(n1985), .Z(ereg_next[576]) );
  AND U2458 ( .A(mul_pow), .B(n1986), .Z(n1985) );
  XOR U2459 ( .A(ein[576]), .B(ein[575]), .Z(n1986) );
  XOR U2460 ( .A(ein[574]), .B(n1987), .Z(ereg_next[575]) );
  AND U2461 ( .A(mul_pow), .B(n1988), .Z(n1987) );
  XOR U2462 ( .A(ein[575]), .B(ein[574]), .Z(n1988) );
  XOR U2463 ( .A(ein[573]), .B(n1989), .Z(ereg_next[574]) );
  AND U2464 ( .A(mul_pow), .B(n1990), .Z(n1989) );
  XOR U2465 ( .A(ein[574]), .B(ein[573]), .Z(n1990) );
  XOR U2466 ( .A(ein[572]), .B(n1991), .Z(ereg_next[573]) );
  AND U2467 ( .A(mul_pow), .B(n1992), .Z(n1991) );
  XOR U2468 ( .A(ein[573]), .B(ein[572]), .Z(n1992) );
  XOR U2469 ( .A(ein[571]), .B(n1993), .Z(ereg_next[572]) );
  AND U2470 ( .A(mul_pow), .B(n1994), .Z(n1993) );
  XOR U2471 ( .A(ein[572]), .B(ein[571]), .Z(n1994) );
  XOR U2472 ( .A(ein[570]), .B(n1995), .Z(ereg_next[571]) );
  AND U2473 ( .A(mul_pow), .B(n1996), .Z(n1995) );
  XOR U2474 ( .A(ein[571]), .B(ein[570]), .Z(n1996) );
  XOR U2475 ( .A(ein[569]), .B(n1997), .Z(ereg_next[570]) );
  AND U2476 ( .A(mul_pow), .B(n1998), .Z(n1997) );
  XOR U2477 ( .A(ein[570]), .B(ein[569]), .Z(n1998) );
  XOR U2478 ( .A(ein[55]), .B(n1999), .Z(ereg_next[56]) );
  AND U2479 ( .A(mul_pow), .B(n2000), .Z(n1999) );
  XOR U2480 ( .A(ein[56]), .B(ein[55]), .Z(n2000) );
  XOR U2481 ( .A(ein[568]), .B(n2001), .Z(ereg_next[569]) );
  AND U2482 ( .A(mul_pow), .B(n2002), .Z(n2001) );
  XOR U2483 ( .A(ein[569]), .B(ein[568]), .Z(n2002) );
  XOR U2484 ( .A(ein[567]), .B(n2003), .Z(ereg_next[568]) );
  AND U2485 ( .A(mul_pow), .B(n2004), .Z(n2003) );
  XOR U2486 ( .A(ein[568]), .B(ein[567]), .Z(n2004) );
  XOR U2487 ( .A(ein[566]), .B(n2005), .Z(ereg_next[567]) );
  AND U2488 ( .A(mul_pow), .B(n2006), .Z(n2005) );
  XOR U2489 ( .A(ein[567]), .B(ein[566]), .Z(n2006) );
  XOR U2490 ( .A(ein[565]), .B(n2007), .Z(ereg_next[566]) );
  AND U2491 ( .A(mul_pow), .B(n2008), .Z(n2007) );
  XOR U2492 ( .A(ein[566]), .B(ein[565]), .Z(n2008) );
  XOR U2493 ( .A(ein[564]), .B(n2009), .Z(ereg_next[565]) );
  AND U2494 ( .A(mul_pow), .B(n2010), .Z(n2009) );
  XOR U2495 ( .A(ein[565]), .B(ein[564]), .Z(n2010) );
  XOR U2496 ( .A(ein[563]), .B(n2011), .Z(ereg_next[564]) );
  AND U2497 ( .A(mul_pow), .B(n2012), .Z(n2011) );
  XOR U2498 ( .A(ein[564]), .B(ein[563]), .Z(n2012) );
  XOR U2499 ( .A(ein[562]), .B(n2013), .Z(ereg_next[563]) );
  AND U2500 ( .A(mul_pow), .B(n2014), .Z(n2013) );
  XOR U2501 ( .A(ein[563]), .B(ein[562]), .Z(n2014) );
  XOR U2502 ( .A(ein[561]), .B(n2015), .Z(ereg_next[562]) );
  AND U2503 ( .A(mul_pow), .B(n2016), .Z(n2015) );
  XOR U2504 ( .A(ein[562]), .B(ein[561]), .Z(n2016) );
  XOR U2505 ( .A(ein[560]), .B(n2017), .Z(ereg_next[561]) );
  AND U2506 ( .A(mul_pow), .B(n2018), .Z(n2017) );
  XOR U2507 ( .A(ein[561]), .B(ein[560]), .Z(n2018) );
  XOR U2508 ( .A(ein[559]), .B(n2019), .Z(ereg_next[560]) );
  AND U2509 ( .A(mul_pow), .B(n2020), .Z(n2019) );
  XOR U2510 ( .A(ein[560]), .B(ein[559]), .Z(n2020) );
  XOR U2511 ( .A(ein[54]), .B(n2021), .Z(ereg_next[55]) );
  AND U2512 ( .A(mul_pow), .B(n2022), .Z(n2021) );
  XOR U2513 ( .A(ein[55]), .B(ein[54]), .Z(n2022) );
  XOR U2514 ( .A(ein[558]), .B(n2023), .Z(ereg_next[559]) );
  AND U2515 ( .A(mul_pow), .B(n2024), .Z(n2023) );
  XOR U2516 ( .A(ein[559]), .B(ein[558]), .Z(n2024) );
  XOR U2517 ( .A(ein[557]), .B(n2025), .Z(ereg_next[558]) );
  AND U2518 ( .A(mul_pow), .B(n2026), .Z(n2025) );
  XOR U2519 ( .A(ein[558]), .B(ein[557]), .Z(n2026) );
  XOR U2520 ( .A(ein[556]), .B(n2027), .Z(ereg_next[557]) );
  AND U2521 ( .A(mul_pow), .B(n2028), .Z(n2027) );
  XOR U2522 ( .A(ein[557]), .B(ein[556]), .Z(n2028) );
  XOR U2523 ( .A(ein[555]), .B(n2029), .Z(ereg_next[556]) );
  AND U2524 ( .A(mul_pow), .B(n2030), .Z(n2029) );
  XOR U2525 ( .A(ein[556]), .B(ein[555]), .Z(n2030) );
  XOR U2526 ( .A(ein[554]), .B(n2031), .Z(ereg_next[555]) );
  AND U2527 ( .A(mul_pow), .B(n2032), .Z(n2031) );
  XOR U2528 ( .A(ein[555]), .B(ein[554]), .Z(n2032) );
  XOR U2529 ( .A(ein[553]), .B(n2033), .Z(ereg_next[554]) );
  AND U2530 ( .A(mul_pow), .B(n2034), .Z(n2033) );
  XOR U2531 ( .A(ein[554]), .B(ein[553]), .Z(n2034) );
  XOR U2532 ( .A(ein[552]), .B(n2035), .Z(ereg_next[553]) );
  AND U2533 ( .A(mul_pow), .B(n2036), .Z(n2035) );
  XOR U2534 ( .A(ein[553]), .B(ein[552]), .Z(n2036) );
  XOR U2535 ( .A(ein[551]), .B(n2037), .Z(ereg_next[552]) );
  AND U2536 ( .A(mul_pow), .B(n2038), .Z(n2037) );
  XOR U2537 ( .A(ein[552]), .B(ein[551]), .Z(n2038) );
  XOR U2538 ( .A(ein[550]), .B(n2039), .Z(ereg_next[551]) );
  AND U2539 ( .A(mul_pow), .B(n2040), .Z(n2039) );
  XOR U2540 ( .A(ein[551]), .B(ein[550]), .Z(n2040) );
  XOR U2541 ( .A(ein[549]), .B(n2041), .Z(ereg_next[550]) );
  AND U2542 ( .A(mul_pow), .B(n2042), .Z(n2041) );
  XOR U2543 ( .A(ein[550]), .B(ein[549]), .Z(n2042) );
  XOR U2544 ( .A(ein[53]), .B(n2043), .Z(ereg_next[54]) );
  AND U2545 ( .A(mul_pow), .B(n2044), .Z(n2043) );
  XOR U2546 ( .A(ein[54]), .B(ein[53]), .Z(n2044) );
  XOR U2547 ( .A(ein[548]), .B(n2045), .Z(ereg_next[549]) );
  AND U2548 ( .A(mul_pow), .B(n2046), .Z(n2045) );
  XOR U2549 ( .A(ein[549]), .B(ein[548]), .Z(n2046) );
  XOR U2550 ( .A(ein[547]), .B(n2047), .Z(ereg_next[548]) );
  AND U2551 ( .A(mul_pow), .B(n2048), .Z(n2047) );
  XOR U2552 ( .A(ein[548]), .B(ein[547]), .Z(n2048) );
  XOR U2553 ( .A(ein[546]), .B(n2049), .Z(ereg_next[547]) );
  AND U2554 ( .A(mul_pow), .B(n2050), .Z(n2049) );
  XOR U2555 ( .A(ein[547]), .B(ein[546]), .Z(n2050) );
  XOR U2556 ( .A(ein[545]), .B(n2051), .Z(ereg_next[546]) );
  AND U2557 ( .A(mul_pow), .B(n2052), .Z(n2051) );
  XOR U2558 ( .A(ein[546]), .B(ein[545]), .Z(n2052) );
  XOR U2559 ( .A(ein[544]), .B(n2053), .Z(ereg_next[545]) );
  AND U2560 ( .A(mul_pow), .B(n2054), .Z(n2053) );
  XOR U2561 ( .A(ein[545]), .B(ein[544]), .Z(n2054) );
  XOR U2562 ( .A(ein[543]), .B(n2055), .Z(ereg_next[544]) );
  AND U2563 ( .A(mul_pow), .B(n2056), .Z(n2055) );
  XOR U2564 ( .A(ein[544]), .B(ein[543]), .Z(n2056) );
  XOR U2565 ( .A(ein[542]), .B(n2057), .Z(ereg_next[543]) );
  AND U2566 ( .A(mul_pow), .B(n2058), .Z(n2057) );
  XOR U2567 ( .A(ein[543]), .B(ein[542]), .Z(n2058) );
  XOR U2568 ( .A(ein[541]), .B(n2059), .Z(ereg_next[542]) );
  AND U2569 ( .A(mul_pow), .B(n2060), .Z(n2059) );
  XOR U2570 ( .A(ein[542]), .B(ein[541]), .Z(n2060) );
  XOR U2571 ( .A(ein[540]), .B(n2061), .Z(ereg_next[541]) );
  AND U2572 ( .A(mul_pow), .B(n2062), .Z(n2061) );
  XOR U2573 ( .A(ein[541]), .B(ein[540]), .Z(n2062) );
  XOR U2574 ( .A(ein[539]), .B(n2063), .Z(ereg_next[540]) );
  AND U2575 ( .A(mul_pow), .B(n2064), .Z(n2063) );
  XOR U2576 ( .A(ein[540]), .B(ein[539]), .Z(n2064) );
  XOR U2577 ( .A(ein[52]), .B(n2065), .Z(ereg_next[53]) );
  AND U2578 ( .A(mul_pow), .B(n2066), .Z(n2065) );
  XOR U2579 ( .A(ein[53]), .B(ein[52]), .Z(n2066) );
  XOR U2580 ( .A(ein[538]), .B(n2067), .Z(ereg_next[539]) );
  AND U2581 ( .A(mul_pow), .B(n2068), .Z(n2067) );
  XOR U2582 ( .A(ein[539]), .B(ein[538]), .Z(n2068) );
  XOR U2583 ( .A(ein[537]), .B(n2069), .Z(ereg_next[538]) );
  AND U2584 ( .A(mul_pow), .B(n2070), .Z(n2069) );
  XOR U2585 ( .A(ein[538]), .B(ein[537]), .Z(n2070) );
  XOR U2586 ( .A(ein[536]), .B(n2071), .Z(ereg_next[537]) );
  AND U2587 ( .A(mul_pow), .B(n2072), .Z(n2071) );
  XOR U2588 ( .A(ein[537]), .B(ein[536]), .Z(n2072) );
  XOR U2589 ( .A(ein[535]), .B(n2073), .Z(ereg_next[536]) );
  AND U2590 ( .A(mul_pow), .B(n2074), .Z(n2073) );
  XOR U2591 ( .A(ein[536]), .B(ein[535]), .Z(n2074) );
  XOR U2592 ( .A(ein[534]), .B(n2075), .Z(ereg_next[535]) );
  AND U2593 ( .A(mul_pow), .B(n2076), .Z(n2075) );
  XOR U2594 ( .A(ein[535]), .B(ein[534]), .Z(n2076) );
  XOR U2595 ( .A(ein[533]), .B(n2077), .Z(ereg_next[534]) );
  AND U2596 ( .A(mul_pow), .B(n2078), .Z(n2077) );
  XOR U2597 ( .A(ein[534]), .B(ein[533]), .Z(n2078) );
  XOR U2598 ( .A(ein[532]), .B(n2079), .Z(ereg_next[533]) );
  AND U2599 ( .A(mul_pow), .B(n2080), .Z(n2079) );
  XOR U2600 ( .A(ein[533]), .B(ein[532]), .Z(n2080) );
  XOR U2601 ( .A(ein[531]), .B(n2081), .Z(ereg_next[532]) );
  AND U2602 ( .A(mul_pow), .B(n2082), .Z(n2081) );
  XOR U2603 ( .A(ein[532]), .B(ein[531]), .Z(n2082) );
  XOR U2604 ( .A(ein[530]), .B(n2083), .Z(ereg_next[531]) );
  AND U2605 ( .A(mul_pow), .B(n2084), .Z(n2083) );
  XOR U2606 ( .A(ein[531]), .B(ein[530]), .Z(n2084) );
  XOR U2607 ( .A(ein[529]), .B(n2085), .Z(ereg_next[530]) );
  AND U2608 ( .A(mul_pow), .B(n2086), .Z(n2085) );
  XOR U2609 ( .A(ein[530]), .B(ein[529]), .Z(n2086) );
  XOR U2610 ( .A(ein[51]), .B(n2087), .Z(ereg_next[52]) );
  AND U2611 ( .A(mul_pow), .B(n2088), .Z(n2087) );
  XOR U2612 ( .A(ein[52]), .B(ein[51]), .Z(n2088) );
  XOR U2613 ( .A(ein[528]), .B(n2089), .Z(ereg_next[529]) );
  AND U2614 ( .A(mul_pow), .B(n2090), .Z(n2089) );
  XOR U2615 ( .A(ein[529]), .B(ein[528]), .Z(n2090) );
  XOR U2616 ( .A(ein[527]), .B(n2091), .Z(ereg_next[528]) );
  AND U2617 ( .A(mul_pow), .B(n2092), .Z(n2091) );
  XOR U2618 ( .A(ein[528]), .B(ein[527]), .Z(n2092) );
  XOR U2619 ( .A(ein[526]), .B(n2093), .Z(ereg_next[527]) );
  AND U2620 ( .A(mul_pow), .B(n2094), .Z(n2093) );
  XOR U2621 ( .A(ein[527]), .B(ein[526]), .Z(n2094) );
  XOR U2622 ( .A(ein[525]), .B(n2095), .Z(ereg_next[526]) );
  AND U2623 ( .A(mul_pow), .B(n2096), .Z(n2095) );
  XOR U2624 ( .A(ein[526]), .B(ein[525]), .Z(n2096) );
  XOR U2625 ( .A(ein[524]), .B(n2097), .Z(ereg_next[525]) );
  AND U2626 ( .A(mul_pow), .B(n2098), .Z(n2097) );
  XOR U2627 ( .A(ein[525]), .B(ein[524]), .Z(n2098) );
  XOR U2628 ( .A(ein[523]), .B(n2099), .Z(ereg_next[524]) );
  AND U2629 ( .A(mul_pow), .B(n2100), .Z(n2099) );
  XOR U2630 ( .A(ein[524]), .B(ein[523]), .Z(n2100) );
  XOR U2631 ( .A(ein[522]), .B(n2101), .Z(ereg_next[523]) );
  AND U2632 ( .A(mul_pow), .B(n2102), .Z(n2101) );
  XOR U2633 ( .A(ein[523]), .B(ein[522]), .Z(n2102) );
  XOR U2634 ( .A(ein[521]), .B(n2103), .Z(ereg_next[522]) );
  AND U2635 ( .A(mul_pow), .B(n2104), .Z(n2103) );
  XOR U2636 ( .A(ein[522]), .B(ein[521]), .Z(n2104) );
  XOR U2637 ( .A(ein[520]), .B(n2105), .Z(ereg_next[521]) );
  AND U2638 ( .A(mul_pow), .B(n2106), .Z(n2105) );
  XOR U2639 ( .A(ein[521]), .B(ein[520]), .Z(n2106) );
  XOR U2640 ( .A(ein[519]), .B(n2107), .Z(ereg_next[520]) );
  AND U2641 ( .A(mul_pow), .B(n2108), .Z(n2107) );
  XOR U2642 ( .A(ein[520]), .B(ein[519]), .Z(n2108) );
  XOR U2643 ( .A(ein[50]), .B(n2109), .Z(ereg_next[51]) );
  AND U2644 ( .A(mul_pow), .B(n2110), .Z(n2109) );
  XOR U2645 ( .A(ein[51]), .B(ein[50]), .Z(n2110) );
  XOR U2646 ( .A(ein[518]), .B(n2111), .Z(ereg_next[519]) );
  AND U2647 ( .A(mul_pow), .B(n2112), .Z(n2111) );
  XOR U2648 ( .A(ein[519]), .B(ein[518]), .Z(n2112) );
  XOR U2649 ( .A(ein[517]), .B(n2113), .Z(ereg_next[518]) );
  AND U2650 ( .A(mul_pow), .B(n2114), .Z(n2113) );
  XOR U2651 ( .A(ein[518]), .B(ein[517]), .Z(n2114) );
  XOR U2652 ( .A(ein[516]), .B(n2115), .Z(ereg_next[517]) );
  AND U2653 ( .A(mul_pow), .B(n2116), .Z(n2115) );
  XOR U2654 ( .A(ein[517]), .B(ein[516]), .Z(n2116) );
  XOR U2655 ( .A(ein[515]), .B(n2117), .Z(ereg_next[516]) );
  AND U2656 ( .A(mul_pow), .B(n2118), .Z(n2117) );
  XOR U2657 ( .A(ein[516]), .B(ein[515]), .Z(n2118) );
  XOR U2658 ( .A(ein[514]), .B(n2119), .Z(ereg_next[515]) );
  AND U2659 ( .A(mul_pow), .B(n2120), .Z(n2119) );
  XOR U2660 ( .A(ein[515]), .B(ein[514]), .Z(n2120) );
  XOR U2661 ( .A(ein[513]), .B(n2121), .Z(ereg_next[514]) );
  AND U2662 ( .A(mul_pow), .B(n2122), .Z(n2121) );
  XOR U2663 ( .A(ein[514]), .B(ein[513]), .Z(n2122) );
  XOR U2664 ( .A(ein[512]), .B(n2123), .Z(ereg_next[513]) );
  AND U2665 ( .A(mul_pow), .B(n2124), .Z(n2123) );
  XOR U2666 ( .A(ein[513]), .B(ein[512]), .Z(n2124) );
  XOR U2667 ( .A(ein[511]), .B(n2125), .Z(ereg_next[512]) );
  AND U2668 ( .A(mul_pow), .B(n2126), .Z(n2125) );
  XOR U2669 ( .A(ein[512]), .B(ein[511]), .Z(n2126) );
  XOR U2670 ( .A(ein[510]), .B(n2127), .Z(ereg_next[511]) );
  AND U2671 ( .A(mul_pow), .B(n2128), .Z(n2127) );
  XOR U2672 ( .A(ein[511]), .B(ein[510]), .Z(n2128) );
  XOR U2673 ( .A(ein[509]), .B(n2129), .Z(ereg_next[510]) );
  AND U2674 ( .A(mul_pow), .B(n2130), .Z(n2129) );
  XOR U2675 ( .A(ein[510]), .B(ein[509]), .Z(n2130) );
  XOR U2676 ( .A(ein[49]), .B(n2131), .Z(ereg_next[50]) );
  AND U2677 ( .A(mul_pow), .B(n2132), .Z(n2131) );
  XOR U2678 ( .A(ein[50]), .B(ein[49]), .Z(n2132) );
  XOR U2679 ( .A(ein[508]), .B(n2133), .Z(ereg_next[509]) );
  AND U2680 ( .A(mul_pow), .B(n2134), .Z(n2133) );
  XOR U2681 ( .A(ein[509]), .B(ein[508]), .Z(n2134) );
  XOR U2682 ( .A(ein[507]), .B(n2135), .Z(ereg_next[508]) );
  AND U2683 ( .A(mul_pow), .B(n2136), .Z(n2135) );
  XOR U2684 ( .A(ein[508]), .B(ein[507]), .Z(n2136) );
  XOR U2685 ( .A(ein[506]), .B(n2137), .Z(ereg_next[507]) );
  AND U2686 ( .A(mul_pow), .B(n2138), .Z(n2137) );
  XOR U2687 ( .A(ein[507]), .B(ein[506]), .Z(n2138) );
  XOR U2688 ( .A(ein[505]), .B(n2139), .Z(ereg_next[506]) );
  AND U2689 ( .A(mul_pow), .B(n2140), .Z(n2139) );
  XOR U2690 ( .A(ein[506]), .B(ein[505]), .Z(n2140) );
  XOR U2691 ( .A(ein[504]), .B(n2141), .Z(ereg_next[505]) );
  AND U2692 ( .A(mul_pow), .B(n2142), .Z(n2141) );
  XOR U2693 ( .A(ein[505]), .B(ein[504]), .Z(n2142) );
  XOR U2694 ( .A(ein[503]), .B(n2143), .Z(ereg_next[504]) );
  AND U2695 ( .A(mul_pow), .B(n2144), .Z(n2143) );
  XOR U2696 ( .A(ein[504]), .B(ein[503]), .Z(n2144) );
  XOR U2697 ( .A(ein[502]), .B(n2145), .Z(ereg_next[503]) );
  AND U2698 ( .A(mul_pow), .B(n2146), .Z(n2145) );
  XOR U2699 ( .A(ein[503]), .B(ein[502]), .Z(n2146) );
  XOR U2700 ( .A(ein[501]), .B(n2147), .Z(ereg_next[502]) );
  AND U2701 ( .A(mul_pow), .B(n2148), .Z(n2147) );
  XOR U2702 ( .A(ein[502]), .B(ein[501]), .Z(n2148) );
  XOR U2703 ( .A(ein[500]), .B(n2149), .Z(ereg_next[501]) );
  AND U2704 ( .A(mul_pow), .B(n2150), .Z(n2149) );
  XOR U2705 ( .A(ein[501]), .B(ein[500]), .Z(n2150) );
  XOR U2706 ( .A(ein[499]), .B(n2151), .Z(ereg_next[500]) );
  AND U2707 ( .A(mul_pow), .B(n2152), .Z(n2151) );
  XOR U2708 ( .A(ein[500]), .B(ein[499]), .Z(n2152) );
  XOR U2709 ( .A(ein[3]), .B(n2153), .Z(ereg_next[4]) );
  AND U2710 ( .A(mul_pow), .B(n2154), .Z(n2153) );
  XOR U2711 ( .A(ein[4]), .B(ein[3]), .Z(n2154) );
  XOR U2712 ( .A(ein[48]), .B(n2155), .Z(ereg_next[49]) );
  AND U2713 ( .A(mul_pow), .B(n2156), .Z(n2155) );
  XOR U2714 ( .A(ein[49]), .B(ein[48]), .Z(n2156) );
  XOR U2715 ( .A(ein[498]), .B(n2157), .Z(ereg_next[499]) );
  AND U2716 ( .A(mul_pow), .B(n2158), .Z(n2157) );
  XOR U2717 ( .A(ein[499]), .B(ein[498]), .Z(n2158) );
  XOR U2718 ( .A(ein[497]), .B(n2159), .Z(ereg_next[498]) );
  AND U2719 ( .A(mul_pow), .B(n2160), .Z(n2159) );
  XOR U2720 ( .A(ein[498]), .B(ein[497]), .Z(n2160) );
  XOR U2721 ( .A(ein[496]), .B(n2161), .Z(ereg_next[497]) );
  AND U2722 ( .A(mul_pow), .B(n2162), .Z(n2161) );
  XOR U2723 ( .A(ein[497]), .B(ein[496]), .Z(n2162) );
  XOR U2724 ( .A(ein[495]), .B(n2163), .Z(ereg_next[496]) );
  AND U2725 ( .A(mul_pow), .B(n2164), .Z(n2163) );
  XOR U2726 ( .A(ein[496]), .B(ein[495]), .Z(n2164) );
  XOR U2727 ( .A(ein[494]), .B(n2165), .Z(ereg_next[495]) );
  AND U2728 ( .A(mul_pow), .B(n2166), .Z(n2165) );
  XOR U2729 ( .A(ein[495]), .B(ein[494]), .Z(n2166) );
  XOR U2730 ( .A(ein[493]), .B(n2167), .Z(ereg_next[494]) );
  AND U2731 ( .A(mul_pow), .B(n2168), .Z(n2167) );
  XOR U2732 ( .A(ein[494]), .B(ein[493]), .Z(n2168) );
  XOR U2733 ( .A(ein[492]), .B(n2169), .Z(ereg_next[493]) );
  AND U2734 ( .A(mul_pow), .B(n2170), .Z(n2169) );
  XOR U2735 ( .A(ein[493]), .B(ein[492]), .Z(n2170) );
  XOR U2736 ( .A(ein[491]), .B(n2171), .Z(ereg_next[492]) );
  AND U2737 ( .A(mul_pow), .B(n2172), .Z(n2171) );
  XOR U2738 ( .A(ein[492]), .B(ein[491]), .Z(n2172) );
  XOR U2739 ( .A(ein[490]), .B(n2173), .Z(ereg_next[491]) );
  AND U2740 ( .A(mul_pow), .B(n2174), .Z(n2173) );
  XOR U2741 ( .A(ein[491]), .B(ein[490]), .Z(n2174) );
  XOR U2742 ( .A(ein[489]), .B(n2175), .Z(ereg_next[490]) );
  AND U2743 ( .A(mul_pow), .B(n2176), .Z(n2175) );
  XOR U2744 ( .A(ein[490]), .B(ein[489]), .Z(n2176) );
  XOR U2745 ( .A(ein[47]), .B(n2177), .Z(ereg_next[48]) );
  AND U2746 ( .A(mul_pow), .B(n2178), .Z(n2177) );
  XOR U2747 ( .A(ein[48]), .B(ein[47]), .Z(n2178) );
  XOR U2748 ( .A(ein[488]), .B(n2179), .Z(ereg_next[489]) );
  AND U2749 ( .A(mul_pow), .B(n2180), .Z(n2179) );
  XOR U2750 ( .A(ein[489]), .B(ein[488]), .Z(n2180) );
  XOR U2751 ( .A(ein[487]), .B(n2181), .Z(ereg_next[488]) );
  AND U2752 ( .A(mul_pow), .B(n2182), .Z(n2181) );
  XOR U2753 ( .A(ein[488]), .B(ein[487]), .Z(n2182) );
  XOR U2754 ( .A(ein[486]), .B(n2183), .Z(ereg_next[487]) );
  AND U2755 ( .A(mul_pow), .B(n2184), .Z(n2183) );
  XOR U2756 ( .A(ein[487]), .B(ein[486]), .Z(n2184) );
  XOR U2757 ( .A(ein[485]), .B(n2185), .Z(ereg_next[486]) );
  AND U2758 ( .A(mul_pow), .B(n2186), .Z(n2185) );
  XOR U2759 ( .A(ein[486]), .B(ein[485]), .Z(n2186) );
  XOR U2760 ( .A(ein[484]), .B(n2187), .Z(ereg_next[485]) );
  AND U2761 ( .A(mul_pow), .B(n2188), .Z(n2187) );
  XOR U2762 ( .A(ein[485]), .B(ein[484]), .Z(n2188) );
  XOR U2763 ( .A(ein[483]), .B(n2189), .Z(ereg_next[484]) );
  AND U2764 ( .A(mul_pow), .B(n2190), .Z(n2189) );
  XOR U2765 ( .A(ein[484]), .B(ein[483]), .Z(n2190) );
  XOR U2766 ( .A(ein[482]), .B(n2191), .Z(ereg_next[483]) );
  AND U2767 ( .A(mul_pow), .B(n2192), .Z(n2191) );
  XOR U2768 ( .A(ein[483]), .B(ein[482]), .Z(n2192) );
  XOR U2769 ( .A(ein[481]), .B(n2193), .Z(ereg_next[482]) );
  AND U2770 ( .A(mul_pow), .B(n2194), .Z(n2193) );
  XOR U2771 ( .A(ein[482]), .B(ein[481]), .Z(n2194) );
  XOR U2772 ( .A(ein[480]), .B(n2195), .Z(ereg_next[481]) );
  AND U2773 ( .A(mul_pow), .B(n2196), .Z(n2195) );
  XOR U2774 ( .A(ein[481]), .B(ein[480]), .Z(n2196) );
  XOR U2775 ( .A(ein[479]), .B(n2197), .Z(ereg_next[480]) );
  AND U2776 ( .A(mul_pow), .B(n2198), .Z(n2197) );
  XOR U2777 ( .A(ein[480]), .B(ein[479]), .Z(n2198) );
  XOR U2778 ( .A(ein[46]), .B(n2199), .Z(ereg_next[47]) );
  AND U2779 ( .A(mul_pow), .B(n2200), .Z(n2199) );
  XOR U2780 ( .A(ein[47]), .B(ein[46]), .Z(n2200) );
  XOR U2781 ( .A(ein[478]), .B(n2201), .Z(ereg_next[479]) );
  AND U2782 ( .A(mul_pow), .B(n2202), .Z(n2201) );
  XOR U2783 ( .A(ein[479]), .B(ein[478]), .Z(n2202) );
  XOR U2784 ( .A(ein[477]), .B(n2203), .Z(ereg_next[478]) );
  AND U2785 ( .A(mul_pow), .B(n2204), .Z(n2203) );
  XOR U2786 ( .A(ein[478]), .B(ein[477]), .Z(n2204) );
  XOR U2787 ( .A(ein[476]), .B(n2205), .Z(ereg_next[477]) );
  AND U2788 ( .A(mul_pow), .B(n2206), .Z(n2205) );
  XOR U2789 ( .A(ein[477]), .B(ein[476]), .Z(n2206) );
  XOR U2790 ( .A(ein[475]), .B(n2207), .Z(ereg_next[476]) );
  AND U2791 ( .A(mul_pow), .B(n2208), .Z(n2207) );
  XOR U2792 ( .A(ein[476]), .B(ein[475]), .Z(n2208) );
  XOR U2793 ( .A(ein[474]), .B(n2209), .Z(ereg_next[475]) );
  AND U2794 ( .A(mul_pow), .B(n2210), .Z(n2209) );
  XOR U2795 ( .A(ein[475]), .B(ein[474]), .Z(n2210) );
  XOR U2796 ( .A(ein[473]), .B(n2211), .Z(ereg_next[474]) );
  AND U2797 ( .A(mul_pow), .B(n2212), .Z(n2211) );
  XOR U2798 ( .A(ein[474]), .B(ein[473]), .Z(n2212) );
  XOR U2799 ( .A(ein[472]), .B(n2213), .Z(ereg_next[473]) );
  AND U2800 ( .A(mul_pow), .B(n2214), .Z(n2213) );
  XOR U2801 ( .A(ein[473]), .B(ein[472]), .Z(n2214) );
  XOR U2802 ( .A(ein[471]), .B(n2215), .Z(ereg_next[472]) );
  AND U2803 ( .A(mul_pow), .B(n2216), .Z(n2215) );
  XOR U2804 ( .A(ein[472]), .B(ein[471]), .Z(n2216) );
  XOR U2805 ( .A(ein[470]), .B(n2217), .Z(ereg_next[471]) );
  AND U2806 ( .A(mul_pow), .B(n2218), .Z(n2217) );
  XOR U2807 ( .A(ein[471]), .B(ein[470]), .Z(n2218) );
  XOR U2808 ( .A(ein[469]), .B(n2219), .Z(ereg_next[470]) );
  AND U2809 ( .A(mul_pow), .B(n2220), .Z(n2219) );
  XOR U2810 ( .A(ein[470]), .B(ein[469]), .Z(n2220) );
  XOR U2811 ( .A(ein[45]), .B(n2221), .Z(ereg_next[46]) );
  AND U2812 ( .A(mul_pow), .B(n2222), .Z(n2221) );
  XOR U2813 ( .A(ein[46]), .B(ein[45]), .Z(n2222) );
  XOR U2814 ( .A(ein[468]), .B(n2223), .Z(ereg_next[469]) );
  AND U2815 ( .A(mul_pow), .B(n2224), .Z(n2223) );
  XOR U2816 ( .A(ein[469]), .B(ein[468]), .Z(n2224) );
  XOR U2817 ( .A(ein[467]), .B(n2225), .Z(ereg_next[468]) );
  AND U2818 ( .A(mul_pow), .B(n2226), .Z(n2225) );
  XOR U2819 ( .A(ein[468]), .B(ein[467]), .Z(n2226) );
  XOR U2820 ( .A(ein[466]), .B(n2227), .Z(ereg_next[467]) );
  AND U2821 ( .A(mul_pow), .B(n2228), .Z(n2227) );
  XOR U2822 ( .A(ein[467]), .B(ein[466]), .Z(n2228) );
  XOR U2823 ( .A(ein[465]), .B(n2229), .Z(ereg_next[466]) );
  AND U2824 ( .A(mul_pow), .B(n2230), .Z(n2229) );
  XOR U2825 ( .A(ein[466]), .B(ein[465]), .Z(n2230) );
  XOR U2826 ( .A(ein[464]), .B(n2231), .Z(ereg_next[465]) );
  AND U2827 ( .A(mul_pow), .B(n2232), .Z(n2231) );
  XOR U2828 ( .A(ein[465]), .B(ein[464]), .Z(n2232) );
  XOR U2829 ( .A(ein[463]), .B(n2233), .Z(ereg_next[464]) );
  AND U2830 ( .A(mul_pow), .B(n2234), .Z(n2233) );
  XOR U2831 ( .A(ein[464]), .B(ein[463]), .Z(n2234) );
  XOR U2832 ( .A(ein[462]), .B(n2235), .Z(ereg_next[463]) );
  AND U2833 ( .A(mul_pow), .B(n2236), .Z(n2235) );
  XOR U2834 ( .A(ein[463]), .B(ein[462]), .Z(n2236) );
  XOR U2835 ( .A(ein[461]), .B(n2237), .Z(ereg_next[462]) );
  AND U2836 ( .A(mul_pow), .B(n2238), .Z(n2237) );
  XOR U2837 ( .A(ein[462]), .B(ein[461]), .Z(n2238) );
  XOR U2838 ( .A(ein[460]), .B(n2239), .Z(ereg_next[461]) );
  AND U2839 ( .A(mul_pow), .B(n2240), .Z(n2239) );
  XOR U2840 ( .A(ein[461]), .B(ein[460]), .Z(n2240) );
  XOR U2841 ( .A(ein[459]), .B(n2241), .Z(ereg_next[460]) );
  AND U2842 ( .A(mul_pow), .B(n2242), .Z(n2241) );
  XOR U2843 ( .A(ein[460]), .B(ein[459]), .Z(n2242) );
  XOR U2844 ( .A(ein[44]), .B(n2243), .Z(ereg_next[45]) );
  AND U2845 ( .A(mul_pow), .B(n2244), .Z(n2243) );
  XOR U2846 ( .A(ein[45]), .B(ein[44]), .Z(n2244) );
  XOR U2847 ( .A(ein[458]), .B(n2245), .Z(ereg_next[459]) );
  AND U2848 ( .A(mul_pow), .B(n2246), .Z(n2245) );
  XOR U2849 ( .A(ein[459]), .B(ein[458]), .Z(n2246) );
  XOR U2850 ( .A(ein[457]), .B(n2247), .Z(ereg_next[458]) );
  AND U2851 ( .A(mul_pow), .B(n2248), .Z(n2247) );
  XOR U2852 ( .A(ein[458]), .B(ein[457]), .Z(n2248) );
  XOR U2853 ( .A(ein[456]), .B(n2249), .Z(ereg_next[457]) );
  AND U2854 ( .A(mul_pow), .B(n2250), .Z(n2249) );
  XOR U2855 ( .A(ein[457]), .B(ein[456]), .Z(n2250) );
  XOR U2856 ( .A(ein[455]), .B(n2251), .Z(ereg_next[456]) );
  AND U2857 ( .A(mul_pow), .B(n2252), .Z(n2251) );
  XOR U2858 ( .A(ein[456]), .B(ein[455]), .Z(n2252) );
  XOR U2859 ( .A(ein[454]), .B(n2253), .Z(ereg_next[455]) );
  AND U2860 ( .A(mul_pow), .B(n2254), .Z(n2253) );
  XOR U2861 ( .A(ein[455]), .B(ein[454]), .Z(n2254) );
  XOR U2862 ( .A(ein[453]), .B(n2255), .Z(ereg_next[454]) );
  AND U2863 ( .A(mul_pow), .B(n2256), .Z(n2255) );
  XOR U2864 ( .A(ein[454]), .B(ein[453]), .Z(n2256) );
  XOR U2865 ( .A(ein[452]), .B(n2257), .Z(ereg_next[453]) );
  AND U2866 ( .A(mul_pow), .B(n2258), .Z(n2257) );
  XOR U2867 ( .A(ein[453]), .B(ein[452]), .Z(n2258) );
  XOR U2868 ( .A(ein[451]), .B(n2259), .Z(ereg_next[452]) );
  AND U2869 ( .A(mul_pow), .B(n2260), .Z(n2259) );
  XOR U2870 ( .A(ein[452]), .B(ein[451]), .Z(n2260) );
  XOR U2871 ( .A(ein[450]), .B(n2261), .Z(ereg_next[451]) );
  AND U2872 ( .A(mul_pow), .B(n2262), .Z(n2261) );
  XOR U2873 ( .A(ein[451]), .B(ein[450]), .Z(n2262) );
  XOR U2874 ( .A(ein[449]), .B(n2263), .Z(ereg_next[450]) );
  AND U2875 ( .A(mul_pow), .B(n2264), .Z(n2263) );
  XOR U2876 ( .A(ein[450]), .B(ein[449]), .Z(n2264) );
  XOR U2877 ( .A(ein[43]), .B(n2265), .Z(ereg_next[44]) );
  AND U2878 ( .A(mul_pow), .B(n2266), .Z(n2265) );
  XOR U2879 ( .A(ein[44]), .B(ein[43]), .Z(n2266) );
  XOR U2880 ( .A(ein[448]), .B(n2267), .Z(ereg_next[449]) );
  AND U2881 ( .A(mul_pow), .B(n2268), .Z(n2267) );
  XOR U2882 ( .A(ein[449]), .B(ein[448]), .Z(n2268) );
  XOR U2883 ( .A(ein[447]), .B(n2269), .Z(ereg_next[448]) );
  AND U2884 ( .A(mul_pow), .B(n2270), .Z(n2269) );
  XOR U2885 ( .A(ein[448]), .B(ein[447]), .Z(n2270) );
  XOR U2886 ( .A(ein[446]), .B(n2271), .Z(ereg_next[447]) );
  AND U2887 ( .A(mul_pow), .B(n2272), .Z(n2271) );
  XOR U2888 ( .A(ein[447]), .B(ein[446]), .Z(n2272) );
  XOR U2889 ( .A(ein[445]), .B(n2273), .Z(ereg_next[446]) );
  AND U2890 ( .A(mul_pow), .B(n2274), .Z(n2273) );
  XOR U2891 ( .A(ein[446]), .B(ein[445]), .Z(n2274) );
  XOR U2892 ( .A(ein[444]), .B(n2275), .Z(ereg_next[445]) );
  AND U2893 ( .A(mul_pow), .B(n2276), .Z(n2275) );
  XOR U2894 ( .A(ein[445]), .B(ein[444]), .Z(n2276) );
  XOR U2895 ( .A(ein[443]), .B(n2277), .Z(ereg_next[444]) );
  AND U2896 ( .A(mul_pow), .B(n2278), .Z(n2277) );
  XOR U2897 ( .A(ein[444]), .B(ein[443]), .Z(n2278) );
  XOR U2898 ( .A(ein[442]), .B(n2279), .Z(ereg_next[443]) );
  AND U2899 ( .A(mul_pow), .B(n2280), .Z(n2279) );
  XOR U2900 ( .A(ein[443]), .B(ein[442]), .Z(n2280) );
  XOR U2901 ( .A(ein[441]), .B(n2281), .Z(ereg_next[442]) );
  AND U2902 ( .A(mul_pow), .B(n2282), .Z(n2281) );
  XOR U2903 ( .A(ein[442]), .B(ein[441]), .Z(n2282) );
  XOR U2904 ( .A(ein[440]), .B(n2283), .Z(ereg_next[441]) );
  AND U2905 ( .A(mul_pow), .B(n2284), .Z(n2283) );
  XOR U2906 ( .A(ein[441]), .B(ein[440]), .Z(n2284) );
  XOR U2907 ( .A(ein[439]), .B(n2285), .Z(ereg_next[440]) );
  AND U2908 ( .A(mul_pow), .B(n2286), .Z(n2285) );
  XOR U2909 ( .A(ein[440]), .B(ein[439]), .Z(n2286) );
  XOR U2910 ( .A(ein[42]), .B(n2287), .Z(ereg_next[43]) );
  AND U2911 ( .A(mul_pow), .B(n2288), .Z(n2287) );
  XOR U2912 ( .A(ein[43]), .B(ein[42]), .Z(n2288) );
  XOR U2913 ( .A(ein[438]), .B(n2289), .Z(ereg_next[439]) );
  AND U2914 ( .A(mul_pow), .B(n2290), .Z(n2289) );
  XOR U2915 ( .A(ein[439]), .B(ein[438]), .Z(n2290) );
  XOR U2916 ( .A(ein[437]), .B(n2291), .Z(ereg_next[438]) );
  AND U2917 ( .A(mul_pow), .B(n2292), .Z(n2291) );
  XOR U2918 ( .A(ein[438]), .B(ein[437]), .Z(n2292) );
  XOR U2919 ( .A(ein[436]), .B(n2293), .Z(ereg_next[437]) );
  AND U2920 ( .A(mul_pow), .B(n2294), .Z(n2293) );
  XOR U2921 ( .A(ein[437]), .B(ein[436]), .Z(n2294) );
  XOR U2922 ( .A(ein[435]), .B(n2295), .Z(ereg_next[436]) );
  AND U2923 ( .A(mul_pow), .B(n2296), .Z(n2295) );
  XOR U2924 ( .A(ein[436]), .B(ein[435]), .Z(n2296) );
  XOR U2925 ( .A(ein[434]), .B(n2297), .Z(ereg_next[435]) );
  AND U2926 ( .A(mul_pow), .B(n2298), .Z(n2297) );
  XOR U2927 ( .A(ein[435]), .B(ein[434]), .Z(n2298) );
  XOR U2928 ( .A(ein[433]), .B(n2299), .Z(ereg_next[434]) );
  AND U2929 ( .A(mul_pow), .B(n2300), .Z(n2299) );
  XOR U2930 ( .A(ein[434]), .B(ein[433]), .Z(n2300) );
  XOR U2931 ( .A(ein[432]), .B(n2301), .Z(ereg_next[433]) );
  AND U2932 ( .A(mul_pow), .B(n2302), .Z(n2301) );
  XOR U2933 ( .A(ein[433]), .B(ein[432]), .Z(n2302) );
  XOR U2934 ( .A(ein[431]), .B(n2303), .Z(ereg_next[432]) );
  AND U2935 ( .A(mul_pow), .B(n2304), .Z(n2303) );
  XOR U2936 ( .A(ein[432]), .B(ein[431]), .Z(n2304) );
  XOR U2937 ( .A(ein[430]), .B(n2305), .Z(ereg_next[431]) );
  AND U2938 ( .A(mul_pow), .B(n2306), .Z(n2305) );
  XOR U2939 ( .A(ein[431]), .B(ein[430]), .Z(n2306) );
  XOR U2940 ( .A(ein[429]), .B(n2307), .Z(ereg_next[430]) );
  AND U2941 ( .A(mul_pow), .B(n2308), .Z(n2307) );
  XOR U2942 ( .A(ein[430]), .B(ein[429]), .Z(n2308) );
  XOR U2943 ( .A(ein[41]), .B(n2309), .Z(ereg_next[42]) );
  AND U2944 ( .A(mul_pow), .B(n2310), .Z(n2309) );
  XOR U2945 ( .A(ein[42]), .B(ein[41]), .Z(n2310) );
  XOR U2946 ( .A(ein[428]), .B(n2311), .Z(ereg_next[429]) );
  AND U2947 ( .A(mul_pow), .B(n2312), .Z(n2311) );
  XOR U2948 ( .A(ein[429]), .B(ein[428]), .Z(n2312) );
  XOR U2949 ( .A(ein[427]), .B(n2313), .Z(ereg_next[428]) );
  AND U2950 ( .A(mul_pow), .B(n2314), .Z(n2313) );
  XOR U2951 ( .A(ein[428]), .B(ein[427]), .Z(n2314) );
  XOR U2952 ( .A(ein[426]), .B(n2315), .Z(ereg_next[427]) );
  AND U2953 ( .A(mul_pow), .B(n2316), .Z(n2315) );
  XOR U2954 ( .A(ein[427]), .B(ein[426]), .Z(n2316) );
  XOR U2955 ( .A(ein[425]), .B(n2317), .Z(ereg_next[426]) );
  AND U2956 ( .A(mul_pow), .B(n2318), .Z(n2317) );
  XOR U2957 ( .A(ein[426]), .B(ein[425]), .Z(n2318) );
  XOR U2958 ( .A(ein[424]), .B(n2319), .Z(ereg_next[425]) );
  AND U2959 ( .A(mul_pow), .B(n2320), .Z(n2319) );
  XOR U2960 ( .A(ein[425]), .B(ein[424]), .Z(n2320) );
  XOR U2961 ( .A(ein[423]), .B(n2321), .Z(ereg_next[424]) );
  AND U2962 ( .A(mul_pow), .B(n2322), .Z(n2321) );
  XOR U2963 ( .A(ein[424]), .B(ein[423]), .Z(n2322) );
  XOR U2964 ( .A(ein[422]), .B(n2323), .Z(ereg_next[423]) );
  AND U2965 ( .A(mul_pow), .B(n2324), .Z(n2323) );
  XOR U2966 ( .A(ein[423]), .B(ein[422]), .Z(n2324) );
  XOR U2967 ( .A(ein[421]), .B(n2325), .Z(ereg_next[422]) );
  AND U2968 ( .A(mul_pow), .B(n2326), .Z(n2325) );
  XOR U2969 ( .A(ein[422]), .B(ein[421]), .Z(n2326) );
  XOR U2970 ( .A(ein[420]), .B(n2327), .Z(ereg_next[421]) );
  AND U2971 ( .A(mul_pow), .B(n2328), .Z(n2327) );
  XOR U2972 ( .A(ein[421]), .B(ein[420]), .Z(n2328) );
  XOR U2973 ( .A(ein[419]), .B(n2329), .Z(ereg_next[420]) );
  AND U2974 ( .A(mul_pow), .B(n2330), .Z(n2329) );
  XOR U2975 ( .A(ein[420]), .B(ein[419]), .Z(n2330) );
  XOR U2976 ( .A(ein[40]), .B(n2331), .Z(ereg_next[41]) );
  AND U2977 ( .A(mul_pow), .B(n2332), .Z(n2331) );
  XOR U2978 ( .A(ein[41]), .B(ein[40]), .Z(n2332) );
  XOR U2979 ( .A(ein[418]), .B(n2333), .Z(ereg_next[419]) );
  AND U2980 ( .A(mul_pow), .B(n2334), .Z(n2333) );
  XOR U2981 ( .A(ein[419]), .B(ein[418]), .Z(n2334) );
  XOR U2982 ( .A(ein[417]), .B(n2335), .Z(ereg_next[418]) );
  AND U2983 ( .A(mul_pow), .B(n2336), .Z(n2335) );
  XOR U2984 ( .A(ein[418]), .B(ein[417]), .Z(n2336) );
  XOR U2985 ( .A(ein[416]), .B(n2337), .Z(ereg_next[417]) );
  AND U2986 ( .A(mul_pow), .B(n2338), .Z(n2337) );
  XOR U2987 ( .A(ein[417]), .B(ein[416]), .Z(n2338) );
  XOR U2988 ( .A(ein[415]), .B(n2339), .Z(ereg_next[416]) );
  AND U2989 ( .A(mul_pow), .B(n2340), .Z(n2339) );
  XOR U2990 ( .A(ein[416]), .B(ein[415]), .Z(n2340) );
  XOR U2991 ( .A(ein[414]), .B(n2341), .Z(ereg_next[415]) );
  AND U2992 ( .A(mul_pow), .B(n2342), .Z(n2341) );
  XOR U2993 ( .A(ein[415]), .B(ein[414]), .Z(n2342) );
  XOR U2994 ( .A(ein[413]), .B(n2343), .Z(ereg_next[414]) );
  AND U2995 ( .A(mul_pow), .B(n2344), .Z(n2343) );
  XOR U2996 ( .A(ein[414]), .B(ein[413]), .Z(n2344) );
  XOR U2997 ( .A(ein[412]), .B(n2345), .Z(ereg_next[413]) );
  AND U2998 ( .A(mul_pow), .B(n2346), .Z(n2345) );
  XOR U2999 ( .A(ein[413]), .B(ein[412]), .Z(n2346) );
  XOR U3000 ( .A(ein[411]), .B(n2347), .Z(ereg_next[412]) );
  AND U3001 ( .A(mul_pow), .B(n2348), .Z(n2347) );
  XOR U3002 ( .A(ein[412]), .B(ein[411]), .Z(n2348) );
  XOR U3003 ( .A(ein[410]), .B(n2349), .Z(ereg_next[411]) );
  AND U3004 ( .A(mul_pow), .B(n2350), .Z(n2349) );
  XOR U3005 ( .A(ein[411]), .B(ein[410]), .Z(n2350) );
  XOR U3006 ( .A(ein[409]), .B(n2351), .Z(ereg_next[410]) );
  AND U3007 ( .A(mul_pow), .B(n2352), .Z(n2351) );
  XOR U3008 ( .A(ein[410]), .B(ein[409]), .Z(n2352) );
  XOR U3009 ( .A(ein[39]), .B(n2353), .Z(ereg_next[40]) );
  AND U3010 ( .A(mul_pow), .B(n2354), .Z(n2353) );
  XOR U3011 ( .A(ein[40]), .B(ein[39]), .Z(n2354) );
  XOR U3012 ( .A(ein[408]), .B(n2355), .Z(ereg_next[409]) );
  AND U3013 ( .A(mul_pow), .B(n2356), .Z(n2355) );
  XOR U3014 ( .A(ein[409]), .B(ein[408]), .Z(n2356) );
  XOR U3015 ( .A(ein[407]), .B(n2357), .Z(ereg_next[408]) );
  AND U3016 ( .A(mul_pow), .B(n2358), .Z(n2357) );
  XOR U3017 ( .A(ein[408]), .B(ein[407]), .Z(n2358) );
  XOR U3018 ( .A(ein[406]), .B(n2359), .Z(ereg_next[407]) );
  AND U3019 ( .A(mul_pow), .B(n2360), .Z(n2359) );
  XOR U3020 ( .A(ein[407]), .B(ein[406]), .Z(n2360) );
  XOR U3021 ( .A(ein[405]), .B(n2361), .Z(ereg_next[406]) );
  AND U3022 ( .A(mul_pow), .B(n2362), .Z(n2361) );
  XOR U3023 ( .A(ein[406]), .B(ein[405]), .Z(n2362) );
  XOR U3024 ( .A(ein[404]), .B(n2363), .Z(ereg_next[405]) );
  AND U3025 ( .A(mul_pow), .B(n2364), .Z(n2363) );
  XOR U3026 ( .A(ein[405]), .B(ein[404]), .Z(n2364) );
  XOR U3027 ( .A(ein[403]), .B(n2365), .Z(ereg_next[404]) );
  AND U3028 ( .A(mul_pow), .B(n2366), .Z(n2365) );
  XOR U3029 ( .A(ein[404]), .B(ein[403]), .Z(n2366) );
  XOR U3030 ( .A(ein[402]), .B(n2367), .Z(ereg_next[403]) );
  AND U3031 ( .A(mul_pow), .B(n2368), .Z(n2367) );
  XOR U3032 ( .A(ein[403]), .B(ein[402]), .Z(n2368) );
  XOR U3033 ( .A(ein[401]), .B(n2369), .Z(ereg_next[402]) );
  AND U3034 ( .A(mul_pow), .B(n2370), .Z(n2369) );
  XOR U3035 ( .A(ein[402]), .B(ein[401]), .Z(n2370) );
  XOR U3036 ( .A(ein[400]), .B(n2371), .Z(ereg_next[401]) );
  AND U3037 ( .A(mul_pow), .B(n2372), .Z(n2371) );
  XOR U3038 ( .A(ein[401]), .B(ein[400]), .Z(n2372) );
  XOR U3039 ( .A(ein[399]), .B(n2373), .Z(ereg_next[400]) );
  AND U3040 ( .A(mul_pow), .B(n2374), .Z(n2373) );
  XOR U3041 ( .A(ein[400]), .B(ein[399]), .Z(n2374) );
  XOR U3042 ( .A(ein[2]), .B(n2375), .Z(ereg_next[3]) );
  AND U3043 ( .A(mul_pow), .B(n2376), .Z(n2375) );
  XOR U3044 ( .A(ein[3]), .B(ein[2]), .Z(n2376) );
  XOR U3045 ( .A(ein[38]), .B(n2377), .Z(ereg_next[39]) );
  AND U3046 ( .A(mul_pow), .B(n2378), .Z(n2377) );
  XOR U3047 ( .A(ein[39]), .B(ein[38]), .Z(n2378) );
  XOR U3048 ( .A(ein[398]), .B(n2379), .Z(ereg_next[399]) );
  AND U3049 ( .A(mul_pow), .B(n2380), .Z(n2379) );
  XOR U3050 ( .A(ein[399]), .B(ein[398]), .Z(n2380) );
  XOR U3051 ( .A(ein[397]), .B(n2381), .Z(ereg_next[398]) );
  AND U3052 ( .A(mul_pow), .B(n2382), .Z(n2381) );
  XOR U3053 ( .A(ein[398]), .B(ein[397]), .Z(n2382) );
  XOR U3054 ( .A(ein[396]), .B(n2383), .Z(ereg_next[397]) );
  AND U3055 ( .A(mul_pow), .B(n2384), .Z(n2383) );
  XOR U3056 ( .A(ein[397]), .B(ein[396]), .Z(n2384) );
  XOR U3057 ( .A(ein[395]), .B(n2385), .Z(ereg_next[396]) );
  AND U3058 ( .A(mul_pow), .B(n2386), .Z(n2385) );
  XOR U3059 ( .A(ein[396]), .B(ein[395]), .Z(n2386) );
  XOR U3060 ( .A(ein[394]), .B(n2387), .Z(ereg_next[395]) );
  AND U3061 ( .A(mul_pow), .B(n2388), .Z(n2387) );
  XOR U3062 ( .A(ein[395]), .B(ein[394]), .Z(n2388) );
  XOR U3063 ( .A(ein[393]), .B(n2389), .Z(ereg_next[394]) );
  AND U3064 ( .A(mul_pow), .B(n2390), .Z(n2389) );
  XOR U3065 ( .A(ein[394]), .B(ein[393]), .Z(n2390) );
  XOR U3066 ( .A(ein[392]), .B(n2391), .Z(ereg_next[393]) );
  AND U3067 ( .A(mul_pow), .B(n2392), .Z(n2391) );
  XOR U3068 ( .A(ein[393]), .B(ein[392]), .Z(n2392) );
  XOR U3069 ( .A(ein[391]), .B(n2393), .Z(ereg_next[392]) );
  AND U3070 ( .A(mul_pow), .B(n2394), .Z(n2393) );
  XOR U3071 ( .A(ein[392]), .B(ein[391]), .Z(n2394) );
  XOR U3072 ( .A(ein[390]), .B(n2395), .Z(ereg_next[391]) );
  AND U3073 ( .A(mul_pow), .B(n2396), .Z(n2395) );
  XOR U3074 ( .A(ein[391]), .B(ein[390]), .Z(n2396) );
  XOR U3075 ( .A(ein[389]), .B(n2397), .Z(ereg_next[390]) );
  AND U3076 ( .A(mul_pow), .B(n2398), .Z(n2397) );
  XOR U3077 ( .A(ein[390]), .B(ein[389]), .Z(n2398) );
  XOR U3078 ( .A(ein[37]), .B(n2399), .Z(ereg_next[38]) );
  AND U3079 ( .A(mul_pow), .B(n2400), .Z(n2399) );
  XOR U3080 ( .A(ein[38]), .B(ein[37]), .Z(n2400) );
  XOR U3081 ( .A(ein[388]), .B(n2401), .Z(ereg_next[389]) );
  AND U3082 ( .A(mul_pow), .B(n2402), .Z(n2401) );
  XOR U3083 ( .A(ein[389]), .B(ein[388]), .Z(n2402) );
  XOR U3084 ( .A(ein[387]), .B(n2403), .Z(ereg_next[388]) );
  AND U3085 ( .A(mul_pow), .B(n2404), .Z(n2403) );
  XOR U3086 ( .A(ein[388]), .B(ein[387]), .Z(n2404) );
  XOR U3087 ( .A(ein[386]), .B(n2405), .Z(ereg_next[387]) );
  AND U3088 ( .A(mul_pow), .B(n2406), .Z(n2405) );
  XOR U3089 ( .A(ein[387]), .B(ein[386]), .Z(n2406) );
  XOR U3090 ( .A(ein[385]), .B(n2407), .Z(ereg_next[386]) );
  AND U3091 ( .A(mul_pow), .B(n2408), .Z(n2407) );
  XOR U3092 ( .A(ein[386]), .B(ein[385]), .Z(n2408) );
  XOR U3093 ( .A(ein[384]), .B(n2409), .Z(ereg_next[385]) );
  AND U3094 ( .A(mul_pow), .B(n2410), .Z(n2409) );
  XOR U3095 ( .A(ein[385]), .B(ein[384]), .Z(n2410) );
  XOR U3096 ( .A(ein[383]), .B(n2411), .Z(ereg_next[384]) );
  AND U3097 ( .A(mul_pow), .B(n2412), .Z(n2411) );
  XOR U3098 ( .A(ein[384]), .B(ein[383]), .Z(n2412) );
  XOR U3099 ( .A(ein[382]), .B(n2413), .Z(ereg_next[383]) );
  AND U3100 ( .A(mul_pow), .B(n2414), .Z(n2413) );
  XOR U3101 ( .A(ein[383]), .B(ein[382]), .Z(n2414) );
  XOR U3102 ( .A(ein[381]), .B(n2415), .Z(ereg_next[382]) );
  AND U3103 ( .A(mul_pow), .B(n2416), .Z(n2415) );
  XOR U3104 ( .A(ein[382]), .B(ein[381]), .Z(n2416) );
  XOR U3105 ( .A(ein[380]), .B(n2417), .Z(ereg_next[381]) );
  AND U3106 ( .A(mul_pow), .B(n2418), .Z(n2417) );
  XOR U3107 ( .A(ein[381]), .B(ein[380]), .Z(n2418) );
  XOR U3108 ( .A(ein[379]), .B(n2419), .Z(ereg_next[380]) );
  AND U3109 ( .A(mul_pow), .B(n2420), .Z(n2419) );
  XOR U3110 ( .A(ein[380]), .B(ein[379]), .Z(n2420) );
  XOR U3111 ( .A(ein[36]), .B(n2421), .Z(ereg_next[37]) );
  AND U3112 ( .A(mul_pow), .B(n2422), .Z(n2421) );
  XOR U3113 ( .A(ein[37]), .B(ein[36]), .Z(n2422) );
  XOR U3114 ( .A(ein[378]), .B(n2423), .Z(ereg_next[379]) );
  AND U3115 ( .A(mul_pow), .B(n2424), .Z(n2423) );
  XOR U3116 ( .A(ein[379]), .B(ein[378]), .Z(n2424) );
  XOR U3117 ( .A(ein[377]), .B(n2425), .Z(ereg_next[378]) );
  AND U3118 ( .A(mul_pow), .B(n2426), .Z(n2425) );
  XOR U3119 ( .A(ein[378]), .B(ein[377]), .Z(n2426) );
  XOR U3120 ( .A(ein[376]), .B(n2427), .Z(ereg_next[377]) );
  AND U3121 ( .A(mul_pow), .B(n2428), .Z(n2427) );
  XOR U3122 ( .A(ein[377]), .B(ein[376]), .Z(n2428) );
  XOR U3123 ( .A(ein[375]), .B(n2429), .Z(ereg_next[376]) );
  AND U3124 ( .A(mul_pow), .B(n2430), .Z(n2429) );
  XOR U3125 ( .A(ein[376]), .B(ein[375]), .Z(n2430) );
  XOR U3126 ( .A(ein[374]), .B(n2431), .Z(ereg_next[375]) );
  AND U3127 ( .A(mul_pow), .B(n2432), .Z(n2431) );
  XOR U3128 ( .A(ein[375]), .B(ein[374]), .Z(n2432) );
  XOR U3129 ( .A(ein[373]), .B(n2433), .Z(ereg_next[374]) );
  AND U3130 ( .A(mul_pow), .B(n2434), .Z(n2433) );
  XOR U3131 ( .A(ein[374]), .B(ein[373]), .Z(n2434) );
  XOR U3132 ( .A(ein[372]), .B(n2435), .Z(ereg_next[373]) );
  AND U3133 ( .A(mul_pow), .B(n2436), .Z(n2435) );
  XOR U3134 ( .A(ein[373]), .B(ein[372]), .Z(n2436) );
  XOR U3135 ( .A(ein[371]), .B(n2437), .Z(ereg_next[372]) );
  AND U3136 ( .A(mul_pow), .B(n2438), .Z(n2437) );
  XOR U3137 ( .A(ein[372]), .B(ein[371]), .Z(n2438) );
  XOR U3138 ( .A(ein[370]), .B(n2439), .Z(ereg_next[371]) );
  AND U3139 ( .A(mul_pow), .B(n2440), .Z(n2439) );
  XOR U3140 ( .A(ein[371]), .B(ein[370]), .Z(n2440) );
  XOR U3141 ( .A(ein[369]), .B(n2441), .Z(ereg_next[370]) );
  AND U3142 ( .A(mul_pow), .B(n2442), .Z(n2441) );
  XOR U3143 ( .A(ein[370]), .B(ein[369]), .Z(n2442) );
  XOR U3144 ( .A(ein[35]), .B(n2443), .Z(ereg_next[36]) );
  AND U3145 ( .A(mul_pow), .B(n2444), .Z(n2443) );
  XOR U3146 ( .A(ein[36]), .B(ein[35]), .Z(n2444) );
  XOR U3147 ( .A(ein[368]), .B(n2445), .Z(ereg_next[369]) );
  AND U3148 ( .A(mul_pow), .B(n2446), .Z(n2445) );
  XOR U3149 ( .A(ein[369]), .B(ein[368]), .Z(n2446) );
  XOR U3150 ( .A(ein[367]), .B(n2447), .Z(ereg_next[368]) );
  AND U3151 ( .A(mul_pow), .B(n2448), .Z(n2447) );
  XOR U3152 ( .A(ein[368]), .B(ein[367]), .Z(n2448) );
  XOR U3153 ( .A(ein[366]), .B(n2449), .Z(ereg_next[367]) );
  AND U3154 ( .A(mul_pow), .B(n2450), .Z(n2449) );
  XOR U3155 ( .A(ein[367]), .B(ein[366]), .Z(n2450) );
  XOR U3156 ( .A(ein[365]), .B(n2451), .Z(ereg_next[366]) );
  AND U3157 ( .A(mul_pow), .B(n2452), .Z(n2451) );
  XOR U3158 ( .A(ein[366]), .B(ein[365]), .Z(n2452) );
  XOR U3159 ( .A(ein[364]), .B(n2453), .Z(ereg_next[365]) );
  AND U3160 ( .A(mul_pow), .B(n2454), .Z(n2453) );
  XOR U3161 ( .A(ein[365]), .B(ein[364]), .Z(n2454) );
  XOR U3162 ( .A(ein[363]), .B(n2455), .Z(ereg_next[364]) );
  AND U3163 ( .A(mul_pow), .B(n2456), .Z(n2455) );
  XOR U3164 ( .A(ein[364]), .B(ein[363]), .Z(n2456) );
  XOR U3165 ( .A(ein[362]), .B(n2457), .Z(ereg_next[363]) );
  AND U3166 ( .A(mul_pow), .B(n2458), .Z(n2457) );
  XOR U3167 ( .A(ein[363]), .B(ein[362]), .Z(n2458) );
  XOR U3168 ( .A(ein[361]), .B(n2459), .Z(ereg_next[362]) );
  AND U3169 ( .A(mul_pow), .B(n2460), .Z(n2459) );
  XOR U3170 ( .A(ein[362]), .B(ein[361]), .Z(n2460) );
  XOR U3171 ( .A(ein[360]), .B(n2461), .Z(ereg_next[361]) );
  AND U3172 ( .A(mul_pow), .B(n2462), .Z(n2461) );
  XOR U3173 ( .A(ein[361]), .B(ein[360]), .Z(n2462) );
  XOR U3174 ( .A(ein[359]), .B(n2463), .Z(ereg_next[360]) );
  AND U3175 ( .A(mul_pow), .B(n2464), .Z(n2463) );
  XOR U3176 ( .A(ein[360]), .B(ein[359]), .Z(n2464) );
  XOR U3177 ( .A(ein[34]), .B(n2465), .Z(ereg_next[35]) );
  AND U3178 ( .A(mul_pow), .B(n2466), .Z(n2465) );
  XOR U3179 ( .A(ein[35]), .B(ein[34]), .Z(n2466) );
  XOR U3180 ( .A(ein[358]), .B(n2467), .Z(ereg_next[359]) );
  AND U3181 ( .A(mul_pow), .B(n2468), .Z(n2467) );
  XOR U3182 ( .A(ein[359]), .B(ein[358]), .Z(n2468) );
  XOR U3183 ( .A(ein[357]), .B(n2469), .Z(ereg_next[358]) );
  AND U3184 ( .A(mul_pow), .B(n2470), .Z(n2469) );
  XOR U3185 ( .A(ein[358]), .B(ein[357]), .Z(n2470) );
  XOR U3186 ( .A(ein[356]), .B(n2471), .Z(ereg_next[357]) );
  AND U3187 ( .A(mul_pow), .B(n2472), .Z(n2471) );
  XOR U3188 ( .A(ein[357]), .B(ein[356]), .Z(n2472) );
  XOR U3189 ( .A(ein[355]), .B(n2473), .Z(ereg_next[356]) );
  AND U3190 ( .A(mul_pow), .B(n2474), .Z(n2473) );
  XOR U3191 ( .A(ein[356]), .B(ein[355]), .Z(n2474) );
  XOR U3192 ( .A(ein[354]), .B(n2475), .Z(ereg_next[355]) );
  AND U3193 ( .A(mul_pow), .B(n2476), .Z(n2475) );
  XOR U3194 ( .A(ein[355]), .B(ein[354]), .Z(n2476) );
  XOR U3195 ( .A(ein[353]), .B(n2477), .Z(ereg_next[354]) );
  AND U3196 ( .A(mul_pow), .B(n2478), .Z(n2477) );
  XOR U3197 ( .A(ein[354]), .B(ein[353]), .Z(n2478) );
  XOR U3198 ( .A(ein[352]), .B(n2479), .Z(ereg_next[353]) );
  AND U3199 ( .A(mul_pow), .B(n2480), .Z(n2479) );
  XOR U3200 ( .A(ein[353]), .B(ein[352]), .Z(n2480) );
  XOR U3201 ( .A(ein[351]), .B(n2481), .Z(ereg_next[352]) );
  AND U3202 ( .A(mul_pow), .B(n2482), .Z(n2481) );
  XOR U3203 ( .A(ein[352]), .B(ein[351]), .Z(n2482) );
  XOR U3204 ( .A(ein[350]), .B(n2483), .Z(ereg_next[351]) );
  AND U3205 ( .A(mul_pow), .B(n2484), .Z(n2483) );
  XOR U3206 ( .A(ein[351]), .B(ein[350]), .Z(n2484) );
  XOR U3207 ( .A(ein[349]), .B(n2485), .Z(ereg_next[350]) );
  AND U3208 ( .A(mul_pow), .B(n2486), .Z(n2485) );
  XOR U3209 ( .A(ein[350]), .B(ein[349]), .Z(n2486) );
  XOR U3210 ( .A(ein[33]), .B(n2487), .Z(ereg_next[34]) );
  AND U3211 ( .A(mul_pow), .B(n2488), .Z(n2487) );
  XOR U3212 ( .A(ein[34]), .B(ein[33]), .Z(n2488) );
  XOR U3213 ( .A(ein[348]), .B(n2489), .Z(ereg_next[349]) );
  AND U3214 ( .A(mul_pow), .B(n2490), .Z(n2489) );
  XOR U3215 ( .A(ein[349]), .B(ein[348]), .Z(n2490) );
  XOR U3216 ( .A(ein[347]), .B(n2491), .Z(ereg_next[348]) );
  AND U3217 ( .A(mul_pow), .B(n2492), .Z(n2491) );
  XOR U3218 ( .A(ein[348]), .B(ein[347]), .Z(n2492) );
  XOR U3219 ( .A(ein[346]), .B(n2493), .Z(ereg_next[347]) );
  AND U3220 ( .A(mul_pow), .B(n2494), .Z(n2493) );
  XOR U3221 ( .A(ein[347]), .B(ein[346]), .Z(n2494) );
  XOR U3222 ( .A(ein[345]), .B(n2495), .Z(ereg_next[346]) );
  AND U3223 ( .A(mul_pow), .B(n2496), .Z(n2495) );
  XOR U3224 ( .A(ein[346]), .B(ein[345]), .Z(n2496) );
  XOR U3225 ( .A(ein[344]), .B(n2497), .Z(ereg_next[345]) );
  AND U3226 ( .A(mul_pow), .B(n2498), .Z(n2497) );
  XOR U3227 ( .A(ein[345]), .B(ein[344]), .Z(n2498) );
  XOR U3228 ( .A(ein[343]), .B(n2499), .Z(ereg_next[344]) );
  AND U3229 ( .A(mul_pow), .B(n2500), .Z(n2499) );
  XOR U3230 ( .A(ein[344]), .B(ein[343]), .Z(n2500) );
  XOR U3231 ( .A(ein[342]), .B(n2501), .Z(ereg_next[343]) );
  AND U3232 ( .A(mul_pow), .B(n2502), .Z(n2501) );
  XOR U3233 ( .A(ein[343]), .B(ein[342]), .Z(n2502) );
  XOR U3234 ( .A(ein[341]), .B(n2503), .Z(ereg_next[342]) );
  AND U3235 ( .A(mul_pow), .B(n2504), .Z(n2503) );
  XOR U3236 ( .A(ein[342]), .B(ein[341]), .Z(n2504) );
  XOR U3237 ( .A(ein[340]), .B(n2505), .Z(ereg_next[341]) );
  AND U3238 ( .A(mul_pow), .B(n2506), .Z(n2505) );
  XOR U3239 ( .A(ein[341]), .B(ein[340]), .Z(n2506) );
  XOR U3240 ( .A(ein[339]), .B(n2507), .Z(ereg_next[340]) );
  AND U3241 ( .A(mul_pow), .B(n2508), .Z(n2507) );
  XOR U3242 ( .A(ein[340]), .B(ein[339]), .Z(n2508) );
  XOR U3243 ( .A(ein[32]), .B(n2509), .Z(ereg_next[33]) );
  AND U3244 ( .A(mul_pow), .B(n2510), .Z(n2509) );
  XOR U3245 ( .A(ein[33]), .B(ein[32]), .Z(n2510) );
  XOR U3246 ( .A(ein[338]), .B(n2511), .Z(ereg_next[339]) );
  AND U3247 ( .A(mul_pow), .B(n2512), .Z(n2511) );
  XOR U3248 ( .A(ein[339]), .B(ein[338]), .Z(n2512) );
  XOR U3249 ( .A(ein[337]), .B(n2513), .Z(ereg_next[338]) );
  AND U3250 ( .A(mul_pow), .B(n2514), .Z(n2513) );
  XOR U3251 ( .A(ein[338]), .B(ein[337]), .Z(n2514) );
  XOR U3252 ( .A(ein[336]), .B(n2515), .Z(ereg_next[337]) );
  AND U3253 ( .A(mul_pow), .B(n2516), .Z(n2515) );
  XOR U3254 ( .A(ein[337]), .B(ein[336]), .Z(n2516) );
  XOR U3255 ( .A(ein[335]), .B(n2517), .Z(ereg_next[336]) );
  AND U3256 ( .A(mul_pow), .B(n2518), .Z(n2517) );
  XOR U3257 ( .A(ein[336]), .B(ein[335]), .Z(n2518) );
  XOR U3258 ( .A(ein[334]), .B(n2519), .Z(ereg_next[335]) );
  AND U3259 ( .A(mul_pow), .B(n2520), .Z(n2519) );
  XOR U3260 ( .A(ein[335]), .B(ein[334]), .Z(n2520) );
  XOR U3261 ( .A(ein[333]), .B(n2521), .Z(ereg_next[334]) );
  AND U3262 ( .A(mul_pow), .B(n2522), .Z(n2521) );
  XOR U3263 ( .A(ein[334]), .B(ein[333]), .Z(n2522) );
  XOR U3264 ( .A(ein[332]), .B(n2523), .Z(ereg_next[333]) );
  AND U3265 ( .A(mul_pow), .B(n2524), .Z(n2523) );
  XOR U3266 ( .A(ein[333]), .B(ein[332]), .Z(n2524) );
  XOR U3267 ( .A(ein[331]), .B(n2525), .Z(ereg_next[332]) );
  AND U3268 ( .A(mul_pow), .B(n2526), .Z(n2525) );
  XOR U3269 ( .A(ein[332]), .B(ein[331]), .Z(n2526) );
  XOR U3270 ( .A(ein[330]), .B(n2527), .Z(ereg_next[331]) );
  AND U3271 ( .A(mul_pow), .B(n2528), .Z(n2527) );
  XOR U3272 ( .A(ein[331]), .B(ein[330]), .Z(n2528) );
  XOR U3273 ( .A(ein[329]), .B(n2529), .Z(ereg_next[330]) );
  AND U3274 ( .A(mul_pow), .B(n2530), .Z(n2529) );
  XOR U3275 ( .A(ein[330]), .B(ein[329]), .Z(n2530) );
  XOR U3276 ( .A(ein[31]), .B(n2531), .Z(ereg_next[32]) );
  AND U3277 ( .A(mul_pow), .B(n2532), .Z(n2531) );
  XOR U3278 ( .A(ein[32]), .B(ein[31]), .Z(n2532) );
  XOR U3279 ( .A(ein[328]), .B(n2533), .Z(ereg_next[329]) );
  AND U3280 ( .A(mul_pow), .B(n2534), .Z(n2533) );
  XOR U3281 ( .A(ein[329]), .B(ein[328]), .Z(n2534) );
  XOR U3282 ( .A(ein[327]), .B(n2535), .Z(ereg_next[328]) );
  AND U3283 ( .A(mul_pow), .B(n2536), .Z(n2535) );
  XOR U3284 ( .A(ein[328]), .B(ein[327]), .Z(n2536) );
  XOR U3285 ( .A(ein[326]), .B(n2537), .Z(ereg_next[327]) );
  AND U3286 ( .A(mul_pow), .B(n2538), .Z(n2537) );
  XOR U3287 ( .A(ein[327]), .B(ein[326]), .Z(n2538) );
  XOR U3288 ( .A(ein[325]), .B(n2539), .Z(ereg_next[326]) );
  AND U3289 ( .A(mul_pow), .B(n2540), .Z(n2539) );
  XOR U3290 ( .A(ein[326]), .B(ein[325]), .Z(n2540) );
  XOR U3291 ( .A(ein[324]), .B(n2541), .Z(ereg_next[325]) );
  AND U3292 ( .A(mul_pow), .B(n2542), .Z(n2541) );
  XOR U3293 ( .A(ein[325]), .B(ein[324]), .Z(n2542) );
  XOR U3294 ( .A(ein[323]), .B(n2543), .Z(ereg_next[324]) );
  AND U3295 ( .A(mul_pow), .B(n2544), .Z(n2543) );
  XOR U3296 ( .A(ein[324]), .B(ein[323]), .Z(n2544) );
  XOR U3297 ( .A(ein[322]), .B(n2545), .Z(ereg_next[323]) );
  AND U3298 ( .A(mul_pow), .B(n2546), .Z(n2545) );
  XOR U3299 ( .A(ein[323]), .B(ein[322]), .Z(n2546) );
  XOR U3300 ( .A(ein[321]), .B(n2547), .Z(ereg_next[322]) );
  AND U3301 ( .A(mul_pow), .B(n2548), .Z(n2547) );
  XOR U3302 ( .A(ein[322]), .B(ein[321]), .Z(n2548) );
  XOR U3303 ( .A(ein[320]), .B(n2549), .Z(ereg_next[321]) );
  AND U3304 ( .A(mul_pow), .B(n2550), .Z(n2549) );
  XOR U3305 ( .A(ein[321]), .B(ein[320]), .Z(n2550) );
  XOR U3306 ( .A(ein[319]), .B(n2551), .Z(ereg_next[320]) );
  AND U3307 ( .A(mul_pow), .B(n2552), .Z(n2551) );
  XOR U3308 ( .A(ein[320]), .B(ein[319]), .Z(n2552) );
  XOR U3309 ( .A(ein[30]), .B(n2553), .Z(ereg_next[31]) );
  AND U3310 ( .A(mul_pow), .B(n2554), .Z(n2553) );
  XOR U3311 ( .A(ein[31]), .B(ein[30]), .Z(n2554) );
  XOR U3312 ( .A(ein[318]), .B(n2555), .Z(ereg_next[319]) );
  AND U3313 ( .A(mul_pow), .B(n2556), .Z(n2555) );
  XOR U3314 ( .A(ein[319]), .B(ein[318]), .Z(n2556) );
  XOR U3315 ( .A(ein[317]), .B(n2557), .Z(ereg_next[318]) );
  AND U3316 ( .A(mul_pow), .B(n2558), .Z(n2557) );
  XOR U3317 ( .A(ein[318]), .B(ein[317]), .Z(n2558) );
  XOR U3318 ( .A(ein[316]), .B(n2559), .Z(ereg_next[317]) );
  AND U3319 ( .A(mul_pow), .B(n2560), .Z(n2559) );
  XOR U3320 ( .A(ein[317]), .B(ein[316]), .Z(n2560) );
  XOR U3321 ( .A(ein[315]), .B(n2561), .Z(ereg_next[316]) );
  AND U3322 ( .A(mul_pow), .B(n2562), .Z(n2561) );
  XOR U3323 ( .A(ein[316]), .B(ein[315]), .Z(n2562) );
  XOR U3324 ( .A(ein[314]), .B(n2563), .Z(ereg_next[315]) );
  AND U3325 ( .A(mul_pow), .B(n2564), .Z(n2563) );
  XOR U3326 ( .A(ein[315]), .B(ein[314]), .Z(n2564) );
  XOR U3327 ( .A(ein[313]), .B(n2565), .Z(ereg_next[314]) );
  AND U3328 ( .A(mul_pow), .B(n2566), .Z(n2565) );
  XOR U3329 ( .A(ein[314]), .B(ein[313]), .Z(n2566) );
  XOR U3330 ( .A(ein[312]), .B(n2567), .Z(ereg_next[313]) );
  AND U3331 ( .A(mul_pow), .B(n2568), .Z(n2567) );
  XOR U3332 ( .A(ein[313]), .B(ein[312]), .Z(n2568) );
  XOR U3333 ( .A(ein[311]), .B(n2569), .Z(ereg_next[312]) );
  AND U3334 ( .A(mul_pow), .B(n2570), .Z(n2569) );
  XOR U3335 ( .A(ein[312]), .B(ein[311]), .Z(n2570) );
  XOR U3336 ( .A(ein[310]), .B(n2571), .Z(ereg_next[311]) );
  AND U3337 ( .A(mul_pow), .B(n2572), .Z(n2571) );
  XOR U3338 ( .A(ein[311]), .B(ein[310]), .Z(n2572) );
  XOR U3339 ( .A(ein[309]), .B(n2573), .Z(ereg_next[310]) );
  AND U3340 ( .A(mul_pow), .B(n2574), .Z(n2573) );
  XOR U3341 ( .A(ein[310]), .B(ein[309]), .Z(n2574) );
  XOR U3342 ( .A(ein[29]), .B(n2575), .Z(ereg_next[30]) );
  AND U3343 ( .A(mul_pow), .B(n2576), .Z(n2575) );
  XOR U3344 ( .A(ein[30]), .B(ein[29]), .Z(n2576) );
  XOR U3345 ( .A(ein[308]), .B(n2577), .Z(ereg_next[309]) );
  AND U3346 ( .A(mul_pow), .B(n2578), .Z(n2577) );
  XOR U3347 ( .A(ein[309]), .B(ein[308]), .Z(n2578) );
  XOR U3348 ( .A(ein[307]), .B(n2579), .Z(ereg_next[308]) );
  AND U3349 ( .A(mul_pow), .B(n2580), .Z(n2579) );
  XOR U3350 ( .A(ein[308]), .B(ein[307]), .Z(n2580) );
  XOR U3351 ( .A(ein[306]), .B(n2581), .Z(ereg_next[307]) );
  AND U3352 ( .A(mul_pow), .B(n2582), .Z(n2581) );
  XOR U3353 ( .A(ein[307]), .B(ein[306]), .Z(n2582) );
  XOR U3354 ( .A(ein[305]), .B(n2583), .Z(ereg_next[306]) );
  AND U3355 ( .A(mul_pow), .B(n2584), .Z(n2583) );
  XOR U3356 ( .A(ein[306]), .B(ein[305]), .Z(n2584) );
  XOR U3357 ( .A(ein[304]), .B(n2585), .Z(ereg_next[305]) );
  AND U3358 ( .A(mul_pow), .B(n2586), .Z(n2585) );
  XOR U3359 ( .A(ein[305]), .B(ein[304]), .Z(n2586) );
  XOR U3360 ( .A(ein[303]), .B(n2587), .Z(ereg_next[304]) );
  AND U3361 ( .A(mul_pow), .B(n2588), .Z(n2587) );
  XOR U3362 ( .A(ein[304]), .B(ein[303]), .Z(n2588) );
  XOR U3363 ( .A(ein[302]), .B(n2589), .Z(ereg_next[303]) );
  AND U3364 ( .A(mul_pow), .B(n2590), .Z(n2589) );
  XOR U3365 ( .A(ein[303]), .B(ein[302]), .Z(n2590) );
  XOR U3366 ( .A(ein[301]), .B(n2591), .Z(ereg_next[302]) );
  AND U3367 ( .A(mul_pow), .B(n2592), .Z(n2591) );
  XOR U3368 ( .A(ein[302]), .B(ein[301]), .Z(n2592) );
  XOR U3369 ( .A(ein[300]), .B(n2593), .Z(ereg_next[301]) );
  AND U3370 ( .A(mul_pow), .B(n2594), .Z(n2593) );
  XOR U3371 ( .A(ein[301]), .B(ein[300]), .Z(n2594) );
  XOR U3372 ( .A(ein[299]), .B(n2595), .Z(ereg_next[300]) );
  AND U3373 ( .A(mul_pow), .B(n2596), .Z(n2595) );
  XOR U3374 ( .A(ein[300]), .B(ein[299]), .Z(n2596) );
  XOR U3375 ( .A(ein[1]), .B(n2597), .Z(ereg_next[2]) );
  AND U3376 ( .A(mul_pow), .B(n2598), .Z(n2597) );
  XOR U3377 ( .A(ein[2]), .B(ein[1]), .Z(n2598) );
  XOR U3378 ( .A(ein[28]), .B(n2599), .Z(ereg_next[29]) );
  AND U3379 ( .A(mul_pow), .B(n2600), .Z(n2599) );
  XOR U3380 ( .A(ein[29]), .B(ein[28]), .Z(n2600) );
  XOR U3381 ( .A(ein[298]), .B(n2601), .Z(ereg_next[299]) );
  AND U3382 ( .A(mul_pow), .B(n2602), .Z(n2601) );
  XOR U3383 ( .A(ein[299]), .B(ein[298]), .Z(n2602) );
  XOR U3384 ( .A(ein[297]), .B(n2603), .Z(ereg_next[298]) );
  AND U3385 ( .A(mul_pow), .B(n2604), .Z(n2603) );
  XOR U3386 ( .A(ein[298]), .B(ein[297]), .Z(n2604) );
  XOR U3387 ( .A(ein[296]), .B(n2605), .Z(ereg_next[297]) );
  AND U3388 ( .A(mul_pow), .B(n2606), .Z(n2605) );
  XOR U3389 ( .A(ein[297]), .B(ein[296]), .Z(n2606) );
  XOR U3390 ( .A(ein[295]), .B(n2607), .Z(ereg_next[296]) );
  AND U3391 ( .A(mul_pow), .B(n2608), .Z(n2607) );
  XOR U3392 ( .A(ein[296]), .B(ein[295]), .Z(n2608) );
  XOR U3393 ( .A(ein[294]), .B(n2609), .Z(ereg_next[295]) );
  AND U3394 ( .A(mul_pow), .B(n2610), .Z(n2609) );
  XOR U3395 ( .A(ein[295]), .B(ein[294]), .Z(n2610) );
  XOR U3396 ( .A(ein[293]), .B(n2611), .Z(ereg_next[294]) );
  AND U3397 ( .A(mul_pow), .B(n2612), .Z(n2611) );
  XOR U3398 ( .A(ein[294]), .B(ein[293]), .Z(n2612) );
  XOR U3399 ( .A(ein[292]), .B(n2613), .Z(ereg_next[293]) );
  AND U3400 ( .A(mul_pow), .B(n2614), .Z(n2613) );
  XOR U3401 ( .A(ein[293]), .B(ein[292]), .Z(n2614) );
  XOR U3402 ( .A(ein[291]), .B(n2615), .Z(ereg_next[292]) );
  AND U3403 ( .A(mul_pow), .B(n2616), .Z(n2615) );
  XOR U3404 ( .A(ein[292]), .B(ein[291]), .Z(n2616) );
  XOR U3405 ( .A(ein[290]), .B(n2617), .Z(ereg_next[291]) );
  AND U3406 ( .A(mul_pow), .B(n2618), .Z(n2617) );
  XOR U3407 ( .A(ein[291]), .B(ein[290]), .Z(n2618) );
  XOR U3408 ( .A(ein[289]), .B(n2619), .Z(ereg_next[290]) );
  AND U3409 ( .A(mul_pow), .B(n2620), .Z(n2619) );
  XOR U3410 ( .A(ein[290]), .B(ein[289]), .Z(n2620) );
  XOR U3411 ( .A(ein[27]), .B(n2621), .Z(ereg_next[28]) );
  AND U3412 ( .A(mul_pow), .B(n2622), .Z(n2621) );
  XOR U3413 ( .A(ein[28]), .B(ein[27]), .Z(n2622) );
  XOR U3414 ( .A(ein[288]), .B(n2623), .Z(ereg_next[289]) );
  AND U3415 ( .A(mul_pow), .B(n2624), .Z(n2623) );
  XOR U3416 ( .A(ein[289]), .B(ein[288]), .Z(n2624) );
  XOR U3417 ( .A(ein[287]), .B(n2625), .Z(ereg_next[288]) );
  AND U3418 ( .A(mul_pow), .B(n2626), .Z(n2625) );
  XOR U3419 ( .A(ein[288]), .B(ein[287]), .Z(n2626) );
  XOR U3420 ( .A(ein[286]), .B(n2627), .Z(ereg_next[287]) );
  AND U3421 ( .A(mul_pow), .B(n2628), .Z(n2627) );
  XOR U3422 ( .A(ein[287]), .B(ein[286]), .Z(n2628) );
  XOR U3423 ( .A(ein[285]), .B(n2629), .Z(ereg_next[286]) );
  AND U3424 ( .A(mul_pow), .B(n2630), .Z(n2629) );
  XOR U3425 ( .A(ein[286]), .B(ein[285]), .Z(n2630) );
  XOR U3426 ( .A(ein[284]), .B(n2631), .Z(ereg_next[285]) );
  AND U3427 ( .A(mul_pow), .B(n2632), .Z(n2631) );
  XOR U3428 ( .A(ein[285]), .B(ein[284]), .Z(n2632) );
  XOR U3429 ( .A(ein[283]), .B(n2633), .Z(ereg_next[284]) );
  AND U3430 ( .A(mul_pow), .B(n2634), .Z(n2633) );
  XOR U3431 ( .A(ein[284]), .B(ein[283]), .Z(n2634) );
  XOR U3432 ( .A(ein[282]), .B(n2635), .Z(ereg_next[283]) );
  AND U3433 ( .A(mul_pow), .B(n2636), .Z(n2635) );
  XOR U3434 ( .A(ein[283]), .B(ein[282]), .Z(n2636) );
  XOR U3435 ( .A(ein[281]), .B(n2637), .Z(ereg_next[282]) );
  AND U3436 ( .A(mul_pow), .B(n2638), .Z(n2637) );
  XOR U3437 ( .A(ein[282]), .B(ein[281]), .Z(n2638) );
  XOR U3438 ( .A(ein[280]), .B(n2639), .Z(ereg_next[281]) );
  AND U3439 ( .A(mul_pow), .B(n2640), .Z(n2639) );
  XOR U3440 ( .A(ein[281]), .B(ein[280]), .Z(n2640) );
  XOR U3441 ( .A(ein[279]), .B(n2641), .Z(ereg_next[280]) );
  AND U3442 ( .A(mul_pow), .B(n2642), .Z(n2641) );
  XOR U3443 ( .A(ein[280]), .B(ein[279]), .Z(n2642) );
  XOR U3444 ( .A(ein[26]), .B(n2643), .Z(ereg_next[27]) );
  AND U3445 ( .A(mul_pow), .B(n2644), .Z(n2643) );
  XOR U3446 ( .A(ein[27]), .B(ein[26]), .Z(n2644) );
  XOR U3447 ( .A(ein[278]), .B(n2645), .Z(ereg_next[279]) );
  AND U3448 ( .A(mul_pow), .B(n2646), .Z(n2645) );
  XOR U3449 ( .A(ein[279]), .B(ein[278]), .Z(n2646) );
  XOR U3450 ( .A(ein[277]), .B(n2647), .Z(ereg_next[278]) );
  AND U3451 ( .A(mul_pow), .B(n2648), .Z(n2647) );
  XOR U3452 ( .A(ein[278]), .B(ein[277]), .Z(n2648) );
  XOR U3453 ( .A(ein[276]), .B(n2649), .Z(ereg_next[277]) );
  AND U3454 ( .A(mul_pow), .B(n2650), .Z(n2649) );
  XOR U3455 ( .A(ein[277]), .B(ein[276]), .Z(n2650) );
  XOR U3456 ( .A(ein[275]), .B(n2651), .Z(ereg_next[276]) );
  AND U3457 ( .A(mul_pow), .B(n2652), .Z(n2651) );
  XOR U3458 ( .A(ein[276]), .B(ein[275]), .Z(n2652) );
  XOR U3459 ( .A(ein[274]), .B(n2653), .Z(ereg_next[275]) );
  AND U3460 ( .A(mul_pow), .B(n2654), .Z(n2653) );
  XOR U3461 ( .A(ein[275]), .B(ein[274]), .Z(n2654) );
  XOR U3462 ( .A(ein[273]), .B(n2655), .Z(ereg_next[274]) );
  AND U3463 ( .A(mul_pow), .B(n2656), .Z(n2655) );
  XOR U3464 ( .A(ein[274]), .B(ein[273]), .Z(n2656) );
  XOR U3465 ( .A(ein[272]), .B(n2657), .Z(ereg_next[273]) );
  AND U3466 ( .A(mul_pow), .B(n2658), .Z(n2657) );
  XOR U3467 ( .A(ein[273]), .B(ein[272]), .Z(n2658) );
  XOR U3468 ( .A(ein[271]), .B(n2659), .Z(ereg_next[272]) );
  AND U3469 ( .A(mul_pow), .B(n2660), .Z(n2659) );
  XOR U3470 ( .A(ein[272]), .B(ein[271]), .Z(n2660) );
  XOR U3471 ( .A(ein[270]), .B(n2661), .Z(ereg_next[271]) );
  AND U3472 ( .A(mul_pow), .B(n2662), .Z(n2661) );
  XOR U3473 ( .A(ein[271]), .B(ein[270]), .Z(n2662) );
  XOR U3474 ( .A(ein[269]), .B(n2663), .Z(ereg_next[270]) );
  AND U3475 ( .A(mul_pow), .B(n2664), .Z(n2663) );
  XOR U3476 ( .A(ein[270]), .B(ein[269]), .Z(n2664) );
  XOR U3477 ( .A(ein[25]), .B(n2665), .Z(ereg_next[26]) );
  AND U3478 ( .A(mul_pow), .B(n2666), .Z(n2665) );
  XOR U3479 ( .A(ein[26]), .B(ein[25]), .Z(n2666) );
  XOR U3480 ( .A(ein[268]), .B(n2667), .Z(ereg_next[269]) );
  AND U3481 ( .A(mul_pow), .B(n2668), .Z(n2667) );
  XOR U3482 ( .A(ein[269]), .B(ein[268]), .Z(n2668) );
  XOR U3483 ( .A(ein[267]), .B(n2669), .Z(ereg_next[268]) );
  AND U3484 ( .A(mul_pow), .B(n2670), .Z(n2669) );
  XOR U3485 ( .A(ein[268]), .B(ein[267]), .Z(n2670) );
  XOR U3486 ( .A(ein[266]), .B(n2671), .Z(ereg_next[267]) );
  AND U3487 ( .A(mul_pow), .B(n2672), .Z(n2671) );
  XOR U3488 ( .A(ein[267]), .B(ein[266]), .Z(n2672) );
  XOR U3489 ( .A(ein[265]), .B(n2673), .Z(ereg_next[266]) );
  AND U3490 ( .A(mul_pow), .B(n2674), .Z(n2673) );
  XOR U3491 ( .A(ein[266]), .B(ein[265]), .Z(n2674) );
  XOR U3492 ( .A(ein[264]), .B(n2675), .Z(ereg_next[265]) );
  AND U3493 ( .A(mul_pow), .B(n2676), .Z(n2675) );
  XOR U3494 ( .A(ein[265]), .B(ein[264]), .Z(n2676) );
  XOR U3495 ( .A(ein[263]), .B(n2677), .Z(ereg_next[264]) );
  AND U3496 ( .A(mul_pow), .B(n2678), .Z(n2677) );
  XOR U3497 ( .A(ein[264]), .B(ein[263]), .Z(n2678) );
  XOR U3498 ( .A(ein[262]), .B(n2679), .Z(ereg_next[263]) );
  AND U3499 ( .A(mul_pow), .B(n2680), .Z(n2679) );
  XOR U3500 ( .A(ein[263]), .B(ein[262]), .Z(n2680) );
  XOR U3501 ( .A(ein[261]), .B(n2681), .Z(ereg_next[262]) );
  AND U3502 ( .A(mul_pow), .B(n2682), .Z(n2681) );
  XOR U3503 ( .A(ein[262]), .B(ein[261]), .Z(n2682) );
  XOR U3504 ( .A(ein[260]), .B(n2683), .Z(ereg_next[261]) );
  AND U3505 ( .A(mul_pow), .B(n2684), .Z(n2683) );
  XOR U3506 ( .A(ein[261]), .B(ein[260]), .Z(n2684) );
  XOR U3507 ( .A(ein[259]), .B(n2685), .Z(ereg_next[260]) );
  AND U3508 ( .A(mul_pow), .B(n2686), .Z(n2685) );
  XOR U3509 ( .A(ein[260]), .B(ein[259]), .Z(n2686) );
  XOR U3510 ( .A(ein[24]), .B(n2687), .Z(ereg_next[25]) );
  AND U3511 ( .A(mul_pow), .B(n2688), .Z(n2687) );
  XOR U3512 ( .A(ein[25]), .B(ein[24]), .Z(n2688) );
  XOR U3513 ( .A(ein[258]), .B(n2689), .Z(ereg_next[259]) );
  AND U3514 ( .A(mul_pow), .B(n2690), .Z(n2689) );
  XOR U3515 ( .A(ein[259]), .B(ein[258]), .Z(n2690) );
  XOR U3516 ( .A(ein[257]), .B(n2691), .Z(ereg_next[258]) );
  AND U3517 ( .A(mul_pow), .B(n2692), .Z(n2691) );
  XOR U3518 ( .A(ein[258]), .B(ein[257]), .Z(n2692) );
  XOR U3519 ( .A(ein[256]), .B(n2693), .Z(ereg_next[257]) );
  AND U3520 ( .A(mul_pow), .B(n2694), .Z(n2693) );
  XOR U3521 ( .A(ein[257]), .B(ein[256]), .Z(n2694) );
  XOR U3522 ( .A(ein[255]), .B(n2695), .Z(ereg_next[256]) );
  AND U3523 ( .A(mul_pow), .B(n2696), .Z(n2695) );
  XOR U3524 ( .A(ein[256]), .B(ein[255]), .Z(n2696) );
  XOR U3525 ( .A(ein[254]), .B(n2697), .Z(ereg_next[255]) );
  AND U3526 ( .A(mul_pow), .B(n2698), .Z(n2697) );
  XOR U3527 ( .A(ein[255]), .B(ein[254]), .Z(n2698) );
  XOR U3528 ( .A(ein[253]), .B(n2699), .Z(ereg_next[254]) );
  AND U3529 ( .A(mul_pow), .B(n2700), .Z(n2699) );
  XOR U3530 ( .A(ein[254]), .B(ein[253]), .Z(n2700) );
  XOR U3531 ( .A(ein[252]), .B(n2701), .Z(ereg_next[253]) );
  AND U3532 ( .A(mul_pow), .B(n2702), .Z(n2701) );
  XOR U3533 ( .A(ein[253]), .B(ein[252]), .Z(n2702) );
  XOR U3534 ( .A(ein[251]), .B(n2703), .Z(ereg_next[252]) );
  AND U3535 ( .A(mul_pow), .B(n2704), .Z(n2703) );
  XOR U3536 ( .A(ein[252]), .B(ein[251]), .Z(n2704) );
  XOR U3537 ( .A(ein[250]), .B(n2705), .Z(ereg_next[251]) );
  AND U3538 ( .A(mul_pow), .B(n2706), .Z(n2705) );
  XOR U3539 ( .A(ein[251]), .B(ein[250]), .Z(n2706) );
  XOR U3540 ( .A(ein[249]), .B(n2707), .Z(ereg_next[250]) );
  AND U3541 ( .A(mul_pow), .B(n2708), .Z(n2707) );
  XOR U3542 ( .A(ein[250]), .B(ein[249]), .Z(n2708) );
  XOR U3543 ( .A(ein[23]), .B(n2709), .Z(ereg_next[24]) );
  AND U3544 ( .A(mul_pow), .B(n2710), .Z(n2709) );
  XOR U3545 ( .A(ein[24]), .B(ein[23]), .Z(n2710) );
  XOR U3546 ( .A(ein[248]), .B(n2711), .Z(ereg_next[249]) );
  AND U3547 ( .A(mul_pow), .B(n2712), .Z(n2711) );
  XOR U3548 ( .A(ein[249]), .B(ein[248]), .Z(n2712) );
  XOR U3549 ( .A(ein[247]), .B(n2713), .Z(ereg_next[248]) );
  AND U3550 ( .A(mul_pow), .B(n2714), .Z(n2713) );
  XOR U3551 ( .A(ein[248]), .B(ein[247]), .Z(n2714) );
  XOR U3552 ( .A(ein[246]), .B(n2715), .Z(ereg_next[247]) );
  AND U3553 ( .A(mul_pow), .B(n2716), .Z(n2715) );
  XOR U3554 ( .A(ein[247]), .B(ein[246]), .Z(n2716) );
  XOR U3555 ( .A(ein[245]), .B(n2717), .Z(ereg_next[246]) );
  AND U3556 ( .A(mul_pow), .B(n2718), .Z(n2717) );
  XOR U3557 ( .A(ein[246]), .B(ein[245]), .Z(n2718) );
  XOR U3558 ( .A(ein[244]), .B(n2719), .Z(ereg_next[245]) );
  AND U3559 ( .A(mul_pow), .B(n2720), .Z(n2719) );
  XOR U3560 ( .A(ein[245]), .B(ein[244]), .Z(n2720) );
  XOR U3561 ( .A(ein[243]), .B(n2721), .Z(ereg_next[244]) );
  AND U3562 ( .A(mul_pow), .B(n2722), .Z(n2721) );
  XOR U3563 ( .A(ein[244]), .B(ein[243]), .Z(n2722) );
  XOR U3564 ( .A(ein[242]), .B(n2723), .Z(ereg_next[243]) );
  AND U3565 ( .A(mul_pow), .B(n2724), .Z(n2723) );
  XOR U3566 ( .A(ein[243]), .B(ein[242]), .Z(n2724) );
  XOR U3567 ( .A(ein[241]), .B(n2725), .Z(ereg_next[242]) );
  AND U3568 ( .A(mul_pow), .B(n2726), .Z(n2725) );
  XOR U3569 ( .A(ein[242]), .B(ein[241]), .Z(n2726) );
  XOR U3570 ( .A(ein[240]), .B(n2727), .Z(ereg_next[241]) );
  AND U3571 ( .A(mul_pow), .B(n2728), .Z(n2727) );
  XOR U3572 ( .A(ein[241]), .B(ein[240]), .Z(n2728) );
  XOR U3573 ( .A(ein[239]), .B(n2729), .Z(ereg_next[240]) );
  AND U3574 ( .A(mul_pow), .B(n2730), .Z(n2729) );
  XOR U3575 ( .A(ein[240]), .B(ein[239]), .Z(n2730) );
  XOR U3576 ( .A(ein[22]), .B(n2731), .Z(ereg_next[23]) );
  AND U3577 ( .A(mul_pow), .B(n2732), .Z(n2731) );
  XOR U3578 ( .A(ein[23]), .B(ein[22]), .Z(n2732) );
  XOR U3579 ( .A(ein[238]), .B(n2733), .Z(ereg_next[239]) );
  AND U3580 ( .A(mul_pow), .B(n2734), .Z(n2733) );
  XOR U3581 ( .A(ein[239]), .B(ein[238]), .Z(n2734) );
  XOR U3582 ( .A(ein[237]), .B(n2735), .Z(ereg_next[238]) );
  AND U3583 ( .A(mul_pow), .B(n2736), .Z(n2735) );
  XOR U3584 ( .A(ein[238]), .B(ein[237]), .Z(n2736) );
  XOR U3585 ( .A(ein[236]), .B(n2737), .Z(ereg_next[237]) );
  AND U3586 ( .A(mul_pow), .B(n2738), .Z(n2737) );
  XOR U3587 ( .A(ein[237]), .B(ein[236]), .Z(n2738) );
  XOR U3588 ( .A(ein[235]), .B(n2739), .Z(ereg_next[236]) );
  AND U3589 ( .A(mul_pow), .B(n2740), .Z(n2739) );
  XOR U3590 ( .A(ein[236]), .B(ein[235]), .Z(n2740) );
  XOR U3591 ( .A(ein[234]), .B(n2741), .Z(ereg_next[235]) );
  AND U3592 ( .A(mul_pow), .B(n2742), .Z(n2741) );
  XOR U3593 ( .A(ein[235]), .B(ein[234]), .Z(n2742) );
  XOR U3594 ( .A(ein[233]), .B(n2743), .Z(ereg_next[234]) );
  AND U3595 ( .A(mul_pow), .B(n2744), .Z(n2743) );
  XOR U3596 ( .A(ein[234]), .B(ein[233]), .Z(n2744) );
  XOR U3597 ( .A(ein[232]), .B(n2745), .Z(ereg_next[233]) );
  AND U3598 ( .A(mul_pow), .B(n2746), .Z(n2745) );
  XOR U3599 ( .A(ein[233]), .B(ein[232]), .Z(n2746) );
  XOR U3600 ( .A(ein[231]), .B(n2747), .Z(ereg_next[232]) );
  AND U3601 ( .A(mul_pow), .B(n2748), .Z(n2747) );
  XOR U3602 ( .A(ein[232]), .B(ein[231]), .Z(n2748) );
  XOR U3603 ( .A(ein[230]), .B(n2749), .Z(ereg_next[231]) );
  AND U3604 ( .A(mul_pow), .B(n2750), .Z(n2749) );
  XOR U3605 ( .A(ein[231]), .B(ein[230]), .Z(n2750) );
  XOR U3606 ( .A(ein[229]), .B(n2751), .Z(ereg_next[230]) );
  AND U3607 ( .A(mul_pow), .B(n2752), .Z(n2751) );
  XOR U3608 ( .A(ein[230]), .B(ein[229]), .Z(n2752) );
  XOR U3609 ( .A(ein[21]), .B(n2753), .Z(ereg_next[22]) );
  AND U3610 ( .A(mul_pow), .B(n2754), .Z(n2753) );
  XOR U3611 ( .A(ein[22]), .B(ein[21]), .Z(n2754) );
  XOR U3612 ( .A(ein[228]), .B(n2755), .Z(ereg_next[229]) );
  AND U3613 ( .A(mul_pow), .B(n2756), .Z(n2755) );
  XOR U3614 ( .A(ein[229]), .B(ein[228]), .Z(n2756) );
  XOR U3615 ( .A(ein[227]), .B(n2757), .Z(ereg_next[228]) );
  AND U3616 ( .A(mul_pow), .B(n2758), .Z(n2757) );
  XOR U3617 ( .A(ein[228]), .B(ein[227]), .Z(n2758) );
  XOR U3618 ( .A(ein[226]), .B(n2759), .Z(ereg_next[227]) );
  AND U3619 ( .A(mul_pow), .B(n2760), .Z(n2759) );
  XOR U3620 ( .A(ein[227]), .B(ein[226]), .Z(n2760) );
  XOR U3621 ( .A(ein[225]), .B(n2761), .Z(ereg_next[226]) );
  AND U3622 ( .A(mul_pow), .B(n2762), .Z(n2761) );
  XOR U3623 ( .A(ein[226]), .B(ein[225]), .Z(n2762) );
  XOR U3624 ( .A(ein[224]), .B(n2763), .Z(ereg_next[225]) );
  AND U3625 ( .A(mul_pow), .B(n2764), .Z(n2763) );
  XOR U3626 ( .A(ein[225]), .B(ein[224]), .Z(n2764) );
  XOR U3627 ( .A(ein[223]), .B(n2765), .Z(ereg_next[224]) );
  AND U3628 ( .A(mul_pow), .B(n2766), .Z(n2765) );
  XOR U3629 ( .A(ein[224]), .B(ein[223]), .Z(n2766) );
  XOR U3630 ( .A(ein[222]), .B(n2767), .Z(ereg_next[223]) );
  AND U3631 ( .A(mul_pow), .B(n2768), .Z(n2767) );
  XOR U3632 ( .A(ein[223]), .B(ein[222]), .Z(n2768) );
  XOR U3633 ( .A(ein[221]), .B(n2769), .Z(ereg_next[222]) );
  AND U3634 ( .A(mul_pow), .B(n2770), .Z(n2769) );
  XOR U3635 ( .A(ein[222]), .B(ein[221]), .Z(n2770) );
  XOR U3636 ( .A(ein[220]), .B(n2771), .Z(ereg_next[221]) );
  AND U3637 ( .A(mul_pow), .B(n2772), .Z(n2771) );
  XOR U3638 ( .A(ein[221]), .B(ein[220]), .Z(n2772) );
  XOR U3639 ( .A(ein[219]), .B(n2773), .Z(ereg_next[220]) );
  AND U3640 ( .A(mul_pow), .B(n2774), .Z(n2773) );
  XOR U3641 ( .A(ein[220]), .B(ein[219]), .Z(n2774) );
  XOR U3642 ( .A(ein[20]), .B(n2775), .Z(ereg_next[21]) );
  AND U3643 ( .A(mul_pow), .B(n2776), .Z(n2775) );
  XOR U3644 ( .A(ein[21]), .B(ein[20]), .Z(n2776) );
  XOR U3645 ( .A(ein[218]), .B(n2777), .Z(ereg_next[219]) );
  AND U3646 ( .A(mul_pow), .B(n2778), .Z(n2777) );
  XOR U3647 ( .A(ein[219]), .B(ein[218]), .Z(n2778) );
  XOR U3648 ( .A(ein[217]), .B(n2779), .Z(ereg_next[218]) );
  AND U3649 ( .A(mul_pow), .B(n2780), .Z(n2779) );
  XOR U3650 ( .A(ein[218]), .B(ein[217]), .Z(n2780) );
  XOR U3651 ( .A(ein[216]), .B(n2781), .Z(ereg_next[217]) );
  AND U3652 ( .A(mul_pow), .B(n2782), .Z(n2781) );
  XOR U3653 ( .A(ein[217]), .B(ein[216]), .Z(n2782) );
  XOR U3654 ( .A(ein[215]), .B(n2783), .Z(ereg_next[216]) );
  AND U3655 ( .A(mul_pow), .B(n2784), .Z(n2783) );
  XOR U3656 ( .A(ein[216]), .B(ein[215]), .Z(n2784) );
  XOR U3657 ( .A(ein[214]), .B(n2785), .Z(ereg_next[215]) );
  AND U3658 ( .A(mul_pow), .B(n2786), .Z(n2785) );
  XOR U3659 ( .A(ein[215]), .B(ein[214]), .Z(n2786) );
  XOR U3660 ( .A(ein[213]), .B(n2787), .Z(ereg_next[214]) );
  AND U3661 ( .A(mul_pow), .B(n2788), .Z(n2787) );
  XOR U3662 ( .A(ein[214]), .B(ein[213]), .Z(n2788) );
  XOR U3663 ( .A(ein[212]), .B(n2789), .Z(ereg_next[213]) );
  AND U3664 ( .A(mul_pow), .B(n2790), .Z(n2789) );
  XOR U3665 ( .A(ein[213]), .B(ein[212]), .Z(n2790) );
  XOR U3666 ( .A(ein[211]), .B(n2791), .Z(ereg_next[212]) );
  AND U3667 ( .A(mul_pow), .B(n2792), .Z(n2791) );
  XOR U3668 ( .A(ein[212]), .B(ein[211]), .Z(n2792) );
  XOR U3669 ( .A(ein[210]), .B(n2793), .Z(ereg_next[211]) );
  AND U3670 ( .A(mul_pow), .B(n2794), .Z(n2793) );
  XOR U3671 ( .A(ein[211]), .B(ein[210]), .Z(n2794) );
  XOR U3672 ( .A(ein[209]), .B(n2795), .Z(ereg_next[210]) );
  AND U3673 ( .A(mul_pow), .B(n2796), .Z(n2795) );
  XOR U3674 ( .A(ein[210]), .B(ein[209]), .Z(n2796) );
  XOR U3675 ( .A(ein[19]), .B(n2797), .Z(ereg_next[20]) );
  AND U3676 ( .A(mul_pow), .B(n2798), .Z(n2797) );
  XOR U3677 ( .A(ein[20]), .B(ein[19]), .Z(n2798) );
  XOR U3678 ( .A(ein[208]), .B(n2799), .Z(ereg_next[209]) );
  AND U3679 ( .A(mul_pow), .B(n2800), .Z(n2799) );
  XOR U3680 ( .A(ein[209]), .B(ein[208]), .Z(n2800) );
  XOR U3681 ( .A(ein[207]), .B(n2801), .Z(ereg_next[208]) );
  AND U3682 ( .A(mul_pow), .B(n2802), .Z(n2801) );
  XOR U3683 ( .A(ein[208]), .B(ein[207]), .Z(n2802) );
  XOR U3684 ( .A(ein[206]), .B(n2803), .Z(ereg_next[207]) );
  AND U3685 ( .A(mul_pow), .B(n2804), .Z(n2803) );
  XOR U3686 ( .A(ein[207]), .B(ein[206]), .Z(n2804) );
  XOR U3687 ( .A(ein[205]), .B(n2805), .Z(ereg_next[206]) );
  AND U3688 ( .A(mul_pow), .B(n2806), .Z(n2805) );
  XOR U3689 ( .A(ein[206]), .B(ein[205]), .Z(n2806) );
  XOR U3690 ( .A(ein[204]), .B(n2807), .Z(ereg_next[205]) );
  AND U3691 ( .A(mul_pow), .B(n2808), .Z(n2807) );
  XOR U3692 ( .A(ein[205]), .B(ein[204]), .Z(n2808) );
  XOR U3693 ( .A(ein[203]), .B(n2809), .Z(ereg_next[204]) );
  AND U3694 ( .A(mul_pow), .B(n2810), .Z(n2809) );
  XOR U3695 ( .A(ein[204]), .B(ein[203]), .Z(n2810) );
  XOR U3696 ( .A(ein[202]), .B(n2811), .Z(ereg_next[203]) );
  AND U3697 ( .A(mul_pow), .B(n2812), .Z(n2811) );
  XOR U3698 ( .A(ein[203]), .B(ein[202]), .Z(n2812) );
  XOR U3699 ( .A(ein[201]), .B(n2813), .Z(ereg_next[202]) );
  AND U3700 ( .A(mul_pow), .B(n2814), .Z(n2813) );
  XOR U3701 ( .A(ein[202]), .B(ein[201]), .Z(n2814) );
  XOR U3702 ( .A(ein[200]), .B(n2815), .Z(ereg_next[201]) );
  AND U3703 ( .A(mul_pow), .B(n2816), .Z(n2815) );
  XOR U3704 ( .A(ein[201]), .B(ein[200]), .Z(n2816) );
  XOR U3705 ( .A(ein[199]), .B(n2817), .Z(ereg_next[200]) );
  AND U3706 ( .A(mul_pow), .B(n2818), .Z(n2817) );
  XOR U3707 ( .A(ein[200]), .B(ein[199]), .Z(n2818) );
  XOR U3708 ( .A(ein[0]), .B(n2819), .Z(ereg_next[1]) );
  AND U3709 ( .A(mul_pow), .B(n2820), .Z(n2819) );
  XOR U3710 ( .A(ein[1]), .B(ein[0]), .Z(n2820) );
  XOR U3711 ( .A(ein[18]), .B(n2821), .Z(ereg_next[19]) );
  AND U3712 ( .A(mul_pow), .B(n2822), .Z(n2821) );
  XOR U3713 ( .A(ein[19]), .B(ein[18]), .Z(n2822) );
  XOR U3714 ( .A(ein[198]), .B(n2823), .Z(ereg_next[199]) );
  AND U3715 ( .A(mul_pow), .B(n2824), .Z(n2823) );
  XOR U3716 ( .A(ein[199]), .B(ein[198]), .Z(n2824) );
  XOR U3717 ( .A(ein[197]), .B(n2825), .Z(ereg_next[198]) );
  AND U3718 ( .A(mul_pow), .B(n2826), .Z(n2825) );
  XOR U3719 ( .A(ein[198]), .B(ein[197]), .Z(n2826) );
  XOR U3720 ( .A(ein[196]), .B(n2827), .Z(ereg_next[197]) );
  AND U3721 ( .A(mul_pow), .B(n2828), .Z(n2827) );
  XOR U3722 ( .A(ein[197]), .B(ein[196]), .Z(n2828) );
  XOR U3723 ( .A(ein[195]), .B(n2829), .Z(ereg_next[196]) );
  AND U3724 ( .A(mul_pow), .B(n2830), .Z(n2829) );
  XOR U3725 ( .A(ein[196]), .B(ein[195]), .Z(n2830) );
  XOR U3726 ( .A(ein[194]), .B(n2831), .Z(ereg_next[195]) );
  AND U3727 ( .A(mul_pow), .B(n2832), .Z(n2831) );
  XOR U3728 ( .A(ein[195]), .B(ein[194]), .Z(n2832) );
  XOR U3729 ( .A(ein[193]), .B(n2833), .Z(ereg_next[194]) );
  AND U3730 ( .A(mul_pow), .B(n2834), .Z(n2833) );
  XOR U3731 ( .A(ein[194]), .B(ein[193]), .Z(n2834) );
  XOR U3732 ( .A(ein[192]), .B(n2835), .Z(ereg_next[193]) );
  AND U3733 ( .A(mul_pow), .B(n2836), .Z(n2835) );
  XOR U3734 ( .A(ein[193]), .B(ein[192]), .Z(n2836) );
  XOR U3735 ( .A(ein[191]), .B(n2837), .Z(ereg_next[192]) );
  AND U3736 ( .A(mul_pow), .B(n2838), .Z(n2837) );
  XOR U3737 ( .A(ein[192]), .B(ein[191]), .Z(n2838) );
  XOR U3738 ( .A(ein[190]), .B(n2839), .Z(ereg_next[191]) );
  AND U3739 ( .A(mul_pow), .B(n2840), .Z(n2839) );
  XOR U3740 ( .A(ein[191]), .B(ein[190]), .Z(n2840) );
  XOR U3741 ( .A(ein[189]), .B(n2841), .Z(ereg_next[190]) );
  AND U3742 ( .A(mul_pow), .B(n2842), .Z(n2841) );
  XOR U3743 ( .A(ein[190]), .B(ein[189]), .Z(n2842) );
  XOR U3744 ( .A(ein[17]), .B(n2843), .Z(ereg_next[18]) );
  AND U3745 ( .A(mul_pow), .B(n2844), .Z(n2843) );
  XOR U3746 ( .A(ein[18]), .B(ein[17]), .Z(n2844) );
  XOR U3747 ( .A(ein[188]), .B(n2845), .Z(ereg_next[189]) );
  AND U3748 ( .A(mul_pow), .B(n2846), .Z(n2845) );
  XOR U3749 ( .A(ein[189]), .B(ein[188]), .Z(n2846) );
  XOR U3750 ( .A(ein[187]), .B(n2847), .Z(ereg_next[188]) );
  AND U3751 ( .A(mul_pow), .B(n2848), .Z(n2847) );
  XOR U3752 ( .A(ein[188]), .B(ein[187]), .Z(n2848) );
  XOR U3753 ( .A(ein[186]), .B(n2849), .Z(ereg_next[187]) );
  AND U3754 ( .A(mul_pow), .B(n2850), .Z(n2849) );
  XOR U3755 ( .A(ein[187]), .B(ein[186]), .Z(n2850) );
  XOR U3756 ( .A(ein[185]), .B(n2851), .Z(ereg_next[186]) );
  AND U3757 ( .A(mul_pow), .B(n2852), .Z(n2851) );
  XOR U3758 ( .A(ein[186]), .B(ein[185]), .Z(n2852) );
  XOR U3759 ( .A(ein[184]), .B(n2853), .Z(ereg_next[185]) );
  AND U3760 ( .A(mul_pow), .B(n2854), .Z(n2853) );
  XOR U3761 ( .A(ein[185]), .B(ein[184]), .Z(n2854) );
  XOR U3762 ( .A(ein[183]), .B(n2855), .Z(ereg_next[184]) );
  AND U3763 ( .A(mul_pow), .B(n2856), .Z(n2855) );
  XOR U3764 ( .A(ein[184]), .B(ein[183]), .Z(n2856) );
  XOR U3765 ( .A(ein[182]), .B(n2857), .Z(ereg_next[183]) );
  AND U3766 ( .A(mul_pow), .B(n2858), .Z(n2857) );
  XOR U3767 ( .A(ein[183]), .B(ein[182]), .Z(n2858) );
  XOR U3768 ( .A(ein[181]), .B(n2859), .Z(ereg_next[182]) );
  AND U3769 ( .A(mul_pow), .B(n2860), .Z(n2859) );
  XOR U3770 ( .A(ein[182]), .B(ein[181]), .Z(n2860) );
  XOR U3771 ( .A(ein[180]), .B(n2861), .Z(ereg_next[181]) );
  AND U3772 ( .A(mul_pow), .B(n2862), .Z(n2861) );
  XOR U3773 ( .A(ein[181]), .B(ein[180]), .Z(n2862) );
  XOR U3774 ( .A(ein[179]), .B(n2863), .Z(ereg_next[180]) );
  AND U3775 ( .A(mul_pow), .B(n2864), .Z(n2863) );
  XOR U3776 ( .A(ein[180]), .B(ein[179]), .Z(n2864) );
  XOR U3777 ( .A(ein[16]), .B(n2865), .Z(ereg_next[17]) );
  AND U3778 ( .A(mul_pow), .B(n2866), .Z(n2865) );
  XOR U3779 ( .A(ein[17]), .B(ein[16]), .Z(n2866) );
  XOR U3780 ( .A(ein[178]), .B(n2867), .Z(ereg_next[179]) );
  AND U3781 ( .A(mul_pow), .B(n2868), .Z(n2867) );
  XOR U3782 ( .A(ein[179]), .B(ein[178]), .Z(n2868) );
  XOR U3783 ( .A(ein[177]), .B(n2869), .Z(ereg_next[178]) );
  AND U3784 ( .A(mul_pow), .B(n2870), .Z(n2869) );
  XOR U3785 ( .A(ein[178]), .B(ein[177]), .Z(n2870) );
  XOR U3786 ( .A(ein[176]), .B(n2871), .Z(ereg_next[177]) );
  AND U3787 ( .A(mul_pow), .B(n2872), .Z(n2871) );
  XOR U3788 ( .A(ein[177]), .B(ein[176]), .Z(n2872) );
  XOR U3789 ( .A(ein[175]), .B(n2873), .Z(ereg_next[176]) );
  AND U3790 ( .A(mul_pow), .B(n2874), .Z(n2873) );
  XOR U3791 ( .A(ein[176]), .B(ein[175]), .Z(n2874) );
  XOR U3792 ( .A(ein[174]), .B(n2875), .Z(ereg_next[175]) );
  AND U3793 ( .A(mul_pow), .B(n2876), .Z(n2875) );
  XOR U3794 ( .A(ein[175]), .B(ein[174]), .Z(n2876) );
  XOR U3795 ( .A(ein[173]), .B(n2877), .Z(ereg_next[174]) );
  AND U3796 ( .A(mul_pow), .B(n2878), .Z(n2877) );
  XOR U3797 ( .A(ein[174]), .B(ein[173]), .Z(n2878) );
  XOR U3798 ( .A(ein[172]), .B(n2879), .Z(ereg_next[173]) );
  AND U3799 ( .A(mul_pow), .B(n2880), .Z(n2879) );
  XOR U3800 ( .A(ein[173]), .B(ein[172]), .Z(n2880) );
  XOR U3801 ( .A(ein[171]), .B(n2881), .Z(ereg_next[172]) );
  AND U3802 ( .A(mul_pow), .B(n2882), .Z(n2881) );
  XOR U3803 ( .A(ein[172]), .B(ein[171]), .Z(n2882) );
  XOR U3804 ( .A(ein[170]), .B(n2883), .Z(ereg_next[171]) );
  AND U3805 ( .A(mul_pow), .B(n2884), .Z(n2883) );
  XOR U3806 ( .A(ein[171]), .B(ein[170]), .Z(n2884) );
  XOR U3807 ( .A(ein[169]), .B(n2885), .Z(ereg_next[170]) );
  AND U3808 ( .A(mul_pow), .B(n2886), .Z(n2885) );
  XOR U3809 ( .A(ein[170]), .B(ein[169]), .Z(n2886) );
  XOR U3810 ( .A(ein[15]), .B(n2887), .Z(ereg_next[16]) );
  AND U3811 ( .A(mul_pow), .B(n2888), .Z(n2887) );
  XOR U3812 ( .A(ein[16]), .B(ein[15]), .Z(n2888) );
  XOR U3813 ( .A(ein[168]), .B(n2889), .Z(ereg_next[169]) );
  AND U3814 ( .A(mul_pow), .B(n2890), .Z(n2889) );
  XOR U3815 ( .A(ein[169]), .B(ein[168]), .Z(n2890) );
  XOR U3816 ( .A(ein[167]), .B(n2891), .Z(ereg_next[168]) );
  AND U3817 ( .A(mul_pow), .B(n2892), .Z(n2891) );
  XOR U3818 ( .A(ein[168]), .B(ein[167]), .Z(n2892) );
  XOR U3819 ( .A(ein[166]), .B(n2893), .Z(ereg_next[167]) );
  AND U3820 ( .A(mul_pow), .B(n2894), .Z(n2893) );
  XOR U3821 ( .A(ein[167]), .B(ein[166]), .Z(n2894) );
  XOR U3822 ( .A(ein[165]), .B(n2895), .Z(ereg_next[166]) );
  AND U3823 ( .A(mul_pow), .B(n2896), .Z(n2895) );
  XOR U3824 ( .A(ein[166]), .B(ein[165]), .Z(n2896) );
  XOR U3825 ( .A(ein[164]), .B(n2897), .Z(ereg_next[165]) );
  AND U3826 ( .A(mul_pow), .B(n2898), .Z(n2897) );
  XOR U3827 ( .A(ein[165]), .B(ein[164]), .Z(n2898) );
  XOR U3828 ( .A(ein[163]), .B(n2899), .Z(ereg_next[164]) );
  AND U3829 ( .A(mul_pow), .B(n2900), .Z(n2899) );
  XOR U3830 ( .A(ein[164]), .B(ein[163]), .Z(n2900) );
  XOR U3831 ( .A(ein[162]), .B(n2901), .Z(ereg_next[163]) );
  AND U3832 ( .A(mul_pow), .B(n2902), .Z(n2901) );
  XOR U3833 ( .A(ein[163]), .B(ein[162]), .Z(n2902) );
  XOR U3834 ( .A(ein[161]), .B(n2903), .Z(ereg_next[162]) );
  AND U3835 ( .A(mul_pow), .B(n2904), .Z(n2903) );
  XOR U3836 ( .A(ein[162]), .B(ein[161]), .Z(n2904) );
  XOR U3837 ( .A(ein[160]), .B(n2905), .Z(ereg_next[161]) );
  AND U3838 ( .A(mul_pow), .B(n2906), .Z(n2905) );
  XOR U3839 ( .A(ein[161]), .B(ein[160]), .Z(n2906) );
  XOR U3840 ( .A(ein[159]), .B(n2907), .Z(ereg_next[160]) );
  AND U3841 ( .A(mul_pow), .B(n2908), .Z(n2907) );
  XOR U3842 ( .A(ein[160]), .B(ein[159]), .Z(n2908) );
  XOR U3843 ( .A(ein[14]), .B(n2909), .Z(ereg_next[15]) );
  AND U3844 ( .A(mul_pow), .B(n2910), .Z(n2909) );
  XOR U3845 ( .A(ein[15]), .B(ein[14]), .Z(n2910) );
  XOR U3846 ( .A(ein[158]), .B(n2911), .Z(ereg_next[159]) );
  AND U3847 ( .A(mul_pow), .B(n2912), .Z(n2911) );
  XOR U3848 ( .A(ein[159]), .B(ein[158]), .Z(n2912) );
  XOR U3849 ( .A(ein[157]), .B(n2913), .Z(ereg_next[158]) );
  AND U3850 ( .A(mul_pow), .B(n2914), .Z(n2913) );
  XOR U3851 ( .A(ein[158]), .B(ein[157]), .Z(n2914) );
  XOR U3852 ( .A(ein[156]), .B(n2915), .Z(ereg_next[157]) );
  AND U3853 ( .A(mul_pow), .B(n2916), .Z(n2915) );
  XOR U3854 ( .A(ein[157]), .B(ein[156]), .Z(n2916) );
  XOR U3855 ( .A(ein[155]), .B(n2917), .Z(ereg_next[156]) );
  AND U3856 ( .A(mul_pow), .B(n2918), .Z(n2917) );
  XOR U3857 ( .A(ein[156]), .B(ein[155]), .Z(n2918) );
  XOR U3858 ( .A(ein[154]), .B(n2919), .Z(ereg_next[155]) );
  AND U3859 ( .A(mul_pow), .B(n2920), .Z(n2919) );
  XOR U3860 ( .A(ein[155]), .B(ein[154]), .Z(n2920) );
  XOR U3861 ( .A(ein[153]), .B(n2921), .Z(ereg_next[154]) );
  AND U3862 ( .A(mul_pow), .B(n2922), .Z(n2921) );
  XOR U3863 ( .A(ein[154]), .B(ein[153]), .Z(n2922) );
  XOR U3864 ( .A(ein[152]), .B(n2923), .Z(ereg_next[153]) );
  AND U3865 ( .A(mul_pow), .B(n2924), .Z(n2923) );
  XOR U3866 ( .A(ein[153]), .B(ein[152]), .Z(n2924) );
  XOR U3867 ( .A(ein[151]), .B(n2925), .Z(ereg_next[152]) );
  AND U3868 ( .A(mul_pow), .B(n2926), .Z(n2925) );
  XOR U3869 ( .A(ein[152]), .B(ein[151]), .Z(n2926) );
  XOR U3870 ( .A(ein[150]), .B(n2927), .Z(ereg_next[151]) );
  AND U3871 ( .A(mul_pow), .B(n2928), .Z(n2927) );
  XOR U3872 ( .A(ein[151]), .B(ein[150]), .Z(n2928) );
  XOR U3873 ( .A(ein[149]), .B(n2929), .Z(ereg_next[150]) );
  AND U3874 ( .A(mul_pow), .B(n2930), .Z(n2929) );
  XOR U3875 ( .A(ein[150]), .B(ein[149]), .Z(n2930) );
  XOR U3876 ( .A(ein[13]), .B(n2931), .Z(ereg_next[14]) );
  AND U3877 ( .A(mul_pow), .B(n2932), .Z(n2931) );
  XOR U3878 ( .A(ein[14]), .B(ein[13]), .Z(n2932) );
  XOR U3879 ( .A(ein[148]), .B(n2933), .Z(ereg_next[149]) );
  AND U3880 ( .A(mul_pow), .B(n2934), .Z(n2933) );
  XOR U3881 ( .A(ein[149]), .B(ein[148]), .Z(n2934) );
  XOR U3882 ( .A(ein[147]), .B(n2935), .Z(ereg_next[148]) );
  AND U3883 ( .A(mul_pow), .B(n2936), .Z(n2935) );
  XOR U3884 ( .A(ein[148]), .B(ein[147]), .Z(n2936) );
  XOR U3885 ( .A(ein[146]), .B(n2937), .Z(ereg_next[147]) );
  AND U3886 ( .A(mul_pow), .B(n2938), .Z(n2937) );
  XOR U3887 ( .A(ein[147]), .B(ein[146]), .Z(n2938) );
  XOR U3888 ( .A(ein[145]), .B(n2939), .Z(ereg_next[146]) );
  AND U3889 ( .A(mul_pow), .B(n2940), .Z(n2939) );
  XOR U3890 ( .A(ein[146]), .B(ein[145]), .Z(n2940) );
  XOR U3891 ( .A(ein[144]), .B(n2941), .Z(ereg_next[145]) );
  AND U3892 ( .A(mul_pow), .B(n2942), .Z(n2941) );
  XOR U3893 ( .A(ein[145]), .B(ein[144]), .Z(n2942) );
  XOR U3894 ( .A(ein[143]), .B(n2943), .Z(ereg_next[144]) );
  AND U3895 ( .A(mul_pow), .B(n2944), .Z(n2943) );
  XOR U3896 ( .A(ein[144]), .B(ein[143]), .Z(n2944) );
  XOR U3897 ( .A(ein[142]), .B(n2945), .Z(ereg_next[143]) );
  AND U3898 ( .A(mul_pow), .B(n2946), .Z(n2945) );
  XOR U3899 ( .A(ein[143]), .B(ein[142]), .Z(n2946) );
  XOR U3900 ( .A(ein[141]), .B(n2947), .Z(ereg_next[142]) );
  AND U3901 ( .A(mul_pow), .B(n2948), .Z(n2947) );
  XOR U3902 ( .A(ein[142]), .B(ein[141]), .Z(n2948) );
  XOR U3903 ( .A(ein[140]), .B(n2949), .Z(ereg_next[141]) );
  AND U3904 ( .A(mul_pow), .B(n2950), .Z(n2949) );
  XOR U3905 ( .A(ein[141]), .B(ein[140]), .Z(n2950) );
  XOR U3906 ( .A(ein[139]), .B(n2951), .Z(ereg_next[140]) );
  AND U3907 ( .A(mul_pow), .B(n2952), .Z(n2951) );
  XOR U3908 ( .A(ein[140]), .B(ein[139]), .Z(n2952) );
  XOR U3909 ( .A(ein[12]), .B(n2953), .Z(ereg_next[13]) );
  AND U3910 ( .A(mul_pow), .B(n2954), .Z(n2953) );
  XOR U3911 ( .A(ein[13]), .B(ein[12]), .Z(n2954) );
  XOR U3912 ( .A(ein[138]), .B(n2955), .Z(ereg_next[139]) );
  AND U3913 ( .A(mul_pow), .B(n2956), .Z(n2955) );
  XOR U3914 ( .A(ein[139]), .B(ein[138]), .Z(n2956) );
  XOR U3915 ( .A(ein[137]), .B(n2957), .Z(ereg_next[138]) );
  AND U3916 ( .A(mul_pow), .B(n2958), .Z(n2957) );
  XOR U3917 ( .A(ein[138]), .B(ein[137]), .Z(n2958) );
  XOR U3918 ( .A(ein[136]), .B(n2959), .Z(ereg_next[137]) );
  AND U3919 ( .A(mul_pow), .B(n2960), .Z(n2959) );
  XOR U3920 ( .A(ein[137]), .B(ein[136]), .Z(n2960) );
  XOR U3921 ( .A(ein[135]), .B(n2961), .Z(ereg_next[136]) );
  AND U3922 ( .A(mul_pow), .B(n2962), .Z(n2961) );
  XOR U3923 ( .A(ein[136]), .B(ein[135]), .Z(n2962) );
  XOR U3924 ( .A(ein[134]), .B(n2963), .Z(ereg_next[135]) );
  AND U3925 ( .A(mul_pow), .B(n2964), .Z(n2963) );
  XOR U3926 ( .A(ein[135]), .B(ein[134]), .Z(n2964) );
  XOR U3927 ( .A(ein[133]), .B(n2965), .Z(ereg_next[134]) );
  AND U3928 ( .A(mul_pow), .B(n2966), .Z(n2965) );
  XOR U3929 ( .A(ein[134]), .B(ein[133]), .Z(n2966) );
  XOR U3930 ( .A(ein[132]), .B(n2967), .Z(ereg_next[133]) );
  AND U3931 ( .A(mul_pow), .B(n2968), .Z(n2967) );
  XOR U3932 ( .A(ein[133]), .B(ein[132]), .Z(n2968) );
  XOR U3933 ( .A(ein[131]), .B(n2969), .Z(ereg_next[132]) );
  AND U3934 ( .A(mul_pow), .B(n2970), .Z(n2969) );
  XOR U3935 ( .A(ein[132]), .B(ein[131]), .Z(n2970) );
  XOR U3936 ( .A(ein[130]), .B(n2971), .Z(ereg_next[131]) );
  AND U3937 ( .A(mul_pow), .B(n2972), .Z(n2971) );
  XOR U3938 ( .A(ein[131]), .B(ein[130]), .Z(n2972) );
  XOR U3939 ( .A(ein[129]), .B(n2973), .Z(ereg_next[130]) );
  AND U3940 ( .A(mul_pow), .B(n2974), .Z(n2973) );
  XOR U3941 ( .A(ein[130]), .B(ein[129]), .Z(n2974) );
  XOR U3942 ( .A(ein[11]), .B(n2975), .Z(ereg_next[12]) );
  AND U3943 ( .A(mul_pow), .B(n2976), .Z(n2975) );
  XOR U3944 ( .A(ein[12]), .B(ein[11]), .Z(n2976) );
  XOR U3945 ( .A(ein[128]), .B(n2977), .Z(ereg_next[129]) );
  AND U3946 ( .A(mul_pow), .B(n2978), .Z(n2977) );
  XOR U3947 ( .A(ein[129]), .B(ein[128]), .Z(n2978) );
  XOR U3948 ( .A(ein[127]), .B(n2979), .Z(ereg_next[128]) );
  AND U3949 ( .A(mul_pow), .B(n2980), .Z(n2979) );
  XOR U3950 ( .A(ein[128]), .B(ein[127]), .Z(n2980) );
  XOR U3951 ( .A(ein[126]), .B(n2981), .Z(ereg_next[127]) );
  AND U3952 ( .A(mul_pow), .B(n2982), .Z(n2981) );
  XOR U3953 ( .A(ein[127]), .B(ein[126]), .Z(n2982) );
  XOR U3954 ( .A(ein[125]), .B(n2983), .Z(ereg_next[126]) );
  AND U3955 ( .A(mul_pow), .B(n2984), .Z(n2983) );
  XOR U3956 ( .A(ein[126]), .B(ein[125]), .Z(n2984) );
  XOR U3957 ( .A(ein[124]), .B(n2985), .Z(ereg_next[125]) );
  AND U3958 ( .A(mul_pow), .B(n2986), .Z(n2985) );
  XOR U3959 ( .A(ein[125]), .B(ein[124]), .Z(n2986) );
  XOR U3960 ( .A(ein[123]), .B(n2987), .Z(ereg_next[124]) );
  AND U3961 ( .A(mul_pow), .B(n2988), .Z(n2987) );
  XOR U3962 ( .A(ein[124]), .B(ein[123]), .Z(n2988) );
  XOR U3963 ( .A(ein[122]), .B(n2989), .Z(ereg_next[123]) );
  AND U3964 ( .A(mul_pow), .B(n2990), .Z(n2989) );
  XOR U3965 ( .A(ein[123]), .B(ein[122]), .Z(n2990) );
  XOR U3966 ( .A(ein[121]), .B(n2991), .Z(ereg_next[122]) );
  AND U3967 ( .A(mul_pow), .B(n2992), .Z(n2991) );
  XOR U3968 ( .A(ein[122]), .B(ein[121]), .Z(n2992) );
  XOR U3969 ( .A(ein[120]), .B(n2993), .Z(ereg_next[121]) );
  AND U3970 ( .A(mul_pow), .B(n2994), .Z(n2993) );
  XOR U3971 ( .A(ein[121]), .B(ein[120]), .Z(n2994) );
  XOR U3972 ( .A(ein[119]), .B(n2995), .Z(ereg_next[120]) );
  AND U3973 ( .A(mul_pow), .B(n2996), .Z(n2995) );
  XOR U3974 ( .A(ein[120]), .B(ein[119]), .Z(n2996) );
  XOR U3975 ( .A(ein[10]), .B(n2997), .Z(ereg_next[11]) );
  AND U3976 ( .A(mul_pow), .B(n2998), .Z(n2997) );
  XOR U3977 ( .A(ein[11]), .B(ein[10]), .Z(n2998) );
  XOR U3978 ( .A(ein[118]), .B(n2999), .Z(ereg_next[119]) );
  AND U3979 ( .A(mul_pow), .B(n3000), .Z(n2999) );
  XOR U3980 ( .A(ein[119]), .B(ein[118]), .Z(n3000) );
  XOR U3981 ( .A(ein[117]), .B(n3001), .Z(ereg_next[118]) );
  AND U3982 ( .A(mul_pow), .B(n3002), .Z(n3001) );
  XOR U3983 ( .A(ein[118]), .B(ein[117]), .Z(n3002) );
  XOR U3984 ( .A(ein[116]), .B(n3003), .Z(ereg_next[117]) );
  AND U3985 ( .A(mul_pow), .B(n3004), .Z(n3003) );
  XOR U3986 ( .A(ein[117]), .B(ein[116]), .Z(n3004) );
  XOR U3987 ( .A(ein[115]), .B(n3005), .Z(ereg_next[116]) );
  AND U3988 ( .A(mul_pow), .B(n3006), .Z(n3005) );
  XOR U3989 ( .A(ein[116]), .B(ein[115]), .Z(n3006) );
  XOR U3990 ( .A(ein[114]), .B(n3007), .Z(ereg_next[115]) );
  AND U3991 ( .A(mul_pow), .B(n3008), .Z(n3007) );
  XOR U3992 ( .A(ein[115]), .B(ein[114]), .Z(n3008) );
  XOR U3993 ( .A(ein[113]), .B(n3009), .Z(ereg_next[114]) );
  AND U3994 ( .A(mul_pow), .B(n3010), .Z(n3009) );
  XOR U3995 ( .A(ein[114]), .B(ein[113]), .Z(n3010) );
  XOR U3996 ( .A(ein[112]), .B(n3011), .Z(ereg_next[113]) );
  AND U3997 ( .A(mul_pow), .B(n3012), .Z(n3011) );
  XOR U3998 ( .A(ein[113]), .B(ein[112]), .Z(n3012) );
  XOR U3999 ( .A(ein[111]), .B(n3013), .Z(ereg_next[112]) );
  AND U4000 ( .A(mul_pow), .B(n3014), .Z(n3013) );
  XOR U4001 ( .A(ein[112]), .B(ein[111]), .Z(n3014) );
  XOR U4002 ( .A(ein[110]), .B(n3015), .Z(ereg_next[111]) );
  AND U4003 ( .A(mul_pow), .B(n3016), .Z(n3015) );
  XOR U4004 ( .A(ein[111]), .B(ein[110]), .Z(n3016) );
  XOR U4005 ( .A(ein[109]), .B(n3017), .Z(ereg_next[110]) );
  AND U4006 ( .A(mul_pow), .B(n3018), .Z(n3017) );
  XOR U4007 ( .A(ein[110]), .B(ein[109]), .Z(n3018) );
  XOR U4008 ( .A(ein[9]), .B(n3019), .Z(ereg_next[10]) );
  AND U4009 ( .A(mul_pow), .B(n3020), .Z(n3019) );
  XOR U4010 ( .A(ein[9]), .B(ein[10]), .Z(n3020) );
  XOR U4011 ( .A(ein[108]), .B(n3021), .Z(ereg_next[109]) );
  AND U4012 ( .A(mul_pow), .B(n3022), .Z(n3021) );
  XOR U4013 ( .A(ein[109]), .B(ein[108]), .Z(n3022) );
  XOR U4014 ( .A(ein[107]), .B(n3023), .Z(ereg_next[108]) );
  AND U4015 ( .A(mul_pow), .B(n3024), .Z(n3023) );
  XOR U4016 ( .A(ein[108]), .B(ein[107]), .Z(n3024) );
  XOR U4017 ( .A(ein[106]), .B(n3025), .Z(ereg_next[107]) );
  AND U4018 ( .A(mul_pow), .B(n3026), .Z(n3025) );
  XOR U4019 ( .A(ein[107]), .B(ein[106]), .Z(n3026) );
  XOR U4020 ( .A(ein[105]), .B(n3027), .Z(ereg_next[106]) );
  AND U4021 ( .A(mul_pow), .B(n3028), .Z(n3027) );
  XOR U4022 ( .A(ein[106]), .B(ein[105]), .Z(n3028) );
  XOR U4023 ( .A(ein[104]), .B(n3029), .Z(ereg_next[105]) );
  AND U4024 ( .A(mul_pow), .B(n3030), .Z(n3029) );
  XOR U4025 ( .A(ein[105]), .B(ein[104]), .Z(n3030) );
  XOR U4026 ( .A(ein[103]), .B(n3031), .Z(ereg_next[104]) );
  AND U4027 ( .A(mul_pow), .B(n3032), .Z(n3031) );
  XOR U4028 ( .A(ein[104]), .B(ein[103]), .Z(n3032) );
  XOR U4029 ( .A(ein[102]), .B(n3033), .Z(ereg_next[103]) );
  AND U4030 ( .A(mul_pow), .B(n3034), .Z(n3033) );
  XOR U4031 ( .A(ein[103]), .B(ein[102]), .Z(n3034) );
  XOR U4032 ( .A(ein[101]), .B(n3035), .Z(ereg_next[102]) );
  AND U4033 ( .A(mul_pow), .B(n3036), .Z(n3035) );
  XOR U4034 ( .A(ein[102]), .B(ein[101]), .Z(n3036) );
  XOR U4035 ( .A(ein[1022]), .B(n3037), .Z(ereg_next[1023]) );
  AND U4036 ( .A(mul_pow), .B(n3038), .Z(n3037) );
  XOR U4037 ( .A(ein[1023]), .B(ein[1022]), .Z(n3038) );
  XOR U4038 ( .A(ein[1021]), .B(n3039), .Z(ereg_next[1022]) );
  AND U4039 ( .A(mul_pow), .B(n3040), .Z(n3039) );
  XOR U4040 ( .A(ein[1022]), .B(ein[1021]), .Z(n3040) );
  XOR U4041 ( .A(ein[1020]), .B(n3041), .Z(ereg_next[1021]) );
  AND U4042 ( .A(mul_pow), .B(n3042), .Z(n3041) );
  XOR U4043 ( .A(ein[1021]), .B(ein[1020]), .Z(n3042) );
  XOR U4044 ( .A(ein[1019]), .B(n3043), .Z(ereg_next[1020]) );
  AND U4045 ( .A(mul_pow), .B(n3044), .Z(n3043) );
  XOR U4046 ( .A(ein[1020]), .B(ein[1019]), .Z(n3044) );
  XOR U4047 ( .A(ein[100]), .B(n3045), .Z(ereg_next[101]) );
  AND U4048 ( .A(mul_pow), .B(n3046), .Z(n3045) );
  XOR U4049 ( .A(ein[101]), .B(ein[100]), .Z(n3046) );
  XOR U4050 ( .A(ein[1018]), .B(n3047), .Z(ereg_next[1019]) );
  AND U4051 ( .A(mul_pow), .B(n3048), .Z(n3047) );
  XOR U4052 ( .A(ein[1019]), .B(ein[1018]), .Z(n3048) );
  XOR U4053 ( .A(ein[1017]), .B(n3049), .Z(ereg_next[1018]) );
  AND U4054 ( .A(mul_pow), .B(n3050), .Z(n3049) );
  XOR U4055 ( .A(ein[1018]), .B(ein[1017]), .Z(n3050) );
  XOR U4056 ( .A(ein[1016]), .B(n3051), .Z(ereg_next[1017]) );
  AND U4057 ( .A(mul_pow), .B(n3052), .Z(n3051) );
  XOR U4058 ( .A(ein[1017]), .B(ein[1016]), .Z(n3052) );
  XOR U4059 ( .A(ein[1015]), .B(n3053), .Z(ereg_next[1016]) );
  AND U4060 ( .A(mul_pow), .B(n3054), .Z(n3053) );
  XOR U4061 ( .A(ein[1016]), .B(ein[1015]), .Z(n3054) );
  XOR U4062 ( .A(ein[1014]), .B(n3055), .Z(ereg_next[1015]) );
  AND U4063 ( .A(mul_pow), .B(n3056), .Z(n3055) );
  XOR U4064 ( .A(ein[1015]), .B(ein[1014]), .Z(n3056) );
  XOR U4065 ( .A(ein[1013]), .B(n3057), .Z(ereg_next[1014]) );
  AND U4066 ( .A(mul_pow), .B(n3058), .Z(n3057) );
  XOR U4067 ( .A(ein[1014]), .B(ein[1013]), .Z(n3058) );
  XOR U4068 ( .A(ein[1012]), .B(n3059), .Z(ereg_next[1013]) );
  AND U4069 ( .A(mul_pow), .B(n3060), .Z(n3059) );
  XOR U4070 ( .A(ein[1013]), .B(ein[1012]), .Z(n3060) );
  XOR U4071 ( .A(ein[1011]), .B(n3061), .Z(ereg_next[1012]) );
  AND U4072 ( .A(mul_pow), .B(n3062), .Z(n3061) );
  XOR U4073 ( .A(ein[1012]), .B(ein[1011]), .Z(n3062) );
  XOR U4074 ( .A(ein[1010]), .B(n3063), .Z(ereg_next[1011]) );
  AND U4075 ( .A(mul_pow), .B(n3064), .Z(n3063) );
  XOR U4076 ( .A(ein[1011]), .B(ein[1010]), .Z(n3064) );
  XOR U4077 ( .A(ein[1009]), .B(n3065), .Z(ereg_next[1010]) );
  AND U4078 ( .A(mul_pow), .B(n3066), .Z(n3065) );
  XOR U4079 ( .A(ein[1010]), .B(ein[1009]), .Z(n3066) );
  XOR U4080 ( .A(ein[99]), .B(n3067), .Z(ereg_next[100]) );
  AND U4081 ( .A(mul_pow), .B(n3068), .Z(n3067) );
  XOR U4082 ( .A(ein[99]), .B(ein[100]), .Z(n3068) );
  XOR U4083 ( .A(ein[1008]), .B(n3069), .Z(ereg_next[1009]) );
  AND U4084 ( .A(mul_pow), .B(n3070), .Z(n3069) );
  XOR U4085 ( .A(ein[1009]), .B(ein[1008]), .Z(n3070) );
  XOR U4086 ( .A(ein[1007]), .B(n3071), .Z(ereg_next[1008]) );
  AND U4087 ( .A(mul_pow), .B(n3072), .Z(n3071) );
  XOR U4088 ( .A(ein[1008]), .B(ein[1007]), .Z(n3072) );
  XOR U4089 ( .A(ein[1006]), .B(n3073), .Z(ereg_next[1007]) );
  AND U4090 ( .A(mul_pow), .B(n3074), .Z(n3073) );
  XOR U4091 ( .A(ein[1007]), .B(ein[1006]), .Z(n3074) );
  XOR U4092 ( .A(ein[1005]), .B(n3075), .Z(ereg_next[1006]) );
  AND U4093 ( .A(mul_pow), .B(n3076), .Z(n3075) );
  XOR U4094 ( .A(ein[1006]), .B(ein[1005]), .Z(n3076) );
  XOR U4095 ( .A(ein[1004]), .B(n3077), .Z(ereg_next[1005]) );
  AND U4096 ( .A(mul_pow), .B(n3078), .Z(n3077) );
  XOR U4097 ( .A(ein[1005]), .B(ein[1004]), .Z(n3078) );
  XOR U4098 ( .A(ein[1003]), .B(n3079), .Z(ereg_next[1004]) );
  AND U4099 ( .A(mul_pow), .B(n3080), .Z(n3079) );
  XOR U4100 ( .A(ein[1004]), .B(ein[1003]), .Z(n3080) );
  XOR U4101 ( .A(ein[1002]), .B(n3081), .Z(ereg_next[1003]) );
  AND U4102 ( .A(mul_pow), .B(n3082), .Z(n3081) );
  XOR U4103 ( .A(ein[1003]), .B(ein[1002]), .Z(n3082) );
  XOR U4104 ( .A(ein[1001]), .B(n3083), .Z(ereg_next[1002]) );
  AND U4105 ( .A(mul_pow), .B(n3084), .Z(n3083) );
  XOR U4106 ( .A(ein[1002]), .B(ein[1001]), .Z(n3084) );
  XOR U4107 ( .A(ein[1000]), .B(n3085), .Z(ereg_next[1001]) );
  AND U4108 ( .A(mul_pow), .B(n3086), .Z(n3085) );
  XOR U4109 ( .A(ein[1001]), .B(ein[1000]), .Z(n3086) );
  XOR U4110 ( .A(ein[999]), .B(n3087), .Z(ereg_next[1000]) );
  AND U4111 ( .A(mul_pow), .B(n3088), .Z(n3087) );
  XOR U4112 ( .A(ein[999]), .B(ein[1000]), .Z(n3088) );
  AND U4113 ( .A(ein[0]), .B(mul_pow), .Z(ereg_next[0]) );
  XOR U4114 ( .A(n3089), .B(o[9]), .Z(creg_next[9]) );
  AND U4115 ( .A(n3090), .B(n3091), .Z(n3089) );
  XNOR U4116 ( .A(c[9]), .B(n3092), .Z(n3091) );
  IV U4117 ( .A(o[9]), .Z(n3092) );
  XNOR U4118 ( .A(n3093), .B(n3094), .Z(o[9]) );
  XOR U4119 ( .A(n3095), .B(o[99]), .Z(creg_next[99]) );
  AND U4120 ( .A(n3090), .B(n3096), .Z(n3095) );
  XNOR U4121 ( .A(c[99]), .B(n3097), .Z(n3096) );
  IV U4122 ( .A(o[99]), .Z(n3097) );
  XNOR U4123 ( .A(n3098), .B(n3099), .Z(o[99]) );
  XOR U4124 ( .A(n3100), .B(o[999]), .Z(creg_next[999]) );
  AND U4125 ( .A(n3090), .B(n3101), .Z(n3100) );
  XNOR U4126 ( .A(c[999]), .B(n3102), .Z(n3101) );
  IV U4127 ( .A(o[999]), .Z(n3102) );
  XNOR U4128 ( .A(n3103), .B(n3104), .Z(o[999]) );
  XOR U4129 ( .A(n3105), .B(o[998]), .Z(creg_next[998]) );
  AND U4130 ( .A(n3090), .B(n3106), .Z(n3105) );
  XNOR U4131 ( .A(c[998]), .B(n3107), .Z(n3106) );
  IV U4132 ( .A(o[998]), .Z(n3107) );
  XNOR U4133 ( .A(n3108), .B(n3109), .Z(o[998]) );
  XOR U4134 ( .A(n3110), .B(o[997]), .Z(creg_next[997]) );
  AND U4135 ( .A(n3090), .B(n3111), .Z(n3110) );
  XNOR U4136 ( .A(c[997]), .B(n3112), .Z(n3111) );
  IV U4137 ( .A(o[997]), .Z(n3112) );
  XNOR U4138 ( .A(n3113), .B(n3114), .Z(o[997]) );
  XOR U4139 ( .A(n3115), .B(o[996]), .Z(creg_next[996]) );
  AND U4140 ( .A(n3090), .B(n3116), .Z(n3115) );
  XNOR U4141 ( .A(c[996]), .B(n3117), .Z(n3116) );
  IV U4142 ( .A(o[996]), .Z(n3117) );
  XNOR U4143 ( .A(n3118), .B(n3119), .Z(o[996]) );
  XOR U4144 ( .A(n3120), .B(o[995]), .Z(creg_next[995]) );
  AND U4145 ( .A(n3090), .B(n3121), .Z(n3120) );
  XNOR U4146 ( .A(c[995]), .B(n3122), .Z(n3121) );
  IV U4147 ( .A(o[995]), .Z(n3122) );
  XNOR U4148 ( .A(n3123), .B(n3124), .Z(o[995]) );
  XOR U4149 ( .A(n3125), .B(o[994]), .Z(creg_next[994]) );
  AND U4150 ( .A(n3090), .B(n3126), .Z(n3125) );
  XNOR U4151 ( .A(c[994]), .B(n3127), .Z(n3126) );
  IV U4152 ( .A(o[994]), .Z(n3127) );
  XNOR U4153 ( .A(n3128), .B(n3129), .Z(o[994]) );
  XOR U4154 ( .A(n3130), .B(o[993]), .Z(creg_next[993]) );
  AND U4155 ( .A(n3090), .B(n3131), .Z(n3130) );
  XNOR U4156 ( .A(c[993]), .B(n3132), .Z(n3131) );
  IV U4157 ( .A(o[993]), .Z(n3132) );
  XNOR U4158 ( .A(n3133), .B(n3134), .Z(o[993]) );
  XOR U4159 ( .A(n3135), .B(o[992]), .Z(creg_next[992]) );
  AND U4160 ( .A(n3090), .B(n3136), .Z(n3135) );
  XNOR U4161 ( .A(c[992]), .B(n3137), .Z(n3136) );
  IV U4162 ( .A(o[992]), .Z(n3137) );
  XNOR U4163 ( .A(n3138), .B(n3139), .Z(o[992]) );
  XOR U4164 ( .A(n3140), .B(o[991]), .Z(creg_next[991]) );
  AND U4165 ( .A(n3090), .B(n3141), .Z(n3140) );
  XNOR U4166 ( .A(c[991]), .B(n3142), .Z(n3141) );
  IV U4167 ( .A(o[991]), .Z(n3142) );
  XNOR U4168 ( .A(n3143), .B(n3144), .Z(o[991]) );
  XOR U4169 ( .A(n3145), .B(o[990]), .Z(creg_next[990]) );
  AND U4170 ( .A(n3090), .B(n3146), .Z(n3145) );
  XNOR U4171 ( .A(c[990]), .B(n3147), .Z(n3146) );
  IV U4172 ( .A(o[990]), .Z(n3147) );
  XNOR U4173 ( .A(n3148), .B(n3149), .Z(o[990]) );
  XOR U4174 ( .A(n3150), .B(o[98]), .Z(creg_next[98]) );
  AND U4175 ( .A(n3090), .B(n3151), .Z(n3150) );
  XNOR U4176 ( .A(c[98]), .B(n3152), .Z(n3151) );
  IV U4177 ( .A(o[98]), .Z(n3152) );
  XNOR U4178 ( .A(n3153), .B(n3154), .Z(o[98]) );
  XOR U4179 ( .A(n3155), .B(o[989]), .Z(creg_next[989]) );
  AND U4180 ( .A(n3090), .B(n3156), .Z(n3155) );
  XNOR U4181 ( .A(c[989]), .B(n3157), .Z(n3156) );
  IV U4182 ( .A(o[989]), .Z(n3157) );
  XNOR U4183 ( .A(n3158), .B(n3159), .Z(o[989]) );
  XOR U4184 ( .A(n3160), .B(o[988]), .Z(creg_next[988]) );
  AND U4185 ( .A(n3090), .B(n3161), .Z(n3160) );
  XNOR U4186 ( .A(c[988]), .B(n3162), .Z(n3161) );
  IV U4187 ( .A(o[988]), .Z(n3162) );
  XNOR U4188 ( .A(n3163), .B(n3164), .Z(o[988]) );
  XOR U4189 ( .A(n3165), .B(o[987]), .Z(creg_next[987]) );
  AND U4190 ( .A(n3090), .B(n3166), .Z(n3165) );
  XNOR U4191 ( .A(c[987]), .B(n3167), .Z(n3166) );
  IV U4192 ( .A(o[987]), .Z(n3167) );
  XNOR U4193 ( .A(n3168), .B(n3169), .Z(o[987]) );
  XOR U4194 ( .A(n3170), .B(o[986]), .Z(creg_next[986]) );
  AND U4195 ( .A(n3090), .B(n3171), .Z(n3170) );
  XNOR U4196 ( .A(c[986]), .B(n3172), .Z(n3171) );
  IV U4197 ( .A(o[986]), .Z(n3172) );
  XNOR U4198 ( .A(n3173), .B(n3174), .Z(o[986]) );
  XOR U4199 ( .A(n3175), .B(o[985]), .Z(creg_next[985]) );
  AND U4200 ( .A(n3090), .B(n3176), .Z(n3175) );
  XNOR U4201 ( .A(c[985]), .B(n3177), .Z(n3176) );
  IV U4202 ( .A(o[985]), .Z(n3177) );
  XNOR U4203 ( .A(n3178), .B(n3179), .Z(o[985]) );
  XOR U4204 ( .A(n3180), .B(o[984]), .Z(creg_next[984]) );
  AND U4205 ( .A(n3090), .B(n3181), .Z(n3180) );
  XNOR U4206 ( .A(c[984]), .B(n3182), .Z(n3181) );
  IV U4207 ( .A(o[984]), .Z(n3182) );
  XNOR U4208 ( .A(n3183), .B(n3184), .Z(o[984]) );
  XOR U4209 ( .A(n3185), .B(o[983]), .Z(creg_next[983]) );
  AND U4210 ( .A(n3090), .B(n3186), .Z(n3185) );
  XNOR U4211 ( .A(c[983]), .B(n3187), .Z(n3186) );
  IV U4212 ( .A(o[983]), .Z(n3187) );
  XNOR U4213 ( .A(n3188), .B(n3189), .Z(o[983]) );
  XOR U4214 ( .A(n3190), .B(o[982]), .Z(creg_next[982]) );
  AND U4215 ( .A(n3090), .B(n3191), .Z(n3190) );
  XNOR U4216 ( .A(c[982]), .B(n3192), .Z(n3191) );
  IV U4217 ( .A(o[982]), .Z(n3192) );
  XNOR U4218 ( .A(n3193), .B(n3194), .Z(o[982]) );
  XOR U4219 ( .A(n3195), .B(o[981]), .Z(creg_next[981]) );
  AND U4220 ( .A(n3090), .B(n3196), .Z(n3195) );
  XNOR U4221 ( .A(c[981]), .B(n3197), .Z(n3196) );
  IV U4222 ( .A(o[981]), .Z(n3197) );
  XNOR U4223 ( .A(n3198), .B(n3199), .Z(o[981]) );
  XOR U4224 ( .A(n3200), .B(o[980]), .Z(creg_next[980]) );
  AND U4225 ( .A(n3090), .B(n3201), .Z(n3200) );
  XNOR U4226 ( .A(c[980]), .B(n3202), .Z(n3201) );
  IV U4227 ( .A(o[980]), .Z(n3202) );
  XNOR U4228 ( .A(n3203), .B(n3204), .Z(o[980]) );
  XOR U4229 ( .A(n3205), .B(o[97]), .Z(creg_next[97]) );
  AND U4230 ( .A(n3090), .B(n3206), .Z(n3205) );
  XNOR U4231 ( .A(c[97]), .B(n3207), .Z(n3206) );
  IV U4232 ( .A(o[97]), .Z(n3207) );
  XNOR U4233 ( .A(n3208), .B(n3209), .Z(o[97]) );
  XOR U4234 ( .A(n3210), .B(o[979]), .Z(creg_next[979]) );
  AND U4235 ( .A(n3090), .B(n3211), .Z(n3210) );
  XNOR U4236 ( .A(c[979]), .B(n3212), .Z(n3211) );
  IV U4237 ( .A(o[979]), .Z(n3212) );
  XNOR U4238 ( .A(n3213), .B(n3214), .Z(o[979]) );
  XOR U4239 ( .A(n3215), .B(o[978]), .Z(creg_next[978]) );
  AND U4240 ( .A(n3090), .B(n3216), .Z(n3215) );
  XNOR U4241 ( .A(c[978]), .B(n3217), .Z(n3216) );
  IV U4242 ( .A(o[978]), .Z(n3217) );
  XNOR U4243 ( .A(n3218), .B(n3219), .Z(o[978]) );
  XOR U4244 ( .A(n3220), .B(o[977]), .Z(creg_next[977]) );
  AND U4245 ( .A(n3090), .B(n3221), .Z(n3220) );
  XNOR U4246 ( .A(c[977]), .B(n3222), .Z(n3221) );
  IV U4247 ( .A(o[977]), .Z(n3222) );
  XNOR U4248 ( .A(n3223), .B(n3224), .Z(o[977]) );
  XOR U4249 ( .A(n3225), .B(o[976]), .Z(creg_next[976]) );
  AND U4250 ( .A(n3090), .B(n3226), .Z(n3225) );
  XNOR U4251 ( .A(c[976]), .B(n3227), .Z(n3226) );
  IV U4252 ( .A(o[976]), .Z(n3227) );
  XNOR U4253 ( .A(n3228), .B(n3229), .Z(o[976]) );
  XOR U4254 ( .A(n3230), .B(o[975]), .Z(creg_next[975]) );
  AND U4255 ( .A(n3090), .B(n3231), .Z(n3230) );
  XNOR U4256 ( .A(c[975]), .B(n3232), .Z(n3231) );
  IV U4257 ( .A(o[975]), .Z(n3232) );
  XNOR U4258 ( .A(n3233), .B(n3234), .Z(o[975]) );
  XOR U4259 ( .A(n3235), .B(o[974]), .Z(creg_next[974]) );
  AND U4260 ( .A(n3090), .B(n3236), .Z(n3235) );
  XNOR U4261 ( .A(c[974]), .B(n3237), .Z(n3236) );
  IV U4262 ( .A(o[974]), .Z(n3237) );
  XNOR U4263 ( .A(n3238), .B(n3239), .Z(o[974]) );
  XOR U4264 ( .A(n3240), .B(o[973]), .Z(creg_next[973]) );
  AND U4265 ( .A(n3090), .B(n3241), .Z(n3240) );
  XNOR U4266 ( .A(c[973]), .B(n3242), .Z(n3241) );
  IV U4267 ( .A(o[973]), .Z(n3242) );
  XNOR U4268 ( .A(n3243), .B(n3244), .Z(o[973]) );
  XOR U4269 ( .A(n3245), .B(o[972]), .Z(creg_next[972]) );
  AND U4270 ( .A(n3090), .B(n3246), .Z(n3245) );
  XNOR U4271 ( .A(c[972]), .B(n3247), .Z(n3246) );
  IV U4272 ( .A(o[972]), .Z(n3247) );
  XNOR U4273 ( .A(n3248), .B(n3249), .Z(o[972]) );
  XOR U4274 ( .A(n3250), .B(o[971]), .Z(creg_next[971]) );
  AND U4275 ( .A(n3090), .B(n3251), .Z(n3250) );
  XNOR U4276 ( .A(c[971]), .B(n3252), .Z(n3251) );
  IV U4277 ( .A(o[971]), .Z(n3252) );
  XNOR U4278 ( .A(n3253), .B(n3254), .Z(o[971]) );
  XOR U4279 ( .A(n3255), .B(o[970]), .Z(creg_next[970]) );
  AND U4280 ( .A(n3090), .B(n3256), .Z(n3255) );
  XNOR U4281 ( .A(c[970]), .B(n3257), .Z(n3256) );
  IV U4282 ( .A(o[970]), .Z(n3257) );
  XNOR U4283 ( .A(n3258), .B(n3259), .Z(o[970]) );
  XOR U4284 ( .A(n3260), .B(o[96]), .Z(creg_next[96]) );
  AND U4285 ( .A(n3090), .B(n3261), .Z(n3260) );
  XNOR U4286 ( .A(c[96]), .B(n3262), .Z(n3261) );
  IV U4287 ( .A(o[96]), .Z(n3262) );
  XNOR U4288 ( .A(n3263), .B(n3264), .Z(o[96]) );
  XOR U4289 ( .A(n3265), .B(o[969]), .Z(creg_next[969]) );
  AND U4290 ( .A(n3090), .B(n3266), .Z(n3265) );
  XNOR U4291 ( .A(c[969]), .B(n3267), .Z(n3266) );
  IV U4292 ( .A(o[969]), .Z(n3267) );
  XNOR U4293 ( .A(n3268), .B(n3269), .Z(o[969]) );
  XOR U4294 ( .A(n3270), .B(o[968]), .Z(creg_next[968]) );
  AND U4295 ( .A(n3090), .B(n3271), .Z(n3270) );
  XNOR U4296 ( .A(c[968]), .B(n3272), .Z(n3271) );
  IV U4297 ( .A(o[968]), .Z(n3272) );
  XNOR U4298 ( .A(n3273), .B(n3274), .Z(o[968]) );
  XOR U4299 ( .A(n3275), .B(o[967]), .Z(creg_next[967]) );
  AND U4300 ( .A(n3090), .B(n3276), .Z(n3275) );
  XNOR U4301 ( .A(c[967]), .B(n3277), .Z(n3276) );
  IV U4302 ( .A(o[967]), .Z(n3277) );
  XNOR U4303 ( .A(n3278), .B(n3279), .Z(o[967]) );
  XOR U4304 ( .A(n3280), .B(o[966]), .Z(creg_next[966]) );
  AND U4305 ( .A(n3090), .B(n3281), .Z(n3280) );
  XNOR U4306 ( .A(c[966]), .B(n3282), .Z(n3281) );
  IV U4307 ( .A(o[966]), .Z(n3282) );
  XNOR U4308 ( .A(n3283), .B(n3284), .Z(o[966]) );
  XOR U4309 ( .A(n3285), .B(o[965]), .Z(creg_next[965]) );
  AND U4310 ( .A(n3090), .B(n3286), .Z(n3285) );
  XNOR U4311 ( .A(c[965]), .B(n3287), .Z(n3286) );
  IV U4312 ( .A(o[965]), .Z(n3287) );
  XNOR U4313 ( .A(n3288), .B(n3289), .Z(o[965]) );
  XOR U4314 ( .A(n3290), .B(o[964]), .Z(creg_next[964]) );
  AND U4315 ( .A(n3090), .B(n3291), .Z(n3290) );
  XNOR U4316 ( .A(c[964]), .B(n3292), .Z(n3291) );
  IV U4317 ( .A(o[964]), .Z(n3292) );
  XNOR U4318 ( .A(n3293), .B(n3294), .Z(o[964]) );
  XOR U4319 ( .A(n3295), .B(o[963]), .Z(creg_next[963]) );
  AND U4320 ( .A(n3090), .B(n3296), .Z(n3295) );
  XNOR U4321 ( .A(c[963]), .B(n3297), .Z(n3296) );
  IV U4322 ( .A(o[963]), .Z(n3297) );
  XNOR U4323 ( .A(n3298), .B(n3299), .Z(o[963]) );
  XOR U4324 ( .A(n3300), .B(o[962]), .Z(creg_next[962]) );
  AND U4325 ( .A(n3090), .B(n3301), .Z(n3300) );
  XNOR U4326 ( .A(c[962]), .B(n3302), .Z(n3301) );
  IV U4327 ( .A(o[962]), .Z(n3302) );
  XNOR U4328 ( .A(n3303), .B(n3304), .Z(o[962]) );
  XOR U4329 ( .A(n3305), .B(o[961]), .Z(creg_next[961]) );
  AND U4330 ( .A(n3090), .B(n3306), .Z(n3305) );
  XNOR U4331 ( .A(c[961]), .B(n3307), .Z(n3306) );
  IV U4332 ( .A(o[961]), .Z(n3307) );
  XNOR U4333 ( .A(n3308), .B(n3309), .Z(o[961]) );
  XOR U4334 ( .A(n3310), .B(o[960]), .Z(creg_next[960]) );
  AND U4335 ( .A(n3090), .B(n3311), .Z(n3310) );
  XNOR U4336 ( .A(c[960]), .B(n3312), .Z(n3311) );
  IV U4337 ( .A(o[960]), .Z(n3312) );
  XNOR U4338 ( .A(n3313), .B(n3314), .Z(o[960]) );
  XOR U4339 ( .A(n3315), .B(o[95]), .Z(creg_next[95]) );
  AND U4340 ( .A(n3090), .B(n3316), .Z(n3315) );
  XNOR U4341 ( .A(c[95]), .B(n3317), .Z(n3316) );
  IV U4342 ( .A(o[95]), .Z(n3317) );
  XNOR U4343 ( .A(n3318), .B(n3319), .Z(o[95]) );
  XOR U4344 ( .A(n3320), .B(o[959]), .Z(creg_next[959]) );
  AND U4345 ( .A(n3090), .B(n3321), .Z(n3320) );
  XNOR U4346 ( .A(c[959]), .B(n3322), .Z(n3321) );
  IV U4347 ( .A(o[959]), .Z(n3322) );
  XNOR U4348 ( .A(n3323), .B(n3324), .Z(o[959]) );
  XOR U4349 ( .A(n3325), .B(o[958]), .Z(creg_next[958]) );
  AND U4350 ( .A(n3090), .B(n3326), .Z(n3325) );
  XNOR U4351 ( .A(c[958]), .B(n3327), .Z(n3326) );
  IV U4352 ( .A(o[958]), .Z(n3327) );
  XNOR U4353 ( .A(n3328), .B(n3329), .Z(o[958]) );
  XOR U4354 ( .A(n3330), .B(o[957]), .Z(creg_next[957]) );
  AND U4355 ( .A(n3090), .B(n3331), .Z(n3330) );
  XNOR U4356 ( .A(c[957]), .B(n3332), .Z(n3331) );
  IV U4357 ( .A(o[957]), .Z(n3332) );
  XNOR U4358 ( .A(n3333), .B(n3334), .Z(o[957]) );
  XOR U4359 ( .A(n3335), .B(o[956]), .Z(creg_next[956]) );
  AND U4360 ( .A(n3090), .B(n3336), .Z(n3335) );
  XNOR U4361 ( .A(c[956]), .B(n3337), .Z(n3336) );
  IV U4362 ( .A(o[956]), .Z(n3337) );
  XNOR U4363 ( .A(n3338), .B(n3339), .Z(o[956]) );
  XOR U4364 ( .A(n3340), .B(o[955]), .Z(creg_next[955]) );
  AND U4365 ( .A(n3090), .B(n3341), .Z(n3340) );
  XNOR U4366 ( .A(c[955]), .B(n3342), .Z(n3341) );
  IV U4367 ( .A(o[955]), .Z(n3342) );
  XNOR U4368 ( .A(n3343), .B(n3344), .Z(o[955]) );
  XOR U4369 ( .A(n3345), .B(o[954]), .Z(creg_next[954]) );
  AND U4370 ( .A(n3090), .B(n3346), .Z(n3345) );
  XNOR U4371 ( .A(c[954]), .B(n3347), .Z(n3346) );
  IV U4372 ( .A(o[954]), .Z(n3347) );
  XNOR U4373 ( .A(n3348), .B(n3349), .Z(o[954]) );
  XOR U4374 ( .A(n3350), .B(o[953]), .Z(creg_next[953]) );
  AND U4375 ( .A(n3090), .B(n3351), .Z(n3350) );
  XNOR U4376 ( .A(c[953]), .B(n3352), .Z(n3351) );
  IV U4377 ( .A(o[953]), .Z(n3352) );
  XNOR U4378 ( .A(n3353), .B(n3354), .Z(o[953]) );
  XOR U4379 ( .A(n3355), .B(o[952]), .Z(creg_next[952]) );
  AND U4380 ( .A(n3090), .B(n3356), .Z(n3355) );
  XNOR U4381 ( .A(c[952]), .B(n3357), .Z(n3356) );
  IV U4382 ( .A(o[952]), .Z(n3357) );
  XNOR U4383 ( .A(n3358), .B(n3359), .Z(o[952]) );
  XOR U4384 ( .A(n3360), .B(o[951]), .Z(creg_next[951]) );
  AND U4385 ( .A(n3090), .B(n3361), .Z(n3360) );
  XNOR U4386 ( .A(c[951]), .B(n3362), .Z(n3361) );
  IV U4387 ( .A(o[951]), .Z(n3362) );
  XNOR U4388 ( .A(n3363), .B(n3364), .Z(o[951]) );
  XOR U4389 ( .A(n3365), .B(o[950]), .Z(creg_next[950]) );
  AND U4390 ( .A(n3090), .B(n3366), .Z(n3365) );
  XNOR U4391 ( .A(c[950]), .B(n3367), .Z(n3366) );
  IV U4392 ( .A(o[950]), .Z(n3367) );
  XNOR U4393 ( .A(n3368), .B(n3369), .Z(o[950]) );
  XOR U4394 ( .A(n3370), .B(o[94]), .Z(creg_next[94]) );
  AND U4395 ( .A(n3090), .B(n3371), .Z(n3370) );
  XNOR U4396 ( .A(c[94]), .B(n3372), .Z(n3371) );
  IV U4397 ( .A(o[94]), .Z(n3372) );
  XNOR U4398 ( .A(n3373), .B(n3374), .Z(o[94]) );
  XOR U4399 ( .A(n3375), .B(o[949]), .Z(creg_next[949]) );
  AND U4400 ( .A(n3090), .B(n3376), .Z(n3375) );
  XNOR U4401 ( .A(c[949]), .B(n3377), .Z(n3376) );
  IV U4402 ( .A(o[949]), .Z(n3377) );
  XNOR U4403 ( .A(n3378), .B(n3379), .Z(o[949]) );
  XOR U4404 ( .A(n3380), .B(o[948]), .Z(creg_next[948]) );
  AND U4405 ( .A(n3090), .B(n3381), .Z(n3380) );
  XNOR U4406 ( .A(c[948]), .B(n3382), .Z(n3381) );
  IV U4407 ( .A(o[948]), .Z(n3382) );
  XNOR U4408 ( .A(n3383), .B(n3384), .Z(o[948]) );
  XOR U4409 ( .A(n3385), .B(o[947]), .Z(creg_next[947]) );
  AND U4410 ( .A(n3090), .B(n3386), .Z(n3385) );
  XNOR U4411 ( .A(c[947]), .B(n3387), .Z(n3386) );
  IV U4412 ( .A(o[947]), .Z(n3387) );
  XNOR U4413 ( .A(n3388), .B(n3389), .Z(o[947]) );
  XOR U4414 ( .A(n3390), .B(o[946]), .Z(creg_next[946]) );
  AND U4415 ( .A(n3090), .B(n3391), .Z(n3390) );
  XNOR U4416 ( .A(c[946]), .B(n3392), .Z(n3391) );
  IV U4417 ( .A(o[946]), .Z(n3392) );
  XNOR U4418 ( .A(n3393), .B(n3394), .Z(o[946]) );
  XOR U4419 ( .A(n3395), .B(o[945]), .Z(creg_next[945]) );
  AND U4420 ( .A(n3090), .B(n3396), .Z(n3395) );
  XNOR U4421 ( .A(c[945]), .B(n3397), .Z(n3396) );
  IV U4422 ( .A(o[945]), .Z(n3397) );
  XNOR U4423 ( .A(n3398), .B(n3399), .Z(o[945]) );
  XOR U4424 ( .A(n3400), .B(o[944]), .Z(creg_next[944]) );
  AND U4425 ( .A(n3090), .B(n3401), .Z(n3400) );
  XNOR U4426 ( .A(c[944]), .B(n3402), .Z(n3401) );
  IV U4427 ( .A(o[944]), .Z(n3402) );
  XNOR U4428 ( .A(n3403), .B(n3404), .Z(o[944]) );
  XOR U4429 ( .A(n3405), .B(o[943]), .Z(creg_next[943]) );
  AND U4430 ( .A(n3090), .B(n3406), .Z(n3405) );
  XNOR U4431 ( .A(c[943]), .B(n3407), .Z(n3406) );
  IV U4432 ( .A(o[943]), .Z(n3407) );
  XNOR U4433 ( .A(n3408), .B(n3409), .Z(o[943]) );
  XOR U4434 ( .A(n3410), .B(o[942]), .Z(creg_next[942]) );
  AND U4435 ( .A(n3090), .B(n3411), .Z(n3410) );
  XNOR U4436 ( .A(c[942]), .B(n3412), .Z(n3411) );
  IV U4437 ( .A(o[942]), .Z(n3412) );
  XNOR U4438 ( .A(n3413), .B(n3414), .Z(o[942]) );
  XOR U4439 ( .A(n3415), .B(o[941]), .Z(creg_next[941]) );
  AND U4440 ( .A(n3090), .B(n3416), .Z(n3415) );
  XNOR U4441 ( .A(c[941]), .B(n3417), .Z(n3416) );
  IV U4442 ( .A(o[941]), .Z(n3417) );
  XNOR U4443 ( .A(n3418), .B(n3419), .Z(o[941]) );
  XOR U4444 ( .A(n3420), .B(o[940]), .Z(creg_next[940]) );
  AND U4445 ( .A(n3090), .B(n3421), .Z(n3420) );
  XNOR U4446 ( .A(c[940]), .B(n3422), .Z(n3421) );
  IV U4447 ( .A(o[940]), .Z(n3422) );
  XNOR U4448 ( .A(n3423), .B(n3424), .Z(o[940]) );
  XOR U4449 ( .A(n3425), .B(o[93]), .Z(creg_next[93]) );
  AND U4450 ( .A(n3090), .B(n3426), .Z(n3425) );
  XNOR U4451 ( .A(c[93]), .B(n3427), .Z(n3426) );
  IV U4452 ( .A(o[93]), .Z(n3427) );
  XNOR U4453 ( .A(n3428), .B(n3429), .Z(o[93]) );
  XOR U4454 ( .A(n3430), .B(o[939]), .Z(creg_next[939]) );
  AND U4455 ( .A(n3090), .B(n3431), .Z(n3430) );
  XNOR U4456 ( .A(c[939]), .B(n3432), .Z(n3431) );
  IV U4457 ( .A(o[939]), .Z(n3432) );
  XNOR U4458 ( .A(n3433), .B(n3434), .Z(o[939]) );
  XOR U4459 ( .A(n3435), .B(o[938]), .Z(creg_next[938]) );
  AND U4460 ( .A(n3090), .B(n3436), .Z(n3435) );
  XNOR U4461 ( .A(c[938]), .B(n3437), .Z(n3436) );
  IV U4462 ( .A(o[938]), .Z(n3437) );
  XNOR U4463 ( .A(n3438), .B(n3439), .Z(o[938]) );
  XOR U4464 ( .A(n3440), .B(o[937]), .Z(creg_next[937]) );
  AND U4465 ( .A(n3090), .B(n3441), .Z(n3440) );
  XNOR U4466 ( .A(c[937]), .B(n3442), .Z(n3441) );
  IV U4467 ( .A(o[937]), .Z(n3442) );
  XNOR U4468 ( .A(n3443), .B(n3444), .Z(o[937]) );
  XOR U4469 ( .A(n3445), .B(o[936]), .Z(creg_next[936]) );
  AND U4470 ( .A(n3090), .B(n3446), .Z(n3445) );
  XNOR U4471 ( .A(c[936]), .B(n3447), .Z(n3446) );
  IV U4472 ( .A(o[936]), .Z(n3447) );
  XNOR U4473 ( .A(n3448), .B(n3449), .Z(o[936]) );
  XOR U4474 ( .A(n3450), .B(o[935]), .Z(creg_next[935]) );
  AND U4475 ( .A(n3090), .B(n3451), .Z(n3450) );
  XNOR U4476 ( .A(c[935]), .B(n3452), .Z(n3451) );
  IV U4477 ( .A(o[935]), .Z(n3452) );
  XNOR U4478 ( .A(n3453), .B(n3454), .Z(o[935]) );
  XOR U4479 ( .A(n3455), .B(o[934]), .Z(creg_next[934]) );
  AND U4480 ( .A(n3090), .B(n3456), .Z(n3455) );
  XNOR U4481 ( .A(c[934]), .B(n3457), .Z(n3456) );
  IV U4482 ( .A(o[934]), .Z(n3457) );
  XNOR U4483 ( .A(n3458), .B(n3459), .Z(o[934]) );
  XOR U4484 ( .A(n3460), .B(o[933]), .Z(creg_next[933]) );
  AND U4485 ( .A(n3090), .B(n3461), .Z(n3460) );
  XNOR U4486 ( .A(c[933]), .B(n3462), .Z(n3461) );
  IV U4487 ( .A(o[933]), .Z(n3462) );
  XNOR U4488 ( .A(n3463), .B(n3464), .Z(o[933]) );
  XOR U4489 ( .A(n3465), .B(o[932]), .Z(creg_next[932]) );
  AND U4490 ( .A(n3090), .B(n3466), .Z(n3465) );
  XNOR U4491 ( .A(c[932]), .B(n3467), .Z(n3466) );
  IV U4492 ( .A(o[932]), .Z(n3467) );
  XNOR U4493 ( .A(n3468), .B(n3469), .Z(o[932]) );
  XOR U4494 ( .A(n3470), .B(o[931]), .Z(creg_next[931]) );
  AND U4495 ( .A(n3090), .B(n3471), .Z(n3470) );
  XNOR U4496 ( .A(c[931]), .B(n3472), .Z(n3471) );
  IV U4497 ( .A(o[931]), .Z(n3472) );
  XNOR U4498 ( .A(n3473), .B(n3474), .Z(o[931]) );
  XOR U4499 ( .A(n3475), .B(o[930]), .Z(creg_next[930]) );
  AND U4500 ( .A(n3090), .B(n3476), .Z(n3475) );
  XNOR U4501 ( .A(c[930]), .B(n3477), .Z(n3476) );
  IV U4502 ( .A(o[930]), .Z(n3477) );
  XNOR U4503 ( .A(n3478), .B(n3479), .Z(o[930]) );
  XOR U4504 ( .A(n3480), .B(o[92]), .Z(creg_next[92]) );
  AND U4505 ( .A(n3090), .B(n3481), .Z(n3480) );
  XNOR U4506 ( .A(c[92]), .B(n3482), .Z(n3481) );
  IV U4507 ( .A(o[92]), .Z(n3482) );
  XNOR U4508 ( .A(n3483), .B(n3484), .Z(o[92]) );
  XOR U4509 ( .A(n3485), .B(o[929]), .Z(creg_next[929]) );
  AND U4510 ( .A(n3090), .B(n3486), .Z(n3485) );
  XNOR U4511 ( .A(c[929]), .B(n3487), .Z(n3486) );
  IV U4512 ( .A(o[929]), .Z(n3487) );
  XNOR U4513 ( .A(n3488), .B(n3489), .Z(o[929]) );
  XOR U4514 ( .A(n3490), .B(o[928]), .Z(creg_next[928]) );
  AND U4515 ( .A(n3090), .B(n3491), .Z(n3490) );
  XNOR U4516 ( .A(c[928]), .B(n3492), .Z(n3491) );
  IV U4517 ( .A(o[928]), .Z(n3492) );
  XNOR U4518 ( .A(n3493), .B(n3494), .Z(o[928]) );
  XOR U4519 ( .A(n3495), .B(o[927]), .Z(creg_next[927]) );
  AND U4520 ( .A(n3090), .B(n3496), .Z(n3495) );
  XNOR U4521 ( .A(c[927]), .B(n3497), .Z(n3496) );
  IV U4522 ( .A(o[927]), .Z(n3497) );
  XNOR U4523 ( .A(n3498), .B(n3499), .Z(o[927]) );
  XOR U4524 ( .A(n3500), .B(o[926]), .Z(creg_next[926]) );
  AND U4525 ( .A(n3090), .B(n3501), .Z(n3500) );
  XNOR U4526 ( .A(c[926]), .B(n3502), .Z(n3501) );
  IV U4527 ( .A(o[926]), .Z(n3502) );
  XNOR U4528 ( .A(n3503), .B(n3504), .Z(o[926]) );
  XOR U4529 ( .A(n3505), .B(o[925]), .Z(creg_next[925]) );
  AND U4530 ( .A(n3090), .B(n3506), .Z(n3505) );
  XNOR U4531 ( .A(c[925]), .B(n3507), .Z(n3506) );
  IV U4532 ( .A(o[925]), .Z(n3507) );
  XNOR U4533 ( .A(n3508), .B(n3509), .Z(o[925]) );
  XOR U4534 ( .A(n3510), .B(o[924]), .Z(creg_next[924]) );
  AND U4535 ( .A(n3090), .B(n3511), .Z(n3510) );
  XNOR U4536 ( .A(c[924]), .B(n3512), .Z(n3511) );
  IV U4537 ( .A(o[924]), .Z(n3512) );
  XNOR U4538 ( .A(n3513), .B(n3514), .Z(o[924]) );
  XOR U4539 ( .A(n3515), .B(o[923]), .Z(creg_next[923]) );
  AND U4540 ( .A(n3090), .B(n3516), .Z(n3515) );
  XNOR U4541 ( .A(c[923]), .B(n3517), .Z(n3516) );
  IV U4542 ( .A(o[923]), .Z(n3517) );
  XNOR U4543 ( .A(n3518), .B(n3519), .Z(o[923]) );
  XOR U4544 ( .A(n3520), .B(o[922]), .Z(creg_next[922]) );
  AND U4545 ( .A(n3090), .B(n3521), .Z(n3520) );
  XNOR U4546 ( .A(c[922]), .B(n3522), .Z(n3521) );
  IV U4547 ( .A(o[922]), .Z(n3522) );
  XNOR U4548 ( .A(n3523), .B(n3524), .Z(o[922]) );
  XOR U4549 ( .A(n3525), .B(o[921]), .Z(creg_next[921]) );
  AND U4550 ( .A(n3090), .B(n3526), .Z(n3525) );
  XNOR U4551 ( .A(c[921]), .B(n3527), .Z(n3526) );
  IV U4552 ( .A(o[921]), .Z(n3527) );
  XNOR U4553 ( .A(n3528), .B(n3529), .Z(o[921]) );
  XOR U4554 ( .A(n3530), .B(o[920]), .Z(creg_next[920]) );
  AND U4555 ( .A(n3090), .B(n3531), .Z(n3530) );
  XNOR U4556 ( .A(c[920]), .B(n3532), .Z(n3531) );
  IV U4557 ( .A(o[920]), .Z(n3532) );
  XNOR U4558 ( .A(n3533), .B(n3534), .Z(o[920]) );
  XOR U4559 ( .A(n3535), .B(o[91]), .Z(creg_next[91]) );
  AND U4560 ( .A(n3090), .B(n3536), .Z(n3535) );
  XNOR U4561 ( .A(c[91]), .B(n3537), .Z(n3536) );
  IV U4562 ( .A(o[91]), .Z(n3537) );
  XNOR U4563 ( .A(n3538), .B(n3539), .Z(o[91]) );
  XOR U4564 ( .A(n3540), .B(o[919]), .Z(creg_next[919]) );
  AND U4565 ( .A(n3090), .B(n3541), .Z(n3540) );
  XNOR U4566 ( .A(c[919]), .B(n3542), .Z(n3541) );
  IV U4567 ( .A(o[919]), .Z(n3542) );
  XNOR U4568 ( .A(n3543), .B(n3544), .Z(o[919]) );
  XOR U4569 ( .A(n3545), .B(o[918]), .Z(creg_next[918]) );
  AND U4570 ( .A(n3090), .B(n3546), .Z(n3545) );
  XNOR U4571 ( .A(c[918]), .B(n3547), .Z(n3546) );
  IV U4572 ( .A(o[918]), .Z(n3547) );
  XNOR U4573 ( .A(n3548), .B(n3549), .Z(o[918]) );
  XOR U4574 ( .A(n3550), .B(o[917]), .Z(creg_next[917]) );
  AND U4575 ( .A(n3090), .B(n3551), .Z(n3550) );
  XNOR U4576 ( .A(c[917]), .B(n3552), .Z(n3551) );
  IV U4577 ( .A(o[917]), .Z(n3552) );
  XNOR U4578 ( .A(n3553), .B(n3554), .Z(o[917]) );
  XOR U4579 ( .A(n3555), .B(o[916]), .Z(creg_next[916]) );
  AND U4580 ( .A(n3090), .B(n3556), .Z(n3555) );
  XNOR U4581 ( .A(c[916]), .B(n3557), .Z(n3556) );
  IV U4582 ( .A(o[916]), .Z(n3557) );
  XNOR U4583 ( .A(n3558), .B(n3559), .Z(o[916]) );
  XOR U4584 ( .A(n3560), .B(o[915]), .Z(creg_next[915]) );
  AND U4585 ( .A(n3090), .B(n3561), .Z(n3560) );
  XNOR U4586 ( .A(c[915]), .B(n3562), .Z(n3561) );
  IV U4587 ( .A(o[915]), .Z(n3562) );
  XNOR U4588 ( .A(n3563), .B(n3564), .Z(o[915]) );
  XOR U4589 ( .A(n3565), .B(o[914]), .Z(creg_next[914]) );
  AND U4590 ( .A(n3090), .B(n3566), .Z(n3565) );
  XNOR U4591 ( .A(c[914]), .B(n3567), .Z(n3566) );
  IV U4592 ( .A(o[914]), .Z(n3567) );
  XNOR U4593 ( .A(n3568), .B(n3569), .Z(o[914]) );
  XOR U4594 ( .A(n3570), .B(o[913]), .Z(creg_next[913]) );
  AND U4595 ( .A(n3090), .B(n3571), .Z(n3570) );
  XNOR U4596 ( .A(c[913]), .B(n3572), .Z(n3571) );
  IV U4597 ( .A(o[913]), .Z(n3572) );
  XNOR U4598 ( .A(n3573), .B(n3574), .Z(o[913]) );
  XOR U4599 ( .A(n3575), .B(o[912]), .Z(creg_next[912]) );
  AND U4600 ( .A(n3090), .B(n3576), .Z(n3575) );
  XNOR U4601 ( .A(c[912]), .B(n3577), .Z(n3576) );
  IV U4602 ( .A(o[912]), .Z(n3577) );
  XNOR U4603 ( .A(n3578), .B(n3579), .Z(o[912]) );
  XOR U4604 ( .A(n3580), .B(o[911]), .Z(creg_next[911]) );
  AND U4605 ( .A(n3090), .B(n3581), .Z(n3580) );
  XNOR U4606 ( .A(c[911]), .B(n3582), .Z(n3581) );
  IV U4607 ( .A(o[911]), .Z(n3582) );
  XNOR U4608 ( .A(n3583), .B(n3584), .Z(o[911]) );
  XOR U4609 ( .A(n3585), .B(o[910]), .Z(creg_next[910]) );
  AND U4610 ( .A(n3090), .B(n3586), .Z(n3585) );
  XNOR U4611 ( .A(c[910]), .B(n3587), .Z(n3586) );
  IV U4612 ( .A(o[910]), .Z(n3587) );
  XNOR U4613 ( .A(n3588), .B(n3589), .Z(o[910]) );
  XOR U4614 ( .A(n3590), .B(o[90]), .Z(creg_next[90]) );
  AND U4615 ( .A(n3090), .B(n3591), .Z(n3590) );
  XNOR U4616 ( .A(c[90]), .B(n3592), .Z(n3591) );
  IV U4617 ( .A(o[90]), .Z(n3592) );
  XNOR U4618 ( .A(n3593), .B(n3594), .Z(o[90]) );
  XOR U4619 ( .A(n3595), .B(o[909]), .Z(creg_next[909]) );
  AND U4620 ( .A(n3090), .B(n3596), .Z(n3595) );
  XNOR U4621 ( .A(c[909]), .B(n3597), .Z(n3596) );
  IV U4622 ( .A(o[909]), .Z(n3597) );
  XNOR U4623 ( .A(n3598), .B(n3599), .Z(o[909]) );
  XOR U4624 ( .A(n3600), .B(o[908]), .Z(creg_next[908]) );
  AND U4625 ( .A(n3090), .B(n3601), .Z(n3600) );
  XNOR U4626 ( .A(c[908]), .B(n3602), .Z(n3601) );
  IV U4627 ( .A(o[908]), .Z(n3602) );
  XNOR U4628 ( .A(n3603), .B(n3604), .Z(o[908]) );
  XOR U4629 ( .A(n3605), .B(o[907]), .Z(creg_next[907]) );
  AND U4630 ( .A(n3090), .B(n3606), .Z(n3605) );
  XNOR U4631 ( .A(c[907]), .B(n3607), .Z(n3606) );
  IV U4632 ( .A(o[907]), .Z(n3607) );
  XNOR U4633 ( .A(n3608), .B(n3609), .Z(o[907]) );
  XOR U4634 ( .A(n3610), .B(o[906]), .Z(creg_next[906]) );
  AND U4635 ( .A(n3090), .B(n3611), .Z(n3610) );
  XNOR U4636 ( .A(c[906]), .B(n3612), .Z(n3611) );
  IV U4637 ( .A(o[906]), .Z(n3612) );
  XNOR U4638 ( .A(n3613), .B(n3614), .Z(o[906]) );
  XOR U4639 ( .A(n3615), .B(o[905]), .Z(creg_next[905]) );
  AND U4640 ( .A(n3090), .B(n3616), .Z(n3615) );
  XNOR U4641 ( .A(c[905]), .B(n3617), .Z(n3616) );
  IV U4642 ( .A(o[905]), .Z(n3617) );
  XNOR U4643 ( .A(n3618), .B(n3619), .Z(o[905]) );
  XOR U4644 ( .A(n3620), .B(o[904]), .Z(creg_next[904]) );
  AND U4645 ( .A(n3090), .B(n3621), .Z(n3620) );
  XNOR U4646 ( .A(c[904]), .B(n3622), .Z(n3621) );
  IV U4647 ( .A(o[904]), .Z(n3622) );
  XNOR U4648 ( .A(n3623), .B(n3624), .Z(o[904]) );
  XOR U4649 ( .A(n3625), .B(o[903]), .Z(creg_next[903]) );
  AND U4650 ( .A(n3090), .B(n3626), .Z(n3625) );
  XNOR U4651 ( .A(c[903]), .B(n3627), .Z(n3626) );
  IV U4652 ( .A(o[903]), .Z(n3627) );
  XNOR U4653 ( .A(n3628), .B(n3629), .Z(o[903]) );
  XOR U4654 ( .A(n3630), .B(o[902]), .Z(creg_next[902]) );
  AND U4655 ( .A(n3090), .B(n3631), .Z(n3630) );
  XNOR U4656 ( .A(c[902]), .B(n3632), .Z(n3631) );
  IV U4657 ( .A(o[902]), .Z(n3632) );
  XNOR U4658 ( .A(n3633), .B(n3634), .Z(o[902]) );
  XOR U4659 ( .A(n3635), .B(o[901]), .Z(creg_next[901]) );
  AND U4660 ( .A(n3090), .B(n3636), .Z(n3635) );
  XNOR U4661 ( .A(c[901]), .B(n3637), .Z(n3636) );
  IV U4662 ( .A(o[901]), .Z(n3637) );
  XNOR U4663 ( .A(n3638), .B(n3639), .Z(o[901]) );
  XOR U4664 ( .A(n3640), .B(o[900]), .Z(creg_next[900]) );
  AND U4665 ( .A(n3090), .B(n3641), .Z(n3640) );
  XNOR U4666 ( .A(c[900]), .B(n3642), .Z(n3641) );
  IV U4667 ( .A(o[900]), .Z(n3642) );
  XNOR U4668 ( .A(n3643), .B(n3644), .Z(o[900]) );
  XOR U4669 ( .A(n3645), .B(o[8]), .Z(creg_next[8]) );
  AND U4670 ( .A(n3090), .B(n3646), .Z(n3645) );
  XNOR U4671 ( .A(c[8]), .B(n3647), .Z(n3646) );
  IV U4672 ( .A(o[8]), .Z(n3647) );
  XNOR U4673 ( .A(n3648), .B(n3649), .Z(o[8]) );
  XOR U4674 ( .A(n3650), .B(o[89]), .Z(creg_next[89]) );
  AND U4675 ( .A(n3090), .B(n3651), .Z(n3650) );
  XNOR U4676 ( .A(c[89]), .B(n3652), .Z(n3651) );
  IV U4677 ( .A(o[89]), .Z(n3652) );
  XNOR U4678 ( .A(n3653), .B(n3654), .Z(o[89]) );
  XOR U4679 ( .A(n3655), .B(o[899]), .Z(creg_next[899]) );
  AND U4680 ( .A(n3090), .B(n3656), .Z(n3655) );
  XNOR U4681 ( .A(c[899]), .B(n3657), .Z(n3656) );
  IV U4682 ( .A(o[899]), .Z(n3657) );
  XNOR U4683 ( .A(n3658), .B(n3659), .Z(o[899]) );
  XOR U4684 ( .A(n3660), .B(o[898]), .Z(creg_next[898]) );
  AND U4685 ( .A(n3090), .B(n3661), .Z(n3660) );
  XNOR U4686 ( .A(c[898]), .B(n3662), .Z(n3661) );
  IV U4687 ( .A(o[898]), .Z(n3662) );
  XNOR U4688 ( .A(n3663), .B(n3664), .Z(o[898]) );
  XOR U4689 ( .A(n3665), .B(o[897]), .Z(creg_next[897]) );
  AND U4690 ( .A(n3090), .B(n3666), .Z(n3665) );
  XNOR U4691 ( .A(c[897]), .B(n3667), .Z(n3666) );
  IV U4692 ( .A(o[897]), .Z(n3667) );
  XNOR U4693 ( .A(n3668), .B(n3669), .Z(o[897]) );
  XOR U4694 ( .A(n3670), .B(o[896]), .Z(creg_next[896]) );
  AND U4695 ( .A(n3090), .B(n3671), .Z(n3670) );
  XNOR U4696 ( .A(c[896]), .B(n3672), .Z(n3671) );
  IV U4697 ( .A(o[896]), .Z(n3672) );
  XNOR U4698 ( .A(n3673), .B(n3674), .Z(o[896]) );
  XOR U4699 ( .A(n3675), .B(o[895]), .Z(creg_next[895]) );
  AND U4700 ( .A(n3090), .B(n3676), .Z(n3675) );
  XNOR U4701 ( .A(c[895]), .B(n3677), .Z(n3676) );
  IV U4702 ( .A(o[895]), .Z(n3677) );
  XNOR U4703 ( .A(n3678), .B(n3679), .Z(o[895]) );
  XOR U4704 ( .A(n3680), .B(o[894]), .Z(creg_next[894]) );
  AND U4705 ( .A(n3090), .B(n3681), .Z(n3680) );
  XNOR U4706 ( .A(c[894]), .B(n3682), .Z(n3681) );
  IV U4707 ( .A(o[894]), .Z(n3682) );
  XNOR U4708 ( .A(n3683), .B(n3684), .Z(o[894]) );
  XOR U4709 ( .A(n3685), .B(o[893]), .Z(creg_next[893]) );
  AND U4710 ( .A(n3090), .B(n3686), .Z(n3685) );
  XNOR U4711 ( .A(c[893]), .B(n3687), .Z(n3686) );
  IV U4712 ( .A(o[893]), .Z(n3687) );
  XNOR U4713 ( .A(n3688), .B(n3689), .Z(o[893]) );
  XOR U4714 ( .A(n3690), .B(o[892]), .Z(creg_next[892]) );
  AND U4715 ( .A(n3090), .B(n3691), .Z(n3690) );
  XNOR U4716 ( .A(c[892]), .B(n3692), .Z(n3691) );
  IV U4717 ( .A(o[892]), .Z(n3692) );
  XNOR U4718 ( .A(n3693), .B(n3694), .Z(o[892]) );
  XOR U4719 ( .A(n3695), .B(o[891]), .Z(creg_next[891]) );
  AND U4720 ( .A(n3090), .B(n3696), .Z(n3695) );
  XNOR U4721 ( .A(c[891]), .B(n3697), .Z(n3696) );
  IV U4722 ( .A(o[891]), .Z(n3697) );
  XNOR U4723 ( .A(n3698), .B(n3699), .Z(o[891]) );
  XOR U4724 ( .A(n3700), .B(o[890]), .Z(creg_next[890]) );
  AND U4725 ( .A(n3090), .B(n3701), .Z(n3700) );
  XNOR U4726 ( .A(c[890]), .B(n3702), .Z(n3701) );
  IV U4727 ( .A(o[890]), .Z(n3702) );
  XNOR U4728 ( .A(n3703), .B(n3704), .Z(o[890]) );
  XOR U4729 ( .A(n3705), .B(o[88]), .Z(creg_next[88]) );
  AND U4730 ( .A(n3090), .B(n3706), .Z(n3705) );
  XNOR U4731 ( .A(c[88]), .B(n3707), .Z(n3706) );
  IV U4732 ( .A(o[88]), .Z(n3707) );
  XNOR U4733 ( .A(n3708), .B(n3709), .Z(o[88]) );
  XOR U4734 ( .A(n3710), .B(o[889]), .Z(creg_next[889]) );
  AND U4735 ( .A(n3090), .B(n3711), .Z(n3710) );
  XNOR U4736 ( .A(c[889]), .B(n3712), .Z(n3711) );
  IV U4737 ( .A(o[889]), .Z(n3712) );
  XNOR U4738 ( .A(n3713), .B(n3714), .Z(o[889]) );
  XOR U4739 ( .A(n3715), .B(o[888]), .Z(creg_next[888]) );
  AND U4740 ( .A(n3090), .B(n3716), .Z(n3715) );
  XNOR U4741 ( .A(c[888]), .B(n3717), .Z(n3716) );
  IV U4742 ( .A(o[888]), .Z(n3717) );
  XNOR U4743 ( .A(n3718), .B(n3719), .Z(o[888]) );
  XOR U4744 ( .A(n3720), .B(o[887]), .Z(creg_next[887]) );
  AND U4745 ( .A(n3090), .B(n3721), .Z(n3720) );
  XNOR U4746 ( .A(c[887]), .B(n3722), .Z(n3721) );
  IV U4747 ( .A(o[887]), .Z(n3722) );
  XNOR U4748 ( .A(n3723), .B(n3724), .Z(o[887]) );
  XOR U4749 ( .A(n3725), .B(o[886]), .Z(creg_next[886]) );
  AND U4750 ( .A(n3090), .B(n3726), .Z(n3725) );
  XNOR U4751 ( .A(c[886]), .B(n3727), .Z(n3726) );
  IV U4752 ( .A(o[886]), .Z(n3727) );
  XNOR U4753 ( .A(n3728), .B(n3729), .Z(o[886]) );
  XOR U4754 ( .A(n3730), .B(o[885]), .Z(creg_next[885]) );
  AND U4755 ( .A(n3090), .B(n3731), .Z(n3730) );
  XNOR U4756 ( .A(c[885]), .B(n3732), .Z(n3731) );
  IV U4757 ( .A(o[885]), .Z(n3732) );
  XNOR U4758 ( .A(n3733), .B(n3734), .Z(o[885]) );
  XOR U4759 ( .A(n3735), .B(o[884]), .Z(creg_next[884]) );
  AND U4760 ( .A(n3090), .B(n3736), .Z(n3735) );
  XNOR U4761 ( .A(c[884]), .B(n3737), .Z(n3736) );
  IV U4762 ( .A(o[884]), .Z(n3737) );
  XNOR U4763 ( .A(n3738), .B(n3739), .Z(o[884]) );
  XOR U4764 ( .A(n3740), .B(o[883]), .Z(creg_next[883]) );
  AND U4765 ( .A(n3090), .B(n3741), .Z(n3740) );
  XNOR U4766 ( .A(c[883]), .B(n3742), .Z(n3741) );
  IV U4767 ( .A(o[883]), .Z(n3742) );
  XNOR U4768 ( .A(n3743), .B(n3744), .Z(o[883]) );
  XOR U4769 ( .A(n3745), .B(o[882]), .Z(creg_next[882]) );
  AND U4770 ( .A(n3090), .B(n3746), .Z(n3745) );
  XNOR U4771 ( .A(c[882]), .B(n3747), .Z(n3746) );
  IV U4772 ( .A(o[882]), .Z(n3747) );
  XNOR U4773 ( .A(n3748), .B(n3749), .Z(o[882]) );
  XOR U4774 ( .A(n3750), .B(o[881]), .Z(creg_next[881]) );
  AND U4775 ( .A(n3090), .B(n3751), .Z(n3750) );
  XNOR U4776 ( .A(c[881]), .B(n3752), .Z(n3751) );
  IV U4777 ( .A(o[881]), .Z(n3752) );
  XNOR U4778 ( .A(n3753), .B(n3754), .Z(o[881]) );
  XOR U4779 ( .A(n3755), .B(o[880]), .Z(creg_next[880]) );
  AND U4780 ( .A(n3090), .B(n3756), .Z(n3755) );
  XNOR U4781 ( .A(c[880]), .B(n3757), .Z(n3756) );
  IV U4782 ( .A(o[880]), .Z(n3757) );
  XNOR U4783 ( .A(n3758), .B(n3759), .Z(o[880]) );
  XOR U4784 ( .A(n3760), .B(o[87]), .Z(creg_next[87]) );
  AND U4785 ( .A(n3090), .B(n3761), .Z(n3760) );
  XNOR U4786 ( .A(c[87]), .B(n3762), .Z(n3761) );
  IV U4787 ( .A(o[87]), .Z(n3762) );
  XNOR U4788 ( .A(n3763), .B(n3764), .Z(o[87]) );
  XOR U4789 ( .A(n3765), .B(o[879]), .Z(creg_next[879]) );
  AND U4790 ( .A(n3090), .B(n3766), .Z(n3765) );
  XNOR U4791 ( .A(c[879]), .B(n3767), .Z(n3766) );
  IV U4792 ( .A(o[879]), .Z(n3767) );
  XNOR U4793 ( .A(n3768), .B(n3769), .Z(o[879]) );
  XOR U4794 ( .A(n3770), .B(o[878]), .Z(creg_next[878]) );
  AND U4795 ( .A(n3090), .B(n3771), .Z(n3770) );
  XNOR U4796 ( .A(c[878]), .B(n3772), .Z(n3771) );
  IV U4797 ( .A(o[878]), .Z(n3772) );
  XNOR U4798 ( .A(n3773), .B(n3774), .Z(o[878]) );
  XOR U4799 ( .A(n3775), .B(o[877]), .Z(creg_next[877]) );
  AND U4800 ( .A(n3090), .B(n3776), .Z(n3775) );
  XNOR U4801 ( .A(c[877]), .B(n3777), .Z(n3776) );
  IV U4802 ( .A(o[877]), .Z(n3777) );
  XNOR U4803 ( .A(n3778), .B(n3779), .Z(o[877]) );
  XOR U4804 ( .A(n3780), .B(o[876]), .Z(creg_next[876]) );
  AND U4805 ( .A(n3090), .B(n3781), .Z(n3780) );
  XNOR U4806 ( .A(c[876]), .B(n3782), .Z(n3781) );
  IV U4807 ( .A(o[876]), .Z(n3782) );
  XNOR U4808 ( .A(n3783), .B(n3784), .Z(o[876]) );
  XOR U4809 ( .A(n3785), .B(o[875]), .Z(creg_next[875]) );
  AND U4810 ( .A(n3090), .B(n3786), .Z(n3785) );
  XNOR U4811 ( .A(c[875]), .B(n3787), .Z(n3786) );
  IV U4812 ( .A(o[875]), .Z(n3787) );
  XNOR U4813 ( .A(n3788), .B(n3789), .Z(o[875]) );
  XOR U4814 ( .A(n3790), .B(o[874]), .Z(creg_next[874]) );
  AND U4815 ( .A(n3090), .B(n3791), .Z(n3790) );
  XNOR U4816 ( .A(c[874]), .B(n3792), .Z(n3791) );
  IV U4817 ( .A(o[874]), .Z(n3792) );
  XNOR U4818 ( .A(n3793), .B(n3794), .Z(o[874]) );
  XOR U4819 ( .A(n3795), .B(o[873]), .Z(creg_next[873]) );
  AND U4820 ( .A(n3090), .B(n3796), .Z(n3795) );
  XNOR U4821 ( .A(c[873]), .B(n3797), .Z(n3796) );
  IV U4822 ( .A(o[873]), .Z(n3797) );
  XNOR U4823 ( .A(n3798), .B(n3799), .Z(o[873]) );
  XOR U4824 ( .A(n3800), .B(o[872]), .Z(creg_next[872]) );
  AND U4825 ( .A(n3090), .B(n3801), .Z(n3800) );
  XNOR U4826 ( .A(c[872]), .B(n3802), .Z(n3801) );
  IV U4827 ( .A(o[872]), .Z(n3802) );
  XNOR U4828 ( .A(n3803), .B(n3804), .Z(o[872]) );
  XOR U4829 ( .A(n3805), .B(o[871]), .Z(creg_next[871]) );
  AND U4830 ( .A(n3090), .B(n3806), .Z(n3805) );
  XNOR U4831 ( .A(c[871]), .B(n3807), .Z(n3806) );
  IV U4832 ( .A(o[871]), .Z(n3807) );
  XNOR U4833 ( .A(n3808), .B(n3809), .Z(o[871]) );
  XOR U4834 ( .A(n3810), .B(o[870]), .Z(creg_next[870]) );
  AND U4835 ( .A(n3090), .B(n3811), .Z(n3810) );
  XNOR U4836 ( .A(c[870]), .B(n3812), .Z(n3811) );
  IV U4837 ( .A(o[870]), .Z(n3812) );
  XNOR U4838 ( .A(n3813), .B(n3814), .Z(o[870]) );
  XOR U4839 ( .A(n3815), .B(o[86]), .Z(creg_next[86]) );
  AND U4840 ( .A(n3090), .B(n3816), .Z(n3815) );
  XNOR U4841 ( .A(c[86]), .B(n3817), .Z(n3816) );
  IV U4842 ( .A(o[86]), .Z(n3817) );
  XNOR U4843 ( .A(n3818), .B(n3819), .Z(o[86]) );
  XOR U4844 ( .A(n3820), .B(o[869]), .Z(creg_next[869]) );
  AND U4845 ( .A(n3090), .B(n3821), .Z(n3820) );
  XNOR U4846 ( .A(c[869]), .B(n3822), .Z(n3821) );
  IV U4847 ( .A(o[869]), .Z(n3822) );
  XNOR U4848 ( .A(n3823), .B(n3824), .Z(o[869]) );
  XOR U4849 ( .A(n3825), .B(o[868]), .Z(creg_next[868]) );
  AND U4850 ( .A(n3090), .B(n3826), .Z(n3825) );
  XNOR U4851 ( .A(c[868]), .B(n3827), .Z(n3826) );
  IV U4852 ( .A(o[868]), .Z(n3827) );
  XNOR U4853 ( .A(n3828), .B(n3829), .Z(o[868]) );
  XOR U4854 ( .A(n3830), .B(o[867]), .Z(creg_next[867]) );
  AND U4855 ( .A(n3090), .B(n3831), .Z(n3830) );
  XNOR U4856 ( .A(c[867]), .B(n3832), .Z(n3831) );
  IV U4857 ( .A(o[867]), .Z(n3832) );
  XNOR U4858 ( .A(n3833), .B(n3834), .Z(o[867]) );
  XOR U4859 ( .A(n3835), .B(o[866]), .Z(creg_next[866]) );
  AND U4860 ( .A(n3090), .B(n3836), .Z(n3835) );
  XNOR U4861 ( .A(c[866]), .B(n3837), .Z(n3836) );
  IV U4862 ( .A(o[866]), .Z(n3837) );
  XNOR U4863 ( .A(n3838), .B(n3839), .Z(o[866]) );
  XOR U4864 ( .A(n3840), .B(o[865]), .Z(creg_next[865]) );
  AND U4865 ( .A(n3090), .B(n3841), .Z(n3840) );
  XNOR U4866 ( .A(c[865]), .B(n3842), .Z(n3841) );
  IV U4867 ( .A(o[865]), .Z(n3842) );
  XNOR U4868 ( .A(n3843), .B(n3844), .Z(o[865]) );
  XOR U4869 ( .A(n3845), .B(o[864]), .Z(creg_next[864]) );
  AND U4870 ( .A(n3090), .B(n3846), .Z(n3845) );
  XNOR U4871 ( .A(c[864]), .B(n3847), .Z(n3846) );
  IV U4872 ( .A(o[864]), .Z(n3847) );
  XNOR U4873 ( .A(n3848), .B(n3849), .Z(o[864]) );
  XOR U4874 ( .A(n3850), .B(o[863]), .Z(creg_next[863]) );
  AND U4875 ( .A(n3090), .B(n3851), .Z(n3850) );
  XNOR U4876 ( .A(c[863]), .B(n3852), .Z(n3851) );
  IV U4877 ( .A(o[863]), .Z(n3852) );
  XNOR U4878 ( .A(n3853), .B(n3854), .Z(o[863]) );
  XOR U4879 ( .A(n3855), .B(o[862]), .Z(creg_next[862]) );
  AND U4880 ( .A(n3090), .B(n3856), .Z(n3855) );
  XNOR U4881 ( .A(c[862]), .B(n3857), .Z(n3856) );
  IV U4882 ( .A(o[862]), .Z(n3857) );
  XNOR U4883 ( .A(n3858), .B(n3859), .Z(o[862]) );
  XOR U4884 ( .A(n3860), .B(o[861]), .Z(creg_next[861]) );
  AND U4885 ( .A(n3090), .B(n3861), .Z(n3860) );
  XNOR U4886 ( .A(c[861]), .B(n3862), .Z(n3861) );
  IV U4887 ( .A(o[861]), .Z(n3862) );
  XNOR U4888 ( .A(n3863), .B(n3864), .Z(o[861]) );
  XOR U4889 ( .A(n3865), .B(o[860]), .Z(creg_next[860]) );
  AND U4890 ( .A(n3090), .B(n3866), .Z(n3865) );
  XNOR U4891 ( .A(c[860]), .B(n3867), .Z(n3866) );
  IV U4892 ( .A(o[860]), .Z(n3867) );
  XNOR U4893 ( .A(n3868), .B(n3869), .Z(o[860]) );
  XOR U4894 ( .A(n3870), .B(o[85]), .Z(creg_next[85]) );
  AND U4895 ( .A(n3090), .B(n3871), .Z(n3870) );
  XNOR U4896 ( .A(c[85]), .B(n3872), .Z(n3871) );
  IV U4897 ( .A(o[85]), .Z(n3872) );
  XNOR U4898 ( .A(n3873), .B(n3874), .Z(o[85]) );
  XOR U4899 ( .A(n3875), .B(o[859]), .Z(creg_next[859]) );
  AND U4900 ( .A(n3090), .B(n3876), .Z(n3875) );
  XNOR U4901 ( .A(c[859]), .B(n3877), .Z(n3876) );
  IV U4902 ( .A(o[859]), .Z(n3877) );
  XNOR U4903 ( .A(n3878), .B(n3879), .Z(o[859]) );
  XOR U4904 ( .A(n3880), .B(o[858]), .Z(creg_next[858]) );
  AND U4905 ( .A(n3090), .B(n3881), .Z(n3880) );
  XNOR U4906 ( .A(c[858]), .B(n3882), .Z(n3881) );
  IV U4907 ( .A(o[858]), .Z(n3882) );
  XNOR U4908 ( .A(n3883), .B(n3884), .Z(o[858]) );
  XOR U4909 ( .A(n3885), .B(o[857]), .Z(creg_next[857]) );
  AND U4910 ( .A(n3090), .B(n3886), .Z(n3885) );
  XNOR U4911 ( .A(c[857]), .B(n3887), .Z(n3886) );
  IV U4912 ( .A(o[857]), .Z(n3887) );
  XNOR U4913 ( .A(n3888), .B(n3889), .Z(o[857]) );
  XOR U4914 ( .A(n3890), .B(o[856]), .Z(creg_next[856]) );
  AND U4915 ( .A(n3090), .B(n3891), .Z(n3890) );
  XNOR U4916 ( .A(c[856]), .B(n3892), .Z(n3891) );
  IV U4917 ( .A(o[856]), .Z(n3892) );
  XNOR U4918 ( .A(n3893), .B(n3894), .Z(o[856]) );
  XOR U4919 ( .A(n3895), .B(o[855]), .Z(creg_next[855]) );
  AND U4920 ( .A(n3090), .B(n3896), .Z(n3895) );
  XNOR U4921 ( .A(c[855]), .B(n3897), .Z(n3896) );
  IV U4922 ( .A(o[855]), .Z(n3897) );
  XNOR U4923 ( .A(n3898), .B(n3899), .Z(o[855]) );
  XOR U4924 ( .A(n3900), .B(o[854]), .Z(creg_next[854]) );
  AND U4925 ( .A(n3090), .B(n3901), .Z(n3900) );
  XNOR U4926 ( .A(c[854]), .B(n3902), .Z(n3901) );
  IV U4927 ( .A(o[854]), .Z(n3902) );
  XNOR U4928 ( .A(n3903), .B(n3904), .Z(o[854]) );
  XOR U4929 ( .A(n3905), .B(o[853]), .Z(creg_next[853]) );
  AND U4930 ( .A(n3090), .B(n3906), .Z(n3905) );
  XNOR U4931 ( .A(c[853]), .B(n3907), .Z(n3906) );
  IV U4932 ( .A(o[853]), .Z(n3907) );
  XNOR U4933 ( .A(n3908), .B(n3909), .Z(o[853]) );
  XOR U4934 ( .A(n3910), .B(o[852]), .Z(creg_next[852]) );
  AND U4935 ( .A(n3090), .B(n3911), .Z(n3910) );
  XNOR U4936 ( .A(c[852]), .B(n3912), .Z(n3911) );
  IV U4937 ( .A(o[852]), .Z(n3912) );
  XNOR U4938 ( .A(n3913), .B(n3914), .Z(o[852]) );
  XOR U4939 ( .A(n3915), .B(o[851]), .Z(creg_next[851]) );
  AND U4940 ( .A(n3090), .B(n3916), .Z(n3915) );
  XNOR U4941 ( .A(c[851]), .B(n3917), .Z(n3916) );
  IV U4942 ( .A(o[851]), .Z(n3917) );
  XNOR U4943 ( .A(n3918), .B(n3919), .Z(o[851]) );
  XOR U4944 ( .A(n3920), .B(o[850]), .Z(creg_next[850]) );
  AND U4945 ( .A(n3090), .B(n3921), .Z(n3920) );
  XNOR U4946 ( .A(c[850]), .B(n3922), .Z(n3921) );
  IV U4947 ( .A(o[850]), .Z(n3922) );
  XNOR U4948 ( .A(n3923), .B(n3924), .Z(o[850]) );
  XOR U4949 ( .A(n3925), .B(o[84]), .Z(creg_next[84]) );
  AND U4950 ( .A(n3090), .B(n3926), .Z(n3925) );
  XNOR U4951 ( .A(c[84]), .B(n3927), .Z(n3926) );
  IV U4952 ( .A(o[84]), .Z(n3927) );
  XNOR U4953 ( .A(n3928), .B(n3929), .Z(o[84]) );
  XOR U4954 ( .A(n3930), .B(o[849]), .Z(creg_next[849]) );
  AND U4955 ( .A(n3090), .B(n3931), .Z(n3930) );
  XNOR U4956 ( .A(c[849]), .B(n3932), .Z(n3931) );
  IV U4957 ( .A(o[849]), .Z(n3932) );
  XNOR U4958 ( .A(n3933), .B(n3934), .Z(o[849]) );
  XOR U4959 ( .A(n3935), .B(o[848]), .Z(creg_next[848]) );
  AND U4960 ( .A(n3090), .B(n3936), .Z(n3935) );
  XNOR U4961 ( .A(c[848]), .B(n3937), .Z(n3936) );
  IV U4962 ( .A(o[848]), .Z(n3937) );
  XNOR U4963 ( .A(n3938), .B(n3939), .Z(o[848]) );
  XOR U4964 ( .A(n3940), .B(o[847]), .Z(creg_next[847]) );
  AND U4965 ( .A(n3090), .B(n3941), .Z(n3940) );
  XNOR U4966 ( .A(c[847]), .B(n3942), .Z(n3941) );
  IV U4967 ( .A(o[847]), .Z(n3942) );
  XNOR U4968 ( .A(n3943), .B(n3944), .Z(o[847]) );
  XOR U4969 ( .A(n3945), .B(o[846]), .Z(creg_next[846]) );
  AND U4970 ( .A(n3090), .B(n3946), .Z(n3945) );
  XNOR U4971 ( .A(c[846]), .B(n3947), .Z(n3946) );
  IV U4972 ( .A(o[846]), .Z(n3947) );
  XNOR U4973 ( .A(n3948), .B(n3949), .Z(o[846]) );
  XOR U4974 ( .A(n3950), .B(o[845]), .Z(creg_next[845]) );
  AND U4975 ( .A(n3090), .B(n3951), .Z(n3950) );
  XNOR U4976 ( .A(c[845]), .B(n3952), .Z(n3951) );
  IV U4977 ( .A(o[845]), .Z(n3952) );
  XNOR U4978 ( .A(n3953), .B(n3954), .Z(o[845]) );
  XOR U4979 ( .A(n3955), .B(o[844]), .Z(creg_next[844]) );
  AND U4980 ( .A(n3090), .B(n3956), .Z(n3955) );
  XNOR U4981 ( .A(c[844]), .B(n3957), .Z(n3956) );
  IV U4982 ( .A(o[844]), .Z(n3957) );
  XNOR U4983 ( .A(n3958), .B(n3959), .Z(o[844]) );
  XOR U4984 ( .A(n3960), .B(o[843]), .Z(creg_next[843]) );
  AND U4985 ( .A(n3090), .B(n3961), .Z(n3960) );
  XNOR U4986 ( .A(c[843]), .B(n3962), .Z(n3961) );
  IV U4987 ( .A(o[843]), .Z(n3962) );
  XNOR U4988 ( .A(n3963), .B(n3964), .Z(o[843]) );
  XOR U4989 ( .A(n3965), .B(o[842]), .Z(creg_next[842]) );
  AND U4990 ( .A(n3090), .B(n3966), .Z(n3965) );
  XNOR U4991 ( .A(c[842]), .B(n3967), .Z(n3966) );
  IV U4992 ( .A(o[842]), .Z(n3967) );
  XNOR U4993 ( .A(n3968), .B(n3969), .Z(o[842]) );
  XOR U4994 ( .A(n3970), .B(o[841]), .Z(creg_next[841]) );
  AND U4995 ( .A(n3090), .B(n3971), .Z(n3970) );
  XNOR U4996 ( .A(c[841]), .B(n3972), .Z(n3971) );
  IV U4997 ( .A(o[841]), .Z(n3972) );
  XNOR U4998 ( .A(n3973), .B(n3974), .Z(o[841]) );
  XOR U4999 ( .A(n3975), .B(o[840]), .Z(creg_next[840]) );
  AND U5000 ( .A(n3090), .B(n3976), .Z(n3975) );
  XNOR U5001 ( .A(c[840]), .B(n3977), .Z(n3976) );
  IV U5002 ( .A(o[840]), .Z(n3977) );
  XNOR U5003 ( .A(n3978), .B(n3979), .Z(o[840]) );
  XOR U5004 ( .A(n3980), .B(o[83]), .Z(creg_next[83]) );
  AND U5005 ( .A(n3090), .B(n3981), .Z(n3980) );
  XNOR U5006 ( .A(c[83]), .B(n3982), .Z(n3981) );
  IV U5007 ( .A(o[83]), .Z(n3982) );
  XNOR U5008 ( .A(n3983), .B(n3984), .Z(o[83]) );
  XOR U5009 ( .A(n3985), .B(o[839]), .Z(creg_next[839]) );
  AND U5010 ( .A(n3090), .B(n3986), .Z(n3985) );
  XNOR U5011 ( .A(c[839]), .B(n3987), .Z(n3986) );
  IV U5012 ( .A(o[839]), .Z(n3987) );
  XNOR U5013 ( .A(n3988), .B(n3989), .Z(o[839]) );
  XOR U5014 ( .A(n3990), .B(o[838]), .Z(creg_next[838]) );
  AND U5015 ( .A(n3090), .B(n3991), .Z(n3990) );
  XNOR U5016 ( .A(c[838]), .B(n3992), .Z(n3991) );
  IV U5017 ( .A(o[838]), .Z(n3992) );
  XNOR U5018 ( .A(n3993), .B(n3994), .Z(o[838]) );
  XOR U5019 ( .A(n3995), .B(o[837]), .Z(creg_next[837]) );
  AND U5020 ( .A(n3090), .B(n3996), .Z(n3995) );
  XNOR U5021 ( .A(c[837]), .B(n3997), .Z(n3996) );
  IV U5022 ( .A(o[837]), .Z(n3997) );
  XNOR U5023 ( .A(n3998), .B(n3999), .Z(o[837]) );
  XOR U5024 ( .A(n4000), .B(o[836]), .Z(creg_next[836]) );
  AND U5025 ( .A(n3090), .B(n4001), .Z(n4000) );
  XNOR U5026 ( .A(c[836]), .B(n4002), .Z(n4001) );
  IV U5027 ( .A(o[836]), .Z(n4002) );
  XNOR U5028 ( .A(n4003), .B(n4004), .Z(o[836]) );
  XOR U5029 ( .A(n4005), .B(o[835]), .Z(creg_next[835]) );
  AND U5030 ( .A(n3090), .B(n4006), .Z(n4005) );
  XNOR U5031 ( .A(c[835]), .B(n4007), .Z(n4006) );
  IV U5032 ( .A(o[835]), .Z(n4007) );
  XNOR U5033 ( .A(n4008), .B(n4009), .Z(o[835]) );
  XOR U5034 ( .A(n4010), .B(o[834]), .Z(creg_next[834]) );
  AND U5035 ( .A(n3090), .B(n4011), .Z(n4010) );
  XNOR U5036 ( .A(c[834]), .B(n4012), .Z(n4011) );
  IV U5037 ( .A(o[834]), .Z(n4012) );
  XNOR U5038 ( .A(n4013), .B(n4014), .Z(o[834]) );
  XOR U5039 ( .A(n4015), .B(o[833]), .Z(creg_next[833]) );
  AND U5040 ( .A(n3090), .B(n4016), .Z(n4015) );
  XNOR U5041 ( .A(c[833]), .B(n4017), .Z(n4016) );
  IV U5042 ( .A(o[833]), .Z(n4017) );
  XNOR U5043 ( .A(n4018), .B(n4019), .Z(o[833]) );
  XOR U5044 ( .A(n4020), .B(o[832]), .Z(creg_next[832]) );
  AND U5045 ( .A(n3090), .B(n4021), .Z(n4020) );
  XNOR U5046 ( .A(c[832]), .B(n4022), .Z(n4021) );
  IV U5047 ( .A(o[832]), .Z(n4022) );
  XNOR U5048 ( .A(n4023), .B(n4024), .Z(o[832]) );
  XOR U5049 ( .A(n4025), .B(o[831]), .Z(creg_next[831]) );
  AND U5050 ( .A(n3090), .B(n4026), .Z(n4025) );
  XNOR U5051 ( .A(c[831]), .B(n4027), .Z(n4026) );
  IV U5052 ( .A(o[831]), .Z(n4027) );
  XNOR U5053 ( .A(n4028), .B(n4029), .Z(o[831]) );
  XOR U5054 ( .A(n4030), .B(o[830]), .Z(creg_next[830]) );
  AND U5055 ( .A(n3090), .B(n4031), .Z(n4030) );
  XNOR U5056 ( .A(c[830]), .B(n4032), .Z(n4031) );
  IV U5057 ( .A(o[830]), .Z(n4032) );
  XNOR U5058 ( .A(n4033), .B(n4034), .Z(o[830]) );
  XOR U5059 ( .A(n4035), .B(o[82]), .Z(creg_next[82]) );
  AND U5060 ( .A(n3090), .B(n4036), .Z(n4035) );
  XNOR U5061 ( .A(c[82]), .B(n4037), .Z(n4036) );
  IV U5062 ( .A(o[82]), .Z(n4037) );
  XNOR U5063 ( .A(n4038), .B(n4039), .Z(o[82]) );
  XOR U5064 ( .A(n4040), .B(o[829]), .Z(creg_next[829]) );
  AND U5065 ( .A(n3090), .B(n4041), .Z(n4040) );
  XNOR U5066 ( .A(c[829]), .B(n4042), .Z(n4041) );
  IV U5067 ( .A(o[829]), .Z(n4042) );
  XNOR U5068 ( .A(n4043), .B(n4044), .Z(o[829]) );
  XOR U5069 ( .A(n4045), .B(o[828]), .Z(creg_next[828]) );
  AND U5070 ( .A(n3090), .B(n4046), .Z(n4045) );
  XNOR U5071 ( .A(c[828]), .B(n4047), .Z(n4046) );
  IV U5072 ( .A(o[828]), .Z(n4047) );
  XNOR U5073 ( .A(n4048), .B(n4049), .Z(o[828]) );
  XOR U5074 ( .A(n4050), .B(o[827]), .Z(creg_next[827]) );
  AND U5075 ( .A(n3090), .B(n4051), .Z(n4050) );
  XNOR U5076 ( .A(c[827]), .B(n4052), .Z(n4051) );
  IV U5077 ( .A(o[827]), .Z(n4052) );
  XNOR U5078 ( .A(n4053), .B(n4054), .Z(o[827]) );
  XOR U5079 ( .A(n4055), .B(o[826]), .Z(creg_next[826]) );
  AND U5080 ( .A(n3090), .B(n4056), .Z(n4055) );
  XNOR U5081 ( .A(c[826]), .B(n4057), .Z(n4056) );
  IV U5082 ( .A(o[826]), .Z(n4057) );
  XNOR U5083 ( .A(n4058), .B(n4059), .Z(o[826]) );
  XOR U5084 ( .A(n4060), .B(o[825]), .Z(creg_next[825]) );
  AND U5085 ( .A(n3090), .B(n4061), .Z(n4060) );
  XNOR U5086 ( .A(c[825]), .B(n4062), .Z(n4061) );
  IV U5087 ( .A(o[825]), .Z(n4062) );
  XNOR U5088 ( .A(n4063), .B(n4064), .Z(o[825]) );
  XOR U5089 ( .A(n4065), .B(o[824]), .Z(creg_next[824]) );
  AND U5090 ( .A(n3090), .B(n4066), .Z(n4065) );
  XNOR U5091 ( .A(c[824]), .B(n4067), .Z(n4066) );
  IV U5092 ( .A(o[824]), .Z(n4067) );
  XNOR U5093 ( .A(n4068), .B(n4069), .Z(o[824]) );
  XOR U5094 ( .A(n4070), .B(o[823]), .Z(creg_next[823]) );
  AND U5095 ( .A(n3090), .B(n4071), .Z(n4070) );
  XNOR U5096 ( .A(c[823]), .B(n4072), .Z(n4071) );
  IV U5097 ( .A(o[823]), .Z(n4072) );
  XNOR U5098 ( .A(n4073), .B(n4074), .Z(o[823]) );
  XOR U5099 ( .A(n4075), .B(o[822]), .Z(creg_next[822]) );
  AND U5100 ( .A(n3090), .B(n4076), .Z(n4075) );
  XNOR U5101 ( .A(c[822]), .B(n4077), .Z(n4076) );
  IV U5102 ( .A(o[822]), .Z(n4077) );
  XNOR U5103 ( .A(n4078), .B(n4079), .Z(o[822]) );
  XOR U5104 ( .A(n4080), .B(o[821]), .Z(creg_next[821]) );
  AND U5105 ( .A(n3090), .B(n4081), .Z(n4080) );
  XNOR U5106 ( .A(c[821]), .B(n4082), .Z(n4081) );
  IV U5107 ( .A(o[821]), .Z(n4082) );
  XNOR U5108 ( .A(n4083), .B(n4084), .Z(o[821]) );
  XOR U5109 ( .A(n4085), .B(o[820]), .Z(creg_next[820]) );
  AND U5110 ( .A(n3090), .B(n4086), .Z(n4085) );
  XNOR U5111 ( .A(c[820]), .B(n4087), .Z(n4086) );
  IV U5112 ( .A(o[820]), .Z(n4087) );
  XNOR U5113 ( .A(n4088), .B(n4089), .Z(o[820]) );
  XOR U5114 ( .A(n4090), .B(o[81]), .Z(creg_next[81]) );
  AND U5115 ( .A(n3090), .B(n4091), .Z(n4090) );
  XNOR U5116 ( .A(c[81]), .B(n4092), .Z(n4091) );
  IV U5117 ( .A(o[81]), .Z(n4092) );
  XNOR U5118 ( .A(n4093), .B(n4094), .Z(o[81]) );
  XOR U5119 ( .A(n4095), .B(o[819]), .Z(creg_next[819]) );
  AND U5120 ( .A(n3090), .B(n4096), .Z(n4095) );
  XNOR U5121 ( .A(c[819]), .B(n4097), .Z(n4096) );
  IV U5122 ( .A(o[819]), .Z(n4097) );
  XNOR U5123 ( .A(n4098), .B(n4099), .Z(o[819]) );
  XOR U5124 ( .A(n4100), .B(o[818]), .Z(creg_next[818]) );
  AND U5125 ( .A(n3090), .B(n4101), .Z(n4100) );
  XNOR U5126 ( .A(c[818]), .B(n4102), .Z(n4101) );
  IV U5127 ( .A(o[818]), .Z(n4102) );
  XNOR U5128 ( .A(n4103), .B(n4104), .Z(o[818]) );
  XOR U5129 ( .A(n4105), .B(o[817]), .Z(creg_next[817]) );
  AND U5130 ( .A(n3090), .B(n4106), .Z(n4105) );
  XNOR U5131 ( .A(c[817]), .B(n4107), .Z(n4106) );
  IV U5132 ( .A(o[817]), .Z(n4107) );
  XNOR U5133 ( .A(n4108), .B(n4109), .Z(o[817]) );
  XOR U5134 ( .A(n4110), .B(o[816]), .Z(creg_next[816]) );
  AND U5135 ( .A(n3090), .B(n4111), .Z(n4110) );
  XNOR U5136 ( .A(c[816]), .B(n4112), .Z(n4111) );
  IV U5137 ( .A(o[816]), .Z(n4112) );
  XNOR U5138 ( .A(n4113), .B(n4114), .Z(o[816]) );
  XOR U5139 ( .A(n4115), .B(o[815]), .Z(creg_next[815]) );
  AND U5140 ( .A(n3090), .B(n4116), .Z(n4115) );
  XNOR U5141 ( .A(c[815]), .B(n4117), .Z(n4116) );
  IV U5142 ( .A(o[815]), .Z(n4117) );
  XNOR U5143 ( .A(n4118), .B(n4119), .Z(o[815]) );
  XOR U5144 ( .A(n4120), .B(o[814]), .Z(creg_next[814]) );
  AND U5145 ( .A(n3090), .B(n4121), .Z(n4120) );
  XNOR U5146 ( .A(c[814]), .B(n4122), .Z(n4121) );
  IV U5147 ( .A(o[814]), .Z(n4122) );
  XNOR U5148 ( .A(n4123), .B(n4124), .Z(o[814]) );
  XOR U5149 ( .A(n4125), .B(o[813]), .Z(creg_next[813]) );
  AND U5150 ( .A(n3090), .B(n4126), .Z(n4125) );
  XNOR U5151 ( .A(c[813]), .B(n4127), .Z(n4126) );
  IV U5152 ( .A(o[813]), .Z(n4127) );
  XNOR U5153 ( .A(n4128), .B(n4129), .Z(o[813]) );
  XOR U5154 ( .A(n4130), .B(o[812]), .Z(creg_next[812]) );
  AND U5155 ( .A(n3090), .B(n4131), .Z(n4130) );
  XNOR U5156 ( .A(c[812]), .B(n4132), .Z(n4131) );
  IV U5157 ( .A(o[812]), .Z(n4132) );
  XNOR U5158 ( .A(n4133), .B(n4134), .Z(o[812]) );
  XOR U5159 ( .A(n4135), .B(o[811]), .Z(creg_next[811]) );
  AND U5160 ( .A(n3090), .B(n4136), .Z(n4135) );
  XNOR U5161 ( .A(c[811]), .B(n4137), .Z(n4136) );
  IV U5162 ( .A(o[811]), .Z(n4137) );
  XNOR U5163 ( .A(n4138), .B(n4139), .Z(o[811]) );
  XOR U5164 ( .A(n4140), .B(o[810]), .Z(creg_next[810]) );
  AND U5165 ( .A(n3090), .B(n4141), .Z(n4140) );
  XNOR U5166 ( .A(c[810]), .B(n4142), .Z(n4141) );
  IV U5167 ( .A(o[810]), .Z(n4142) );
  XNOR U5168 ( .A(n4143), .B(n4144), .Z(o[810]) );
  XOR U5169 ( .A(n4145), .B(o[80]), .Z(creg_next[80]) );
  AND U5170 ( .A(n3090), .B(n4146), .Z(n4145) );
  XNOR U5171 ( .A(c[80]), .B(n4147), .Z(n4146) );
  IV U5172 ( .A(o[80]), .Z(n4147) );
  XNOR U5173 ( .A(n4148), .B(n4149), .Z(o[80]) );
  XOR U5174 ( .A(n4150), .B(o[809]), .Z(creg_next[809]) );
  AND U5175 ( .A(n3090), .B(n4151), .Z(n4150) );
  XNOR U5176 ( .A(c[809]), .B(n4152), .Z(n4151) );
  IV U5177 ( .A(o[809]), .Z(n4152) );
  XNOR U5178 ( .A(n4153), .B(n4154), .Z(o[809]) );
  XOR U5179 ( .A(n4155), .B(o[808]), .Z(creg_next[808]) );
  AND U5180 ( .A(n3090), .B(n4156), .Z(n4155) );
  XNOR U5181 ( .A(c[808]), .B(n4157), .Z(n4156) );
  IV U5182 ( .A(o[808]), .Z(n4157) );
  XNOR U5183 ( .A(n4158), .B(n4159), .Z(o[808]) );
  XOR U5184 ( .A(n4160), .B(o[807]), .Z(creg_next[807]) );
  AND U5185 ( .A(n3090), .B(n4161), .Z(n4160) );
  XNOR U5186 ( .A(c[807]), .B(n4162), .Z(n4161) );
  IV U5187 ( .A(o[807]), .Z(n4162) );
  XNOR U5188 ( .A(n4163), .B(n4164), .Z(o[807]) );
  XOR U5189 ( .A(n4165), .B(o[806]), .Z(creg_next[806]) );
  AND U5190 ( .A(n3090), .B(n4166), .Z(n4165) );
  XNOR U5191 ( .A(c[806]), .B(n4167), .Z(n4166) );
  IV U5192 ( .A(o[806]), .Z(n4167) );
  XNOR U5193 ( .A(n4168), .B(n4169), .Z(o[806]) );
  XOR U5194 ( .A(n4170), .B(o[805]), .Z(creg_next[805]) );
  AND U5195 ( .A(n3090), .B(n4171), .Z(n4170) );
  XNOR U5196 ( .A(c[805]), .B(n4172), .Z(n4171) );
  IV U5197 ( .A(o[805]), .Z(n4172) );
  XNOR U5198 ( .A(n4173), .B(n4174), .Z(o[805]) );
  XOR U5199 ( .A(n4175), .B(o[804]), .Z(creg_next[804]) );
  AND U5200 ( .A(n3090), .B(n4176), .Z(n4175) );
  XNOR U5201 ( .A(c[804]), .B(n4177), .Z(n4176) );
  IV U5202 ( .A(o[804]), .Z(n4177) );
  XNOR U5203 ( .A(n4178), .B(n4179), .Z(o[804]) );
  XOR U5204 ( .A(n4180), .B(o[803]), .Z(creg_next[803]) );
  AND U5205 ( .A(n3090), .B(n4181), .Z(n4180) );
  XNOR U5206 ( .A(c[803]), .B(n4182), .Z(n4181) );
  IV U5207 ( .A(o[803]), .Z(n4182) );
  XNOR U5208 ( .A(n4183), .B(n4184), .Z(o[803]) );
  XOR U5209 ( .A(n4185), .B(o[802]), .Z(creg_next[802]) );
  AND U5210 ( .A(n3090), .B(n4186), .Z(n4185) );
  XNOR U5211 ( .A(c[802]), .B(n4187), .Z(n4186) );
  IV U5212 ( .A(o[802]), .Z(n4187) );
  XNOR U5213 ( .A(n4188), .B(n4189), .Z(o[802]) );
  XOR U5214 ( .A(n4190), .B(o[801]), .Z(creg_next[801]) );
  AND U5215 ( .A(n3090), .B(n4191), .Z(n4190) );
  XNOR U5216 ( .A(c[801]), .B(n4192), .Z(n4191) );
  IV U5217 ( .A(o[801]), .Z(n4192) );
  XNOR U5218 ( .A(n4193), .B(n4194), .Z(o[801]) );
  XOR U5219 ( .A(n4195), .B(o[800]), .Z(creg_next[800]) );
  AND U5220 ( .A(n3090), .B(n4196), .Z(n4195) );
  XNOR U5221 ( .A(c[800]), .B(n4197), .Z(n4196) );
  IV U5222 ( .A(o[800]), .Z(n4197) );
  XNOR U5223 ( .A(n4198), .B(n4199), .Z(o[800]) );
  XOR U5224 ( .A(n4200), .B(o[7]), .Z(creg_next[7]) );
  AND U5225 ( .A(n3090), .B(n4201), .Z(n4200) );
  XNOR U5226 ( .A(c[7]), .B(n4202), .Z(n4201) );
  IV U5227 ( .A(o[7]), .Z(n4202) );
  XNOR U5228 ( .A(n4203), .B(n4204), .Z(o[7]) );
  XOR U5229 ( .A(n4205), .B(o[79]), .Z(creg_next[79]) );
  AND U5230 ( .A(n3090), .B(n4206), .Z(n4205) );
  XNOR U5231 ( .A(c[79]), .B(n4207), .Z(n4206) );
  IV U5232 ( .A(o[79]), .Z(n4207) );
  XNOR U5233 ( .A(n4208), .B(n4209), .Z(o[79]) );
  XOR U5234 ( .A(n4210), .B(o[799]), .Z(creg_next[799]) );
  AND U5235 ( .A(n3090), .B(n4211), .Z(n4210) );
  XNOR U5236 ( .A(c[799]), .B(n4212), .Z(n4211) );
  IV U5237 ( .A(o[799]), .Z(n4212) );
  XNOR U5238 ( .A(n4213), .B(n4214), .Z(o[799]) );
  XOR U5239 ( .A(n4215), .B(o[798]), .Z(creg_next[798]) );
  AND U5240 ( .A(n3090), .B(n4216), .Z(n4215) );
  XNOR U5241 ( .A(c[798]), .B(n4217), .Z(n4216) );
  IV U5242 ( .A(o[798]), .Z(n4217) );
  XNOR U5243 ( .A(n4218), .B(n4219), .Z(o[798]) );
  XOR U5244 ( .A(n4220), .B(o[797]), .Z(creg_next[797]) );
  AND U5245 ( .A(n3090), .B(n4221), .Z(n4220) );
  XNOR U5246 ( .A(c[797]), .B(n4222), .Z(n4221) );
  IV U5247 ( .A(o[797]), .Z(n4222) );
  XNOR U5248 ( .A(n4223), .B(n4224), .Z(o[797]) );
  XOR U5249 ( .A(n4225), .B(o[796]), .Z(creg_next[796]) );
  AND U5250 ( .A(n3090), .B(n4226), .Z(n4225) );
  XNOR U5251 ( .A(c[796]), .B(n4227), .Z(n4226) );
  IV U5252 ( .A(o[796]), .Z(n4227) );
  XNOR U5253 ( .A(n4228), .B(n4229), .Z(o[796]) );
  XOR U5254 ( .A(n4230), .B(o[795]), .Z(creg_next[795]) );
  AND U5255 ( .A(n3090), .B(n4231), .Z(n4230) );
  XNOR U5256 ( .A(c[795]), .B(n4232), .Z(n4231) );
  IV U5257 ( .A(o[795]), .Z(n4232) );
  XNOR U5258 ( .A(n4233), .B(n4234), .Z(o[795]) );
  XOR U5259 ( .A(n4235), .B(o[794]), .Z(creg_next[794]) );
  AND U5260 ( .A(n3090), .B(n4236), .Z(n4235) );
  XNOR U5261 ( .A(c[794]), .B(n4237), .Z(n4236) );
  IV U5262 ( .A(o[794]), .Z(n4237) );
  XNOR U5263 ( .A(n4238), .B(n4239), .Z(o[794]) );
  XOR U5264 ( .A(n4240), .B(o[793]), .Z(creg_next[793]) );
  AND U5265 ( .A(n3090), .B(n4241), .Z(n4240) );
  XNOR U5266 ( .A(c[793]), .B(n4242), .Z(n4241) );
  IV U5267 ( .A(o[793]), .Z(n4242) );
  XNOR U5268 ( .A(n4243), .B(n4244), .Z(o[793]) );
  XOR U5269 ( .A(n4245), .B(o[792]), .Z(creg_next[792]) );
  AND U5270 ( .A(n3090), .B(n4246), .Z(n4245) );
  XNOR U5271 ( .A(c[792]), .B(n4247), .Z(n4246) );
  IV U5272 ( .A(o[792]), .Z(n4247) );
  XNOR U5273 ( .A(n4248), .B(n4249), .Z(o[792]) );
  XOR U5274 ( .A(n4250), .B(o[791]), .Z(creg_next[791]) );
  AND U5275 ( .A(n3090), .B(n4251), .Z(n4250) );
  XNOR U5276 ( .A(c[791]), .B(n4252), .Z(n4251) );
  IV U5277 ( .A(o[791]), .Z(n4252) );
  XNOR U5278 ( .A(n4253), .B(n4254), .Z(o[791]) );
  XOR U5279 ( .A(n4255), .B(o[790]), .Z(creg_next[790]) );
  AND U5280 ( .A(n3090), .B(n4256), .Z(n4255) );
  XNOR U5281 ( .A(c[790]), .B(n4257), .Z(n4256) );
  IV U5282 ( .A(o[790]), .Z(n4257) );
  XNOR U5283 ( .A(n4258), .B(n4259), .Z(o[790]) );
  XOR U5284 ( .A(n4260), .B(o[78]), .Z(creg_next[78]) );
  AND U5285 ( .A(n3090), .B(n4261), .Z(n4260) );
  XNOR U5286 ( .A(c[78]), .B(n4262), .Z(n4261) );
  IV U5287 ( .A(o[78]), .Z(n4262) );
  XNOR U5288 ( .A(n4263), .B(n4264), .Z(o[78]) );
  XOR U5289 ( .A(n4265), .B(o[789]), .Z(creg_next[789]) );
  AND U5290 ( .A(n3090), .B(n4266), .Z(n4265) );
  XNOR U5291 ( .A(c[789]), .B(n4267), .Z(n4266) );
  IV U5292 ( .A(o[789]), .Z(n4267) );
  XNOR U5293 ( .A(n4268), .B(n4269), .Z(o[789]) );
  XOR U5294 ( .A(n4270), .B(o[788]), .Z(creg_next[788]) );
  AND U5295 ( .A(n3090), .B(n4271), .Z(n4270) );
  XNOR U5296 ( .A(c[788]), .B(n4272), .Z(n4271) );
  IV U5297 ( .A(o[788]), .Z(n4272) );
  XNOR U5298 ( .A(n4273), .B(n4274), .Z(o[788]) );
  XOR U5299 ( .A(n4275), .B(o[787]), .Z(creg_next[787]) );
  AND U5300 ( .A(n3090), .B(n4276), .Z(n4275) );
  XNOR U5301 ( .A(c[787]), .B(n4277), .Z(n4276) );
  IV U5302 ( .A(o[787]), .Z(n4277) );
  XNOR U5303 ( .A(n4278), .B(n4279), .Z(o[787]) );
  XOR U5304 ( .A(n4280), .B(o[786]), .Z(creg_next[786]) );
  AND U5305 ( .A(n3090), .B(n4281), .Z(n4280) );
  XNOR U5306 ( .A(c[786]), .B(n4282), .Z(n4281) );
  IV U5307 ( .A(o[786]), .Z(n4282) );
  XNOR U5308 ( .A(n4283), .B(n4284), .Z(o[786]) );
  XOR U5309 ( .A(n4285), .B(o[785]), .Z(creg_next[785]) );
  AND U5310 ( .A(n3090), .B(n4286), .Z(n4285) );
  XNOR U5311 ( .A(c[785]), .B(n4287), .Z(n4286) );
  IV U5312 ( .A(o[785]), .Z(n4287) );
  XNOR U5313 ( .A(n4288), .B(n4289), .Z(o[785]) );
  XOR U5314 ( .A(n4290), .B(o[784]), .Z(creg_next[784]) );
  AND U5315 ( .A(n3090), .B(n4291), .Z(n4290) );
  XNOR U5316 ( .A(c[784]), .B(n4292), .Z(n4291) );
  IV U5317 ( .A(o[784]), .Z(n4292) );
  XNOR U5318 ( .A(n4293), .B(n4294), .Z(o[784]) );
  XOR U5319 ( .A(n4295), .B(o[783]), .Z(creg_next[783]) );
  AND U5320 ( .A(n3090), .B(n4296), .Z(n4295) );
  XNOR U5321 ( .A(c[783]), .B(n4297), .Z(n4296) );
  IV U5322 ( .A(o[783]), .Z(n4297) );
  XNOR U5323 ( .A(n4298), .B(n4299), .Z(o[783]) );
  XOR U5324 ( .A(n4300), .B(o[782]), .Z(creg_next[782]) );
  AND U5325 ( .A(n3090), .B(n4301), .Z(n4300) );
  XNOR U5326 ( .A(c[782]), .B(n4302), .Z(n4301) );
  IV U5327 ( .A(o[782]), .Z(n4302) );
  XNOR U5328 ( .A(n4303), .B(n4304), .Z(o[782]) );
  XOR U5329 ( .A(n4305), .B(o[781]), .Z(creg_next[781]) );
  AND U5330 ( .A(n3090), .B(n4306), .Z(n4305) );
  XNOR U5331 ( .A(c[781]), .B(n4307), .Z(n4306) );
  IV U5332 ( .A(o[781]), .Z(n4307) );
  XNOR U5333 ( .A(n4308), .B(n4309), .Z(o[781]) );
  XOR U5334 ( .A(n4310), .B(o[780]), .Z(creg_next[780]) );
  AND U5335 ( .A(n3090), .B(n4311), .Z(n4310) );
  XNOR U5336 ( .A(c[780]), .B(n4312), .Z(n4311) );
  IV U5337 ( .A(o[780]), .Z(n4312) );
  XNOR U5338 ( .A(n4313), .B(n4314), .Z(o[780]) );
  XOR U5339 ( .A(n4315), .B(o[77]), .Z(creg_next[77]) );
  AND U5340 ( .A(n3090), .B(n4316), .Z(n4315) );
  XNOR U5341 ( .A(c[77]), .B(n4317), .Z(n4316) );
  IV U5342 ( .A(o[77]), .Z(n4317) );
  XNOR U5343 ( .A(n4318), .B(n4319), .Z(o[77]) );
  XOR U5344 ( .A(n4320), .B(o[779]), .Z(creg_next[779]) );
  AND U5345 ( .A(n3090), .B(n4321), .Z(n4320) );
  XNOR U5346 ( .A(c[779]), .B(n4322), .Z(n4321) );
  IV U5347 ( .A(o[779]), .Z(n4322) );
  XNOR U5348 ( .A(n4323), .B(n4324), .Z(o[779]) );
  XOR U5349 ( .A(n4325), .B(o[778]), .Z(creg_next[778]) );
  AND U5350 ( .A(n3090), .B(n4326), .Z(n4325) );
  XNOR U5351 ( .A(c[778]), .B(n4327), .Z(n4326) );
  IV U5352 ( .A(o[778]), .Z(n4327) );
  XNOR U5353 ( .A(n4328), .B(n4329), .Z(o[778]) );
  XOR U5354 ( .A(n4330), .B(o[777]), .Z(creg_next[777]) );
  AND U5355 ( .A(n3090), .B(n4331), .Z(n4330) );
  XNOR U5356 ( .A(c[777]), .B(n4332), .Z(n4331) );
  IV U5357 ( .A(o[777]), .Z(n4332) );
  XNOR U5358 ( .A(n4333), .B(n4334), .Z(o[777]) );
  XOR U5359 ( .A(n4335), .B(o[776]), .Z(creg_next[776]) );
  AND U5360 ( .A(n3090), .B(n4336), .Z(n4335) );
  XNOR U5361 ( .A(c[776]), .B(n4337), .Z(n4336) );
  IV U5362 ( .A(o[776]), .Z(n4337) );
  XNOR U5363 ( .A(n4338), .B(n4339), .Z(o[776]) );
  XOR U5364 ( .A(n4340), .B(o[775]), .Z(creg_next[775]) );
  AND U5365 ( .A(n3090), .B(n4341), .Z(n4340) );
  XNOR U5366 ( .A(c[775]), .B(n4342), .Z(n4341) );
  IV U5367 ( .A(o[775]), .Z(n4342) );
  XNOR U5368 ( .A(n4343), .B(n4344), .Z(o[775]) );
  XOR U5369 ( .A(n4345), .B(o[774]), .Z(creg_next[774]) );
  AND U5370 ( .A(n3090), .B(n4346), .Z(n4345) );
  XNOR U5371 ( .A(c[774]), .B(n4347), .Z(n4346) );
  IV U5372 ( .A(o[774]), .Z(n4347) );
  XNOR U5373 ( .A(n4348), .B(n4349), .Z(o[774]) );
  XOR U5374 ( .A(n4350), .B(o[773]), .Z(creg_next[773]) );
  AND U5375 ( .A(n3090), .B(n4351), .Z(n4350) );
  XNOR U5376 ( .A(c[773]), .B(n4352), .Z(n4351) );
  IV U5377 ( .A(o[773]), .Z(n4352) );
  XNOR U5378 ( .A(n4353), .B(n4354), .Z(o[773]) );
  XOR U5379 ( .A(n4355), .B(o[772]), .Z(creg_next[772]) );
  AND U5380 ( .A(n3090), .B(n4356), .Z(n4355) );
  XNOR U5381 ( .A(c[772]), .B(n4357), .Z(n4356) );
  IV U5382 ( .A(o[772]), .Z(n4357) );
  XNOR U5383 ( .A(n4358), .B(n4359), .Z(o[772]) );
  XOR U5384 ( .A(n4360), .B(o[771]), .Z(creg_next[771]) );
  AND U5385 ( .A(n3090), .B(n4361), .Z(n4360) );
  XNOR U5386 ( .A(c[771]), .B(n4362), .Z(n4361) );
  IV U5387 ( .A(o[771]), .Z(n4362) );
  XNOR U5388 ( .A(n4363), .B(n4364), .Z(o[771]) );
  XOR U5389 ( .A(n4365), .B(o[770]), .Z(creg_next[770]) );
  AND U5390 ( .A(n3090), .B(n4366), .Z(n4365) );
  XNOR U5391 ( .A(c[770]), .B(n4367), .Z(n4366) );
  IV U5392 ( .A(o[770]), .Z(n4367) );
  XNOR U5393 ( .A(n4368), .B(n4369), .Z(o[770]) );
  XOR U5394 ( .A(n4370), .B(o[76]), .Z(creg_next[76]) );
  AND U5395 ( .A(n3090), .B(n4371), .Z(n4370) );
  XNOR U5396 ( .A(c[76]), .B(n4372), .Z(n4371) );
  IV U5397 ( .A(o[76]), .Z(n4372) );
  XNOR U5398 ( .A(n4373), .B(n4374), .Z(o[76]) );
  XOR U5399 ( .A(n4375), .B(o[769]), .Z(creg_next[769]) );
  AND U5400 ( .A(n3090), .B(n4376), .Z(n4375) );
  XNOR U5401 ( .A(c[769]), .B(n4377), .Z(n4376) );
  IV U5402 ( .A(o[769]), .Z(n4377) );
  XNOR U5403 ( .A(n4378), .B(n4379), .Z(o[769]) );
  XOR U5404 ( .A(n4380), .B(o[768]), .Z(creg_next[768]) );
  AND U5405 ( .A(n3090), .B(n4381), .Z(n4380) );
  XNOR U5406 ( .A(c[768]), .B(n4382), .Z(n4381) );
  IV U5407 ( .A(o[768]), .Z(n4382) );
  XNOR U5408 ( .A(n4383), .B(n4384), .Z(o[768]) );
  XOR U5409 ( .A(n4385), .B(o[767]), .Z(creg_next[767]) );
  AND U5410 ( .A(n3090), .B(n4386), .Z(n4385) );
  XNOR U5411 ( .A(c[767]), .B(n4387), .Z(n4386) );
  IV U5412 ( .A(o[767]), .Z(n4387) );
  XNOR U5413 ( .A(n4388), .B(n4389), .Z(o[767]) );
  XOR U5414 ( .A(n4390), .B(o[766]), .Z(creg_next[766]) );
  AND U5415 ( .A(n3090), .B(n4391), .Z(n4390) );
  XNOR U5416 ( .A(c[766]), .B(n4392), .Z(n4391) );
  IV U5417 ( .A(o[766]), .Z(n4392) );
  XNOR U5418 ( .A(n4393), .B(n4394), .Z(o[766]) );
  XOR U5419 ( .A(n4395), .B(o[765]), .Z(creg_next[765]) );
  AND U5420 ( .A(n3090), .B(n4396), .Z(n4395) );
  XNOR U5421 ( .A(c[765]), .B(n4397), .Z(n4396) );
  IV U5422 ( .A(o[765]), .Z(n4397) );
  XNOR U5423 ( .A(n4398), .B(n4399), .Z(o[765]) );
  XOR U5424 ( .A(n4400), .B(o[764]), .Z(creg_next[764]) );
  AND U5425 ( .A(n3090), .B(n4401), .Z(n4400) );
  XNOR U5426 ( .A(c[764]), .B(n4402), .Z(n4401) );
  IV U5427 ( .A(o[764]), .Z(n4402) );
  XNOR U5428 ( .A(n4403), .B(n4404), .Z(o[764]) );
  XOR U5429 ( .A(n4405), .B(o[763]), .Z(creg_next[763]) );
  AND U5430 ( .A(n3090), .B(n4406), .Z(n4405) );
  XNOR U5431 ( .A(c[763]), .B(n4407), .Z(n4406) );
  IV U5432 ( .A(o[763]), .Z(n4407) );
  XNOR U5433 ( .A(n4408), .B(n4409), .Z(o[763]) );
  XOR U5434 ( .A(n4410), .B(o[762]), .Z(creg_next[762]) );
  AND U5435 ( .A(n3090), .B(n4411), .Z(n4410) );
  XNOR U5436 ( .A(c[762]), .B(n4412), .Z(n4411) );
  IV U5437 ( .A(o[762]), .Z(n4412) );
  XNOR U5438 ( .A(n4413), .B(n4414), .Z(o[762]) );
  XOR U5439 ( .A(n4415), .B(o[761]), .Z(creg_next[761]) );
  AND U5440 ( .A(n3090), .B(n4416), .Z(n4415) );
  XNOR U5441 ( .A(c[761]), .B(n4417), .Z(n4416) );
  IV U5442 ( .A(o[761]), .Z(n4417) );
  XNOR U5443 ( .A(n4418), .B(n4419), .Z(o[761]) );
  XOR U5444 ( .A(n4420), .B(o[760]), .Z(creg_next[760]) );
  AND U5445 ( .A(n3090), .B(n4421), .Z(n4420) );
  XNOR U5446 ( .A(c[760]), .B(n4422), .Z(n4421) );
  IV U5447 ( .A(o[760]), .Z(n4422) );
  XNOR U5448 ( .A(n4423), .B(n4424), .Z(o[760]) );
  XOR U5449 ( .A(n4425), .B(o[75]), .Z(creg_next[75]) );
  AND U5450 ( .A(n3090), .B(n4426), .Z(n4425) );
  XNOR U5451 ( .A(c[75]), .B(n4427), .Z(n4426) );
  IV U5452 ( .A(o[75]), .Z(n4427) );
  XNOR U5453 ( .A(n4428), .B(n4429), .Z(o[75]) );
  XOR U5454 ( .A(n4430), .B(o[759]), .Z(creg_next[759]) );
  AND U5455 ( .A(n3090), .B(n4431), .Z(n4430) );
  XNOR U5456 ( .A(c[759]), .B(n4432), .Z(n4431) );
  IV U5457 ( .A(o[759]), .Z(n4432) );
  XNOR U5458 ( .A(n4433), .B(n4434), .Z(o[759]) );
  XOR U5459 ( .A(n4435), .B(o[758]), .Z(creg_next[758]) );
  AND U5460 ( .A(n3090), .B(n4436), .Z(n4435) );
  XNOR U5461 ( .A(c[758]), .B(n4437), .Z(n4436) );
  IV U5462 ( .A(o[758]), .Z(n4437) );
  XNOR U5463 ( .A(n4438), .B(n4439), .Z(o[758]) );
  XOR U5464 ( .A(n4440), .B(o[757]), .Z(creg_next[757]) );
  AND U5465 ( .A(n3090), .B(n4441), .Z(n4440) );
  XNOR U5466 ( .A(c[757]), .B(n4442), .Z(n4441) );
  IV U5467 ( .A(o[757]), .Z(n4442) );
  XNOR U5468 ( .A(n4443), .B(n4444), .Z(o[757]) );
  XOR U5469 ( .A(n4445), .B(o[756]), .Z(creg_next[756]) );
  AND U5470 ( .A(n3090), .B(n4446), .Z(n4445) );
  XNOR U5471 ( .A(c[756]), .B(n4447), .Z(n4446) );
  IV U5472 ( .A(o[756]), .Z(n4447) );
  XNOR U5473 ( .A(n4448), .B(n4449), .Z(o[756]) );
  XOR U5474 ( .A(n4450), .B(o[755]), .Z(creg_next[755]) );
  AND U5475 ( .A(n3090), .B(n4451), .Z(n4450) );
  XNOR U5476 ( .A(c[755]), .B(n4452), .Z(n4451) );
  IV U5477 ( .A(o[755]), .Z(n4452) );
  XNOR U5478 ( .A(n4453), .B(n4454), .Z(o[755]) );
  XOR U5479 ( .A(n4455), .B(o[754]), .Z(creg_next[754]) );
  AND U5480 ( .A(n3090), .B(n4456), .Z(n4455) );
  XNOR U5481 ( .A(c[754]), .B(n4457), .Z(n4456) );
  IV U5482 ( .A(o[754]), .Z(n4457) );
  XNOR U5483 ( .A(n4458), .B(n4459), .Z(o[754]) );
  XOR U5484 ( .A(n4460), .B(o[753]), .Z(creg_next[753]) );
  AND U5485 ( .A(n3090), .B(n4461), .Z(n4460) );
  XNOR U5486 ( .A(c[753]), .B(n4462), .Z(n4461) );
  IV U5487 ( .A(o[753]), .Z(n4462) );
  XNOR U5488 ( .A(n4463), .B(n4464), .Z(o[753]) );
  XOR U5489 ( .A(n4465), .B(o[752]), .Z(creg_next[752]) );
  AND U5490 ( .A(n3090), .B(n4466), .Z(n4465) );
  XNOR U5491 ( .A(c[752]), .B(n4467), .Z(n4466) );
  IV U5492 ( .A(o[752]), .Z(n4467) );
  XNOR U5493 ( .A(n4468), .B(n4469), .Z(o[752]) );
  XOR U5494 ( .A(n4470), .B(o[751]), .Z(creg_next[751]) );
  AND U5495 ( .A(n3090), .B(n4471), .Z(n4470) );
  XNOR U5496 ( .A(c[751]), .B(n4472), .Z(n4471) );
  IV U5497 ( .A(o[751]), .Z(n4472) );
  XNOR U5498 ( .A(n4473), .B(n4474), .Z(o[751]) );
  XOR U5499 ( .A(n4475), .B(o[750]), .Z(creg_next[750]) );
  AND U5500 ( .A(n3090), .B(n4476), .Z(n4475) );
  XNOR U5501 ( .A(c[750]), .B(n4477), .Z(n4476) );
  IV U5502 ( .A(o[750]), .Z(n4477) );
  XNOR U5503 ( .A(n4478), .B(n4479), .Z(o[750]) );
  XOR U5504 ( .A(n4480), .B(o[74]), .Z(creg_next[74]) );
  AND U5505 ( .A(n3090), .B(n4481), .Z(n4480) );
  XNOR U5506 ( .A(c[74]), .B(n4482), .Z(n4481) );
  IV U5507 ( .A(o[74]), .Z(n4482) );
  XNOR U5508 ( .A(n4483), .B(n4484), .Z(o[74]) );
  XOR U5509 ( .A(n4485), .B(o[749]), .Z(creg_next[749]) );
  AND U5510 ( .A(n3090), .B(n4486), .Z(n4485) );
  XNOR U5511 ( .A(c[749]), .B(n4487), .Z(n4486) );
  IV U5512 ( .A(o[749]), .Z(n4487) );
  XNOR U5513 ( .A(n4488), .B(n4489), .Z(o[749]) );
  XOR U5514 ( .A(n4490), .B(o[748]), .Z(creg_next[748]) );
  AND U5515 ( .A(n3090), .B(n4491), .Z(n4490) );
  XNOR U5516 ( .A(c[748]), .B(n4492), .Z(n4491) );
  IV U5517 ( .A(o[748]), .Z(n4492) );
  XNOR U5518 ( .A(n4493), .B(n4494), .Z(o[748]) );
  XOR U5519 ( .A(n4495), .B(o[747]), .Z(creg_next[747]) );
  AND U5520 ( .A(n3090), .B(n4496), .Z(n4495) );
  XNOR U5521 ( .A(c[747]), .B(n4497), .Z(n4496) );
  IV U5522 ( .A(o[747]), .Z(n4497) );
  XNOR U5523 ( .A(n4498), .B(n4499), .Z(o[747]) );
  XOR U5524 ( .A(n4500), .B(o[746]), .Z(creg_next[746]) );
  AND U5525 ( .A(n3090), .B(n4501), .Z(n4500) );
  XNOR U5526 ( .A(c[746]), .B(n4502), .Z(n4501) );
  IV U5527 ( .A(o[746]), .Z(n4502) );
  XNOR U5528 ( .A(n4503), .B(n4504), .Z(o[746]) );
  XOR U5529 ( .A(n4505), .B(o[745]), .Z(creg_next[745]) );
  AND U5530 ( .A(n3090), .B(n4506), .Z(n4505) );
  XNOR U5531 ( .A(c[745]), .B(n4507), .Z(n4506) );
  IV U5532 ( .A(o[745]), .Z(n4507) );
  XNOR U5533 ( .A(n4508), .B(n4509), .Z(o[745]) );
  XOR U5534 ( .A(n4510), .B(o[744]), .Z(creg_next[744]) );
  AND U5535 ( .A(n3090), .B(n4511), .Z(n4510) );
  XNOR U5536 ( .A(c[744]), .B(n4512), .Z(n4511) );
  IV U5537 ( .A(o[744]), .Z(n4512) );
  XNOR U5538 ( .A(n4513), .B(n4514), .Z(o[744]) );
  XOR U5539 ( .A(n4515), .B(o[743]), .Z(creg_next[743]) );
  AND U5540 ( .A(n3090), .B(n4516), .Z(n4515) );
  XNOR U5541 ( .A(c[743]), .B(n4517), .Z(n4516) );
  IV U5542 ( .A(o[743]), .Z(n4517) );
  XNOR U5543 ( .A(n4518), .B(n4519), .Z(o[743]) );
  XOR U5544 ( .A(n4520), .B(o[742]), .Z(creg_next[742]) );
  AND U5545 ( .A(n3090), .B(n4521), .Z(n4520) );
  XNOR U5546 ( .A(c[742]), .B(n4522), .Z(n4521) );
  IV U5547 ( .A(o[742]), .Z(n4522) );
  XNOR U5548 ( .A(n4523), .B(n4524), .Z(o[742]) );
  XOR U5549 ( .A(n4525), .B(o[741]), .Z(creg_next[741]) );
  AND U5550 ( .A(n3090), .B(n4526), .Z(n4525) );
  XNOR U5551 ( .A(c[741]), .B(n4527), .Z(n4526) );
  IV U5552 ( .A(o[741]), .Z(n4527) );
  XNOR U5553 ( .A(n4528), .B(n4529), .Z(o[741]) );
  XOR U5554 ( .A(n4530), .B(o[740]), .Z(creg_next[740]) );
  AND U5555 ( .A(n3090), .B(n4531), .Z(n4530) );
  XNOR U5556 ( .A(c[740]), .B(n4532), .Z(n4531) );
  IV U5557 ( .A(o[740]), .Z(n4532) );
  XNOR U5558 ( .A(n4533), .B(n4534), .Z(o[740]) );
  XOR U5559 ( .A(n4535), .B(o[73]), .Z(creg_next[73]) );
  AND U5560 ( .A(n3090), .B(n4536), .Z(n4535) );
  XNOR U5561 ( .A(c[73]), .B(n4537), .Z(n4536) );
  IV U5562 ( .A(o[73]), .Z(n4537) );
  XNOR U5563 ( .A(n4538), .B(n4539), .Z(o[73]) );
  XOR U5564 ( .A(n4540), .B(o[739]), .Z(creg_next[739]) );
  AND U5565 ( .A(n3090), .B(n4541), .Z(n4540) );
  XNOR U5566 ( .A(c[739]), .B(n4542), .Z(n4541) );
  IV U5567 ( .A(o[739]), .Z(n4542) );
  XNOR U5568 ( .A(n4543), .B(n4544), .Z(o[739]) );
  XOR U5569 ( .A(n4545), .B(o[738]), .Z(creg_next[738]) );
  AND U5570 ( .A(n3090), .B(n4546), .Z(n4545) );
  XNOR U5571 ( .A(c[738]), .B(n4547), .Z(n4546) );
  IV U5572 ( .A(o[738]), .Z(n4547) );
  XNOR U5573 ( .A(n4548), .B(n4549), .Z(o[738]) );
  XOR U5574 ( .A(n4550), .B(o[737]), .Z(creg_next[737]) );
  AND U5575 ( .A(n3090), .B(n4551), .Z(n4550) );
  XNOR U5576 ( .A(c[737]), .B(n4552), .Z(n4551) );
  IV U5577 ( .A(o[737]), .Z(n4552) );
  XNOR U5578 ( .A(n4553), .B(n4554), .Z(o[737]) );
  XOR U5579 ( .A(n4555), .B(o[736]), .Z(creg_next[736]) );
  AND U5580 ( .A(n3090), .B(n4556), .Z(n4555) );
  XNOR U5581 ( .A(c[736]), .B(n4557), .Z(n4556) );
  IV U5582 ( .A(o[736]), .Z(n4557) );
  XNOR U5583 ( .A(n4558), .B(n4559), .Z(o[736]) );
  XOR U5584 ( .A(n4560), .B(o[735]), .Z(creg_next[735]) );
  AND U5585 ( .A(n3090), .B(n4561), .Z(n4560) );
  XNOR U5586 ( .A(c[735]), .B(n4562), .Z(n4561) );
  IV U5587 ( .A(o[735]), .Z(n4562) );
  XNOR U5588 ( .A(n4563), .B(n4564), .Z(o[735]) );
  XOR U5589 ( .A(n4565), .B(o[734]), .Z(creg_next[734]) );
  AND U5590 ( .A(n3090), .B(n4566), .Z(n4565) );
  XNOR U5591 ( .A(c[734]), .B(n4567), .Z(n4566) );
  IV U5592 ( .A(o[734]), .Z(n4567) );
  XNOR U5593 ( .A(n4568), .B(n4569), .Z(o[734]) );
  XOR U5594 ( .A(n4570), .B(o[733]), .Z(creg_next[733]) );
  AND U5595 ( .A(n3090), .B(n4571), .Z(n4570) );
  XNOR U5596 ( .A(c[733]), .B(n4572), .Z(n4571) );
  IV U5597 ( .A(o[733]), .Z(n4572) );
  XNOR U5598 ( .A(n4573), .B(n4574), .Z(o[733]) );
  XOR U5599 ( .A(n4575), .B(o[732]), .Z(creg_next[732]) );
  AND U5600 ( .A(n3090), .B(n4576), .Z(n4575) );
  XNOR U5601 ( .A(c[732]), .B(n4577), .Z(n4576) );
  IV U5602 ( .A(o[732]), .Z(n4577) );
  XNOR U5603 ( .A(n4578), .B(n4579), .Z(o[732]) );
  XOR U5604 ( .A(n4580), .B(o[731]), .Z(creg_next[731]) );
  AND U5605 ( .A(n3090), .B(n4581), .Z(n4580) );
  XNOR U5606 ( .A(c[731]), .B(n4582), .Z(n4581) );
  IV U5607 ( .A(o[731]), .Z(n4582) );
  XNOR U5608 ( .A(n4583), .B(n4584), .Z(o[731]) );
  XOR U5609 ( .A(n4585), .B(o[730]), .Z(creg_next[730]) );
  AND U5610 ( .A(n3090), .B(n4586), .Z(n4585) );
  XNOR U5611 ( .A(c[730]), .B(n4587), .Z(n4586) );
  IV U5612 ( .A(o[730]), .Z(n4587) );
  XNOR U5613 ( .A(n4588), .B(n4589), .Z(o[730]) );
  XOR U5614 ( .A(n4590), .B(o[72]), .Z(creg_next[72]) );
  AND U5615 ( .A(n3090), .B(n4591), .Z(n4590) );
  XNOR U5616 ( .A(c[72]), .B(n4592), .Z(n4591) );
  IV U5617 ( .A(o[72]), .Z(n4592) );
  XNOR U5618 ( .A(n4593), .B(n4594), .Z(o[72]) );
  XOR U5619 ( .A(n4595), .B(o[729]), .Z(creg_next[729]) );
  AND U5620 ( .A(n3090), .B(n4596), .Z(n4595) );
  XNOR U5621 ( .A(c[729]), .B(n4597), .Z(n4596) );
  IV U5622 ( .A(o[729]), .Z(n4597) );
  XNOR U5623 ( .A(n4598), .B(n4599), .Z(o[729]) );
  XOR U5624 ( .A(n4600), .B(o[728]), .Z(creg_next[728]) );
  AND U5625 ( .A(n3090), .B(n4601), .Z(n4600) );
  XNOR U5626 ( .A(c[728]), .B(n4602), .Z(n4601) );
  IV U5627 ( .A(o[728]), .Z(n4602) );
  XNOR U5628 ( .A(n4603), .B(n4604), .Z(o[728]) );
  XOR U5629 ( .A(n4605), .B(o[727]), .Z(creg_next[727]) );
  AND U5630 ( .A(n3090), .B(n4606), .Z(n4605) );
  XNOR U5631 ( .A(c[727]), .B(n4607), .Z(n4606) );
  IV U5632 ( .A(o[727]), .Z(n4607) );
  XNOR U5633 ( .A(n4608), .B(n4609), .Z(o[727]) );
  XOR U5634 ( .A(n4610), .B(o[726]), .Z(creg_next[726]) );
  AND U5635 ( .A(n3090), .B(n4611), .Z(n4610) );
  XNOR U5636 ( .A(c[726]), .B(n4612), .Z(n4611) );
  IV U5637 ( .A(o[726]), .Z(n4612) );
  XNOR U5638 ( .A(n4613), .B(n4614), .Z(o[726]) );
  XOR U5639 ( .A(n4615), .B(o[725]), .Z(creg_next[725]) );
  AND U5640 ( .A(n3090), .B(n4616), .Z(n4615) );
  XNOR U5641 ( .A(c[725]), .B(n4617), .Z(n4616) );
  IV U5642 ( .A(o[725]), .Z(n4617) );
  XNOR U5643 ( .A(n4618), .B(n4619), .Z(o[725]) );
  XOR U5644 ( .A(n4620), .B(o[724]), .Z(creg_next[724]) );
  AND U5645 ( .A(n3090), .B(n4621), .Z(n4620) );
  XNOR U5646 ( .A(c[724]), .B(n4622), .Z(n4621) );
  IV U5647 ( .A(o[724]), .Z(n4622) );
  XNOR U5648 ( .A(n4623), .B(n4624), .Z(o[724]) );
  XOR U5649 ( .A(n4625), .B(o[723]), .Z(creg_next[723]) );
  AND U5650 ( .A(n3090), .B(n4626), .Z(n4625) );
  XNOR U5651 ( .A(c[723]), .B(n4627), .Z(n4626) );
  IV U5652 ( .A(o[723]), .Z(n4627) );
  XNOR U5653 ( .A(n4628), .B(n4629), .Z(o[723]) );
  XOR U5654 ( .A(n4630), .B(o[722]), .Z(creg_next[722]) );
  AND U5655 ( .A(n3090), .B(n4631), .Z(n4630) );
  XNOR U5656 ( .A(c[722]), .B(n4632), .Z(n4631) );
  IV U5657 ( .A(o[722]), .Z(n4632) );
  XNOR U5658 ( .A(n4633), .B(n4634), .Z(o[722]) );
  XOR U5659 ( .A(n4635), .B(o[721]), .Z(creg_next[721]) );
  AND U5660 ( .A(n3090), .B(n4636), .Z(n4635) );
  XNOR U5661 ( .A(c[721]), .B(n4637), .Z(n4636) );
  IV U5662 ( .A(o[721]), .Z(n4637) );
  XNOR U5663 ( .A(n4638), .B(n4639), .Z(o[721]) );
  XOR U5664 ( .A(n4640), .B(o[720]), .Z(creg_next[720]) );
  AND U5665 ( .A(n3090), .B(n4641), .Z(n4640) );
  XNOR U5666 ( .A(c[720]), .B(n4642), .Z(n4641) );
  IV U5667 ( .A(o[720]), .Z(n4642) );
  XNOR U5668 ( .A(n4643), .B(n4644), .Z(o[720]) );
  XOR U5669 ( .A(n4645), .B(o[71]), .Z(creg_next[71]) );
  AND U5670 ( .A(n3090), .B(n4646), .Z(n4645) );
  XNOR U5671 ( .A(c[71]), .B(n4647), .Z(n4646) );
  IV U5672 ( .A(o[71]), .Z(n4647) );
  XNOR U5673 ( .A(n4648), .B(n4649), .Z(o[71]) );
  XOR U5674 ( .A(n4650), .B(o[719]), .Z(creg_next[719]) );
  AND U5675 ( .A(n3090), .B(n4651), .Z(n4650) );
  XNOR U5676 ( .A(c[719]), .B(n4652), .Z(n4651) );
  IV U5677 ( .A(o[719]), .Z(n4652) );
  XNOR U5678 ( .A(n4653), .B(n4654), .Z(o[719]) );
  XOR U5679 ( .A(n4655), .B(o[718]), .Z(creg_next[718]) );
  AND U5680 ( .A(n3090), .B(n4656), .Z(n4655) );
  XNOR U5681 ( .A(c[718]), .B(n4657), .Z(n4656) );
  IV U5682 ( .A(o[718]), .Z(n4657) );
  XNOR U5683 ( .A(n4658), .B(n4659), .Z(o[718]) );
  XOR U5684 ( .A(n4660), .B(o[717]), .Z(creg_next[717]) );
  AND U5685 ( .A(n3090), .B(n4661), .Z(n4660) );
  XNOR U5686 ( .A(c[717]), .B(n4662), .Z(n4661) );
  IV U5687 ( .A(o[717]), .Z(n4662) );
  XNOR U5688 ( .A(n4663), .B(n4664), .Z(o[717]) );
  XOR U5689 ( .A(n4665), .B(o[716]), .Z(creg_next[716]) );
  AND U5690 ( .A(n3090), .B(n4666), .Z(n4665) );
  XNOR U5691 ( .A(c[716]), .B(n4667), .Z(n4666) );
  IV U5692 ( .A(o[716]), .Z(n4667) );
  XNOR U5693 ( .A(n4668), .B(n4669), .Z(o[716]) );
  XOR U5694 ( .A(n4670), .B(o[715]), .Z(creg_next[715]) );
  AND U5695 ( .A(n3090), .B(n4671), .Z(n4670) );
  XNOR U5696 ( .A(c[715]), .B(n4672), .Z(n4671) );
  IV U5697 ( .A(o[715]), .Z(n4672) );
  XNOR U5698 ( .A(n4673), .B(n4674), .Z(o[715]) );
  XOR U5699 ( .A(n4675), .B(o[714]), .Z(creg_next[714]) );
  AND U5700 ( .A(n3090), .B(n4676), .Z(n4675) );
  XNOR U5701 ( .A(c[714]), .B(n4677), .Z(n4676) );
  IV U5702 ( .A(o[714]), .Z(n4677) );
  XNOR U5703 ( .A(n4678), .B(n4679), .Z(o[714]) );
  XOR U5704 ( .A(n4680), .B(o[713]), .Z(creg_next[713]) );
  AND U5705 ( .A(n3090), .B(n4681), .Z(n4680) );
  XNOR U5706 ( .A(c[713]), .B(n4682), .Z(n4681) );
  IV U5707 ( .A(o[713]), .Z(n4682) );
  XNOR U5708 ( .A(n4683), .B(n4684), .Z(o[713]) );
  XOR U5709 ( .A(n4685), .B(o[712]), .Z(creg_next[712]) );
  AND U5710 ( .A(n3090), .B(n4686), .Z(n4685) );
  XNOR U5711 ( .A(c[712]), .B(n4687), .Z(n4686) );
  IV U5712 ( .A(o[712]), .Z(n4687) );
  XNOR U5713 ( .A(n4688), .B(n4689), .Z(o[712]) );
  XOR U5714 ( .A(n4690), .B(o[711]), .Z(creg_next[711]) );
  AND U5715 ( .A(n3090), .B(n4691), .Z(n4690) );
  XNOR U5716 ( .A(c[711]), .B(n4692), .Z(n4691) );
  IV U5717 ( .A(o[711]), .Z(n4692) );
  XNOR U5718 ( .A(n4693), .B(n4694), .Z(o[711]) );
  XOR U5719 ( .A(n4695), .B(o[710]), .Z(creg_next[710]) );
  AND U5720 ( .A(n3090), .B(n4696), .Z(n4695) );
  XNOR U5721 ( .A(c[710]), .B(n4697), .Z(n4696) );
  IV U5722 ( .A(o[710]), .Z(n4697) );
  XNOR U5723 ( .A(n4698), .B(n4699), .Z(o[710]) );
  XOR U5724 ( .A(n4700), .B(o[70]), .Z(creg_next[70]) );
  AND U5725 ( .A(n3090), .B(n4701), .Z(n4700) );
  XNOR U5726 ( .A(c[70]), .B(n4702), .Z(n4701) );
  IV U5727 ( .A(o[70]), .Z(n4702) );
  XNOR U5728 ( .A(n4703), .B(n4704), .Z(o[70]) );
  XOR U5729 ( .A(n4705), .B(o[709]), .Z(creg_next[709]) );
  AND U5730 ( .A(n3090), .B(n4706), .Z(n4705) );
  XNOR U5731 ( .A(c[709]), .B(n4707), .Z(n4706) );
  IV U5732 ( .A(o[709]), .Z(n4707) );
  XNOR U5733 ( .A(n4708), .B(n4709), .Z(o[709]) );
  XOR U5734 ( .A(n4710), .B(o[708]), .Z(creg_next[708]) );
  AND U5735 ( .A(n3090), .B(n4711), .Z(n4710) );
  XNOR U5736 ( .A(c[708]), .B(n4712), .Z(n4711) );
  IV U5737 ( .A(o[708]), .Z(n4712) );
  XNOR U5738 ( .A(n4713), .B(n4714), .Z(o[708]) );
  XOR U5739 ( .A(n4715), .B(o[707]), .Z(creg_next[707]) );
  AND U5740 ( .A(n3090), .B(n4716), .Z(n4715) );
  XNOR U5741 ( .A(c[707]), .B(n4717), .Z(n4716) );
  IV U5742 ( .A(o[707]), .Z(n4717) );
  XNOR U5743 ( .A(n4718), .B(n4719), .Z(o[707]) );
  XOR U5744 ( .A(n4720), .B(o[706]), .Z(creg_next[706]) );
  AND U5745 ( .A(n3090), .B(n4721), .Z(n4720) );
  XNOR U5746 ( .A(c[706]), .B(n4722), .Z(n4721) );
  IV U5747 ( .A(o[706]), .Z(n4722) );
  XNOR U5748 ( .A(n4723), .B(n4724), .Z(o[706]) );
  XOR U5749 ( .A(n4725), .B(o[705]), .Z(creg_next[705]) );
  AND U5750 ( .A(n3090), .B(n4726), .Z(n4725) );
  XNOR U5751 ( .A(c[705]), .B(n4727), .Z(n4726) );
  IV U5752 ( .A(o[705]), .Z(n4727) );
  XNOR U5753 ( .A(n4728), .B(n4729), .Z(o[705]) );
  XOR U5754 ( .A(n4730), .B(o[704]), .Z(creg_next[704]) );
  AND U5755 ( .A(n3090), .B(n4731), .Z(n4730) );
  XNOR U5756 ( .A(c[704]), .B(n4732), .Z(n4731) );
  IV U5757 ( .A(o[704]), .Z(n4732) );
  XNOR U5758 ( .A(n4733), .B(n4734), .Z(o[704]) );
  XOR U5759 ( .A(n4735), .B(o[703]), .Z(creg_next[703]) );
  AND U5760 ( .A(n3090), .B(n4736), .Z(n4735) );
  XNOR U5761 ( .A(c[703]), .B(n4737), .Z(n4736) );
  IV U5762 ( .A(o[703]), .Z(n4737) );
  XNOR U5763 ( .A(n4738), .B(n4739), .Z(o[703]) );
  XOR U5764 ( .A(n4740), .B(o[702]), .Z(creg_next[702]) );
  AND U5765 ( .A(n3090), .B(n4741), .Z(n4740) );
  XNOR U5766 ( .A(c[702]), .B(n4742), .Z(n4741) );
  IV U5767 ( .A(o[702]), .Z(n4742) );
  XNOR U5768 ( .A(n4743), .B(n4744), .Z(o[702]) );
  XOR U5769 ( .A(n4745), .B(o[701]), .Z(creg_next[701]) );
  AND U5770 ( .A(n3090), .B(n4746), .Z(n4745) );
  XNOR U5771 ( .A(c[701]), .B(n4747), .Z(n4746) );
  IV U5772 ( .A(o[701]), .Z(n4747) );
  XNOR U5773 ( .A(n4748), .B(n4749), .Z(o[701]) );
  XOR U5774 ( .A(n4750), .B(o[700]), .Z(creg_next[700]) );
  AND U5775 ( .A(n3090), .B(n4751), .Z(n4750) );
  XNOR U5776 ( .A(c[700]), .B(n4752), .Z(n4751) );
  IV U5777 ( .A(o[700]), .Z(n4752) );
  XNOR U5778 ( .A(n4753), .B(n4754), .Z(o[700]) );
  XOR U5779 ( .A(n4755), .B(o[6]), .Z(creg_next[6]) );
  AND U5780 ( .A(n3090), .B(n4756), .Z(n4755) );
  XNOR U5781 ( .A(c[6]), .B(n4757), .Z(n4756) );
  IV U5782 ( .A(o[6]), .Z(n4757) );
  XNOR U5783 ( .A(n4758), .B(n4759), .Z(o[6]) );
  XOR U5784 ( .A(n4760), .B(o[69]), .Z(creg_next[69]) );
  AND U5785 ( .A(n3090), .B(n4761), .Z(n4760) );
  XNOR U5786 ( .A(c[69]), .B(n4762), .Z(n4761) );
  IV U5787 ( .A(o[69]), .Z(n4762) );
  XNOR U5788 ( .A(n4763), .B(n4764), .Z(o[69]) );
  XOR U5789 ( .A(n4765), .B(o[699]), .Z(creg_next[699]) );
  AND U5790 ( .A(n3090), .B(n4766), .Z(n4765) );
  XNOR U5791 ( .A(c[699]), .B(n4767), .Z(n4766) );
  IV U5792 ( .A(o[699]), .Z(n4767) );
  XNOR U5793 ( .A(n4768), .B(n4769), .Z(o[699]) );
  XOR U5794 ( .A(n4770), .B(o[698]), .Z(creg_next[698]) );
  AND U5795 ( .A(n3090), .B(n4771), .Z(n4770) );
  XNOR U5796 ( .A(c[698]), .B(n4772), .Z(n4771) );
  IV U5797 ( .A(o[698]), .Z(n4772) );
  XNOR U5798 ( .A(n4773), .B(n4774), .Z(o[698]) );
  XOR U5799 ( .A(n4775), .B(o[697]), .Z(creg_next[697]) );
  AND U5800 ( .A(n3090), .B(n4776), .Z(n4775) );
  XNOR U5801 ( .A(c[697]), .B(n4777), .Z(n4776) );
  IV U5802 ( .A(o[697]), .Z(n4777) );
  XNOR U5803 ( .A(n4778), .B(n4779), .Z(o[697]) );
  XOR U5804 ( .A(n4780), .B(o[696]), .Z(creg_next[696]) );
  AND U5805 ( .A(n3090), .B(n4781), .Z(n4780) );
  XNOR U5806 ( .A(c[696]), .B(n4782), .Z(n4781) );
  IV U5807 ( .A(o[696]), .Z(n4782) );
  XNOR U5808 ( .A(n4783), .B(n4784), .Z(o[696]) );
  XOR U5809 ( .A(n4785), .B(o[695]), .Z(creg_next[695]) );
  AND U5810 ( .A(n3090), .B(n4786), .Z(n4785) );
  XNOR U5811 ( .A(c[695]), .B(n4787), .Z(n4786) );
  IV U5812 ( .A(o[695]), .Z(n4787) );
  XNOR U5813 ( .A(n4788), .B(n4789), .Z(o[695]) );
  XOR U5814 ( .A(n4790), .B(o[694]), .Z(creg_next[694]) );
  AND U5815 ( .A(n3090), .B(n4791), .Z(n4790) );
  XNOR U5816 ( .A(c[694]), .B(n4792), .Z(n4791) );
  IV U5817 ( .A(o[694]), .Z(n4792) );
  XNOR U5818 ( .A(n4793), .B(n4794), .Z(o[694]) );
  XOR U5819 ( .A(n4795), .B(o[693]), .Z(creg_next[693]) );
  AND U5820 ( .A(n3090), .B(n4796), .Z(n4795) );
  XNOR U5821 ( .A(c[693]), .B(n4797), .Z(n4796) );
  IV U5822 ( .A(o[693]), .Z(n4797) );
  XNOR U5823 ( .A(n4798), .B(n4799), .Z(o[693]) );
  XOR U5824 ( .A(n4800), .B(o[692]), .Z(creg_next[692]) );
  AND U5825 ( .A(n3090), .B(n4801), .Z(n4800) );
  XNOR U5826 ( .A(c[692]), .B(n4802), .Z(n4801) );
  IV U5827 ( .A(o[692]), .Z(n4802) );
  XNOR U5828 ( .A(n4803), .B(n4804), .Z(o[692]) );
  XOR U5829 ( .A(n4805), .B(o[691]), .Z(creg_next[691]) );
  AND U5830 ( .A(n3090), .B(n4806), .Z(n4805) );
  XNOR U5831 ( .A(c[691]), .B(n4807), .Z(n4806) );
  IV U5832 ( .A(o[691]), .Z(n4807) );
  XNOR U5833 ( .A(n4808), .B(n4809), .Z(o[691]) );
  XOR U5834 ( .A(n4810), .B(o[690]), .Z(creg_next[690]) );
  AND U5835 ( .A(n3090), .B(n4811), .Z(n4810) );
  XNOR U5836 ( .A(c[690]), .B(n4812), .Z(n4811) );
  IV U5837 ( .A(o[690]), .Z(n4812) );
  XNOR U5838 ( .A(n4813), .B(n4814), .Z(o[690]) );
  XOR U5839 ( .A(n4815), .B(o[68]), .Z(creg_next[68]) );
  AND U5840 ( .A(n3090), .B(n4816), .Z(n4815) );
  XNOR U5841 ( .A(c[68]), .B(n4817), .Z(n4816) );
  IV U5842 ( .A(o[68]), .Z(n4817) );
  XNOR U5843 ( .A(n4818), .B(n4819), .Z(o[68]) );
  XOR U5844 ( .A(n4820), .B(o[689]), .Z(creg_next[689]) );
  AND U5845 ( .A(n3090), .B(n4821), .Z(n4820) );
  XNOR U5846 ( .A(c[689]), .B(n4822), .Z(n4821) );
  IV U5847 ( .A(o[689]), .Z(n4822) );
  XNOR U5848 ( .A(n4823), .B(n4824), .Z(o[689]) );
  XOR U5849 ( .A(n4825), .B(o[688]), .Z(creg_next[688]) );
  AND U5850 ( .A(n3090), .B(n4826), .Z(n4825) );
  XNOR U5851 ( .A(c[688]), .B(n4827), .Z(n4826) );
  IV U5852 ( .A(o[688]), .Z(n4827) );
  XNOR U5853 ( .A(n4828), .B(n4829), .Z(o[688]) );
  XOR U5854 ( .A(n4830), .B(o[687]), .Z(creg_next[687]) );
  AND U5855 ( .A(n3090), .B(n4831), .Z(n4830) );
  XNOR U5856 ( .A(c[687]), .B(n4832), .Z(n4831) );
  IV U5857 ( .A(o[687]), .Z(n4832) );
  XNOR U5858 ( .A(n4833), .B(n4834), .Z(o[687]) );
  XOR U5859 ( .A(n4835), .B(o[686]), .Z(creg_next[686]) );
  AND U5860 ( .A(n3090), .B(n4836), .Z(n4835) );
  XNOR U5861 ( .A(c[686]), .B(n4837), .Z(n4836) );
  IV U5862 ( .A(o[686]), .Z(n4837) );
  XNOR U5863 ( .A(n4838), .B(n4839), .Z(o[686]) );
  XOR U5864 ( .A(n4840), .B(o[685]), .Z(creg_next[685]) );
  AND U5865 ( .A(n3090), .B(n4841), .Z(n4840) );
  XNOR U5866 ( .A(c[685]), .B(n4842), .Z(n4841) );
  IV U5867 ( .A(o[685]), .Z(n4842) );
  XNOR U5868 ( .A(n4843), .B(n4844), .Z(o[685]) );
  XOR U5869 ( .A(n4845), .B(o[684]), .Z(creg_next[684]) );
  AND U5870 ( .A(n3090), .B(n4846), .Z(n4845) );
  XNOR U5871 ( .A(c[684]), .B(n4847), .Z(n4846) );
  IV U5872 ( .A(o[684]), .Z(n4847) );
  XNOR U5873 ( .A(n4848), .B(n4849), .Z(o[684]) );
  XOR U5874 ( .A(n4850), .B(o[683]), .Z(creg_next[683]) );
  AND U5875 ( .A(n3090), .B(n4851), .Z(n4850) );
  XNOR U5876 ( .A(c[683]), .B(n4852), .Z(n4851) );
  IV U5877 ( .A(o[683]), .Z(n4852) );
  XNOR U5878 ( .A(n4853), .B(n4854), .Z(o[683]) );
  XOR U5879 ( .A(n4855), .B(o[682]), .Z(creg_next[682]) );
  AND U5880 ( .A(n3090), .B(n4856), .Z(n4855) );
  XNOR U5881 ( .A(c[682]), .B(n4857), .Z(n4856) );
  IV U5882 ( .A(o[682]), .Z(n4857) );
  XNOR U5883 ( .A(n4858), .B(n4859), .Z(o[682]) );
  XOR U5884 ( .A(n4860), .B(o[681]), .Z(creg_next[681]) );
  AND U5885 ( .A(n3090), .B(n4861), .Z(n4860) );
  XNOR U5886 ( .A(c[681]), .B(n4862), .Z(n4861) );
  IV U5887 ( .A(o[681]), .Z(n4862) );
  XNOR U5888 ( .A(n4863), .B(n4864), .Z(o[681]) );
  XOR U5889 ( .A(n4865), .B(o[680]), .Z(creg_next[680]) );
  AND U5890 ( .A(n3090), .B(n4866), .Z(n4865) );
  XNOR U5891 ( .A(c[680]), .B(n4867), .Z(n4866) );
  IV U5892 ( .A(o[680]), .Z(n4867) );
  XNOR U5893 ( .A(n4868), .B(n4869), .Z(o[680]) );
  XOR U5894 ( .A(n4870), .B(o[67]), .Z(creg_next[67]) );
  AND U5895 ( .A(n3090), .B(n4871), .Z(n4870) );
  XNOR U5896 ( .A(c[67]), .B(n4872), .Z(n4871) );
  IV U5897 ( .A(o[67]), .Z(n4872) );
  XNOR U5898 ( .A(n4873), .B(n4874), .Z(o[67]) );
  XOR U5899 ( .A(n4875), .B(o[679]), .Z(creg_next[679]) );
  AND U5900 ( .A(n3090), .B(n4876), .Z(n4875) );
  XNOR U5901 ( .A(c[679]), .B(n4877), .Z(n4876) );
  IV U5902 ( .A(o[679]), .Z(n4877) );
  XNOR U5903 ( .A(n4878), .B(n4879), .Z(o[679]) );
  XOR U5904 ( .A(n4880), .B(o[678]), .Z(creg_next[678]) );
  AND U5905 ( .A(n3090), .B(n4881), .Z(n4880) );
  XNOR U5906 ( .A(c[678]), .B(n4882), .Z(n4881) );
  IV U5907 ( .A(o[678]), .Z(n4882) );
  XNOR U5908 ( .A(n4883), .B(n4884), .Z(o[678]) );
  XOR U5909 ( .A(n4885), .B(o[677]), .Z(creg_next[677]) );
  AND U5910 ( .A(n3090), .B(n4886), .Z(n4885) );
  XNOR U5911 ( .A(c[677]), .B(n4887), .Z(n4886) );
  IV U5912 ( .A(o[677]), .Z(n4887) );
  XNOR U5913 ( .A(n4888), .B(n4889), .Z(o[677]) );
  XOR U5914 ( .A(n4890), .B(o[676]), .Z(creg_next[676]) );
  AND U5915 ( .A(n3090), .B(n4891), .Z(n4890) );
  XNOR U5916 ( .A(c[676]), .B(n4892), .Z(n4891) );
  IV U5917 ( .A(o[676]), .Z(n4892) );
  XNOR U5918 ( .A(n4893), .B(n4894), .Z(o[676]) );
  XOR U5919 ( .A(n4895), .B(o[675]), .Z(creg_next[675]) );
  AND U5920 ( .A(n3090), .B(n4896), .Z(n4895) );
  XNOR U5921 ( .A(c[675]), .B(n4897), .Z(n4896) );
  IV U5922 ( .A(o[675]), .Z(n4897) );
  XNOR U5923 ( .A(n4898), .B(n4899), .Z(o[675]) );
  XOR U5924 ( .A(n4900), .B(o[674]), .Z(creg_next[674]) );
  AND U5925 ( .A(n3090), .B(n4901), .Z(n4900) );
  XNOR U5926 ( .A(c[674]), .B(n4902), .Z(n4901) );
  IV U5927 ( .A(o[674]), .Z(n4902) );
  XNOR U5928 ( .A(n4903), .B(n4904), .Z(o[674]) );
  XOR U5929 ( .A(n4905), .B(o[673]), .Z(creg_next[673]) );
  AND U5930 ( .A(n3090), .B(n4906), .Z(n4905) );
  XNOR U5931 ( .A(c[673]), .B(n4907), .Z(n4906) );
  IV U5932 ( .A(o[673]), .Z(n4907) );
  XNOR U5933 ( .A(n4908), .B(n4909), .Z(o[673]) );
  XOR U5934 ( .A(n4910), .B(o[672]), .Z(creg_next[672]) );
  AND U5935 ( .A(n3090), .B(n4911), .Z(n4910) );
  XNOR U5936 ( .A(c[672]), .B(n4912), .Z(n4911) );
  IV U5937 ( .A(o[672]), .Z(n4912) );
  XNOR U5938 ( .A(n4913), .B(n4914), .Z(o[672]) );
  XOR U5939 ( .A(n4915), .B(o[671]), .Z(creg_next[671]) );
  AND U5940 ( .A(n3090), .B(n4916), .Z(n4915) );
  XNOR U5941 ( .A(c[671]), .B(n4917), .Z(n4916) );
  IV U5942 ( .A(o[671]), .Z(n4917) );
  XNOR U5943 ( .A(n4918), .B(n4919), .Z(o[671]) );
  XOR U5944 ( .A(n4920), .B(o[670]), .Z(creg_next[670]) );
  AND U5945 ( .A(n3090), .B(n4921), .Z(n4920) );
  XNOR U5946 ( .A(c[670]), .B(n4922), .Z(n4921) );
  IV U5947 ( .A(o[670]), .Z(n4922) );
  XNOR U5948 ( .A(n4923), .B(n4924), .Z(o[670]) );
  XOR U5949 ( .A(n4925), .B(o[66]), .Z(creg_next[66]) );
  AND U5950 ( .A(n3090), .B(n4926), .Z(n4925) );
  XNOR U5951 ( .A(c[66]), .B(n4927), .Z(n4926) );
  IV U5952 ( .A(o[66]), .Z(n4927) );
  XNOR U5953 ( .A(n4928), .B(n4929), .Z(o[66]) );
  XOR U5954 ( .A(n4930), .B(o[669]), .Z(creg_next[669]) );
  AND U5955 ( .A(n3090), .B(n4931), .Z(n4930) );
  XNOR U5956 ( .A(c[669]), .B(n4932), .Z(n4931) );
  IV U5957 ( .A(o[669]), .Z(n4932) );
  XNOR U5958 ( .A(n4933), .B(n4934), .Z(o[669]) );
  XOR U5959 ( .A(n4935), .B(o[668]), .Z(creg_next[668]) );
  AND U5960 ( .A(n3090), .B(n4936), .Z(n4935) );
  XNOR U5961 ( .A(c[668]), .B(n4937), .Z(n4936) );
  IV U5962 ( .A(o[668]), .Z(n4937) );
  XNOR U5963 ( .A(n4938), .B(n4939), .Z(o[668]) );
  XOR U5964 ( .A(n4940), .B(o[667]), .Z(creg_next[667]) );
  AND U5965 ( .A(n3090), .B(n4941), .Z(n4940) );
  XNOR U5966 ( .A(c[667]), .B(n4942), .Z(n4941) );
  IV U5967 ( .A(o[667]), .Z(n4942) );
  XNOR U5968 ( .A(n4943), .B(n4944), .Z(o[667]) );
  XOR U5969 ( .A(n4945), .B(o[666]), .Z(creg_next[666]) );
  AND U5970 ( .A(n3090), .B(n4946), .Z(n4945) );
  XNOR U5971 ( .A(c[666]), .B(n4947), .Z(n4946) );
  IV U5972 ( .A(o[666]), .Z(n4947) );
  XNOR U5973 ( .A(n4948), .B(n4949), .Z(o[666]) );
  XOR U5974 ( .A(n4950), .B(o[665]), .Z(creg_next[665]) );
  AND U5975 ( .A(n3090), .B(n4951), .Z(n4950) );
  XNOR U5976 ( .A(c[665]), .B(n4952), .Z(n4951) );
  IV U5977 ( .A(o[665]), .Z(n4952) );
  XNOR U5978 ( .A(n4953), .B(n4954), .Z(o[665]) );
  XOR U5979 ( .A(n4955), .B(o[664]), .Z(creg_next[664]) );
  AND U5980 ( .A(n3090), .B(n4956), .Z(n4955) );
  XNOR U5981 ( .A(c[664]), .B(n4957), .Z(n4956) );
  IV U5982 ( .A(o[664]), .Z(n4957) );
  XNOR U5983 ( .A(n4958), .B(n4959), .Z(o[664]) );
  XOR U5984 ( .A(n4960), .B(o[663]), .Z(creg_next[663]) );
  AND U5985 ( .A(n3090), .B(n4961), .Z(n4960) );
  XNOR U5986 ( .A(c[663]), .B(n4962), .Z(n4961) );
  IV U5987 ( .A(o[663]), .Z(n4962) );
  XNOR U5988 ( .A(n4963), .B(n4964), .Z(o[663]) );
  XOR U5989 ( .A(n4965), .B(o[662]), .Z(creg_next[662]) );
  AND U5990 ( .A(n3090), .B(n4966), .Z(n4965) );
  XNOR U5991 ( .A(c[662]), .B(n4967), .Z(n4966) );
  IV U5992 ( .A(o[662]), .Z(n4967) );
  XNOR U5993 ( .A(n4968), .B(n4969), .Z(o[662]) );
  XOR U5994 ( .A(n4970), .B(o[661]), .Z(creg_next[661]) );
  AND U5995 ( .A(n3090), .B(n4971), .Z(n4970) );
  XNOR U5996 ( .A(c[661]), .B(n4972), .Z(n4971) );
  IV U5997 ( .A(o[661]), .Z(n4972) );
  XNOR U5998 ( .A(n4973), .B(n4974), .Z(o[661]) );
  XOR U5999 ( .A(n4975), .B(o[660]), .Z(creg_next[660]) );
  AND U6000 ( .A(n3090), .B(n4976), .Z(n4975) );
  XNOR U6001 ( .A(c[660]), .B(n4977), .Z(n4976) );
  IV U6002 ( .A(o[660]), .Z(n4977) );
  XNOR U6003 ( .A(n4978), .B(n4979), .Z(o[660]) );
  XOR U6004 ( .A(n4980), .B(o[65]), .Z(creg_next[65]) );
  AND U6005 ( .A(n3090), .B(n4981), .Z(n4980) );
  XNOR U6006 ( .A(c[65]), .B(n4982), .Z(n4981) );
  IV U6007 ( .A(o[65]), .Z(n4982) );
  XNOR U6008 ( .A(n4983), .B(n4984), .Z(o[65]) );
  XOR U6009 ( .A(n4985), .B(o[659]), .Z(creg_next[659]) );
  AND U6010 ( .A(n3090), .B(n4986), .Z(n4985) );
  XNOR U6011 ( .A(c[659]), .B(n4987), .Z(n4986) );
  IV U6012 ( .A(o[659]), .Z(n4987) );
  XNOR U6013 ( .A(n4988), .B(n4989), .Z(o[659]) );
  XOR U6014 ( .A(n4990), .B(o[658]), .Z(creg_next[658]) );
  AND U6015 ( .A(n3090), .B(n4991), .Z(n4990) );
  XNOR U6016 ( .A(c[658]), .B(n4992), .Z(n4991) );
  IV U6017 ( .A(o[658]), .Z(n4992) );
  XNOR U6018 ( .A(n4993), .B(n4994), .Z(o[658]) );
  XOR U6019 ( .A(n4995), .B(o[657]), .Z(creg_next[657]) );
  AND U6020 ( .A(n3090), .B(n4996), .Z(n4995) );
  XNOR U6021 ( .A(c[657]), .B(n4997), .Z(n4996) );
  IV U6022 ( .A(o[657]), .Z(n4997) );
  XNOR U6023 ( .A(n4998), .B(n4999), .Z(o[657]) );
  XOR U6024 ( .A(n5000), .B(o[656]), .Z(creg_next[656]) );
  AND U6025 ( .A(n3090), .B(n5001), .Z(n5000) );
  XNOR U6026 ( .A(c[656]), .B(n5002), .Z(n5001) );
  IV U6027 ( .A(o[656]), .Z(n5002) );
  XNOR U6028 ( .A(n5003), .B(n5004), .Z(o[656]) );
  XOR U6029 ( .A(n5005), .B(o[655]), .Z(creg_next[655]) );
  AND U6030 ( .A(n3090), .B(n5006), .Z(n5005) );
  XNOR U6031 ( .A(c[655]), .B(n5007), .Z(n5006) );
  IV U6032 ( .A(o[655]), .Z(n5007) );
  XNOR U6033 ( .A(n5008), .B(n5009), .Z(o[655]) );
  XOR U6034 ( .A(n5010), .B(o[654]), .Z(creg_next[654]) );
  AND U6035 ( .A(n3090), .B(n5011), .Z(n5010) );
  XNOR U6036 ( .A(c[654]), .B(n5012), .Z(n5011) );
  IV U6037 ( .A(o[654]), .Z(n5012) );
  XNOR U6038 ( .A(n5013), .B(n5014), .Z(o[654]) );
  XOR U6039 ( .A(n5015), .B(o[653]), .Z(creg_next[653]) );
  AND U6040 ( .A(n3090), .B(n5016), .Z(n5015) );
  XNOR U6041 ( .A(c[653]), .B(n5017), .Z(n5016) );
  IV U6042 ( .A(o[653]), .Z(n5017) );
  XNOR U6043 ( .A(n5018), .B(n5019), .Z(o[653]) );
  XOR U6044 ( .A(n5020), .B(o[652]), .Z(creg_next[652]) );
  AND U6045 ( .A(n3090), .B(n5021), .Z(n5020) );
  XNOR U6046 ( .A(c[652]), .B(n5022), .Z(n5021) );
  IV U6047 ( .A(o[652]), .Z(n5022) );
  XNOR U6048 ( .A(n5023), .B(n5024), .Z(o[652]) );
  XOR U6049 ( .A(n5025), .B(o[651]), .Z(creg_next[651]) );
  AND U6050 ( .A(n3090), .B(n5026), .Z(n5025) );
  XNOR U6051 ( .A(c[651]), .B(n5027), .Z(n5026) );
  IV U6052 ( .A(o[651]), .Z(n5027) );
  XNOR U6053 ( .A(n5028), .B(n5029), .Z(o[651]) );
  XOR U6054 ( .A(n5030), .B(o[650]), .Z(creg_next[650]) );
  AND U6055 ( .A(n3090), .B(n5031), .Z(n5030) );
  XNOR U6056 ( .A(c[650]), .B(n5032), .Z(n5031) );
  IV U6057 ( .A(o[650]), .Z(n5032) );
  XNOR U6058 ( .A(n5033), .B(n5034), .Z(o[650]) );
  XOR U6059 ( .A(n5035), .B(o[64]), .Z(creg_next[64]) );
  AND U6060 ( .A(n3090), .B(n5036), .Z(n5035) );
  XNOR U6061 ( .A(c[64]), .B(n5037), .Z(n5036) );
  IV U6062 ( .A(o[64]), .Z(n5037) );
  XNOR U6063 ( .A(n5038), .B(n5039), .Z(o[64]) );
  XOR U6064 ( .A(n5040), .B(o[649]), .Z(creg_next[649]) );
  AND U6065 ( .A(n3090), .B(n5041), .Z(n5040) );
  XNOR U6066 ( .A(c[649]), .B(n5042), .Z(n5041) );
  IV U6067 ( .A(o[649]), .Z(n5042) );
  XNOR U6068 ( .A(n5043), .B(n5044), .Z(o[649]) );
  XOR U6069 ( .A(n5045), .B(o[648]), .Z(creg_next[648]) );
  AND U6070 ( .A(n3090), .B(n5046), .Z(n5045) );
  XNOR U6071 ( .A(c[648]), .B(n5047), .Z(n5046) );
  IV U6072 ( .A(o[648]), .Z(n5047) );
  XNOR U6073 ( .A(n5048), .B(n5049), .Z(o[648]) );
  XOR U6074 ( .A(n5050), .B(o[647]), .Z(creg_next[647]) );
  AND U6075 ( .A(n3090), .B(n5051), .Z(n5050) );
  XNOR U6076 ( .A(c[647]), .B(n5052), .Z(n5051) );
  IV U6077 ( .A(o[647]), .Z(n5052) );
  XNOR U6078 ( .A(n5053), .B(n5054), .Z(o[647]) );
  XOR U6079 ( .A(n5055), .B(o[646]), .Z(creg_next[646]) );
  AND U6080 ( .A(n3090), .B(n5056), .Z(n5055) );
  XNOR U6081 ( .A(c[646]), .B(n5057), .Z(n5056) );
  IV U6082 ( .A(o[646]), .Z(n5057) );
  XNOR U6083 ( .A(n5058), .B(n5059), .Z(o[646]) );
  XOR U6084 ( .A(n5060), .B(o[645]), .Z(creg_next[645]) );
  AND U6085 ( .A(n3090), .B(n5061), .Z(n5060) );
  XNOR U6086 ( .A(c[645]), .B(n5062), .Z(n5061) );
  IV U6087 ( .A(o[645]), .Z(n5062) );
  XNOR U6088 ( .A(n5063), .B(n5064), .Z(o[645]) );
  XOR U6089 ( .A(n5065), .B(o[644]), .Z(creg_next[644]) );
  AND U6090 ( .A(n3090), .B(n5066), .Z(n5065) );
  XNOR U6091 ( .A(c[644]), .B(n5067), .Z(n5066) );
  IV U6092 ( .A(o[644]), .Z(n5067) );
  XNOR U6093 ( .A(n5068), .B(n5069), .Z(o[644]) );
  XOR U6094 ( .A(n5070), .B(o[643]), .Z(creg_next[643]) );
  AND U6095 ( .A(n3090), .B(n5071), .Z(n5070) );
  XNOR U6096 ( .A(c[643]), .B(n5072), .Z(n5071) );
  IV U6097 ( .A(o[643]), .Z(n5072) );
  XNOR U6098 ( .A(n5073), .B(n5074), .Z(o[643]) );
  XOR U6099 ( .A(n5075), .B(o[642]), .Z(creg_next[642]) );
  AND U6100 ( .A(n3090), .B(n5076), .Z(n5075) );
  XNOR U6101 ( .A(c[642]), .B(n5077), .Z(n5076) );
  IV U6102 ( .A(o[642]), .Z(n5077) );
  XNOR U6103 ( .A(n5078), .B(n5079), .Z(o[642]) );
  XOR U6104 ( .A(n5080), .B(o[641]), .Z(creg_next[641]) );
  AND U6105 ( .A(n3090), .B(n5081), .Z(n5080) );
  XNOR U6106 ( .A(c[641]), .B(n5082), .Z(n5081) );
  IV U6107 ( .A(o[641]), .Z(n5082) );
  XNOR U6108 ( .A(n5083), .B(n5084), .Z(o[641]) );
  XOR U6109 ( .A(n5085), .B(o[640]), .Z(creg_next[640]) );
  AND U6110 ( .A(n3090), .B(n5086), .Z(n5085) );
  XNOR U6111 ( .A(c[640]), .B(n5087), .Z(n5086) );
  IV U6112 ( .A(o[640]), .Z(n5087) );
  XNOR U6113 ( .A(n5088), .B(n5089), .Z(o[640]) );
  XOR U6114 ( .A(n5090), .B(o[63]), .Z(creg_next[63]) );
  AND U6115 ( .A(n3090), .B(n5091), .Z(n5090) );
  XNOR U6116 ( .A(c[63]), .B(n5092), .Z(n5091) );
  IV U6117 ( .A(o[63]), .Z(n5092) );
  XNOR U6118 ( .A(n5093), .B(n5094), .Z(o[63]) );
  XOR U6119 ( .A(n5095), .B(o[639]), .Z(creg_next[639]) );
  AND U6120 ( .A(n3090), .B(n5096), .Z(n5095) );
  XNOR U6121 ( .A(c[639]), .B(n5097), .Z(n5096) );
  IV U6122 ( .A(o[639]), .Z(n5097) );
  XNOR U6123 ( .A(n5098), .B(n5099), .Z(o[639]) );
  XOR U6124 ( .A(n5100), .B(o[638]), .Z(creg_next[638]) );
  AND U6125 ( .A(n3090), .B(n5101), .Z(n5100) );
  XNOR U6126 ( .A(c[638]), .B(n5102), .Z(n5101) );
  IV U6127 ( .A(o[638]), .Z(n5102) );
  XNOR U6128 ( .A(n5103), .B(n5104), .Z(o[638]) );
  XOR U6129 ( .A(n5105), .B(o[637]), .Z(creg_next[637]) );
  AND U6130 ( .A(n3090), .B(n5106), .Z(n5105) );
  XNOR U6131 ( .A(c[637]), .B(n5107), .Z(n5106) );
  IV U6132 ( .A(o[637]), .Z(n5107) );
  XNOR U6133 ( .A(n5108), .B(n5109), .Z(o[637]) );
  XOR U6134 ( .A(n5110), .B(o[636]), .Z(creg_next[636]) );
  AND U6135 ( .A(n3090), .B(n5111), .Z(n5110) );
  XNOR U6136 ( .A(c[636]), .B(n5112), .Z(n5111) );
  IV U6137 ( .A(o[636]), .Z(n5112) );
  XNOR U6138 ( .A(n5113), .B(n5114), .Z(o[636]) );
  XOR U6139 ( .A(n5115), .B(o[635]), .Z(creg_next[635]) );
  AND U6140 ( .A(n3090), .B(n5116), .Z(n5115) );
  XNOR U6141 ( .A(c[635]), .B(n5117), .Z(n5116) );
  IV U6142 ( .A(o[635]), .Z(n5117) );
  XNOR U6143 ( .A(n5118), .B(n5119), .Z(o[635]) );
  XOR U6144 ( .A(n5120), .B(o[634]), .Z(creg_next[634]) );
  AND U6145 ( .A(n3090), .B(n5121), .Z(n5120) );
  XNOR U6146 ( .A(c[634]), .B(n5122), .Z(n5121) );
  IV U6147 ( .A(o[634]), .Z(n5122) );
  XNOR U6148 ( .A(n5123), .B(n5124), .Z(o[634]) );
  XOR U6149 ( .A(n5125), .B(o[633]), .Z(creg_next[633]) );
  AND U6150 ( .A(n3090), .B(n5126), .Z(n5125) );
  XNOR U6151 ( .A(c[633]), .B(n5127), .Z(n5126) );
  IV U6152 ( .A(o[633]), .Z(n5127) );
  XNOR U6153 ( .A(n5128), .B(n5129), .Z(o[633]) );
  XOR U6154 ( .A(n5130), .B(o[632]), .Z(creg_next[632]) );
  AND U6155 ( .A(n3090), .B(n5131), .Z(n5130) );
  XNOR U6156 ( .A(c[632]), .B(n5132), .Z(n5131) );
  IV U6157 ( .A(o[632]), .Z(n5132) );
  XNOR U6158 ( .A(n5133), .B(n5134), .Z(o[632]) );
  XOR U6159 ( .A(n5135), .B(o[631]), .Z(creg_next[631]) );
  AND U6160 ( .A(n3090), .B(n5136), .Z(n5135) );
  XNOR U6161 ( .A(c[631]), .B(n5137), .Z(n5136) );
  IV U6162 ( .A(o[631]), .Z(n5137) );
  XNOR U6163 ( .A(n5138), .B(n5139), .Z(o[631]) );
  XOR U6164 ( .A(n5140), .B(o[630]), .Z(creg_next[630]) );
  AND U6165 ( .A(n3090), .B(n5141), .Z(n5140) );
  XNOR U6166 ( .A(c[630]), .B(n5142), .Z(n5141) );
  IV U6167 ( .A(o[630]), .Z(n5142) );
  XNOR U6168 ( .A(n5143), .B(n5144), .Z(o[630]) );
  XOR U6169 ( .A(n5145), .B(o[62]), .Z(creg_next[62]) );
  AND U6170 ( .A(n3090), .B(n5146), .Z(n5145) );
  XNOR U6171 ( .A(c[62]), .B(n5147), .Z(n5146) );
  IV U6172 ( .A(o[62]), .Z(n5147) );
  XNOR U6173 ( .A(n5148), .B(n5149), .Z(o[62]) );
  XOR U6174 ( .A(n5150), .B(o[629]), .Z(creg_next[629]) );
  AND U6175 ( .A(n3090), .B(n5151), .Z(n5150) );
  XNOR U6176 ( .A(c[629]), .B(n5152), .Z(n5151) );
  IV U6177 ( .A(o[629]), .Z(n5152) );
  XNOR U6178 ( .A(n5153), .B(n5154), .Z(o[629]) );
  XOR U6179 ( .A(n5155), .B(o[628]), .Z(creg_next[628]) );
  AND U6180 ( .A(n3090), .B(n5156), .Z(n5155) );
  XNOR U6181 ( .A(c[628]), .B(n5157), .Z(n5156) );
  IV U6182 ( .A(o[628]), .Z(n5157) );
  XNOR U6183 ( .A(n5158), .B(n5159), .Z(o[628]) );
  XOR U6184 ( .A(n5160), .B(o[627]), .Z(creg_next[627]) );
  AND U6185 ( .A(n3090), .B(n5161), .Z(n5160) );
  XNOR U6186 ( .A(c[627]), .B(n5162), .Z(n5161) );
  IV U6187 ( .A(o[627]), .Z(n5162) );
  XNOR U6188 ( .A(n5163), .B(n5164), .Z(o[627]) );
  XOR U6189 ( .A(n5165), .B(o[626]), .Z(creg_next[626]) );
  AND U6190 ( .A(n3090), .B(n5166), .Z(n5165) );
  XNOR U6191 ( .A(c[626]), .B(n5167), .Z(n5166) );
  IV U6192 ( .A(o[626]), .Z(n5167) );
  XNOR U6193 ( .A(n5168), .B(n5169), .Z(o[626]) );
  XOR U6194 ( .A(n5170), .B(o[625]), .Z(creg_next[625]) );
  AND U6195 ( .A(n3090), .B(n5171), .Z(n5170) );
  XNOR U6196 ( .A(c[625]), .B(n5172), .Z(n5171) );
  IV U6197 ( .A(o[625]), .Z(n5172) );
  XNOR U6198 ( .A(n5173), .B(n5174), .Z(o[625]) );
  XOR U6199 ( .A(n5175), .B(o[624]), .Z(creg_next[624]) );
  AND U6200 ( .A(n3090), .B(n5176), .Z(n5175) );
  XNOR U6201 ( .A(c[624]), .B(n5177), .Z(n5176) );
  IV U6202 ( .A(o[624]), .Z(n5177) );
  XNOR U6203 ( .A(n5178), .B(n5179), .Z(o[624]) );
  XOR U6204 ( .A(n5180), .B(o[623]), .Z(creg_next[623]) );
  AND U6205 ( .A(n3090), .B(n5181), .Z(n5180) );
  XNOR U6206 ( .A(c[623]), .B(n5182), .Z(n5181) );
  IV U6207 ( .A(o[623]), .Z(n5182) );
  XNOR U6208 ( .A(n5183), .B(n5184), .Z(o[623]) );
  XOR U6209 ( .A(n5185), .B(o[622]), .Z(creg_next[622]) );
  AND U6210 ( .A(n3090), .B(n5186), .Z(n5185) );
  XNOR U6211 ( .A(c[622]), .B(n5187), .Z(n5186) );
  IV U6212 ( .A(o[622]), .Z(n5187) );
  XNOR U6213 ( .A(n5188), .B(n5189), .Z(o[622]) );
  XOR U6214 ( .A(n5190), .B(o[621]), .Z(creg_next[621]) );
  AND U6215 ( .A(n3090), .B(n5191), .Z(n5190) );
  XNOR U6216 ( .A(c[621]), .B(n5192), .Z(n5191) );
  IV U6217 ( .A(o[621]), .Z(n5192) );
  XNOR U6218 ( .A(n5193), .B(n5194), .Z(o[621]) );
  XOR U6219 ( .A(n5195), .B(o[620]), .Z(creg_next[620]) );
  AND U6220 ( .A(n3090), .B(n5196), .Z(n5195) );
  XNOR U6221 ( .A(c[620]), .B(n5197), .Z(n5196) );
  IV U6222 ( .A(o[620]), .Z(n5197) );
  XNOR U6223 ( .A(n5198), .B(n5199), .Z(o[620]) );
  XOR U6224 ( .A(n5200), .B(o[61]), .Z(creg_next[61]) );
  AND U6225 ( .A(n3090), .B(n5201), .Z(n5200) );
  XNOR U6226 ( .A(c[61]), .B(n5202), .Z(n5201) );
  IV U6227 ( .A(o[61]), .Z(n5202) );
  XNOR U6228 ( .A(n5203), .B(n5204), .Z(o[61]) );
  XOR U6229 ( .A(n5205), .B(o[619]), .Z(creg_next[619]) );
  AND U6230 ( .A(n3090), .B(n5206), .Z(n5205) );
  XNOR U6231 ( .A(c[619]), .B(n5207), .Z(n5206) );
  IV U6232 ( .A(o[619]), .Z(n5207) );
  XNOR U6233 ( .A(n5208), .B(n5209), .Z(o[619]) );
  XOR U6234 ( .A(n5210), .B(o[618]), .Z(creg_next[618]) );
  AND U6235 ( .A(n3090), .B(n5211), .Z(n5210) );
  XNOR U6236 ( .A(c[618]), .B(n5212), .Z(n5211) );
  IV U6237 ( .A(o[618]), .Z(n5212) );
  XNOR U6238 ( .A(n5213), .B(n5214), .Z(o[618]) );
  XOR U6239 ( .A(n5215), .B(o[617]), .Z(creg_next[617]) );
  AND U6240 ( .A(n3090), .B(n5216), .Z(n5215) );
  XNOR U6241 ( .A(c[617]), .B(n5217), .Z(n5216) );
  IV U6242 ( .A(o[617]), .Z(n5217) );
  XNOR U6243 ( .A(n5218), .B(n5219), .Z(o[617]) );
  XOR U6244 ( .A(n5220), .B(o[616]), .Z(creg_next[616]) );
  AND U6245 ( .A(n3090), .B(n5221), .Z(n5220) );
  XNOR U6246 ( .A(c[616]), .B(n5222), .Z(n5221) );
  IV U6247 ( .A(o[616]), .Z(n5222) );
  XNOR U6248 ( .A(n5223), .B(n5224), .Z(o[616]) );
  XOR U6249 ( .A(n5225), .B(o[615]), .Z(creg_next[615]) );
  AND U6250 ( .A(n3090), .B(n5226), .Z(n5225) );
  XNOR U6251 ( .A(c[615]), .B(n5227), .Z(n5226) );
  IV U6252 ( .A(o[615]), .Z(n5227) );
  XNOR U6253 ( .A(n5228), .B(n5229), .Z(o[615]) );
  XOR U6254 ( .A(n5230), .B(o[614]), .Z(creg_next[614]) );
  AND U6255 ( .A(n3090), .B(n5231), .Z(n5230) );
  XNOR U6256 ( .A(c[614]), .B(n5232), .Z(n5231) );
  IV U6257 ( .A(o[614]), .Z(n5232) );
  XNOR U6258 ( .A(n5233), .B(n5234), .Z(o[614]) );
  XOR U6259 ( .A(n5235), .B(o[613]), .Z(creg_next[613]) );
  AND U6260 ( .A(n3090), .B(n5236), .Z(n5235) );
  XNOR U6261 ( .A(c[613]), .B(n5237), .Z(n5236) );
  IV U6262 ( .A(o[613]), .Z(n5237) );
  XNOR U6263 ( .A(n5238), .B(n5239), .Z(o[613]) );
  XOR U6264 ( .A(n5240), .B(o[612]), .Z(creg_next[612]) );
  AND U6265 ( .A(n3090), .B(n5241), .Z(n5240) );
  XNOR U6266 ( .A(c[612]), .B(n5242), .Z(n5241) );
  IV U6267 ( .A(o[612]), .Z(n5242) );
  XNOR U6268 ( .A(n5243), .B(n5244), .Z(o[612]) );
  XOR U6269 ( .A(n5245), .B(o[611]), .Z(creg_next[611]) );
  AND U6270 ( .A(n3090), .B(n5246), .Z(n5245) );
  XNOR U6271 ( .A(c[611]), .B(n5247), .Z(n5246) );
  IV U6272 ( .A(o[611]), .Z(n5247) );
  XNOR U6273 ( .A(n5248), .B(n5249), .Z(o[611]) );
  XOR U6274 ( .A(n5250), .B(o[610]), .Z(creg_next[610]) );
  AND U6275 ( .A(n3090), .B(n5251), .Z(n5250) );
  XNOR U6276 ( .A(c[610]), .B(n5252), .Z(n5251) );
  IV U6277 ( .A(o[610]), .Z(n5252) );
  XNOR U6278 ( .A(n5253), .B(n5254), .Z(o[610]) );
  XOR U6279 ( .A(n5255), .B(o[60]), .Z(creg_next[60]) );
  AND U6280 ( .A(n3090), .B(n5256), .Z(n5255) );
  XNOR U6281 ( .A(c[60]), .B(n5257), .Z(n5256) );
  IV U6282 ( .A(o[60]), .Z(n5257) );
  XNOR U6283 ( .A(n5258), .B(n5259), .Z(o[60]) );
  XOR U6284 ( .A(n5260), .B(o[609]), .Z(creg_next[609]) );
  AND U6285 ( .A(n3090), .B(n5261), .Z(n5260) );
  XNOR U6286 ( .A(c[609]), .B(n5262), .Z(n5261) );
  IV U6287 ( .A(o[609]), .Z(n5262) );
  XNOR U6288 ( .A(n5263), .B(n5264), .Z(o[609]) );
  XOR U6289 ( .A(n5265), .B(o[608]), .Z(creg_next[608]) );
  AND U6290 ( .A(n3090), .B(n5266), .Z(n5265) );
  XNOR U6291 ( .A(c[608]), .B(n5267), .Z(n5266) );
  IV U6292 ( .A(o[608]), .Z(n5267) );
  XNOR U6293 ( .A(n5268), .B(n5269), .Z(o[608]) );
  XOR U6294 ( .A(n5270), .B(o[607]), .Z(creg_next[607]) );
  AND U6295 ( .A(n3090), .B(n5271), .Z(n5270) );
  XNOR U6296 ( .A(c[607]), .B(n5272), .Z(n5271) );
  IV U6297 ( .A(o[607]), .Z(n5272) );
  XNOR U6298 ( .A(n5273), .B(n5274), .Z(o[607]) );
  XOR U6299 ( .A(n5275), .B(o[606]), .Z(creg_next[606]) );
  AND U6300 ( .A(n3090), .B(n5276), .Z(n5275) );
  XNOR U6301 ( .A(c[606]), .B(n5277), .Z(n5276) );
  IV U6302 ( .A(o[606]), .Z(n5277) );
  XNOR U6303 ( .A(n5278), .B(n5279), .Z(o[606]) );
  XOR U6304 ( .A(n5280), .B(o[605]), .Z(creg_next[605]) );
  AND U6305 ( .A(n3090), .B(n5281), .Z(n5280) );
  XNOR U6306 ( .A(c[605]), .B(n5282), .Z(n5281) );
  IV U6307 ( .A(o[605]), .Z(n5282) );
  XNOR U6308 ( .A(n5283), .B(n5284), .Z(o[605]) );
  XOR U6309 ( .A(n5285), .B(o[604]), .Z(creg_next[604]) );
  AND U6310 ( .A(n3090), .B(n5286), .Z(n5285) );
  XNOR U6311 ( .A(c[604]), .B(n5287), .Z(n5286) );
  IV U6312 ( .A(o[604]), .Z(n5287) );
  XNOR U6313 ( .A(n5288), .B(n5289), .Z(o[604]) );
  XOR U6314 ( .A(n5290), .B(o[603]), .Z(creg_next[603]) );
  AND U6315 ( .A(n3090), .B(n5291), .Z(n5290) );
  XNOR U6316 ( .A(c[603]), .B(n5292), .Z(n5291) );
  IV U6317 ( .A(o[603]), .Z(n5292) );
  XNOR U6318 ( .A(n5293), .B(n5294), .Z(o[603]) );
  XOR U6319 ( .A(n5295), .B(o[602]), .Z(creg_next[602]) );
  AND U6320 ( .A(n3090), .B(n5296), .Z(n5295) );
  XNOR U6321 ( .A(c[602]), .B(n5297), .Z(n5296) );
  IV U6322 ( .A(o[602]), .Z(n5297) );
  XNOR U6323 ( .A(n5298), .B(n5299), .Z(o[602]) );
  XOR U6324 ( .A(n5300), .B(o[601]), .Z(creg_next[601]) );
  AND U6325 ( .A(n3090), .B(n5301), .Z(n5300) );
  XNOR U6326 ( .A(c[601]), .B(n5302), .Z(n5301) );
  IV U6327 ( .A(o[601]), .Z(n5302) );
  XNOR U6328 ( .A(n5303), .B(n5304), .Z(o[601]) );
  XOR U6329 ( .A(n5305), .B(o[600]), .Z(creg_next[600]) );
  AND U6330 ( .A(n3090), .B(n5306), .Z(n5305) );
  XNOR U6331 ( .A(c[600]), .B(n5307), .Z(n5306) );
  IV U6332 ( .A(o[600]), .Z(n5307) );
  XNOR U6333 ( .A(n5308), .B(n5309), .Z(o[600]) );
  XOR U6334 ( .A(n5310), .B(o[5]), .Z(creg_next[5]) );
  AND U6335 ( .A(n3090), .B(n5311), .Z(n5310) );
  XNOR U6336 ( .A(c[5]), .B(n5312), .Z(n5311) );
  IV U6337 ( .A(o[5]), .Z(n5312) );
  XNOR U6338 ( .A(n5313), .B(n5314), .Z(o[5]) );
  XOR U6339 ( .A(n5315), .B(o[59]), .Z(creg_next[59]) );
  AND U6340 ( .A(n3090), .B(n5316), .Z(n5315) );
  XNOR U6341 ( .A(c[59]), .B(n5317), .Z(n5316) );
  IV U6342 ( .A(o[59]), .Z(n5317) );
  XNOR U6343 ( .A(n5318), .B(n5319), .Z(o[59]) );
  XOR U6344 ( .A(n5320), .B(o[599]), .Z(creg_next[599]) );
  AND U6345 ( .A(n3090), .B(n5321), .Z(n5320) );
  XNOR U6346 ( .A(c[599]), .B(n5322), .Z(n5321) );
  IV U6347 ( .A(o[599]), .Z(n5322) );
  XNOR U6348 ( .A(n5323), .B(n5324), .Z(o[599]) );
  XOR U6349 ( .A(n5325), .B(o[598]), .Z(creg_next[598]) );
  AND U6350 ( .A(n3090), .B(n5326), .Z(n5325) );
  XNOR U6351 ( .A(c[598]), .B(n5327), .Z(n5326) );
  IV U6352 ( .A(o[598]), .Z(n5327) );
  XNOR U6353 ( .A(n5328), .B(n5329), .Z(o[598]) );
  XOR U6354 ( .A(n5330), .B(o[597]), .Z(creg_next[597]) );
  AND U6355 ( .A(n3090), .B(n5331), .Z(n5330) );
  XNOR U6356 ( .A(c[597]), .B(n5332), .Z(n5331) );
  IV U6357 ( .A(o[597]), .Z(n5332) );
  XNOR U6358 ( .A(n5333), .B(n5334), .Z(o[597]) );
  XOR U6359 ( .A(n5335), .B(o[596]), .Z(creg_next[596]) );
  AND U6360 ( .A(n3090), .B(n5336), .Z(n5335) );
  XNOR U6361 ( .A(c[596]), .B(n5337), .Z(n5336) );
  IV U6362 ( .A(o[596]), .Z(n5337) );
  XNOR U6363 ( .A(n5338), .B(n5339), .Z(o[596]) );
  XOR U6364 ( .A(n5340), .B(o[595]), .Z(creg_next[595]) );
  AND U6365 ( .A(n3090), .B(n5341), .Z(n5340) );
  XNOR U6366 ( .A(c[595]), .B(n5342), .Z(n5341) );
  IV U6367 ( .A(o[595]), .Z(n5342) );
  XNOR U6368 ( .A(n5343), .B(n5344), .Z(o[595]) );
  XOR U6369 ( .A(n5345), .B(o[594]), .Z(creg_next[594]) );
  AND U6370 ( .A(n3090), .B(n5346), .Z(n5345) );
  XNOR U6371 ( .A(c[594]), .B(n5347), .Z(n5346) );
  IV U6372 ( .A(o[594]), .Z(n5347) );
  XNOR U6373 ( .A(n5348), .B(n5349), .Z(o[594]) );
  XOR U6374 ( .A(n5350), .B(o[593]), .Z(creg_next[593]) );
  AND U6375 ( .A(n3090), .B(n5351), .Z(n5350) );
  XNOR U6376 ( .A(c[593]), .B(n5352), .Z(n5351) );
  IV U6377 ( .A(o[593]), .Z(n5352) );
  XNOR U6378 ( .A(n5353), .B(n5354), .Z(o[593]) );
  XOR U6379 ( .A(n5355), .B(o[592]), .Z(creg_next[592]) );
  AND U6380 ( .A(n3090), .B(n5356), .Z(n5355) );
  XNOR U6381 ( .A(c[592]), .B(n5357), .Z(n5356) );
  IV U6382 ( .A(o[592]), .Z(n5357) );
  XNOR U6383 ( .A(n5358), .B(n5359), .Z(o[592]) );
  XOR U6384 ( .A(n5360), .B(o[591]), .Z(creg_next[591]) );
  AND U6385 ( .A(n3090), .B(n5361), .Z(n5360) );
  XNOR U6386 ( .A(c[591]), .B(n5362), .Z(n5361) );
  IV U6387 ( .A(o[591]), .Z(n5362) );
  XNOR U6388 ( .A(n5363), .B(n5364), .Z(o[591]) );
  XOR U6389 ( .A(n5365), .B(o[590]), .Z(creg_next[590]) );
  AND U6390 ( .A(n3090), .B(n5366), .Z(n5365) );
  XNOR U6391 ( .A(c[590]), .B(n5367), .Z(n5366) );
  IV U6392 ( .A(o[590]), .Z(n5367) );
  XNOR U6393 ( .A(n5368), .B(n5369), .Z(o[590]) );
  XOR U6394 ( .A(n5370), .B(o[58]), .Z(creg_next[58]) );
  AND U6395 ( .A(n3090), .B(n5371), .Z(n5370) );
  XNOR U6396 ( .A(c[58]), .B(n5372), .Z(n5371) );
  IV U6397 ( .A(o[58]), .Z(n5372) );
  XNOR U6398 ( .A(n5373), .B(n5374), .Z(o[58]) );
  XOR U6399 ( .A(n5375), .B(o[589]), .Z(creg_next[589]) );
  AND U6400 ( .A(n3090), .B(n5376), .Z(n5375) );
  XNOR U6401 ( .A(c[589]), .B(n5377), .Z(n5376) );
  IV U6402 ( .A(o[589]), .Z(n5377) );
  XNOR U6403 ( .A(n5378), .B(n5379), .Z(o[589]) );
  XOR U6404 ( .A(n5380), .B(o[588]), .Z(creg_next[588]) );
  AND U6405 ( .A(n3090), .B(n5381), .Z(n5380) );
  XNOR U6406 ( .A(c[588]), .B(n5382), .Z(n5381) );
  IV U6407 ( .A(o[588]), .Z(n5382) );
  XNOR U6408 ( .A(n5383), .B(n5384), .Z(o[588]) );
  XOR U6409 ( .A(n5385), .B(o[587]), .Z(creg_next[587]) );
  AND U6410 ( .A(n3090), .B(n5386), .Z(n5385) );
  XNOR U6411 ( .A(c[587]), .B(n5387), .Z(n5386) );
  IV U6412 ( .A(o[587]), .Z(n5387) );
  XNOR U6413 ( .A(n5388), .B(n5389), .Z(o[587]) );
  XOR U6414 ( .A(n5390), .B(o[586]), .Z(creg_next[586]) );
  AND U6415 ( .A(n3090), .B(n5391), .Z(n5390) );
  XNOR U6416 ( .A(c[586]), .B(n5392), .Z(n5391) );
  IV U6417 ( .A(o[586]), .Z(n5392) );
  XNOR U6418 ( .A(n5393), .B(n5394), .Z(o[586]) );
  XOR U6419 ( .A(n5395), .B(o[585]), .Z(creg_next[585]) );
  AND U6420 ( .A(n3090), .B(n5396), .Z(n5395) );
  XNOR U6421 ( .A(c[585]), .B(n5397), .Z(n5396) );
  IV U6422 ( .A(o[585]), .Z(n5397) );
  XNOR U6423 ( .A(n5398), .B(n5399), .Z(o[585]) );
  XOR U6424 ( .A(n5400), .B(o[584]), .Z(creg_next[584]) );
  AND U6425 ( .A(n3090), .B(n5401), .Z(n5400) );
  XNOR U6426 ( .A(c[584]), .B(n5402), .Z(n5401) );
  IV U6427 ( .A(o[584]), .Z(n5402) );
  XNOR U6428 ( .A(n5403), .B(n5404), .Z(o[584]) );
  XOR U6429 ( .A(n5405), .B(o[583]), .Z(creg_next[583]) );
  AND U6430 ( .A(n3090), .B(n5406), .Z(n5405) );
  XNOR U6431 ( .A(c[583]), .B(n5407), .Z(n5406) );
  IV U6432 ( .A(o[583]), .Z(n5407) );
  XNOR U6433 ( .A(n5408), .B(n5409), .Z(o[583]) );
  XOR U6434 ( .A(n5410), .B(o[582]), .Z(creg_next[582]) );
  AND U6435 ( .A(n3090), .B(n5411), .Z(n5410) );
  XNOR U6436 ( .A(c[582]), .B(n5412), .Z(n5411) );
  IV U6437 ( .A(o[582]), .Z(n5412) );
  XNOR U6438 ( .A(n5413), .B(n5414), .Z(o[582]) );
  XOR U6439 ( .A(n5415), .B(o[581]), .Z(creg_next[581]) );
  AND U6440 ( .A(n3090), .B(n5416), .Z(n5415) );
  XNOR U6441 ( .A(c[581]), .B(n5417), .Z(n5416) );
  IV U6442 ( .A(o[581]), .Z(n5417) );
  XNOR U6443 ( .A(n5418), .B(n5419), .Z(o[581]) );
  XOR U6444 ( .A(n5420), .B(o[580]), .Z(creg_next[580]) );
  AND U6445 ( .A(n3090), .B(n5421), .Z(n5420) );
  XNOR U6446 ( .A(c[580]), .B(n5422), .Z(n5421) );
  IV U6447 ( .A(o[580]), .Z(n5422) );
  XNOR U6448 ( .A(n5423), .B(n5424), .Z(o[580]) );
  XOR U6449 ( .A(n5425), .B(o[57]), .Z(creg_next[57]) );
  AND U6450 ( .A(n3090), .B(n5426), .Z(n5425) );
  XNOR U6451 ( .A(c[57]), .B(n5427), .Z(n5426) );
  IV U6452 ( .A(o[57]), .Z(n5427) );
  XNOR U6453 ( .A(n5428), .B(n5429), .Z(o[57]) );
  XOR U6454 ( .A(n5430), .B(o[579]), .Z(creg_next[579]) );
  AND U6455 ( .A(n3090), .B(n5431), .Z(n5430) );
  XNOR U6456 ( .A(c[579]), .B(n5432), .Z(n5431) );
  IV U6457 ( .A(o[579]), .Z(n5432) );
  XNOR U6458 ( .A(n5433), .B(n5434), .Z(o[579]) );
  XOR U6459 ( .A(n5435), .B(o[578]), .Z(creg_next[578]) );
  AND U6460 ( .A(n3090), .B(n5436), .Z(n5435) );
  XNOR U6461 ( .A(c[578]), .B(n5437), .Z(n5436) );
  IV U6462 ( .A(o[578]), .Z(n5437) );
  XNOR U6463 ( .A(n5438), .B(n5439), .Z(o[578]) );
  XOR U6464 ( .A(n5440), .B(o[577]), .Z(creg_next[577]) );
  AND U6465 ( .A(n3090), .B(n5441), .Z(n5440) );
  XNOR U6466 ( .A(c[577]), .B(n5442), .Z(n5441) );
  IV U6467 ( .A(o[577]), .Z(n5442) );
  XNOR U6468 ( .A(n5443), .B(n5444), .Z(o[577]) );
  XOR U6469 ( .A(n5445), .B(o[576]), .Z(creg_next[576]) );
  AND U6470 ( .A(n3090), .B(n5446), .Z(n5445) );
  XNOR U6471 ( .A(c[576]), .B(n5447), .Z(n5446) );
  IV U6472 ( .A(o[576]), .Z(n5447) );
  XNOR U6473 ( .A(n5448), .B(n5449), .Z(o[576]) );
  XOR U6474 ( .A(n5450), .B(o[575]), .Z(creg_next[575]) );
  AND U6475 ( .A(n3090), .B(n5451), .Z(n5450) );
  XNOR U6476 ( .A(c[575]), .B(n5452), .Z(n5451) );
  IV U6477 ( .A(o[575]), .Z(n5452) );
  XNOR U6478 ( .A(n5453), .B(n5454), .Z(o[575]) );
  XOR U6479 ( .A(n5455), .B(o[574]), .Z(creg_next[574]) );
  AND U6480 ( .A(n3090), .B(n5456), .Z(n5455) );
  XNOR U6481 ( .A(c[574]), .B(n5457), .Z(n5456) );
  IV U6482 ( .A(o[574]), .Z(n5457) );
  XNOR U6483 ( .A(n5458), .B(n5459), .Z(o[574]) );
  XOR U6484 ( .A(n5460), .B(o[573]), .Z(creg_next[573]) );
  AND U6485 ( .A(n3090), .B(n5461), .Z(n5460) );
  XNOR U6486 ( .A(c[573]), .B(n5462), .Z(n5461) );
  IV U6487 ( .A(o[573]), .Z(n5462) );
  XNOR U6488 ( .A(n5463), .B(n5464), .Z(o[573]) );
  XOR U6489 ( .A(n5465), .B(o[572]), .Z(creg_next[572]) );
  AND U6490 ( .A(n3090), .B(n5466), .Z(n5465) );
  XNOR U6491 ( .A(c[572]), .B(n5467), .Z(n5466) );
  IV U6492 ( .A(o[572]), .Z(n5467) );
  XNOR U6493 ( .A(n5468), .B(n5469), .Z(o[572]) );
  XOR U6494 ( .A(n5470), .B(o[571]), .Z(creg_next[571]) );
  AND U6495 ( .A(n3090), .B(n5471), .Z(n5470) );
  XNOR U6496 ( .A(c[571]), .B(n5472), .Z(n5471) );
  IV U6497 ( .A(o[571]), .Z(n5472) );
  XNOR U6498 ( .A(n5473), .B(n5474), .Z(o[571]) );
  XOR U6499 ( .A(n5475), .B(o[570]), .Z(creg_next[570]) );
  AND U6500 ( .A(n3090), .B(n5476), .Z(n5475) );
  XNOR U6501 ( .A(c[570]), .B(n5477), .Z(n5476) );
  IV U6502 ( .A(o[570]), .Z(n5477) );
  XNOR U6503 ( .A(n5478), .B(n5479), .Z(o[570]) );
  XOR U6504 ( .A(n5480), .B(o[56]), .Z(creg_next[56]) );
  AND U6505 ( .A(n3090), .B(n5481), .Z(n5480) );
  XNOR U6506 ( .A(c[56]), .B(n5482), .Z(n5481) );
  IV U6507 ( .A(o[56]), .Z(n5482) );
  XNOR U6508 ( .A(n5483), .B(n5484), .Z(o[56]) );
  XOR U6509 ( .A(n5485), .B(o[569]), .Z(creg_next[569]) );
  AND U6510 ( .A(n3090), .B(n5486), .Z(n5485) );
  XNOR U6511 ( .A(c[569]), .B(n5487), .Z(n5486) );
  IV U6512 ( .A(o[569]), .Z(n5487) );
  XNOR U6513 ( .A(n5488), .B(n5489), .Z(o[569]) );
  XOR U6514 ( .A(n5490), .B(o[568]), .Z(creg_next[568]) );
  AND U6515 ( .A(n3090), .B(n5491), .Z(n5490) );
  XNOR U6516 ( .A(c[568]), .B(n5492), .Z(n5491) );
  IV U6517 ( .A(o[568]), .Z(n5492) );
  XNOR U6518 ( .A(n5493), .B(n5494), .Z(o[568]) );
  XOR U6519 ( .A(n5495), .B(o[567]), .Z(creg_next[567]) );
  AND U6520 ( .A(n3090), .B(n5496), .Z(n5495) );
  XNOR U6521 ( .A(c[567]), .B(n5497), .Z(n5496) );
  IV U6522 ( .A(o[567]), .Z(n5497) );
  XNOR U6523 ( .A(n5498), .B(n5499), .Z(o[567]) );
  XOR U6524 ( .A(n5500), .B(o[566]), .Z(creg_next[566]) );
  AND U6525 ( .A(n3090), .B(n5501), .Z(n5500) );
  XNOR U6526 ( .A(c[566]), .B(n5502), .Z(n5501) );
  IV U6527 ( .A(o[566]), .Z(n5502) );
  XNOR U6528 ( .A(n5503), .B(n5504), .Z(o[566]) );
  XOR U6529 ( .A(n5505), .B(o[565]), .Z(creg_next[565]) );
  AND U6530 ( .A(n3090), .B(n5506), .Z(n5505) );
  XNOR U6531 ( .A(c[565]), .B(n5507), .Z(n5506) );
  IV U6532 ( .A(o[565]), .Z(n5507) );
  XNOR U6533 ( .A(n5508), .B(n5509), .Z(o[565]) );
  XOR U6534 ( .A(n5510), .B(o[564]), .Z(creg_next[564]) );
  AND U6535 ( .A(n3090), .B(n5511), .Z(n5510) );
  XNOR U6536 ( .A(c[564]), .B(n5512), .Z(n5511) );
  IV U6537 ( .A(o[564]), .Z(n5512) );
  XNOR U6538 ( .A(n5513), .B(n5514), .Z(o[564]) );
  XOR U6539 ( .A(n5515), .B(o[563]), .Z(creg_next[563]) );
  AND U6540 ( .A(n3090), .B(n5516), .Z(n5515) );
  XNOR U6541 ( .A(c[563]), .B(n5517), .Z(n5516) );
  IV U6542 ( .A(o[563]), .Z(n5517) );
  XNOR U6543 ( .A(n5518), .B(n5519), .Z(o[563]) );
  XOR U6544 ( .A(n5520), .B(o[562]), .Z(creg_next[562]) );
  AND U6545 ( .A(n3090), .B(n5521), .Z(n5520) );
  XNOR U6546 ( .A(c[562]), .B(n5522), .Z(n5521) );
  IV U6547 ( .A(o[562]), .Z(n5522) );
  XNOR U6548 ( .A(n5523), .B(n5524), .Z(o[562]) );
  XOR U6549 ( .A(n5525), .B(o[561]), .Z(creg_next[561]) );
  AND U6550 ( .A(n3090), .B(n5526), .Z(n5525) );
  XNOR U6551 ( .A(c[561]), .B(n5527), .Z(n5526) );
  IV U6552 ( .A(o[561]), .Z(n5527) );
  XNOR U6553 ( .A(n5528), .B(n5529), .Z(o[561]) );
  XOR U6554 ( .A(n5530), .B(o[560]), .Z(creg_next[560]) );
  AND U6555 ( .A(n3090), .B(n5531), .Z(n5530) );
  XNOR U6556 ( .A(c[560]), .B(n5532), .Z(n5531) );
  IV U6557 ( .A(o[560]), .Z(n5532) );
  XNOR U6558 ( .A(n5533), .B(n5534), .Z(o[560]) );
  XOR U6559 ( .A(n5535), .B(o[55]), .Z(creg_next[55]) );
  AND U6560 ( .A(n3090), .B(n5536), .Z(n5535) );
  XNOR U6561 ( .A(c[55]), .B(n5537), .Z(n5536) );
  IV U6562 ( .A(o[55]), .Z(n5537) );
  XNOR U6563 ( .A(n5538), .B(n5539), .Z(o[55]) );
  XOR U6564 ( .A(n5540), .B(o[559]), .Z(creg_next[559]) );
  AND U6565 ( .A(n3090), .B(n5541), .Z(n5540) );
  XNOR U6566 ( .A(c[559]), .B(n5542), .Z(n5541) );
  IV U6567 ( .A(o[559]), .Z(n5542) );
  XNOR U6568 ( .A(n5543), .B(n5544), .Z(o[559]) );
  XOR U6569 ( .A(n5545), .B(o[558]), .Z(creg_next[558]) );
  AND U6570 ( .A(n3090), .B(n5546), .Z(n5545) );
  XNOR U6571 ( .A(c[558]), .B(n5547), .Z(n5546) );
  IV U6572 ( .A(o[558]), .Z(n5547) );
  XNOR U6573 ( .A(n5548), .B(n5549), .Z(o[558]) );
  XOR U6574 ( .A(n5550), .B(o[557]), .Z(creg_next[557]) );
  AND U6575 ( .A(n3090), .B(n5551), .Z(n5550) );
  XNOR U6576 ( .A(c[557]), .B(n5552), .Z(n5551) );
  IV U6577 ( .A(o[557]), .Z(n5552) );
  XNOR U6578 ( .A(n5553), .B(n5554), .Z(o[557]) );
  XOR U6579 ( .A(n5555), .B(o[556]), .Z(creg_next[556]) );
  AND U6580 ( .A(n3090), .B(n5556), .Z(n5555) );
  XNOR U6581 ( .A(c[556]), .B(n5557), .Z(n5556) );
  IV U6582 ( .A(o[556]), .Z(n5557) );
  XNOR U6583 ( .A(n5558), .B(n5559), .Z(o[556]) );
  XOR U6584 ( .A(n5560), .B(o[555]), .Z(creg_next[555]) );
  AND U6585 ( .A(n3090), .B(n5561), .Z(n5560) );
  XNOR U6586 ( .A(c[555]), .B(n5562), .Z(n5561) );
  IV U6587 ( .A(o[555]), .Z(n5562) );
  XNOR U6588 ( .A(n5563), .B(n5564), .Z(o[555]) );
  XOR U6589 ( .A(n5565), .B(o[554]), .Z(creg_next[554]) );
  AND U6590 ( .A(n3090), .B(n5566), .Z(n5565) );
  XNOR U6591 ( .A(c[554]), .B(n5567), .Z(n5566) );
  IV U6592 ( .A(o[554]), .Z(n5567) );
  XNOR U6593 ( .A(n5568), .B(n5569), .Z(o[554]) );
  XOR U6594 ( .A(n5570), .B(o[553]), .Z(creg_next[553]) );
  AND U6595 ( .A(n3090), .B(n5571), .Z(n5570) );
  XNOR U6596 ( .A(c[553]), .B(n5572), .Z(n5571) );
  IV U6597 ( .A(o[553]), .Z(n5572) );
  XNOR U6598 ( .A(n5573), .B(n5574), .Z(o[553]) );
  XOR U6599 ( .A(n5575), .B(o[552]), .Z(creg_next[552]) );
  AND U6600 ( .A(n3090), .B(n5576), .Z(n5575) );
  XNOR U6601 ( .A(c[552]), .B(n5577), .Z(n5576) );
  IV U6602 ( .A(o[552]), .Z(n5577) );
  XNOR U6603 ( .A(n5578), .B(n5579), .Z(o[552]) );
  XOR U6604 ( .A(n5580), .B(o[551]), .Z(creg_next[551]) );
  AND U6605 ( .A(n3090), .B(n5581), .Z(n5580) );
  XNOR U6606 ( .A(c[551]), .B(n5582), .Z(n5581) );
  IV U6607 ( .A(o[551]), .Z(n5582) );
  XNOR U6608 ( .A(n5583), .B(n5584), .Z(o[551]) );
  XOR U6609 ( .A(n5585), .B(o[550]), .Z(creg_next[550]) );
  AND U6610 ( .A(n3090), .B(n5586), .Z(n5585) );
  XNOR U6611 ( .A(c[550]), .B(n5587), .Z(n5586) );
  IV U6612 ( .A(o[550]), .Z(n5587) );
  XNOR U6613 ( .A(n5588), .B(n5589), .Z(o[550]) );
  XOR U6614 ( .A(n5590), .B(o[54]), .Z(creg_next[54]) );
  AND U6615 ( .A(n3090), .B(n5591), .Z(n5590) );
  XNOR U6616 ( .A(c[54]), .B(n5592), .Z(n5591) );
  IV U6617 ( .A(o[54]), .Z(n5592) );
  XNOR U6618 ( .A(n5593), .B(n5594), .Z(o[54]) );
  XOR U6619 ( .A(n5595), .B(o[549]), .Z(creg_next[549]) );
  AND U6620 ( .A(n3090), .B(n5596), .Z(n5595) );
  XNOR U6621 ( .A(c[549]), .B(n5597), .Z(n5596) );
  IV U6622 ( .A(o[549]), .Z(n5597) );
  XNOR U6623 ( .A(n5598), .B(n5599), .Z(o[549]) );
  XOR U6624 ( .A(n5600), .B(o[548]), .Z(creg_next[548]) );
  AND U6625 ( .A(n3090), .B(n5601), .Z(n5600) );
  XNOR U6626 ( .A(c[548]), .B(n5602), .Z(n5601) );
  IV U6627 ( .A(o[548]), .Z(n5602) );
  XNOR U6628 ( .A(n5603), .B(n5604), .Z(o[548]) );
  XOR U6629 ( .A(n5605), .B(o[547]), .Z(creg_next[547]) );
  AND U6630 ( .A(n3090), .B(n5606), .Z(n5605) );
  XNOR U6631 ( .A(c[547]), .B(n5607), .Z(n5606) );
  IV U6632 ( .A(o[547]), .Z(n5607) );
  XNOR U6633 ( .A(n5608), .B(n5609), .Z(o[547]) );
  XOR U6634 ( .A(n5610), .B(o[546]), .Z(creg_next[546]) );
  AND U6635 ( .A(n3090), .B(n5611), .Z(n5610) );
  XNOR U6636 ( .A(c[546]), .B(n5612), .Z(n5611) );
  IV U6637 ( .A(o[546]), .Z(n5612) );
  XNOR U6638 ( .A(n5613), .B(n5614), .Z(o[546]) );
  XOR U6639 ( .A(n5615), .B(o[545]), .Z(creg_next[545]) );
  AND U6640 ( .A(n3090), .B(n5616), .Z(n5615) );
  XNOR U6641 ( .A(c[545]), .B(n5617), .Z(n5616) );
  IV U6642 ( .A(o[545]), .Z(n5617) );
  XNOR U6643 ( .A(n5618), .B(n5619), .Z(o[545]) );
  XOR U6644 ( .A(n5620), .B(o[544]), .Z(creg_next[544]) );
  AND U6645 ( .A(n3090), .B(n5621), .Z(n5620) );
  XNOR U6646 ( .A(c[544]), .B(n5622), .Z(n5621) );
  IV U6647 ( .A(o[544]), .Z(n5622) );
  XNOR U6648 ( .A(n5623), .B(n5624), .Z(o[544]) );
  XOR U6649 ( .A(n5625), .B(o[543]), .Z(creg_next[543]) );
  AND U6650 ( .A(n3090), .B(n5626), .Z(n5625) );
  XNOR U6651 ( .A(c[543]), .B(n5627), .Z(n5626) );
  IV U6652 ( .A(o[543]), .Z(n5627) );
  XNOR U6653 ( .A(n5628), .B(n5629), .Z(o[543]) );
  XOR U6654 ( .A(n5630), .B(o[542]), .Z(creg_next[542]) );
  AND U6655 ( .A(n3090), .B(n5631), .Z(n5630) );
  XNOR U6656 ( .A(c[542]), .B(n5632), .Z(n5631) );
  IV U6657 ( .A(o[542]), .Z(n5632) );
  XNOR U6658 ( .A(n5633), .B(n5634), .Z(o[542]) );
  XOR U6659 ( .A(n5635), .B(o[541]), .Z(creg_next[541]) );
  AND U6660 ( .A(n3090), .B(n5636), .Z(n5635) );
  XNOR U6661 ( .A(c[541]), .B(n5637), .Z(n5636) );
  IV U6662 ( .A(o[541]), .Z(n5637) );
  XNOR U6663 ( .A(n5638), .B(n5639), .Z(o[541]) );
  XOR U6664 ( .A(n5640), .B(o[540]), .Z(creg_next[540]) );
  AND U6665 ( .A(n3090), .B(n5641), .Z(n5640) );
  XNOR U6666 ( .A(c[540]), .B(n5642), .Z(n5641) );
  IV U6667 ( .A(o[540]), .Z(n5642) );
  XNOR U6668 ( .A(n5643), .B(n5644), .Z(o[540]) );
  XOR U6669 ( .A(n5645), .B(o[53]), .Z(creg_next[53]) );
  AND U6670 ( .A(n3090), .B(n5646), .Z(n5645) );
  XNOR U6671 ( .A(c[53]), .B(n5647), .Z(n5646) );
  IV U6672 ( .A(o[53]), .Z(n5647) );
  XNOR U6673 ( .A(n5648), .B(n5649), .Z(o[53]) );
  XOR U6674 ( .A(n5650), .B(o[539]), .Z(creg_next[539]) );
  AND U6675 ( .A(n3090), .B(n5651), .Z(n5650) );
  XNOR U6676 ( .A(c[539]), .B(n5652), .Z(n5651) );
  IV U6677 ( .A(o[539]), .Z(n5652) );
  XNOR U6678 ( .A(n5653), .B(n5654), .Z(o[539]) );
  XOR U6679 ( .A(n5655), .B(o[538]), .Z(creg_next[538]) );
  AND U6680 ( .A(n3090), .B(n5656), .Z(n5655) );
  XNOR U6681 ( .A(c[538]), .B(n5657), .Z(n5656) );
  IV U6682 ( .A(o[538]), .Z(n5657) );
  XNOR U6683 ( .A(n5658), .B(n5659), .Z(o[538]) );
  XOR U6684 ( .A(n5660), .B(o[537]), .Z(creg_next[537]) );
  AND U6685 ( .A(n3090), .B(n5661), .Z(n5660) );
  XNOR U6686 ( .A(c[537]), .B(n5662), .Z(n5661) );
  IV U6687 ( .A(o[537]), .Z(n5662) );
  XNOR U6688 ( .A(n5663), .B(n5664), .Z(o[537]) );
  XOR U6689 ( .A(n5665), .B(o[536]), .Z(creg_next[536]) );
  AND U6690 ( .A(n3090), .B(n5666), .Z(n5665) );
  XNOR U6691 ( .A(c[536]), .B(n5667), .Z(n5666) );
  IV U6692 ( .A(o[536]), .Z(n5667) );
  XNOR U6693 ( .A(n5668), .B(n5669), .Z(o[536]) );
  XOR U6694 ( .A(n5670), .B(o[535]), .Z(creg_next[535]) );
  AND U6695 ( .A(n3090), .B(n5671), .Z(n5670) );
  XNOR U6696 ( .A(c[535]), .B(n5672), .Z(n5671) );
  IV U6697 ( .A(o[535]), .Z(n5672) );
  XNOR U6698 ( .A(n5673), .B(n5674), .Z(o[535]) );
  XOR U6699 ( .A(n5675), .B(o[534]), .Z(creg_next[534]) );
  AND U6700 ( .A(n3090), .B(n5676), .Z(n5675) );
  XNOR U6701 ( .A(c[534]), .B(n5677), .Z(n5676) );
  IV U6702 ( .A(o[534]), .Z(n5677) );
  XNOR U6703 ( .A(n5678), .B(n5679), .Z(o[534]) );
  XOR U6704 ( .A(n5680), .B(o[533]), .Z(creg_next[533]) );
  AND U6705 ( .A(n3090), .B(n5681), .Z(n5680) );
  XNOR U6706 ( .A(c[533]), .B(n5682), .Z(n5681) );
  IV U6707 ( .A(o[533]), .Z(n5682) );
  XNOR U6708 ( .A(n5683), .B(n5684), .Z(o[533]) );
  XOR U6709 ( .A(n5685), .B(o[532]), .Z(creg_next[532]) );
  AND U6710 ( .A(n3090), .B(n5686), .Z(n5685) );
  XNOR U6711 ( .A(c[532]), .B(n5687), .Z(n5686) );
  IV U6712 ( .A(o[532]), .Z(n5687) );
  XNOR U6713 ( .A(n5688), .B(n5689), .Z(o[532]) );
  XOR U6714 ( .A(n5690), .B(o[531]), .Z(creg_next[531]) );
  AND U6715 ( .A(n3090), .B(n5691), .Z(n5690) );
  XNOR U6716 ( .A(c[531]), .B(n5692), .Z(n5691) );
  IV U6717 ( .A(o[531]), .Z(n5692) );
  XNOR U6718 ( .A(n5693), .B(n5694), .Z(o[531]) );
  XOR U6719 ( .A(n5695), .B(o[530]), .Z(creg_next[530]) );
  AND U6720 ( .A(n3090), .B(n5696), .Z(n5695) );
  XNOR U6721 ( .A(c[530]), .B(n5697), .Z(n5696) );
  IV U6722 ( .A(o[530]), .Z(n5697) );
  XNOR U6723 ( .A(n5698), .B(n5699), .Z(o[530]) );
  XOR U6724 ( .A(n5700), .B(o[52]), .Z(creg_next[52]) );
  AND U6725 ( .A(n3090), .B(n5701), .Z(n5700) );
  XNOR U6726 ( .A(c[52]), .B(n5702), .Z(n5701) );
  IV U6727 ( .A(o[52]), .Z(n5702) );
  XNOR U6728 ( .A(n5703), .B(n5704), .Z(o[52]) );
  XOR U6729 ( .A(n5705), .B(o[529]), .Z(creg_next[529]) );
  AND U6730 ( .A(n3090), .B(n5706), .Z(n5705) );
  XNOR U6731 ( .A(c[529]), .B(n5707), .Z(n5706) );
  IV U6732 ( .A(o[529]), .Z(n5707) );
  XNOR U6733 ( .A(n5708), .B(n5709), .Z(o[529]) );
  XOR U6734 ( .A(n5710), .B(o[528]), .Z(creg_next[528]) );
  AND U6735 ( .A(n3090), .B(n5711), .Z(n5710) );
  XNOR U6736 ( .A(c[528]), .B(n5712), .Z(n5711) );
  IV U6737 ( .A(o[528]), .Z(n5712) );
  XNOR U6738 ( .A(n5713), .B(n5714), .Z(o[528]) );
  XOR U6739 ( .A(n5715), .B(o[527]), .Z(creg_next[527]) );
  AND U6740 ( .A(n3090), .B(n5716), .Z(n5715) );
  XNOR U6741 ( .A(c[527]), .B(n5717), .Z(n5716) );
  IV U6742 ( .A(o[527]), .Z(n5717) );
  XNOR U6743 ( .A(n5718), .B(n5719), .Z(o[527]) );
  XOR U6744 ( .A(n5720), .B(o[526]), .Z(creg_next[526]) );
  AND U6745 ( .A(n3090), .B(n5721), .Z(n5720) );
  XNOR U6746 ( .A(c[526]), .B(n5722), .Z(n5721) );
  IV U6747 ( .A(o[526]), .Z(n5722) );
  XNOR U6748 ( .A(n5723), .B(n5724), .Z(o[526]) );
  XOR U6749 ( .A(n5725), .B(o[525]), .Z(creg_next[525]) );
  AND U6750 ( .A(n3090), .B(n5726), .Z(n5725) );
  XNOR U6751 ( .A(c[525]), .B(n5727), .Z(n5726) );
  IV U6752 ( .A(o[525]), .Z(n5727) );
  XNOR U6753 ( .A(n5728), .B(n5729), .Z(o[525]) );
  XOR U6754 ( .A(n5730), .B(o[524]), .Z(creg_next[524]) );
  AND U6755 ( .A(n3090), .B(n5731), .Z(n5730) );
  XNOR U6756 ( .A(c[524]), .B(n5732), .Z(n5731) );
  IV U6757 ( .A(o[524]), .Z(n5732) );
  XNOR U6758 ( .A(n5733), .B(n5734), .Z(o[524]) );
  XOR U6759 ( .A(n5735), .B(o[523]), .Z(creg_next[523]) );
  AND U6760 ( .A(n3090), .B(n5736), .Z(n5735) );
  XNOR U6761 ( .A(c[523]), .B(n5737), .Z(n5736) );
  IV U6762 ( .A(o[523]), .Z(n5737) );
  XNOR U6763 ( .A(n5738), .B(n5739), .Z(o[523]) );
  XOR U6764 ( .A(n5740), .B(o[522]), .Z(creg_next[522]) );
  AND U6765 ( .A(n3090), .B(n5741), .Z(n5740) );
  XNOR U6766 ( .A(c[522]), .B(n5742), .Z(n5741) );
  IV U6767 ( .A(o[522]), .Z(n5742) );
  XNOR U6768 ( .A(n5743), .B(n5744), .Z(o[522]) );
  XOR U6769 ( .A(n5745), .B(o[521]), .Z(creg_next[521]) );
  AND U6770 ( .A(n3090), .B(n5746), .Z(n5745) );
  XNOR U6771 ( .A(c[521]), .B(n5747), .Z(n5746) );
  IV U6772 ( .A(o[521]), .Z(n5747) );
  XNOR U6773 ( .A(n5748), .B(n5749), .Z(o[521]) );
  XOR U6774 ( .A(n5750), .B(o[520]), .Z(creg_next[520]) );
  AND U6775 ( .A(n3090), .B(n5751), .Z(n5750) );
  XNOR U6776 ( .A(c[520]), .B(n5752), .Z(n5751) );
  IV U6777 ( .A(o[520]), .Z(n5752) );
  XNOR U6778 ( .A(n5753), .B(n5754), .Z(o[520]) );
  XOR U6779 ( .A(n5755), .B(o[51]), .Z(creg_next[51]) );
  AND U6780 ( .A(n3090), .B(n5756), .Z(n5755) );
  XNOR U6781 ( .A(c[51]), .B(n5757), .Z(n5756) );
  IV U6782 ( .A(o[51]), .Z(n5757) );
  XNOR U6783 ( .A(n5758), .B(n5759), .Z(o[51]) );
  XOR U6784 ( .A(n5760), .B(o[519]), .Z(creg_next[519]) );
  AND U6785 ( .A(n3090), .B(n5761), .Z(n5760) );
  XNOR U6786 ( .A(c[519]), .B(n5762), .Z(n5761) );
  IV U6787 ( .A(o[519]), .Z(n5762) );
  XNOR U6788 ( .A(n5763), .B(n5764), .Z(o[519]) );
  XOR U6789 ( .A(n5765), .B(o[518]), .Z(creg_next[518]) );
  AND U6790 ( .A(n3090), .B(n5766), .Z(n5765) );
  XNOR U6791 ( .A(c[518]), .B(n5767), .Z(n5766) );
  IV U6792 ( .A(o[518]), .Z(n5767) );
  XNOR U6793 ( .A(n5768), .B(n5769), .Z(o[518]) );
  XOR U6794 ( .A(n5770), .B(o[517]), .Z(creg_next[517]) );
  AND U6795 ( .A(n3090), .B(n5771), .Z(n5770) );
  XNOR U6796 ( .A(c[517]), .B(n5772), .Z(n5771) );
  IV U6797 ( .A(o[517]), .Z(n5772) );
  XNOR U6798 ( .A(n5773), .B(n5774), .Z(o[517]) );
  XOR U6799 ( .A(n5775), .B(o[516]), .Z(creg_next[516]) );
  AND U6800 ( .A(n3090), .B(n5776), .Z(n5775) );
  XNOR U6801 ( .A(c[516]), .B(n5777), .Z(n5776) );
  IV U6802 ( .A(o[516]), .Z(n5777) );
  XNOR U6803 ( .A(n5778), .B(n5779), .Z(o[516]) );
  XOR U6804 ( .A(n5780), .B(o[515]), .Z(creg_next[515]) );
  AND U6805 ( .A(n3090), .B(n5781), .Z(n5780) );
  XNOR U6806 ( .A(c[515]), .B(n5782), .Z(n5781) );
  IV U6807 ( .A(o[515]), .Z(n5782) );
  XNOR U6808 ( .A(n5783), .B(n5784), .Z(o[515]) );
  XOR U6809 ( .A(n5785), .B(o[514]), .Z(creg_next[514]) );
  AND U6810 ( .A(n3090), .B(n5786), .Z(n5785) );
  XNOR U6811 ( .A(c[514]), .B(n5787), .Z(n5786) );
  IV U6812 ( .A(o[514]), .Z(n5787) );
  XNOR U6813 ( .A(n5788), .B(n5789), .Z(o[514]) );
  XOR U6814 ( .A(n5790), .B(o[513]), .Z(creg_next[513]) );
  AND U6815 ( .A(n3090), .B(n5791), .Z(n5790) );
  XNOR U6816 ( .A(c[513]), .B(n5792), .Z(n5791) );
  IV U6817 ( .A(o[513]), .Z(n5792) );
  XNOR U6818 ( .A(n5793), .B(n5794), .Z(o[513]) );
  XOR U6819 ( .A(n5795), .B(o[512]), .Z(creg_next[512]) );
  AND U6820 ( .A(n3090), .B(n5796), .Z(n5795) );
  XNOR U6821 ( .A(c[512]), .B(n5797), .Z(n5796) );
  IV U6822 ( .A(o[512]), .Z(n5797) );
  XNOR U6823 ( .A(n5798), .B(n5799), .Z(o[512]) );
  XOR U6824 ( .A(n5800), .B(o[511]), .Z(creg_next[511]) );
  AND U6825 ( .A(n3090), .B(n5801), .Z(n5800) );
  XNOR U6826 ( .A(c[511]), .B(n5802), .Z(n5801) );
  IV U6827 ( .A(o[511]), .Z(n5802) );
  XNOR U6828 ( .A(n5803), .B(n5804), .Z(o[511]) );
  XOR U6829 ( .A(n5805), .B(o[510]), .Z(creg_next[510]) );
  AND U6830 ( .A(n3090), .B(n5806), .Z(n5805) );
  XNOR U6831 ( .A(c[510]), .B(n5807), .Z(n5806) );
  IV U6832 ( .A(o[510]), .Z(n5807) );
  XNOR U6833 ( .A(n5808), .B(n5809), .Z(o[510]) );
  XOR U6834 ( .A(n5810), .B(o[50]), .Z(creg_next[50]) );
  AND U6835 ( .A(n3090), .B(n5811), .Z(n5810) );
  XNOR U6836 ( .A(c[50]), .B(n5812), .Z(n5811) );
  IV U6837 ( .A(o[50]), .Z(n5812) );
  XNOR U6838 ( .A(n5813), .B(n5814), .Z(o[50]) );
  XOR U6839 ( .A(n5815), .B(o[509]), .Z(creg_next[509]) );
  AND U6840 ( .A(n3090), .B(n5816), .Z(n5815) );
  XNOR U6841 ( .A(c[509]), .B(n5817), .Z(n5816) );
  IV U6842 ( .A(o[509]), .Z(n5817) );
  XNOR U6843 ( .A(n5818), .B(n5819), .Z(o[509]) );
  XOR U6844 ( .A(n5820), .B(o[508]), .Z(creg_next[508]) );
  AND U6845 ( .A(n3090), .B(n5821), .Z(n5820) );
  XNOR U6846 ( .A(c[508]), .B(n5822), .Z(n5821) );
  IV U6847 ( .A(o[508]), .Z(n5822) );
  XNOR U6848 ( .A(n5823), .B(n5824), .Z(o[508]) );
  XOR U6849 ( .A(n5825), .B(o[507]), .Z(creg_next[507]) );
  AND U6850 ( .A(n3090), .B(n5826), .Z(n5825) );
  XNOR U6851 ( .A(c[507]), .B(n5827), .Z(n5826) );
  IV U6852 ( .A(o[507]), .Z(n5827) );
  XNOR U6853 ( .A(n5828), .B(n5829), .Z(o[507]) );
  XOR U6854 ( .A(n5830), .B(o[506]), .Z(creg_next[506]) );
  AND U6855 ( .A(n3090), .B(n5831), .Z(n5830) );
  XNOR U6856 ( .A(c[506]), .B(n5832), .Z(n5831) );
  IV U6857 ( .A(o[506]), .Z(n5832) );
  XNOR U6858 ( .A(n5833), .B(n5834), .Z(o[506]) );
  XOR U6859 ( .A(n5835), .B(o[505]), .Z(creg_next[505]) );
  AND U6860 ( .A(n3090), .B(n5836), .Z(n5835) );
  XNOR U6861 ( .A(c[505]), .B(n5837), .Z(n5836) );
  IV U6862 ( .A(o[505]), .Z(n5837) );
  XNOR U6863 ( .A(n5838), .B(n5839), .Z(o[505]) );
  XOR U6864 ( .A(n5840), .B(o[504]), .Z(creg_next[504]) );
  AND U6865 ( .A(n3090), .B(n5841), .Z(n5840) );
  XNOR U6866 ( .A(c[504]), .B(n5842), .Z(n5841) );
  IV U6867 ( .A(o[504]), .Z(n5842) );
  XNOR U6868 ( .A(n5843), .B(n5844), .Z(o[504]) );
  XOR U6869 ( .A(n5845), .B(o[503]), .Z(creg_next[503]) );
  AND U6870 ( .A(n3090), .B(n5846), .Z(n5845) );
  XNOR U6871 ( .A(c[503]), .B(n5847), .Z(n5846) );
  IV U6872 ( .A(o[503]), .Z(n5847) );
  XNOR U6873 ( .A(n5848), .B(n5849), .Z(o[503]) );
  XOR U6874 ( .A(n5850), .B(o[502]), .Z(creg_next[502]) );
  AND U6875 ( .A(n3090), .B(n5851), .Z(n5850) );
  XNOR U6876 ( .A(c[502]), .B(n5852), .Z(n5851) );
  IV U6877 ( .A(o[502]), .Z(n5852) );
  XNOR U6878 ( .A(n5853), .B(n5854), .Z(o[502]) );
  XOR U6879 ( .A(n5855), .B(o[501]), .Z(creg_next[501]) );
  AND U6880 ( .A(n3090), .B(n5856), .Z(n5855) );
  XNOR U6881 ( .A(c[501]), .B(n5857), .Z(n5856) );
  IV U6882 ( .A(o[501]), .Z(n5857) );
  XNOR U6883 ( .A(n5858), .B(n5859), .Z(o[501]) );
  XOR U6884 ( .A(n5860), .B(o[500]), .Z(creg_next[500]) );
  AND U6885 ( .A(n3090), .B(n5861), .Z(n5860) );
  XNOR U6886 ( .A(c[500]), .B(n5862), .Z(n5861) );
  IV U6887 ( .A(o[500]), .Z(n5862) );
  XNOR U6888 ( .A(n5863), .B(n5864), .Z(o[500]) );
  XOR U6889 ( .A(n5865), .B(o[4]), .Z(creg_next[4]) );
  AND U6890 ( .A(n3090), .B(n5866), .Z(n5865) );
  XNOR U6891 ( .A(c[4]), .B(n5867), .Z(n5866) );
  IV U6892 ( .A(o[4]), .Z(n5867) );
  XNOR U6893 ( .A(n5868), .B(n5869), .Z(o[4]) );
  XOR U6894 ( .A(n5870), .B(o[49]), .Z(creg_next[49]) );
  AND U6895 ( .A(n3090), .B(n5871), .Z(n5870) );
  XNOR U6896 ( .A(c[49]), .B(n5872), .Z(n5871) );
  IV U6897 ( .A(o[49]), .Z(n5872) );
  XNOR U6898 ( .A(n5873), .B(n5874), .Z(o[49]) );
  XOR U6899 ( .A(n5875), .B(o[499]), .Z(creg_next[499]) );
  AND U6900 ( .A(n3090), .B(n5876), .Z(n5875) );
  XNOR U6901 ( .A(c[499]), .B(n5877), .Z(n5876) );
  IV U6902 ( .A(o[499]), .Z(n5877) );
  XNOR U6903 ( .A(n5878), .B(n5879), .Z(o[499]) );
  XOR U6904 ( .A(n5880), .B(o[498]), .Z(creg_next[498]) );
  AND U6905 ( .A(n3090), .B(n5881), .Z(n5880) );
  XNOR U6906 ( .A(c[498]), .B(n5882), .Z(n5881) );
  IV U6907 ( .A(o[498]), .Z(n5882) );
  XNOR U6908 ( .A(n5883), .B(n5884), .Z(o[498]) );
  XOR U6909 ( .A(n5885), .B(o[497]), .Z(creg_next[497]) );
  AND U6910 ( .A(n3090), .B(n5886), .Z(n5885) );
  XNOR U6911 ( .A(c[497]), .B(n5887), .Z(n5886) );
  IV U6912 ( .A(o[497]), .Z(n5887) );
  XNOR U6913 ( .A(n5888), .B(n5889), .Z(o[497]) );
  XOR U6914 ( .A(n5890), .B(o[496]), .Z(creg_next[496]) );
  AND U6915 ( .A(n3090), .B(n5891), .Z(n5890) );
  XNOR U6916 ( .A(c[496]), .B(n5892), .Z(n5891) );
  IV U6917 ( .A(o[496]), .Z(n5892) );
  XNOR U6918 ( .A(n5893), .B(n5894), .Z(o[496]) );
  XOR U6919 ( .A(n5895), .B(o[495]), .Z(creg_next[495]) );
  AND U6920 ( .A(n3090), .B(n5896), .Z(n5895) );
  XNOR U6921 ( .A(c[495]), .B(n5897), .Z(n5896) );
  IV U6922 ( .A(o[495]), .Z(n5897) );
  XNOR U6923 ( .A(n5898), .B(n5899), .Z(o[495]) );
  XOR U6924 ( .A(n5900), .B(o[494]), .Z(creg_next[494]) );
  AND U6925 ( .A(n3090), .B(n5901), .Z(n5900) );
  XNOR U6926 ( .A(c[494]), .B(n5902), .Z(n5901) );
  IV U6927 ( .A(o[494]), .Z(n5902) );
  XNOR U6928 ( .A(n5903), .B(n5904), .Z(o[494]) );
  XOR U6929 ( .A(n5905), .B(o[493]), .Z(creg_next[493]) );
  AND U6930 ( .A(n3090), .B(n5906), .Z(n5905) );
  XNOR U6931 ( .A(c[493]), .B(n5907), .Z(n5906) );
  IV U6932 ( .A(o[493]), .Z(n5907) );
  XNOR U6933 ( .A(n5908), .B(n5909), .Z(o[493]) );
  XOR U6934 ( .A(n5910), .B(o[492]), .Z(creg_next[492]) );
  AND U6935 ( .A(n3090), .B(n5911), .Z(n5910) );
  XNOR U6936 ( .A(c[492]), .B(n5912), .Z(n5911) );
  IV U6937 ( .A(o[492]), .Z(n5912) );
  XNOR U6938 ( .A(n5913), .B(n5914), .Z(o[492]) );
  XOR U6939 ( .A(n5915), .B(o[491]), .Z(creg_next[491]) );
  AND U6940 ( .A(n3090), .B(n5916), .Z(n5915) );
  XNOR U6941 ( .A(c[491]), .B(n5917), .Z(n5916) );
  IV U6942 ( .A(o[491]), .Z(n5917) );
  XNOR U6943 ( .A(n5918), .B(n5919), .Z(o[491]) );
  XOR U6944 ( .A(n5920), .B(o[490]), .Z(creg_next[490]) );
  AND U6945 ( .A(n3090), .B(n5921), .Z(n5920) );
  XNOR U6946 ( .A(c[490]), .B(n5922), .Z(n5921) );
  IV U6947 ( .A(o[490]), .Z(n5922) );
  XNOR U6948 ( .A(n5923), .B(n5924), .Z(o[490]) );
  XOR U6949 ( .A(n5925), .B(o[48]), .Z(creg_next[48]) );
  AND U6950 ( .A(n3090), .B(n5926), .Z(n5925) );
  XNOR U6951 ( .A(c[48]), .B(n5927), .Z(n5926) );
  IV U6952 ( .A(o[48]), .Z(n5927) );
  XNOR U6953 ( .A(n5928), .B(n5929), .Z(o[48]) );
  XOR U6954 ( .A(n5930), .B(o[489]), .Z(creg_next[489]) );
  AND U6955 ( .A(n3090), .B(n5931), .Z(n5930) );
  XNOR U6956 ( .A(c[489]), .B(n5932), .Z(n5931) );
  IV U6957 ( .A(o[489]), .Z(n5932) );
  XNOR U6958 ( .A(n5933), .B(n5934), .Z(o[489]) );
  XOR U6959 ( .A(n5935), .B(o[488]), .Z(creg_next[488]) );
  AND U6960 ( .A(n3090), .B(n5936), .Z(n5935) );
  XNOR U6961 ( .A(c[488]), .B(n5937), .Z(n5936) );
  IV U6962 ( .A(o[488]), .Z(n5937) );
  XNOR U6963 ( .A(n5938), .B(n5939), .Z(o[488]) );
  XOR U6964 ( .A(n5940), .B(o[487]), .Z(creg_next[487]) );
  AND U6965 ( .A(n3090), .B(n5941), .Z(n5940) );
  XNOR U6966 ( .A(c[487]), .B(n5942), .Z(n5941) );
  IV U6967 ( .A(o[487]), .Z(n5942) );
  XNOR U6968 ( .A(n5943), .B(n5944), .Z(o[487]) );
  XOR U6969 ( .A(n5945), .B(o[486]), .Z(creg_next[486]) );
  AND U6970 ( .A(n3090), .B(n5946), .Z(n5945) );
  XNOR U6971 ( .A(c[486]), .B(n5947), .Z(n5946) );
  IV U6972 ( .A(o[486]), .Z(n5947) );
  XNOR U6973 ( .A(n5948), .B(n5949), .Z(o[486]) );
  XOR U6974 ( .A(n5950), .B(o[485]), .Z(creg_next[485]) );
  AND U6975 ( .A(n3090), .B(n5951), .Z(n5950) );
  XNOR U6976 ( .A(c[485]), .B(n5952), .Z(n5951) );
  IV U6977 ( .A(o[485]), .Z(n5952) );
  XNOR U6978 ( .A(n5953), .B(n5954), .Z(o[485]) );
  XOR U6979 ( .A(n5955), .B(o[484]), .Z(creg_next[484]) );
  AND U6980 ( .A(n3090), .B(n5956), .Z(n5955) );
  XNOR U6981 ( .A(c[484]), .B(n5957), .Z(n5956) );
  IV U6982 ( .A(o[484]), .Z(n5957) );
  XNOR U6983 ( .A(n5958), .B(n5959), .Z(o[484]) );
  XOR U6984 ( .A(n5960), .B(o[483]), .Z(creg_next[483]) );
  AND U6985 ( .A(n3090), .B(n5961), .Z(n5960) );
  XNOR U6986 ( .A(c[483]), .B(n5962), .Z(n5961) );
  IV U6987 ( .A(o[483]), .Z(n5962) );
  XNOR U6988 ( .A(n5963), .B(n5964), .Z(o[483]) );
  XOR U6989 ( .A(n5965), .B(o[482]), .Z(creg_next[482]) );
  AND U6990 ( .A(n3090), .B(n5966), .Z(n5965) );
  XNOR U6991 ( .A(c[482]), .B(n5967), .Z(n5966) );
  IV U6992 ( .A(o[482]), .Z(n5967) );
  XNOR U6993 ( .A(n5968), .B(n5969), .Z(o[482]) );
  XOR U6994 ( .A(n5970), .B(o[481]), .Z(creg_next[481]) );
  AND U6995 ( .A(n3090), .B(n5971), .Z(n5970) );
  XNOR U6996 ( .A(c[481]), .B(n5972), .Z(n5971) );
  IV U6997 ( .A(o[481]), .Z(n5972) );
  XNOR U6998 ( .A(n5973), .B(n5974), .Z(o[481]) );
  XOR U6999 ( .A(n5975), .B(o[480]), .Z(creg_next[480]) );
  AND U7000 ( .A(n3090), .B(n5976), .Z(n5975) );
  XNOR U7001 ( .A(c[480]), .B(n5977), .Z(n5976) );
  IV U7002 ( .A(o[480]), .Z(n5977) );
  XNOR U7003 ( .A(n5978), .B(n5979), .Z(o[480]) );
  XOR U7004 ( .A(n5980), .B(o[47]), .Z(creg_next[47]) );
  AND U7005 ( .A(n3090), .B(n5981), .Z(n5980) );
  XNOR U7006 ( .A(c[47]), .B(n5982), .Z(n5981) );
  IV U7007 ( .A(o[47]), .Z(n5982) );
  XNOR U7008 ( .A(n5983), .B(n5984), .Z(o[47]) );
  XOR U7009 ( .A(n5985), .B(o[479]), .Z(creg_next[479]) );
  AND U7010 ( .A(n3090), .B(n5986), .Z(n5985) );
  XNOR U7011 ( .A(c[479]), .B(n5987), .Z(n5986) );
  IV U7012 ( .A(o[479]), .Z(n5987) );
  XNOR U7013 ( .A(n5988), .B(n5989), .Z(o[479]) );
  XOR U7014 ( .A(n5990), .B(o[478]), .Z(creg_next[478]) );
  AND U7015 ( .A(n3090), .B(n5991), .Z(n5990) );
  XNOR U7016 ( .A(c[478]), .B(n5992), .Z(n5991) );
  IV U7017 ( .A(o[478]), .Z(n5992) );
  XNOR U7018 ( .A(n5993), .B(n5994), .Z(o[478]) );
  XOR U7019 ( .A(n5995), .B(o[477]), .Z(creg_next[477]) );
  AND U7020 ( .A(n3090), .B(n5996), .Z(n5995) );
  XNOR U7021 ( .A(c[477]), .B(n5997), .Z(n5996) );
  IV U7022 ( .A(o[477]), .Z(n5997) );
  XNOR U7023 ( .A(n5998), .B(n5999), .Z(o[477]) );
  XOR U7024 ( .A(n6000), .B(o[476]), .Z(creg_next[476]) );
  AND U7025 ( .A(n3090), .B(n6001), .Z(n6000) );
  XNOR U7026 ( .A(c[476]), .B(n6002), .Z(n6001) );
  IV U7027 ( .A(o[476]), .Z(n6002) );
  XNOR U7028 ( .A(n6003), .B(n6004), .Z(o[476]) );
  XOR U7029 ( .A(n6005), .B(o[475]), .Z(creg_next[475]) );
  AND U7030 ( .A(n3090), .B(n6006), .Z(n6005) );
  XNOR U7031 ( .A(c[475]), .B(n6007), .Z(n6006) );
  IV U7032 ( .A(o[475]), .Z(n6007) );
  XNOR U7033 ( .A(n6008), .B(n6009), .Z(o[475]) );
  XOR U7034 ( .A(n6010), .B(o[474]), .Z(creg_next[474]) );
  AND U7035 ( .A(n3090), .B(n6011), .Z(n6010) );
  XNOR U7036 ( .A(c[474]), .B(n6012), .Z(n6011) );
  IV U7037 ( .A(o[474]), .Z(n6012) );
  XNOR U7038 ( .A(n6013), .B(n6014), .Z(o[474]) );
  XOR U7039 ( .A(n6015), .B(o[473]), .Z(creg_next[473]) );
  AND U7040 ( .A(n3090), .B(n6016), .Z(n6015) );
  XNOR U7041 ( .A(c[473]), .B(n6017), .Z(n6016) );
  IV U7042 ( .A(o[473]), .Z(n6017) );
  XNOR U7043 ( .A(n6018), .B(n6019), .Z(o[473]) );
  XOR U7044 ( .A(n6020), .B(o[472]), .Z(creg_next[472]) );
  AND U7045 ( .A(n3090), .B(n6021), .Z(n6020) );
  XNOR U7046 ( .A(c[472]), .B(n6022), .Z(n6021) );
  IV U7047 ( .A(o[472]), .Z(n6022) );
  XNOR U7048 ( .A(n6023), .B(n6024), .Z(o[472]) );
  XOR U7049 ( .A(n6025), .B(o[471]), .Z(creg_next[471]) );
  AND U7050 ( .A(n3090), .B(n6026), .Z(n6025) );
  XNOR U7051 ( .A(c[471]), .B(n6027), .Z(n6026) );
  IV U7052 ( .A(o[471]), .Z(n6027) );
  XNOR U7053 ( .A(n6028), .B(n6029), .Z(o[471]) );
  XOR U7054 ( .A(n6030), .B(o[470]), .Z(creg_next[470]) );
  AND U7055 ( .A(n3090), .B(n6031), .Z(n6030) );
  XNOR U7056 ( .A(c[470]), .B(n6032), .Z(n6031) );
  IV U7057 ( .A(o[470]), .Z(n6032) );
  XNOR U7058 ( .A(n6033), .B(n6034), .Z(o[470]) );
  XOR U7059 ( .A(n6035), .B(o[46]), .Z(creg_next[46]) );
  AND U7060 ( .A(n3090), .B(n6036), .Z(n6035) );
  XNOR U7061 ( .A(c[46]), .B(n6037), .Z(n6036) );
  IV U7062 ( .A(o[46]), .Z(n6037) );
  XNOR U7063 ( .A(n6038), .B(n6039), .Z(o[46]) );
  XOR U7064 ( .A(n6040), .B(o[469]), .Z(creg_next[469]) );
  AND U7065 ( .A(n3090), .B(n6041), .Z(n6040) );
  XNOR U7066 ( .A(c[469]), .B(n6042), .Z(n6041) );
  IV U7067 ( .A(o[469]), .Z(n6042) );
  XNOR U7068 ( .A(n6043), .B(n6044), .Z(o[469]) );
  XOR U7069 ( .A(n6045), .B(o[468]), .Z(creg_next[468]) );
  AND U7070 ( .A(n3090), .B(n6046), .Z(n6045) );
  XNOR U7071 ( .A(c[468]), .B(n6047), .Z(n6046) );
  IV U7072 ( .A(o[468]), .Z(n6047) );
  XNOR U7073 ( .A(n6048), .B(n6049), .Z(o[468]) );
  XOR U7074 ( .A(n6050), .B(o[467]), .Z(creg_next[467]) );
  AND U7075 ( .A(n3090), .B(n6051), .Z(n6050) );
  XNOR U7076 ( .A(c[467]), .B(n6052), .Z(n6051) );
  IV U7077 ( .A(o[467]), .Z(n6052) );
  XNOR U7078 ( .A(n6053), .B(n6054), .Z(o[467]) );
  XOR U7079 ( .A(n6055), .B(o[466]), .Z(creg_next[466]) );
  AND U7080 ( .A(n3090), .B(n6056), .Z(n6055) );
  XNOR U7081 ( .A(c[466]), .B(n6057), .Z(n6056) );
  IV U7082 ( .A(o[466]), .Z(n6057) );
  XNOR U7083 ( .A(n6058), .B(n6059), .Z(o[466]) );
  XOR U7084 ( .A(n6060), .B(o[465]), .Z(creg_next[465]) );
  AND U7085 ( .A(n3090), .B(n6061), .Z(n6060) );
  XNOR U7086 ( .A(c[465]), .B(n6062), .Z(n6061) );
  IV U7087 ( .A(o[465]), .Z(n6062) );
  XNOR U7088 ( .A(n6063), .B(n6064), .Z(o[465]) );
  XOR U7089 ( .A(n6065), .B(o[464]), .Z(creg_next[464]) );
  AND U7090 ( .A(n3090), .B(n6066), .Z(n6065) );
  XNOR U7091 ( .A(c[464]), .B(n6067), .Z(n6066) );
  IV U7092 ( .A(o[464]), .Z(n6067) );
  XNOR U7093 ( .A(n6068), .B(n6069), .Z(o[464]) );
  XOR U7094 ( .A(n6070), .B(o[463]), .Z(creg_next[463]) );
  AND U7095 ( .A(n3090), .B(n6071), .Z(n6070) );
  XNOR U7096 ( .A(c[463]), .B(n6072), .Z(n6071) );
  IV U7097 ( .A(o[463]), .Z(n6072) );
  XNOR U7098 ( .A(n6073), .B(n6074), .Z(o[463]) );
  XOR U7099 ( .A(n6075), .B(o[462]), .Z(creg_next[462]) );
  AND U7100 ( .A(n3090), .B(n6076), .Z(n6075) );
  XNOR U7101 ( .A(c[462]), .B(n6077), .Z(n6076) );
  IV U7102 ( .A(o[462]), .Z(n6077) );
  XNOR U7103 ( .A(n6078), .B(n6079), .Z(o[462]) );
  XOR U7104 ( .A(n6080), .B(o[461]), .Z(creg_next[461]) );
  AND U7105 ( .A(n3090), .B(n6081), .Z(n6080) );
  XNOR U7106 ( .A(c[461]), .B(n6082), .Z(n6081) );
  IV U7107 ( .A(o[461]), .Z(n6082) );
  XNOR U7108 ( .A(n6083), .B(n6084), .Z(o[461]) );
  XOR U7109 ( .A(n6085), .B(o[460]), .Z(creg_next[460]) );
  AND U7110 ( .A(n3090), .B(n6086), .Z(n6085) );
  XNOR U7111 ( .A(c[460]), .B(n6087), .Z(n6086) );
  IV U7112 ( .A(o[460]), .Z(n6087) );
  XNOR U7113 ( .A(n6088), .B(n6089), .Z(o[460]) );
  XOR U7114 ( .A(n6090), .B(o[45]), .Z(creg_next[45]) );
  AND U7115 ( .A(n3090), .B(n6091), .Z(n6090) );
  XNOR U7116 ( .A(c[45]), .B(n6092), .Z(n6091) );
  IV U7117 ( .A(o[45]), .Z(n6092) );
  XNOR U7118 ( .A(n6093), .B(n6094), .Z(o[45]) );
  XOR U7119 ( .A(n6095), .B(o[459]), .Z(creg_next[459]) );
  AND U7120 ( .A(n3090), .B(n6096), .Z(n6095) );
  XNOR U7121 ( .A(c[459]), .B(n6097), .Z(n6096) );
  IV U7122 ( .A(o[459]), .Z(n6097) );
  XNOR U7123 ( .A(n6098), .B(n6099), .Z(o[459]) );
  XOR U7124 ( .A(n6100), .B(o[458]), .Z(creg_next[458]) );
  AND U7125 ( .A(n3090), .B(n6101), .Z(n6100) );
  XNOR U7126 ( .A(c[458]), .B(n6102), .Z(n6101) );
  IV U7127 ( .A(o[458]), .Z(n6102) );
  XNOR U7128 ( .A(n6103), .B(n6104), .Z(o[458]) );
  XOR U7129 ( .A(n6105), .B(o[457]), .Z(creg_next[457]) );
  AND U7130 ( .A(n3090), .B(n6106), .Z(n6105) );
  XNOR U7131 ( .A(c[457]), .B(n6107), .Z(n6106) );
  IV U7132 ( .A(o[457]), .Z(n6107) );
  XNOR U7133 ( .A(n6108), .B(n6109), .Z(o[457]) );
  XOR U7134 ( .A(n6110), .B(o[456]), .Z(creg_next[456]) );
  AND U7135 ( .A(n3090), .B(n6111), .Z(n6110) );
  XNOR U7136 ( .A(c[456]), .B(n6112), .Z(n6111) );
  IV U7137 ( .A(o[456]), .Z(n6112) );
  XNOR U7138 ( .A(n6113), .B(n6114), .Z(o[456]) );
  XOR U7139 ( .A(n6115), .B(o[455]), .Z(creg_next[455]) );
  AND U7140 ( .A(n3090), .B(n6116), .Z(n6115) );
  XNOR U7141 ( .A(c[455]), .B(n6117), .Z(n6116) );
  IV U7142 ( .A(o[455]), .Z(n6117) );
  XNOR U7143 ( .A(n6118), .B(n6119), .Z(o[455]) );
  XOR U7144 ( .A(n6120), .B(o[454]), .Z(creg_next[454]) );
  AND U7145 ( .A(n3090), .B(n6121), .Z(n6120) );
  XNOR U7146 ( .A(c[454]), .B(n6122), .Z(n6121) );
  IV U7147 ( .A(o[454]), .Z(n6122) );
  XNOR U7148 ( .A(n6123), .B(n6124), .Z(o[454]) );
  XOR U7149 ( .A(n6125), .B(o[453]), .Z(creg_next[453]) );
  AND U7150 ( .A(n3090), .B(n6126), .Z(n6125) );
  XNOR U7151 ( .A(c[453]), .B(n6127), .Z(n6126) );
  IV U7152 ( .A(o[453]), .Z(n6127) );
  XNOR U7153 ( .A(n6128), .B(n6129), .Z(o[453]) );
  XOR U7154 ( .A(n6130), .B(o[452]), .Z(creg_next[452]) );
  AND U7155 ( .A(n3090), .B(n6131), .Z(n6130) );
  XNOR U7156 ( .A(c[452]), .B(n6132), .Z(n6131) );
  IV U7157 ( .A(o[452]), .Z(n6132) );
  XNOR U7158 ( .A(n6133), .B(n6134), .Z(o[452]) );
  XOR U7159 ( .A(n6135), .B(o[451]), .Z(creg_next[451]) );
  AND U7160 ( .A(n3090), .B(n6136), .Z(n6135) );
  XNOR U7161 ( .A(c[451]), .B(n6137), .Z(n6136) );
  IV U7162 ( .A(o[451]), .Z(n6137) );
  XNOR U7163 ( .A(n6138), .B(n6139), .Z(o[451]) );
  XOR U7164 ( .A(n6140), .B(o[450]), .Z(creg_next[450]) );
  AND U7165 ( .A(n3090), .B(n6141), .Z(n6140) );
  XNOR U7166 ( .A(c[450]), .B(n6142), .Z(n6141) );
  IV U7167 ( .A(o[450]), .Z(n6142) );
  XNOR U7168 ( .A(n6143), .B(n6144), .Z(o[450]) );
  XOR U7169 ( .A(n6145), .B(o[44]), .Z(creg_next[44]) );
  AND U7170 ( .A(n3090), .B(n6146), .Z(n6145) );
  XNOR U7171 ( .A(c[44]), .B(n6147), .Z(n6146) );
  IV U7172 ( .A(o[44]), .Z(n6147) );
  XNOR U7173 ( .A(n6148), .B(n6149), .Z(o[44]) );
  XOR U7174 ( .A(n6150), .B(o[449]), .Z(creg_next[449]) );
  AND U7175 ( .A(n3090), .B(n6151), .Z(n6150) );
  XNOR U7176 ( .A(c[449]), .B(n6152), .Z(n6151) );
  IV U7177 ( .A(o[449]), .Z(n6152) );
  XNOR U7178 ( .A(n6153), .B(n6154), .Z(o[449]) );
  XOR U7179 ( .A(n6155), .B(o[448]), .Z(creg_next[448]) );
  AND U7180 ( .A(n3090), .B(n6156), .Z(n6155) );
  XNOR U7181 ( .A(c[448]), .B(n6157), .Z(n6156) );
  IV U7182 ( .A(o[448]), .Z(n6157) );
  XNOR U7183 ( .A(n6158), .B(n6159), .Z(o[448]) );
  XOR U7184 ( .A(n6160), .B(o[447]), .Z(creg_next[447]) );
  AND U7185 ( .A(n3090), .B(n6161), .Z(n6160) );
  XNOR U7186 ( .A(c[447]), .B(n6162), .Z(n6161) );
  IV U7187 ( .A(o[447]), .Z(n6162) );
  XNOR U7188 ( .A(n6163), .B(n6164), .Z(o[447]) );
  XOR U7189 ( .A(n6165), .B(o[446]), .Z(creg_next[446]) );
  AND U7190 ( .A(n3090), .B(n6166), .Z(n6165) );
  XNOR U7191 ( .A(c[446]), .B(n6167), .Z(n6166) );
  IV U7192 ( .A(o[446]), .Z(n6167) );
  XNOR U7193 ( .A(n6168), .B(n6169), .Z(o[446]) );
  XOR U7194 ( .A(n6170), .B(o[445]), .Z(creg_next[445]) );
  AND U7195 ( .A(n3090), .B(n6171), .Z(n6170) );
  XNOR U7196 ( .A(c[445]), .B(n6172), .Z(n6171) );
  IV U7197 ( .A(o[445]), .Z(n6172) );
  XNOR U7198 ( .A(n6173), .B(n6174), .Z(o[445]) );
  XOR U7199 ( .A(n6175), .B(o[444]), .Z(creg_next[444]) );
  AND U7200 ( .A(n3090), .B(n6176), .Z(n6175) );
  XNOR U7201 ( .A(c[444]), .B(n6177), .Z(n6176) );
  IV U7202 ( .A(o[444]), .Z(n6177) );
  XNOR U7203 ( .A(n6178), .B(n6179), .Z(o[444]) );
  XOR U7204 ( .A(n6180), .B(o[443]), .Z(creg_next[443]) );
  AND U7205 ( .A(n3090), .B(n6181), .Z(n6180) );
  XNOR U7206 ( .A(c[443]), .B(n6182), .Z(n6181) );
  IV U7207 ( .A(o[443]), .Z(n6182) );
  XNOR U7208 ( .A(n6183), .B(n6184), .Z(o[443]) );
  XOR U7209 ( .A(n6185), .B(o[442]), .Z(creg_next[442]) );
  AND U7210 ( .A(n3090), .B(n6186), .Z(n6185) );
  XNOR U7211 ( .A(c[442]), .B(n6187), .Z(n6186) );
  IV U7212 ( .A(o[442]), .Z(n6187) );
  XNOR U7213 ( .A(n6188), .B(n6189), .Z(o[442]) );
  XOR U7214 ( .A(n6190), .B(o[441]), .Z(creg_next[441]) );
  AND U7215 ( .A(n3090), .B(n6191), .Z(n6190) );
  XNOR U7216 ( .A(c[441]), .B(n6192), .Z(n6191) );
  IV U7217 ( .A(o[441]), .Z(n6192) );
  XNOR U7218 ( .A(n6193), .B(n6194), .Z(o[441]) );
  XOR U7219 ( .A(n6195), .B(o[440]), .Z(creg_next[440]) );
  AND U7220 ( .A(n3090), .B(n6196), .Z(n6195) );
  XNOR U7221 ( .A(c[440]), .B(n6197), .Z(n6196) );
  IV U7222 ( .A(o[440]), .Z(n6197) );
  XNOR U7223 ( .A(n6198), .B(n6199), .Z(o[440]) );
  XOR U7224 ( .A(n6200), .B(o[43]), .Z(creg_next[43]) );
  AND U7225 ( .A(n3090), .B(n6201), .Z(n6200) );
  XNOR U7226 ( .A(c[43]), .B(n6202), .Z(n6201) );
  IV U7227 ( .A(o[43]), .Z(n6202) );
  XNOR U7228 ( .A(n6203), .B(n6204), .Z(o[43]) );
  XOR U7229 ( .A(n6205), .B(o[439]), .Z(creg_next[439]) );
  AND U7230 ( .A(n3090), .B(n6206), .Z(n6205) );
  XNOR U7231 ( .A(c[439]), .B(n6207), .Z(n6206) );
  IV U7232 ( .A(o[439]), .Z(n6207) );
  XNOR U7233 ( .A(n6208), .B(n6209), .Z(o[439]) );
  XOR U7234 ( .A(n6210), .B(o[438]), .Z(creg_next[438]) );
  AND U7235 ( .A(n3090), .B(n6211), .Z(n6210) );
  XNOR U7236 ( .A(c[438]), .B(n6212), .Z(n6211) );
  IV U7237 ( .A(o[438]), .Z(n6212) );
  XNOR U7238 ( .A(n6213), .B(n6214), .Z(o[438]) );
  XOR U7239 ( .A(n6215), .B(o[437]), .Z(creg_next[437]) );
  AND U7240 ( .A(n3090), .B(n6216), .Z(n6215) );
  XNOR U7241 ( .A(c[437]), .B(n6217), .Z(n6216) );
  IV U7242 ( .A(o[437]), .Z(n6217) );
  XNOR U7243 ( .A(n6218), .B(n6219), .Z(o[437]) );
  XOR U7244 ( .A(n6220), .B(o[436]), .Z(creg_next[436]) );
  AND U7245 ( .A(n3090), .B(n6221), .Z(n6220) );
  XNOR U7246 ( .A(c[436]), .B(n6222), .Z(n6221) );
  IV U7247 ( .A(o[436]), .Z(n6222) );
  XNOR U7248 ( .A(n6223), .B(n6224), .Z(o[436]) );
  XOR U7249 ( .A(n6225), .B(o[435]), .Z(creg_next[435]) );
  AND U7250 ( .A(n3090), .B(n6226), .Z(n6225) );
  XNOR U7251 ( .A(c[435]), .B(n6227), .Z(n6226) );
  IV U7252 ( .A(o[435]), .Z(n6227) );
  XNOR U7253 ( .A(n6228), .B(n6229), .Z(o[435]) );
  XOR U7254 ( .A(n6230), .B(o[434]), .Z(creg_next[434]) );
  AND U7255 ( .A(n3090), .B(n6231), .Z(n6230) );
  XNOR U7256 ( .A(c[434]), .B(n6232), .Z(n6231) );
  IV U7257 ( .A(o[434]), .Z(n6232) );
  XNOR U7258 ( .A(n6233), .B(n6234), .Z(o[434]) );
  XOR U7259 ( .A(n6235), .B(o[433]), .Z(creg_next[433]) );
  AND U7260 ( .A(n3090), .B(n6236), .Z(n6235) );
  XNOR U7261 ( .A(c[433]), .B(n6237), .Z(n6236) );
  IV U7262 ( .A(o[433]), .Z(n6237) );
  XNOR U7263 ( .A(n6238), .B(n6239), .Z(o[433]) );
  XOR U7264 ( .A(n6240), .B(o[432]), .Z(creg_next[432]) );
  AND U7265 ( .A(n3090), .B(n6241), .Z(n6240) );
  XNOR U7266 ( .A(c[432]), .B(n6242), .Z(n6241) );
  IV U7267 ( .A(o[432]), .Z(n6242) );
  XNOR U7268 ( .A(n6243), .B(n6244), .Z(o[432]) );
  XOR U7269 ( .A(n6245), .B(o[431]), .Z(creg_next[431]) );
  AND U7270 ( .A(n3090), .B(n6246), .Z(n6245) );
  XNOR U7271 ( .A(c[431]), .B(n6247), .Z(n6246) );
  IV U7272 ( .A(o[431]), .Z(n6247) );
  XNOR U7273 ( .A(n6248), .B(n6249), .Z(o[431]) );
  XOR U7274 ( .A(n6250), .B(o[430]), .Z(creg_next[430]) );
  AND U7275 ( .A(n3090), .B(n6251), .Z(n6250) );
  XNOR U7276 ( .A(c[430]), .B(n6252), .Z(n6251) );
  IV U7277 ( .A(o[430]), .Z(n6252) );
  XNOR U7278 ( .A(n6253), .B(n6254), .Z(o[430]) );
  XOR U7279 ( .A(n6255), .B(o[42]), .Z(creg_next[42]) );
  AND U7280 ( .A(n3090), .B(n6256), .Z(n6255) );
  XNOR U7281 ( .A(c[42]), .B(n6257), .Z(n6256) );
  IV U7282 ( .A(o[42]), .Z(n6257) );
  XNOR U7283 ( .A(n6258), .B(n6259), .Z(o[42]) );
  XOR U7284 ( .A(n6260), .B(o[429]), .Z(creg_next[429]) );
  AND U7285 ( .A(n3090), .B(n6261), .Z(n6260) );
  XNOR U7286 ( .A(c[429]), .B(n6262), .Z(n6261) );
  IV U7287 ( .A(o[429]), .Z(n6262) );
  XNOR U7288 ( .A(n6263), .B(n6264), .Z(o[429]) );
  XOR U7289 ( .A(n6265), .B(o[428]), .Z(creg_next[428]) );
  AND U7290 ( .A(n3090), .B(n6266), .Z(n6265) );
  XNOR U7291 ( .A(c[428]), .B(n6267), .Z(n6266) );
  IV U7292 ( .A(o[428]), .Z(n6267) );
  XNOR U7293 ( .A(n6268), .B(n6269), .Z(o[428]) );
  XOR U7294 ( .A(n6270), .B(o[427]), .Z(creg_next[427]) );
  AND U7295 ( .A(n3090), .B(n6271), .Z(n6270) );
  XNOR U7296 ( .A(c[427]), .B(n6272), .Z(n6271) );
  IV U7297 ( .A(o[427]), .Z(n6272) );
  XNOR U7298 ( .A(n6273), .B(n6274), .Z(o[427]) );
  XOR U7299 ( .A(n6275), .B(o[426]), .Z(creg_next[426]) );
  AND U7300 ( .A(n3090), .B(n6276), .Z(n6275) );
  XNOR U7301 ( .A(c[426]), .B(n6277), .Z(n6276) );
  IV U7302 ( .A(o[426]), .Z(n6277) );
  XNOR U7303 ( .A(n6278), .B(n6279), .Z(o[426]) );
  XOR U7304 ( .A(n6280), .B(o[425]), .Z(creg_next[425]) );
  AND U7305 ( .A(n3090), .B(n6281), .Z(n6280) );
  XNOR U7306 ( .A(c[425]), .B(n6282), .Z(n6281) );
  IV U7307 ( .A(o[425]), .Z(n6282) );
  XNOR U7308 ( .A(n6283), .B(n6284), .Z(o[425]) );
  XOR U7309 ( .A(n6285), .B(o[424]), .Z(creg_next[424]) );
  AND U7310 ( .A(n3090), .B(n6286), .Z(n6285) );
  XNOR U7311 ( .A(c[424]), .B(n6287), .Z(n6286) );
  IV U7312 ( .A(o[424]), .Z(n6287) );
  XNOR U7313 ( .A(n6288), .B(n6289), .Z(o[424]) );
  XOR U7314 ( .A(n6290), .B(o[423]), .Z(creg_next[423]) );
  AND U7315 ( .A(n3090), .B(n6291), .Z(n6290) );
  XNOR U7316 ( .A(c[423]), .B(n6292), .Z(n6291) );
  IV U7317 ( .A(o[423]), .Z(n6292) );
  XNOR U7318 ( .A(n6293), .B(n6294), .Z(o[423]) );
  XOR U7319 ( .A(n6295), .B(o[422]), .Z(creg_next[422]) );
  AND U7320 ( .A(n3090), .B(n6296), .Z(n6295) );
  XNOR U7321 ( .A(c[422]), .B(n6297), .Z(n6296) );
  IV U7322 ( .A(o[422]), .Z(n6297) );
  XNOR U7323 ( .A(n6298), .B(n6299), .Z(o[422]) );
  XOR U7324 ( .A(n6300), .B(o[421]), .Z(creg_next[421]) );
  AND U7325 ( .A(n3090), .B(n6301), .Z(n6300) );
  XNOR U7326 ( .A(c[421]), .B(n6302), .Z(n6301) );
  IV U7327 ( .A(o[421]), .Z(n6302) );
  XNOR U7328 ( .A(n6303), .B(n6304), .Z(o[421]) );
  XOR U7329 ( .A(n6305), .B(o[420]), .Z(creg_next[420]) );
  AND U7330 ( .A(n3090), .B(n6306), .Z(n6305) );
  XNOR U7331 ( .A(c[420]), .B(n6307), .Z(n6306) );
  IV U7332 ( .A(o[420]), .Z(n6307) );
  XNOR U7333 ( .A(n6308), .B(n6309), .Z(o[420]) );
  XOR U7334 ( .A(n6310), .B(o[41]), .Z(creg_next[41]) );
  AND U7335 ( .A(n3090), .B(n6311), .Z(n6310) );
  XNOR U7336 ( .A(c[41]), .B(n6312), .Z(n6311) );
  IV U7337 ( .A(o[41]), .Z(n6312) );
  XNOR U7338 ( .A(n6313), .B(n6314), .Z(o[41]) );
  XOR U7339 ( .A(n6315), .B(o[419]), .Z(creg_next[419]) );
  AND U7340 ( .A(n3090), .B(n6316), .Z(n6315) );
  XNOR U7341 ( .A(c[419]), .B(n6317), .Z(n6316) );
  IV U7342 ( .A(o[419]), .Z(n6317) );
  XNOR U7343 ( .A(n6318), .B(n6319), .Z(o[419]) );
  XOR U7344 ( .A(n6320), .B(o[418]), .Z(creg_next[418]) );
  AND U7345 ( .A(n3090), .B(n6321), .Z(n6320) );
  XNOR U7346 ( .A(c[418]), .B(n6322), .Z(n6321) );
  IV U7347 ( .A(o[418]), .Z(n6322) );
  XNOR U7348 ( .A(n6323), .B(n6324), .Z(o[418]) );
  XOR U7349 ( .A(n6325), .B(o[417]), .Z(creg_next[417]) );
  AND U7350 ( .A(n3090), .B(n6326), .Z(n6325) );
  XNOR U7351 ( .A(c[417]), .B(n6327), .Z(n6326) );
  IV U7352 ( .A(o[417]), .Z(n6327) );
  XNOR U7353 ( .A(n6328), .B(n6329), .Z(o[417]) );
  XOR U7354 ( .A(n6330), .B(o[416]), .Z(creg_next[416]) );
  AND U7355 ( .A(n3090), .B(n6331), .Z(n6330) );
  XNOR U7356 ( .A(c[416]), .B(n6332), .Z(n6331) );
  IV U7357 ( .A(o[416]), .Z(n6332) );
  XNOR U7358 ( .A(n6333), .B(n6334), .Z(o[416]) );
  XOR U7359 ( .A(n6335), .B(o[415]), .Z(creg_next[415]) );
  AND U7360 ( .A(n3090), .B(n6336), .Z(n6335) );
  XNOR U7361 ( .A(c[415]), .B(n6337), .Z(n6336) );
  IV U7362 ( .A(o[415]), .Z(n6337) );
  XNOR U7363 ( .A(n6338), .B(n6339), .Z(o[415]) );
  XOR U7364 ( .A(n6340), .B(o[414]), .Z(creg_next[414]) );
  AND U7365 ( .A(n3090), .B(n6341), .Z(n6340) );
  XNOR U7366 ( .A(c[414]), .B(n6342), .Z(n6341) );
  IV U7367 ( .A(o[414]), .Z(n6342) );
  XNOR U7368 ( .A(n6343), .B(n6344), .Z(o[414]) );
  XOR U7369 ( .A(n6345), .B(o[413]), .Z(creg_next[413]) );
  AND U7370 ( .A(n3090), .B(n6346), .Z(n6345) );
  XNOR U7371 ( .A(c[413]), .B(n6347), .Z(n6346) );
  IV U7372 ( .A(o[413]), .Z(n6347) );
  XNOR U7373 ( .A(n6348), .B(n6349), .Z(o[413]) );
  XOR U7374 ( .A(n6350), .B(o[412]), .Z(creg_next[412]) );
  AND U7375 ( .A(n3090), .B(n6351), .Z(n6350) );
  XNOR U7376 ( .A(c[412]), .B(n6352), .Z(n6351) );
  IV U7377 ( .A(o[412]), .Z(n6352) );
  XNOR U7378 ( .A(n6353), .B(n6354), .Z(o[412]) );
  XOR U7379 ( .A(n6355), .B(o[411]), .Z(creg_next[411]) );
  AND U7380 ( .A(n3090), .B(n6356), .Z(n6355) );
  XNOR U7381 ( .A(c[411]), .B(n6357), .Z(n6356) );
  IV U7382 ( .A(o[411]), .Z(n6357) );
  XNOR U7383 ( .A(n6358), .B(n6359), .Z(o[411]) );
  XOR U7384 ( .A(n6360), .B(o[410]), .Z(creg_next[410]) );
  AND U7385 ( .A(n3090), .B(n6361), .Z(n6360) );
  XNOR U7386 ( .A(c[410]), .B(n6362), .Z(n6361) );
  IV U7387 ( .A(o[410]), .Z(n6362) );
  XNOR U7388 ( .A(n6363), .B(n6364), .Z(o[410]) );
  XOR U7389 ( .A(n6365), .B(o[40]), .Z(creg_next[40]) );
  AND U7390 ( .A(n3090), .B(n6366), .Z(n6365) );
  XNOR U7391 ( .A(c[40]), .B(n6367), .Z(n6366) );
  IV U7392 ( .A(o[40]), .Z(n6367) );
  XNOR U7393 ( .A(n6368), .B(n6369), .Z(o[40]) );
  XOR U7394 ( .A(n6370), .B(o[409]), .Z(creg_next[409]) );
  AND U7395 ( .A(n3090), .B(n6371), .Z(n6370) );
  XNOR U7396 ( .A(c[409]), .B(n6372), .Z(n6371) );
  IV U7397 ( .A(o[409]), .Z(n6372) );
  XNOR U7398 ( .A(n6373), .B(n6374), .Z(o[409]) );
  XOR U7399 ( .A(n6375), .B(o[408]), .Z(creg_next[408]) );
  AND U7400 ( .A(n3090), .B(n6376), .Z(n6375) );
  XNOR U7401 ( .A(c[408]), .B(n6377), .Z(n6376) );
  IV U7402 ( .A(o[408]), .Z(n6377) );
  XNOR U7403 ( .A(n6378), .B(n6379), .Z(o[408]) );
  XOR U7404 ( .A(n6380), .B(o[407]), .Z(creg_next[407]) );
  AND U7405 ( .A(n3090), .B(n6381), .Z(n6380) );
  XNOR U7406 ( .A(c[407]), .B(n6382), .Z(n6381) );
  IV U7407 ( .A(o[407]), .Z(n6382) );
  XNOR U7408 ( .A(n6383), .B(n6384), .Z(o[407]) );
  XOR U7409 ( .A(n6385), .B(o[406]), .Z(creg_next[406]) );
  AND U7410 ( .A(n3090), .B(n6386), .Z(n6385) );
  XNOR U7411 ( .A(c[406]), .B(n6387), .Z(n6386) );
  IV U7412 ( .A(o[406]), .Z(n6387) );
  XNOR U7413 ( .A(n6388), .B(n6389), .Z(o[406]) );
  XOR U7414 ( .A(n6390), .B(o[405]), .Z(creg_next[405]) );
  AND U7415 ( .A(n3090), .B(n6391), .Z(n6390) );
  XNOR U7416 ( .A(c[405]), .B(n6392), .Z(n6391) );
  IV U7417 ( .A(o[405]), .Z(n6392) );
  XNOR U7418 ( .A(n6393), .B(n6394), .Z(o[405]) );
  XOR U7419 ( .A(n6395), .B(o[404]), .Z(creg_next[404]) );
  AND U7420 ( .A(n3090), .B(n6396), .Z(n6395) );
  XNOR U7421 ( .A(c[404]), .B(n6397), .Z(n6396) );
  IV U7422 ( .A(o[404]), .Z(n6397) );
  XNOR U7423 ( .A(n6398), .B(n6399), .Z(o[404]) );
  XOR U7424 ( .A(n6400), .B(o[403]), .Z(creg_next[403]) );
  AND U7425 ( .A(n3090), .B(n6401), .Z(n6400) );
  XNOR U7426 ( .A(c[403]), .B(n6402), .Z(n6401) );
  IV U7427 ( .A(o[403]), .Z(n6402) );
  XNOR U7428 ( .A(n6403), .B(n6404), .Z(o[403]) );
  XOR U7429 ( .A(n6405), .B(o[402]), .Z(creg_next[402]) );
  AND U7430 ( .A(n3090), .B(n6406), .Z(n6405) );
  XNOR U7431 ( .A(c[402]), .B(n6407), .Z(n6406) );
  IV U7432 ( .A(o[402]), .Z(n6407) );
  XNOR U7433 ( .A(n6408), .B(n6409), .Z(o[402]) );
  XOR U7434 ( .A(n6410), .B(o[401]), .Z(creg_next[401]) );
  AND U7435 ( .A(n3090), .B(n6411), .Z(n6410) );
  XNOR U7436 ( .A(c[401]), .B(n6412), .Z(n6411) );
  IV U7437 ( .A(o[401]), .Z(n6412) );
  XNOR U7438 ( .A(n6413), .B(n6414), .Z(o[401]) );
  XOR U7439 ( .A(n6415), .B(o[400]), .Z(creg_next[400]) );
  AND U7440 ( .A(n3090), .B(n6416), .Z(n6415) );
  XNOR U7441 ( .A(c[400]), .B(n6417), .Z(n6416) );
  IV U7442 ( .A(o[400]), .Z(n6417) );
  XNOR U7443 ( .A(n6418), .B(n6419), .Z(o[400]) );
  XOR U7444 ( .A(n6420), .B(o[3]), .Z(creg_next[3]) );
  AND U7445 ( .A(n3090), .B(n6421), .Z(n6420) );
  XNOR U7446 ( .A(c[3]), .B(n6422), .Z(n6421) );
  IV U7447 ( .A(o[3]), .Z(n6422) );
  XNOR U7448 ( .A(n6423), .B(n6424), .Z(o[3]) );
  XOR U7449 ( .A(n6425), .B(o[39]), .Z(creg_next[39]) );
  AND U7450 ( .A(n3090), .B(n6426), .Z(n6425) );
  XNOR U7451 ( .A(c[39]), .B(n6427), .Z(n6426) );
  IV U7452 ( .A(o[39]), .Z(n6427) );
  XNOR U7453 ( .A(n6428), .B(n6429), .Z(o[39]) );
  XOR U7454 ( .A(n6430), .B(o[399]), .Z(creg_next[399]) );
  AND U7455 ( .A(n3090), .B(n6431), .Z(n6430) );
  XNOR U7456 ( .A(c[399]), .B(n6432), .Z(n6431) );
  IV U7457 ( .A(o[399]), .Z(n6432) );
  XNOR U7458 ( .A(n6433), .B(n6434), .Z(o[399]) );
  XOR U7459 ( .A(n6435), .B(o[398]), .Z(creg_next[398]) );
  AND U7460 ( .A(n3090), .B(n6436), .Z(n6435) );
  XNOR U7461 ( .A(c[398]), .B(n6437), .Z(n6436) );
  IV U7462 ( .A(o[398]), .Z(n6437) );
  XNOR U7463 ( .A(n6438), .B(n6439), .Z(o[398]) );
  XOR U7464 ( .A(n6440), .B(o[397]), .Z(creg_next[397]) );
  AND U7465 ( .A(n3090), .B(n6441), .Z(n6440) );
  XNOR U7466 ( .A(c[397]), .B(n6442), .Z(n6441) );
  IV U7467 ( .A(o[397]), .Z(n6442) );
  XNOR U7468 ( .A(n6443), .B(n6444), .Z(o[397]) );
  XOR U7469 ( .A(n6445), .B(o[396]), .Z(creg_next[396]) );
  AND U7470 ( .A(n3090), .B(n6446), .Z(n6445) );
  XNOR U7471 ( .A(c[396]), .B(n6447), .Z(n6446) );
  IV U7472 ( .A(o[396]), .Z(n6447) );
  XNOR U7473 ( .A(n6448), .B(n6449), .Z(o[396]) );
  XOR U7474 ( .A(n6450), .B(o[395]), .Z(creg_next[395]) );
  AND U7475 ( .A(n3090), .B(n6451), .Z(n6450) );
  XNOR U7476 ( .A(c[395]), .B(n6452), .Z(n6451) );
  IV U7477 ( .A(o[395]), .Z(n6452) );
  XNOR U7478 ( .A(n6453), .B(n6454), .Z(o[395]) );
  XOR U7479 ( .A(n6455), .B(o[394]), .Z(creg_next[394]) );
  AND U7480 ( .A(n3090), .B(n6456), .Z(n6455) );
  XNOR U7481 ( .A(c[394]), .B(n6457), .Z(n6456) );
  IV U7482 ( .A(o[394]), .Z(n6457) );
  XNOR U7483 ( .A(n6458), .B(n6459), .Z(o[394]) );
  XOR U7484 ( .A(n6460), .B(o[393]), .Z(creg_next[393]) );
  AND U7485 ( .A(n3090), .B(n6461), .Z(n6460) );
  XNOR U7486 ( .A(c[393]), .B(n6462), .Z(n6461) );
  IV U7487 ( .A(o[393]), .Z(n6462) );
  XNOR U7488 ( .A(n6463), .B(n6464), .Z(o[393]) );
  XOR U7489 ( .A(n6465), .B(o[392]), .Z(creg_next[392]) );
  AND U7490 ( .A(n3090), .B(n6466), .Z(n6465) );
  XNOR U7491 ( .A(c[392]), .B(n6467), .Z(n6466) );
  IV U7492 ( .A(o[392]), .Z(n6467) );
  XNOR U7493 ( .A(n6468), .B(n6469), .Z(o[392]) );
  XOR U7494 ( .A(n6470), .B(o[391]), .Z(creg_next[391]) );
  AND U7495 ( .A(n3090), .B(n6471), .Z(n6470) );
  XNOR U7496 ( .A(c[391]), .B(n6472), .Z(n6471) );
  IV U7497 ( .A(o[391]), .Z(n6472) );
  XNOR U7498 ( .A(n6473), .B(n6474), .Z(o[391]) );
  XOR U7499 ( .A(n6475), .B(o[390]), .Z(creg_next[390]) );
  AND U7500 ( .A(n3090), .B(n6476), .Z(n6475) );
  XNOR U7501 ( .A(c[390]), .B(n6477), .Z(n6476) );
  IV U7502 ( .A(o[390]), .Z(n6477) );
  XNOR U7503 ( .A(n6478), .B(n6479), .Z(o[390]) );
  XOR U7504 ( .A(n6480), .B(o[38]), .Z(creg_next[38]) );
  AND U7505 ( .A(n3090), .B(n6481), .Z(n6480) );
  XNOR U7506 ( .A(c[38]), .B(n6482), .Z(n6481) );
  IV U7507 ( .A(o[38]), .Z(n6482) );
  XNOR U7508 ( .A(n6483), .B(n6484), .Z(o[38]) );
  XOR U7509 ( .A(n6485), .B(o[389]), .Z(creg_next[389]) );
  AND U7510 ( .A(n3090), .B(n6486), .Z(n6485) );
  XNOR U7511 ( .A(c[389]), .B(n6487), .Z(n6486) );
  IV U7512 ( .A(o[389]), .Z(n6487) );
  XNOR U7513 ( .A(n6488), .B(n6489), .Z(o[389]) );
  XOR U7514 ( .A(n6490), .B(o[388]), .Z(creg_next[388]) );
  AND U7515 ( .A(n3090), .B(n6491), .Z(n6490) );
  XNOR U7516 ( .A(c[388]), .B(n6492), .Z(n6491) );
  IV U7517 ( .A(o[388]), .Z(n6492) );
  XNOR U7518 ( .A(n6493), .B(n6494), .Z(o[388]) );
  XOR U7519 ( .A(n6495), .B(o[387]), .Z(creg_next[387]) );
  AND U7520 ( .A(n3090), .B(n6496), .Z(n6495) );
  XNOR U7521 ( .A(c[387]), .B(n6497), .Z(n6496) );
  IV U7522 ( .A(o[387]), .Z(n6497) );
  XNOR U7523 ( .A(n6498), .B(n6499), .Z(o[387]) );
  XOR U7524 ( .A(n6500), .B(o[386]), .Z(creg_next[386]) );
  AND U7525 ( .A(n3090), .B(n6501), .Z(n6500) );
  XNOR U7526 ( .A(c[386]), .B(n6502), .Z(n6501) );
  IV U7527 ( .A(o[386]), .Z(n6502) );
  XNOR U7528 ( .A(n6503), .B(n6504), .Z(o[386]) );
  XOR U7529 ( .A(n6505), .B(o[385]), .Z(creg_next[385]) );
  AND U7530 ( .A(n3090), .B(n6506), .Z(n6505) );
  XNOR U7531 ( .A(c[385]), .B(n6507), .Z(n6506) );
  IV U7532 ( .A(o[385]), .Z(n6507) );
  XNOR U7533 ( .A(n6508), .B(n6509), .Z(o[385]) );
  XOR U7534 ( .A(n6510), .B(o[384]), .Z(creg_next[384]) );
  AND U7535 ( .A(n3090), .B(n6511), .Z(n6510) );
  XNOR U7536 ( .A(c[384]), .B(n6512), .Z(n6511) );
  IV U7537 ( .A(o[384]), .Z(n6512) );
  XNOR U7538 ( .A(n6513), .B(n6514), .Z(o[384]) );
  XOR U7539 ( .A(n6515), .B(o[383]), .Z(creg_next[383]) );
  AND U7540 ( .A(n3090), .B(n6516), .Z(n6515) );
  XNOR U7541 ( .A(c[383]), .B(n6517), .Z(n6516) );
  IV U7542 ( .A(o[383]), .Z(n6517) );
  XNOR U7543 ( .A(n6518), .B(n6519), .Z(o[383]) );
  XOR U7544 ( .A(n6520), .B(o[382]), .Z(creg_next[382]) );
  AND U7545 ( .A(n3090), .B(n6521), .Z(n6520) );
  XNOR U7546 ( .A(c[382]), .B(n6522), .Z(n6521) );
  IV U7547 ( .A(o[382]), .Z(n6522) );
  XNOR U7548 ( .A(n6523), .B(n6524), .Z(o[382]) );
  XOR U7549 ( .A(n6525), .B(o[381]), .Z(creg_next[381]) );
  AND U7550 ( .A(n3090), .B(n6526), .Z(n6525) );
  XNOR U7551 ( .A(c[381]), .B(n6527), .Z(n6526) );
  IV U7552 ( .A(o[381]), .Z(n6527) );
  XNOR U7553 ( .A(n6528), .B(n6529), .Z(o[381]) );
  XOR U7554 ( .A(n6530), .B(o[380]), .Z(creg_next[380]) );
  AND U7555 ( .A(n3090), .B(n6531), .Z(n6530) );
  XNOR U7556 ( .A(c[380]), .B(n6532), .Z(n6531) );
  IV U7557 ( .A(o[380]), .Z(n6532) );
  XNOR U7558 ( .A(n6533), .B(n6534), .Z(o[380]) );
  XOR U7559 ( .A(n6535), .B(o[37]), .Z(creg_next[37]) );
  AND U7560 ( .A(n3090), .B(n6536), .Z(n6535) );
  XNOR U7561 ( .A(c[37]), .B(n6537), .Z(n6536) );
  IV U7562 ( .A(o[37]), .Z(n6537) );
  XNOR U7563 ( .A(n6538), .B(n6539), .Z(o[37]) );
  XOR U7564 ( .A(n6540), .B(o[379]), .Z(creg_next[379]) );
  AND U7565 ( .A(n3090), .B(n6541), .Z(n6540) );
  XNOR U7566 ( .A(c[379]), .B(n6542), .Z(n6541) );
  IV U7567 ( .A(o[379]), .Z(n6542) );
  XNOR U7568 ( .A(n6543), .B(n6544), .Z(o[379]) );
  XOR U7569 ( .A(n6545), .B(o[378]), .Z(creg_next[378]) );
  AND U7570 ( .A(n3090), .B(n6546), .Z(n6545) );
  XNOR U7571 ( .A(c[378]), .B(n6547), .Z(n6546) );
  IV U7572 ( .A(o[378]), .Z(n6547) );
  XNOR U7573 ( .A(n6548), .B(n6549), .Z(o[378]) );
  XOR U7574 ( .A(n6550), .B(o[377]), .Z(creg_next[377]) );
  AND U7575 ( .A(n3090), .B(n6551), .Z(n6550) );
  XNOR U7576 ( .A(c[377]), .B(n6552), .Z(n6551) );
  IV U7577 ( .A(o[377]), .Z(n6552) );
  XNOR U7578 ( .A(n6553), .B(n6554), .Z(o[377]) );
  XOR U7579 ( .A(n6555), .B(o[376]), .Z(creg_next[376]) );
  AND U7580 ( .A(n3090), .B(n6556), .Z(n6555) );
  XNOR U7581 ( .A(c[376]), .B(n6557), .Z(n6556) );
  IV U7582 ( .A(o[376]), .Z(n6557) );
  XNOR U7583 ( .A(n6558), .B(n6559), .Z(o[376]) );
  XOR U7584 ( .A(n6560), .B(o[375]), .Z(creg_next[375]) );
  AND U7585 ( .A(n3090), .B(n6561), .Z(n6560) );
  XNOR U7586 ( .A(c[375]), .B(n6562), .Z(n6561) );
  IV U7587 ( .A(o[375]), .Z(n6562) );
  XNOR U7588 ( .A(n6563), .B(n6564), .Z(o[375]) );
  XOR U7589 ( .A(n6565), .B(o[374]), .Z(creg_next[374]) );
  AND U7590 ( .A(n3090), .B(n6566), .Z(n6565) );
  XNOR U7591 ( .A(c[374]), .B(n6567), .Z(n6566) );
  IV U7592 ( .A(o[374]), .Z(n6567) );
  XNOR U7593 ( .A(n6568), .B(n6569), .Z(o[374]) );
  XOR U7594 ( .A(n6570), .B(o[373]), .Z(creg_next[373]) );
  AND U7595 ( .A(n3090), .B(n6571), .Z(n6570) );
  XNOR U7596 ( .A(c[373]), .B(n6572), .Z(n6571) );
  IV U7597 ( .A(o[373]), .Z(n6572) );
  XNOR U7598 ( .A(n6573), .B(n6574), .Z(o[373]) );
  XOR U7599 ( .A(n6575), .B(o[372]), .Z(creg_next[372]) );
  AND U7600 ( .A(n3090), .B(n6576), .Z(n6575) );
  XNOR U7601 ( .A(c[372]), .B(n6577), .Z(n6576) );
  IV U7602 ( .A(o[372]), .Z(n6577) );
  XNOR U7603 ( .A(n6578), .B(n6579), .Z(o[372]) );
  XOR U7604 ( .A(n6580), .B(o[371]), .Z(creg_next[371]) );
  AND U7605 ( .A(n3090), .B(n6581), .Z(n6580) );
  XNOR U7606 ( .A(c[371]), .B(n6582), .Z(n6581) );
  IV U7607 ( .A(o[371]), .Z(n6582) );
  XNOR U7608 ( .A(n6583), .B(n6584), .Z(o[371]) );
  XOR U7609 ( .A(n6585), .B(o[370]), .Z(creg_next[370]) );
  AND U7610 ( .A(n3090), .B(n6586), .Z(n6585) );
  XNOR U7611 ( .A(c[370]), .B(n6587), .Z(n6586) );
  IV U7612 ( .A(o[370]), .Z(n6587) );
  XNOR U7613 ( .A(n6588), .B(n6589), .Z(o[370]) );
  XOR U7614 ( .A(n6590), .B(o[36]), .Z(creg_next[36]) );
  AND U7615 ( .A(n3090), .B(n6591), .Z(n6590) );
  XNOR U7616 ( .A(c[36]), .B(n6592), .Z(n6591) );
  IV U7617 ( .A(o[36]), .Z(n6592) );
  XNOR U7618 ( .A(n6593), .B(n6594), .Z(o[36]) );
  XOR U7619 ( .A(n6595), .B(o[369]), .Z(creg_next[369]) );
  AND U7620 ( .A(n3090), .B(n6596), .Z(n6595) );
  XNOR U7621 ( .A(c[369]), .B(n6597), .Z(n6596) );
  IV U7622 ( .A(o[369]), .Z(n6597) );
  XNOR U7623 ( .A(n6598), .B(n6599), .Z(o[369]) );
  XOR U7624 ( .A(n6600), .B(o[368]), .Z(creg_next[368]) );
  AND U7625 ( .A(n3090), .B(n6601), .Z(n6600) );
  XNOR U7626 ( .A(c[368]), .B(n6602), .Z(n6601) );
  IV U7627 ( .A(o[368]), .Z(n6602) );
  XNOR U7628 ( .A(n6603), .B(n6604), .Z(o[368]) );
  XOR U7629 ( .A(n6605), .B(o[367]), .Z(creg_next[367]) );
  AND U7630 ( .A(n3090), .B(n6606), .Z(n6605) );
  XNOR U7631 ( .A(c[367]), .B(n6607), .Z(n6606) );
  IV U7632 ( .A(o[367]), .Z(n6607) );
  XNOR U7633 ( .A(n6608), .B(n6609), .Z(o[367]) );
  XOR U7634 ( .A(n6610), .B(o[366]), .Z(creg_next[366]) );
  AND U7635 ( .A(n3090), .B(n6611), .Z(n6610) );
  XNOR U7636 ( .A(c[366]), .B(n6612), .Z(n6611) );
  IV U7637 ( .A(o[366]), .Z(n6612) );
  XNOR U7638 ( .A(n6613), .B(n6614), .Z(o[366]) );
  XOR U7639 ( .A(n6615), .B(o[365]), .Z(creg_next[365]) );
  AND U7640 ( .A(n3090), .B(n6616), .Z(n6615) );
  XNOR U7641 ( .A(c[365]), .B(n6617), .Z(n6616) );
  IV U7642 ( .A(o[365]), .Z(n6617) );
  XNOR U7643 ( .A(n6618), .B(n6619), .Z(o[365]) );
  XOR U7644 ( .A(n6620), .B(o[364]), .Z(creg_next[364]) );
  AND U7645 ( .A(n3090), .B(n6621), .Z(n6620) );
  XNOR U7646 ( .A(c[364]), .B(n6622), .Z(n6621) );
  IV U7647 ( .A(o[364]), .Z(n6622) );
  XNOR U7648 ( .A(n6623), .B(n6624), .Z(o[364]) );
  XOR U7649 ( .A(n6625), .B(o[363]), .Z(creg_next[363]) );
  AND U7650 ( .A(n3090), .B(n6626), .Z(n6625) );
  XNOR U7651 ( .A(c[363]), .B(n6627), .Z(n6626) );
  IV U7652 ( .A(o[363]), .Z(n6627) );
  XNOR U7653 ( .A(n6628), .B(n6629), .Z(o[363]) );
  XOR U7654 ( .A(n6630), .B(o[362]), .Z(creg_next[362]) );
  AND U7655 ( .A(n3090), .B(n6631), .Z(n6630) );
  XNOR U7656 ( .A(c[362]), .B(n6632), .Z(n6631) );
  IV U7657 ( .A(o[362]), .Z(n6632) );
  XNOR U7658 ( .A(n6633), .B(n6634), .Z(o[362]) );
  XOR U7659 ( .A(n6635), .B(o[361]), .Z(creg_next[361]) );
  AND U7660 ( .A(n3090), .B(n6636), .Z(n6635) );
  XNOR U7661 ( .A(c[361]), .B(n6637), .Z(n6636) );
  IV U7662 ( .A(o[361]), .Z(n6637) );
  XNOR U7663 ( .A(n6638), .B(n6639), .Z(o[361]) );
  XOR U7664 ( .A(n6640), .B(o[360]), .Z(creg_next[360]) );
  AND U7665 ( .A(n3090), .B(n6641), .Z(n6640) );
  XNOR U7666 ( .A(c[360]), .B(n6642), .Z(n6641) );
  IV U7667 ( .A(o[360]), .Z(n6642) );
  XNOR U7668 ( .A(n6643), .B(n6644), .Z(o[360]) );
  XOR U7669 ( .A(n6645), .B(o[35]), .Z(creg_next[35]) );
  AND U7670 ( .A(n3090), .B(n6646), .Z(n6645) );
  XNOR U7671 ( .A(c[35]), .B(n6647), .Z(n6646) );
  IV U7672 ( .A(o[35]), .Z(n6647) );
  XNOR U7673 ( .A(n6648), .B(n6649), .Z(o[35]) );
  XOR U7674 ( .A(n6650), .B(o[359]), .Z(creg_next[359]) );
  AND U7675 ( .A(n3090), .B(n6651), .Z(n6650) );
  XNOR U7676 ( .A(c[359]), .B(n6652), .Z(n6651) );
  IV U7677 ( .A(o[359]), .Z(n6652) );
  XNOR U7678 ( .A(n6653), .B(n6654), .Z(o[359]) );
  XOR U7679 ( .A(n6655), .B(o[358]), .Z(creg_next[358]) );
  AND U7680 ( .A(n3090), .B(n6656), .Z(n6655) );
  XNOR U7681 ( .A(c[358]), .B(n6657), .Z(n6656) );
  IV U7682 ( .A(o[358]), .Z(n6657) );
  XNOR U7683 ( .A(n6658), .B(n6659), .Z(o[358]) );
  XOR U7684 ( .A(n6660), .B(o[357]), .Z(creg_next[357]) );
  AND U7685 ( .A(n3090), .B(n6661), .Z(n6660) );
  XNOR U7686 ( .A(c[357]), .B(n6662), .Z(n6661) );
  IV U7687 ( .A(o[357]), .Z(n6662) );
  XNOR U7688 ( .A(n6663), .B(n6664), .Z(o[357]) );
  XOR U7689 ( .A(n6665), .B(o[356]), .Z(creg_next[356]) );
  AND U7690 ( .A(n3090), .B(n6666), .Z(n6665) );
  XNOR U7691 ( .A(c[356]), .B(n6667), .Z(n6666) );
  IV U7692 ( .A(o[356]), .Z(n6667) );
  XNOR U7693 ( .A(n6668), .B(n6669), .Z(o[356]) );
  XOR U7694 ( .A(n6670), .B(o[355]), .Z(creg_next[355]) );
  AND U7695 ( .A(n3090), .B(n6671), .Z(n6670) );
  XNOR U7696 ( .A(c[355]), .B(n6672), .Z(n6671) );
  IV U7697 ( .A(o[355]), .Z(n6672) );
  XNOR U7698 ( .A(n6673), .B(n6674), .Z(o[355]) );
  XOR U7699 ( .A(n6675), .B(o[354]), .Z(creg_next[354]) );
  AND U7700 ( .A(n3090), .B(n6676), .Z(n6675) );
  XNOR U7701 ( .A(c[354]), .B(n6677), .Z(n6676) );
  IV U7702 ( .A(o[354]), .Z(n6677) );
  XNOR U7703 ( .A(n6678), .B(n6679), .Z(o[354]) );
  XOR U7704 ( .A(n6680), .B(o[353]), .Z(creg_next[353]) );
  AND U7705 ( .A(n3090), .B(n6681), .Z(n6680) );
  XNOR U7706 ( .A(c[353]), .B(n6682), .Z(n6681) );
  IV U7707 ( .A(o[353]), .Z(n6682) );
  XNOR U7708 ( .A(n6683), .B(n6684), .Z(o[353]) );
  XOR U7709 ( .A(n6685), .B(o[352]), .Z(creg_next[352]) );
  AND U7710 ( .A(n3090), .B(n6686), .Z(n6685) );
  XNOR U7711 ( .A(c[352]), .B(n6687), .Z(n6686) );
  IV U7712 ( .A(o[352]), .Z(n6687) );
  XNOR U7713 ( .A(n6688), .B(n6689), .Z(o[352]) );
  XOR U7714 ( .A(n6690), .B(o[351]), .Z(creg_next[351]) );
  AND U7715 ( .A(n3090), .B(n6691), .Z(n6690) );
  XNOR U7716 ( .A(c[351]), .B(n6692), .Z(n6691) );
  IV U7717 ( .A(o[351]), .Z(n6692) );
  XNOR U7718 ( .A(n6693), .B(n6694), .Z(o[351]) );
  XOR U7719 ( .A(n6695), .B(o[350]), .Z(creg_next[350]) );
  AND U7720 ( .A(n3090), .B(n6696), .Z(n6695) );
  XNOR U7721 ( .A(c[350]), .B(n6697), .Z(n6696) );
  IV U7722 ( .A(o[350]), .Z(n6697) );
  XNOR U7723 ( .A(n6698), .B(n6699), .Z(o[350]) );
  XOR U7724 ( .A(n6700), .B(o[34]), .Z(creg_next[34]) );
  AND U7725 ( .A(n3090), .B(n6701), .Z(n6700) );
  XNOR U7726 ( .A(c[34]), .B(n6702), .Z(n6701) );
  IV U7727 ( .A(o[34]), .Z(n6702) );
  XNOR U7728 ( .A(n6703), .B(n6704), .Z(o[34]) );
  XOR U7729 ( .A(n6705), .B(o[349]), .Z(creg_next[349]) );
  AND U7730 ( .A(n3090), .B(n6706), .Z(n6705) );
  XNOR U7731 ( .A(c[349]), .B(n6707), .Z(n6706) );
  IV U7732 ( .A(o[349]), .Z(n6707) );
  XNOR U7733 ( .A(n6708), .B(n6709), .Z(o[349]) );
  XOR U7734 ( .A(n6710), .B(o[348]), .Z(creg_next[348]) );
  AND U7735 ( .A(n3090), .B(n6711), .Z(n6710) );
  XNOR U7736 ( .A(c[348]), .B(n6712), .Z(n6711) );
  IV U7737 ( .A(o[348]), .Z(n6712) );
  XNOR U7738 ( .A(n6713), .B(n6714), .Z(o[348]) );
  XOR U7739 ( .A(n6715), .B(o[347]), .Z(creg_next[347]) );
  AND U7740 ( .A(n3090), .B(n6716), .Z(n6715) );
  XNOR U7741 ( .A(c[347]), .B(n6717), .Z(n6716) );
  IV U7742 ( .A(o[347]), .Z(n6717) );
  XNOR U7743 ( .A(n6718), .B(n6719), .Z(o[347]) );
  XOR U7744 ( .A(n6720), .B(o[346]), .Z(creg_next[346]) );
  AND U7745 ( .A(n3090), .B(n6721), .Z(n6720) );
  XNOR U7746 ( .A(c[346]), .B(n6722), .Z(n6721) );
  IV U7747 ( .A(o[346]), .Z(n6722) );
  XNOR U7748 ( .A(n6723), .B(n6724), .Z(o[346]) );
  XOR U7749 ( .A(n6725), .B(o[345]), .Z(creg_next[345]) );
  AND U7750 ( .A(n3090), .B(n6726), .Z(n6725) );
  XNOR U7751 ( .A(c[345]), .B(n6727), .Z(n6726) );
  IV U7752 ( .A(o[345]), .Z(n6727) );
  XNOR U7753 ( .A(n6728), .B(n6729), .Z(o[345]) );
  XOR U7754 ( .A(n6730), .B(o[344]), .Z(creg_next[344]) );
  AND U7755 ( .A(n3090), .B(n6731), .Z(n6730) );
  XNOR U7756 ( .A(c[344]), .B(n6732), .Z(n6731) );
  IV U7757 ( .A(o[344]), .Z(n6732) );
  XNOR U7758 ( .A(n6733), .B(n6734), .Z(o[344]) );
  XOR U7759 ( .A(n6735), .B(o[343]), .Z(creg_next[343]) );
  AND U7760 ( .A(n3090), .B(n6736), .Z(n6735) );
  XNOR U7761 ( .A(c[343]), .B(n6737), .Z(n6736) );
  IV U7762 ( .A(o[343]), .Z(n6737) );
  XNOR U7763 ( .A(n6738), .B(n6739), .Z(o[343]) );
  XOR U7764 ( .A(n6740), .B(o[342]), .Z(creg_next[342]) );
  AND U7765 ( .A(n3090), .B(n6741), .Z(n6740) );
  XNOR U7766 ( .A(c[342]), .B(n6742), .Z(n6741) );
  IV U7767 ( .A(o[342]), .Z(n6742) );
  XNOR U7768 ( .A(n6743), .B(n6744), .Z(o[342]) );
  XOR U7769 ( .A(n6745), .B(o[341]), .Z(creg_next[341]) );
  AND U7770 ( .A(n3090), .B(n6746), .Z(n6745) );
  XNOR U7771 ( .A(c[341]), .B(n6747), .Z(n6746) );
  IV U7772 ( .A(o[341]), .Z(n6747) );
  XNOR U7773 ( .A(n6748), .B(n6749), .Z(o[341]) );
  XOR U7774 ( .A(n6750), .B(o[340]), .Z(creg_next[340]) );
  AND U7775 ( .A(n3090), .B(n6751), .Z(n6750) );
  XNOR U7776 ( .A(c[340]), .B(n6752), .Z(n6751) );
  IV U7777 ( .A(o[340]), .Z(n6752) );
  XNOR U7778 ( .A(n6753), .B(n6754), .Z(o[340]) );
  XOR U7779 ( .A(n6755), .B(o[33]), .Z(creg_next[33]) );
  AND U7780 ( .A(n3090), .B(n6756), .Z(n6755) );
  XNOR U7781 ( .A(c[33]), .B(n6757), .Z(n6756) );
  IV U7782 ( .A(o[33]), .Z(n6757) );
  XNOR U7783 ( .A(n6758), .B(n6759), .Z(o[33]) );
  XOR U7784 ( .A(n6760), .B(o[339]), .Z(creg_next[339]) );
  AND U7785 ( .A(n3090), .B(n6761), .Z(n6760) );
  XNOR U7786 ( .A(c[339]), .B(n6762), .Z(n6761) );
  IV U7787 ( .A(o[339]), .Z(n6762) );
  XNOR U7788 ( .A(n6763), .B(n6764), .Z(o[339]) );
  XOR U7789 ( .A(n6765), .B(o[338]), .Z(creg_next[338]) );
  AND U7790 ( .A(n3090), .B(n6766), .Z(n6765) );
  XNOR U7791 ( .A(c[338]), .B(n6767), .Z(n6766) );
  IV U7792 ( .A(o[338]), .Z(n6767) );
  XNOR U7793 ( .A(n6768), .B(n6769), .Z(o[338]) );
  XOR U7794 ( .A(n6770), .B(o[337]), .Z(creg_next[337]) );
  AND U7795 ( .A(n3090), .B(n6771), .Z(n6770) );
  XNOR U7796 ( .A(c[337]), .B(n6772), .Z(n6771) );
  IV U7797 ( .A(o[337]), .Z(n6772) );
  XNOR U7798 ( .A(n6773), .B(n6774), .Z(o[337]) );
  XOR U7799 ( .A(n6775), .B(o[336]), .Z(creg_next[336]) );
  AND U7800 ( .A(n3090), .B(n6776), .Z(n6775) );
  XNOR U7801 ( .A(c[336]), .B(n6777), .Z(n6776) );
  IV U7802 ( .A(o[336]), .Z(n6777) );
  XNOR U7803 ( .A(n6778), .B(n6779), .Z(o[336]) );
  XOR U7804 ( .A(n6780), .B(o[335]), .Z(creg_next[335]) );
  AND U7805 ( .A(n3090), .B(n6781), .Z(n6780) );
  XNOR U7806 ( .A(c[335]), .B(n6782), .Z(n6781) );
  IV U7807 ( .A(o[335]), .Z(n6782) );
  XNOR U7808 ( .A(n6783), .B(n6784), .Z(o[335]) );
  XOR U7809 ( .A(n6785), .B(o[334]), .Z(creg_next[334]) );
  AND U7810 ( .A(n3090), .B(n6786), .Z(n6785) );
  XNOR U7811 ( .A(c[334]), .B(n6787), .Z(n6786) );
  IV U7812 ( .A(o[334]), .Z(n6787) );
  XNOR U7813 ( .A(n6788), .B(n6789), .Z(o[334]) );
  XOR U7814 ( .A(n6790), .B(o[333]), .Z(creg_next[333]) );
  AND U7815 ( .A(n3090), .B(n6791), .Z(n6790) );
  XNOR U7816 ( .A(c[333]), .B(n6792), .Z(n6791) );
  IV U7817 ( .A(o[333]), .Z(n6792) );
  XNOR U7818 ( .A(n6793), .B(n6794), .Z(o[333]) );
  XOR U7819 ( .A(n6795), .B(o[332]), .Z(creg_next[332]) );
  AND U7820 ( .A(n3090), .B(n6796), .Z(n6795) );
  XNOR U7821 ( .A(c[332]), .B(n6797), .Z(n6796) );
  IV U7822 ( .A(o[332]), .Z(n6797) );
  XNOR U7823 ( .A(n6798), .B(n6799), .Z(o[332]) );
  XOR U7824 ( .A(n6800), .B(o[331]), .Z(creg_next[331]) );
  AND U7825 ( .A(n3090), .B(n6801), .Z(n6800) );
  XNOR U7826 ( .A(c[331]), .B(n6802), .Z(n6801) );
  IV U7827 ( .A(o[331]), .Z(n6802) );
  XNOR U7828 ( .A(n6803), .B(n6804), .Z(o[331]) );
  XOR U7829 ( .A(n6805), .B(o[330]), .Z(creg_next[330]) );
  AND U7830 ( .A(n3090), .B(n6806), .Z(n6805) );
  XNOR U7831 ( .A(c[330]), .B(n6807), .Z(n6806) );
  IV U7832 ( .A(o[330]), .Z(n6807) );
  XNOR U7833 ( .A(n6808), .B(n6809), .Z(o[330]) );
  XOR U7834 ( .A(n6810), .B(o[32]), .Z(creg_next[32]) );
  AND U7835 ( .A(n3090), .B(n6811), .Z(n6810) );
  XNOR U7836 ( .A(c[32]), .B(n6812), .Z(n6811) );
  IV U7837 ( .A(o[32]), .Z(n6812) );
  XNOR U7838 ( .A(n6813), .B(n6814), .Z(o[32]) );
  XOR U7839 ( .A(n6815), .B(o[329]), .Z(creg_next[329]) );
  AND U7840 ( .A(n3090), .B(n6816), .Z(n6815) );
  XNOR U7841 ( .A(c[329]), .B(n6817), .Z(n6816) );
  IV U7842 ( .A(o[329]), .Z(n6817) );
  XNOR U7843 ( .A(n6818), .B(n6819), .Z(o[329]) );
  XOR U7844 ( .A(n6820), .B(o[328]), .Z(creg_next[328]) );
  AND U7845 ( .A(n3090), .B(n6821), .Z(n6820) );
  XNOR U7846 ( .A(c[328]), .B(n6822), .Z(n6821) );
  IV U7847 ( .A(o[328]), .Z(n6822) );
  XNOR U7848 ( .A(n6823), .B(n6824), .Z(o[328]) );
  XOR U7849 ( .A(n6825), .B(o[327]), .Z(creg_next[327]) );
  AND U7850 ( .A(n3090), .B(n6826), .Z(n6825) );
  XNOR U7851 ( .A(c[327]), .B(n6827), .Z(n6826) );
  IV U7852 ( .A(o[327]), .Z(n6827) );
  XNOR U7853 ( .A(n6828), .B(n6829), .Z(o[327]) );
  XOR U7854 ( .A(n6830), .B(o[326]), .Z(creg_next[326]) );
  AND U7855 ( .A(n3090), .B(n6831), .Z(n6830) );
  XNOR U7856 ( .A(c[326]), .B(n6832), .Z(n6831) );
  IV U7857 ( .A(o[326]), .Z(n6832) );
  XNOR U7858 ( .A(n6833), .B(n6834), .Z(o[326]) );
  XOR U7859 ( .A(n6835), .B(o[325]), .Z(creg_next[325]) );
  AND U7860 ( .A(n3090), .B(n6836), .Z(n6835) );
  XNOR U7861 ( .A(c[325]), .B(n6837), .Z(n6836) );
  IV U7862 ( .A(o[325]), .Z(n6837) );
  XNOR U7863 ( .A(n6838), .B(n6839), .Z(o[325]) );
  XOR U7864 ( .A(n6840), .B(o[324]), .Z(creg_next[324]) );
  AND U7865 ( .A(n3090), .B(n6841), .Z(n6840) );
  XNOR U7866 ( .A(c[324]), .B(n6842), .Z(n6841) );
  IV U7867 ( .A(o[324]), .Z(n6842) );
  XNOR U7868 ( .A(n6843), .B(n6844), .Z(o[324]) );
  XOR U7869 ( .A(n6845), .B(o[323]), .Z(creg_next[323]) );
  AND U7870 ( .A(n3090), .B(n6846), .Z(n6845) );
  XNOR U7871 ( .A(c[323]), .B(n6847), .Z(n6846) );
  IV U7872 ( .A(o[323]), .Z(n6847) );
  XNOR U7873 ( .A(n6848), .B(n6849), .Z(o[323]) );
  XOR U7874 ( .A(n6850), .B(o[322]), .Z(creg_next[322]) );
  AND U7875 ( .A(n3090), .B(n6851), .Z(n6850) );
  XNOR U7876 ( .A(c[322]), .B(n6852), .Z(n6851) );
  IV U7877 ( .A(o[322]), .Z(n6852) );
  XNOR U7878 ( .A(n6853), .B(n6854), .Z(o[322]) );
  XOR U7879 ( .A(n6855), .B(o[321]), .Z(creg_next[321]) );
  AND U7880 ( .A(n3090), .B(n6856), .Z(n6855) );
  XNOR U7881 ( .A(c[321]), .B(n6857), .Z(n6856) );
  IV U7882 ( .A(o[321]), .Z(n6857) );
  XNOR U7883 ( .A(n6858), .B(n6859), .Z(o[321]) );
  XOR U7884 ( .A(n6860), .B(o[320]), .Z(creg_next[320]) );
  AND U7885 ( .A(n3090), .B(n6861), .Z(n6860) );
  XNOR U7886 ( .A(c[320]), .B(n6862), .Z(n6861) );
  IV U7887 ( .A(o[320]), .Z(n6862) );
  XNOR U7888 ( .A(n6863), .B(n6864), .Z(o[320]) );
  XOR U7889 ( .A(n6865), .B(o[31]), .Z(creg_next[31]) );
  AND U7890 ( .A(n3090), .B(n6866), .Z(n6865) );
  XNOR U7891 ( .A(c[31]), .B(n6867), .Z(n6866) );
  IV U7892 ( .A(o[31]), .Z(n6867) );
  XNOR U7893 ( .A(n6868), .B(n6869), .Z(o[31]) );
  XOR U7894 ( .A(n6870), .B(o[319]), .Z(creg_next[319]) );
  AND U7895 ( .A(n3090), .B(n6871), .Z(n6870) );
  XNOR U7896 ( .A(c[319]), .B(n6872), .Z(n6871) );
  IV U7897 ( .A(o[319]), .Z(n6872) );
  XNOR U7898 ( .A(n6873), .B(n6874), .Z(o[319]) );
  XOR U7899 ( .A(n6875), .B(o[318]), .Z(creg_next[318]) );
  AND U7900 ( .A(n3090), .B(n6876), .Z(n6875) );
  XNOR U7901 ( .A(c[318]), .B(n6877), .Z(n6876) );
  IV U7902 ( .A(o[318]), .Z(n6877) );
  XNOR U7903 ( .A(n6878), .B(n6879), .Z(o[318]) );
  XOR U7904 ( .A(n6880), .B(o[317]), .Z(creg_next[317]) );
  AND U7905 ( .A(n3090), .B(n6881), .Z(n6880) );
  XNOR U7906 ( .A(c[317]), .B(n6882), .Z(n6881) );
  IV U7907 ( .A(o[317]), .Z(n6882) );
  XNOR U7908 ( .A(n6883), .B(n6884), .Z(o[317]) );
  XOR U7909 ( .A(n6885), .B(o[316]), .Z(creg_next[316]) );
  AND U7910 ( .A(n3090), .B(n6886), .Z(n6885) );
  XNOR U7911 ( .A(c[316]), .B(n6887), .Z(n6886) );
  IV U7912 ( .A(o[316]), .Z(n6887) );
  XNOR U7913 ( .A(n6888), .B(n6889), .Z(o[316]) );
  XOR U7914 ( .A(n6890), .B(o[315]), .Z(creg_next[315]) );
  AND U7915 ( .A(n3090), .B(n6891), .Z(n6890) );
  XNOR U7916 ( .A(c[315]), .B(n6892), .Z(n6891) );
  IV U7917 ( .A(o[315]), .Z(n6892) );
  XNOR U7918 ( .A(n6893), .B(n6894), .Z(o[315]) );
  XOR U7919 ( .A(n6895), .B(o[314]), .Z(creg_next[314]) );
  AND U7920 ( .A(n3090), .B(n6896), .Z(n6895) );
  XNOR U7921 ( .A(c[314]), .B(n6897), .Z(n6896) );
  IV U7922 ( .A(o[314]), .Z(n6897) );
  XNOR U7923 ( .A(n6898), .B(n6899), .Z(o[314]) );
  XOR U7924 ( .A(n6900), .B(o[313]), .Z(creg_next[313]) );
  AND U7925 ( .A(n3090), .B(n6901), .Z(n6900) );
  XNOR U7926 ( .A(c[313]), .B(n6902), .Z(n6901) );
  IV U7927 ( .A(o[313]), .Z(n6902) );
  XNOR U7928 ( .A(n6903), .B(n6904), .Z(o[313]) );
  XOR U7929 ( .A(n6905), .B(o[312]), .Z(creg_next[312]) );
  AND U7930 ( .A(n3090), .B(n6906), .Z(n6905) );
  XNOR U7931 ( .A(c[312]), .B(n6907), .Z(n6906) );
  IV U7932 ( .A(o[312]), .Z(n6907) );
  XNOR U7933 ( .A(n6908), .B(n6909), .Z(o[312]) );
  XOR U7934 ( .A(n6910), .B(o[311]), .Z(creg_next[311]) );
  AND U7935 ( .A(n3090), .B(n6911), .Z(n6910) );
  XNOR U7936 ( .A(c[311]), .B(n6912), .Z(n6911) );
  IV U7937 ( .A(o[311]), .Z(n6912) );
  XNOR U7938 ( .A(n6913), .B(n6914), .Z(o[311]) );
  XOR U7939 ( .A(n6915), .B(o[310]), .Z(creg_next[310]) );
  AND U7940 ( .A(n3090), .B(n6916), .Z(n6915) );
  XNOR U7941 ( .A(c[310]), .B(n6917), .Z(n6916) );
  IV U7942 ( .A(o[310]), .Z(n6917) );
  XNOR U7943 ( .A(n6918), .B(n6919), .Z(o[310]) );
  XOR U7944 ( .A(n6920), .B(o[30]), .Z(creg_next[30]) );
  AND U7945 ( .A(n3090), .B(n6921), .Z(n6920) );
  XNOR U7946 ( .A(c[30]), .B(n6922), .Z(n6921) );
  IV U7947 ( .A(o[30]), .Z(n6922) );
  XNOR U7948 ( .A(n6923), .B(n6924), .Z(o[30]) );
  XOR U7949 ( .A(n6925), .B(o[309]), .Z(creg_next[309]) );
  AND U7950 ( .A(n3090), .B(n6926), .Z(n6925) );
  XNOR U7951 ( .A(c[309]), .B(n6927), .Z(n6926) );
  IV U7952 ( .A(o[309]), .Z(n6927) );
  XNOR U7953 ( .A(n6928), .B(n6929), .Z(o[309]) );
  XOR U7954 ( .A(n6930), .B(o[308]), .Z(creg_next[308]) );
  AND U7955 ( .A(n3090), .B(n6931), .Z(n6930) );
  XNOR U7956 ( .A(c[308]), .B(n6932), .Z(n6931) );
  IV U7957 ( .A(o[308]), .Z(n6932) );
  XNOR U7958 ( .A(n6933), .B(n6934), .Z(o[308]) );
  XOR U7959 ( .A(n6935), .B(o[307]), .Z(creg_next[307]) );
  AND U7960 ( .A(n3090), .B(n6936), .Z(n6935) );
  XNOR U7961 ( .A(c[307]), .B(n6937), .Z(n6936) );
  IV U7962 ( .A(o[307]), .Z(n6937) );
  XNOR U7963 ( .A(n6938), .B(n6939), .Z(o[307]) );
  XOR U7964 ( .A(n6940), .B(o[306]), .Z(creg_next[306]) );
  AND U7965 ( .A(n3090), .B(n6941), .Z(n6940) );
  XNOR U7966 ( .A(c[306]), .B(n6942), .Z(n6941) );
  IV U7967 ( .A(o[306]), .Z(n6942) );
  XNOR U7968 ( .A(n6943), .B(n6944), .Z(o[306]) );
  XOR U7969 ( .A(n6945), .B(o[305]), .Z(creg_next[305]) );
  AND U7970 ( .A(n3090), .B(n6946), .Z(n6945) );
  XNOR U7971 ( .A(c[305]), .B(n6947), .Z(n6946) );
  IV U7972 ( .A(o[305]), .Z(n6947) );
  XNOR U7973 ( .A(n6948), .B(n6949), .Z(o[305]) );
  XOR U7974 ( .A(n6950), .B(o[304]), .Z(creg_next[304]) );
  AND U7975 ( .A(n3090), .B(n6951), .Z(n6950) );
  XNOR U7976 ( .A(c[304]), .B(n6952), .Z(n6951) );
  IV U7977 ( .A(o[304]), .Z(n6952) );
  XNOR U7978 ( .A(n6953), .B(n6954), .Z(o[304]) );
  XOR U7979 ( .A(n6955), .B(o[303]), .Z(creg_next[303]) );
  AND U7980 ( .A(n3090), .B(n6956), .Z(n6955) );
  XNOR U7981 ( .A(c[303]), .B(n6957), .Z(n6956) );
  IV U7982 ( .A(o[303]), .Z(n6957) );
  XNOR U7983 ( .A(n6958), .B(n6959), .Z(o[303]) );
  XOR U7984 ( .A(n6960), .B(o[302]), .Z(creg_next[302]) );
  AND U7985 ( .A(n3090), .B(n6961), .Z(n6960) );
  XNOR U7986 ( .A(c[302]), .B(n6962), .Z(n6961) );
  IV U7987 ( .A(o[302]), .Z(n6962) );
  XNOR U7988 ( .A(n6963), .B(n6964), .Z(o[302]) );
  XOR U7989 ( .A(n6965), .B(o[301]), .Z(creg_next[301]) );
  AND U7990 ( .A(n3090), .B(n6966), .Z(n6965) );
  XNOR U7991 ( .A(c[301]), .B(n6967), .Z(n6966) );
  IV U7992 ( .A(o[301]), .Z(n6967) );
  XNOR U7993 ( .A(n6968), .B(n6969), .Z(o[301]) );
  XOR U7994 ( .A(n6970), .B(o[300]), .Z(creg_next[300]) );
  AND U7995 ( .A(n3090), .B(n6971), .Z(n6970) );
  XNOR U7996 ( .A(c[300]), .B(n6972), .Z(n6971) );
  IV U7997 ( .A(o[300]), .Z(n6972) );
  XNOR U7998 ( .A(n6973), .B(n6974), .Z(o[300]) );
  XOR U7999 ( .A(n6975), .B(o[2]), .Z(creg_next[2]) );
  AND U8000 ( .A(n3090), .B(n6976), .Z(n6975) );
  XNOR U8001 ( .A(c[2]), .B(n6977), .Z(n6976) );
  IV U8002 ( .A(o[2]), .Z(n6977) );
  XNOR U8003 ( .A(n6978), .B(n6979), .Z(o[2]) );
  XOR U8004 ( .A(n6980), .B(o[29]), .Z(creg_next[29]) );
  AND U8005 ( .A(n3090), .B(n6981), .Z(n6980) );
  XNOR U8006 ( .A(c[29]), .B(n6982), .Z(n6981) );
  IV U8007 ( .A(o[29]), .Z(n6982) );
  XNOR U8008 ( .A(n6983), .B(n6984), .Z(o[29]) );
  XOR U8009 ( .A(n6985), .B(o[299]), .Z(creg_next[299]) );
  AND U8010 ( .A(n3090), .B(n6986), .Z(n6985) );
  XNOR U8011 ( .A(c[299]), .B(n6987), .Z(n6986) );
  IV U8012 ( .A(o[299]), .Z(n6987) );
  XNOR U8013 ( .A(n6988), .B(n6989), .Z(o[299]) );
  XOR U8014 ( .A(n6990), .B(o[298]), .Z(creg_next[298]) );
  AND U8015 ( .A(n3090), .B(n6991), .Z(n6990) );
  XNOR U8016 ( .A(c[298]), .B(n6992), .Z(n6991) );
  IV U8017 ( .A(o[298]), .Z(n6992) );
  XNOR U8018 ( .A(n6993), .B(n6994), .Z(o[298]) );
  XOR U8019 ( .A(n6995), .B(o[297]), .Z(creg_next[297]) );
  AND U8020 ( .A(n3090), .B(n6996), .Z(n6995) );
  XNOR U8021 ( .A(c[297]), .B(n6997), .Z(n6996) );
  IV U8022 ( .A(o[297]), .Z(n6997) );
  XNOR U8023 ( .A(n6998), .B(n6999), .Z(o[297]) );
  XOR U8024 ( .A(n7000), .B(o[296]), .Z(creg_next[296]) );
  AND U8025 ( .A(n3090), .B(n7001), .Z(n7000) );
  XNOR U8026 ( .A(c[296]), .B(n7002), .Z(n7001) );
  IV U8027 ( .A(o[296]), .Z(n7002) );
  XNOR U8028 ( .A(n7003), .B(n7004), .Z(o[296]) );
  XOR U8029 ( .A(n7005), .B(o[295]), .Z(creg_next[295]) );
  AND U8030 ( .A(n3090), .B(n7006), .Z(n7005) );
  XNOR U8031 ( .A(c[295]), .B(n7007), .Z(n7006) );
  IV U8032 ( .A(o[295]), .Z(n7007) );
  XNOR U8033 ( .A(n7008), .B(n7009), .Z(o[295]) );
  XOR U8034 ( .A(n7010), .B(o[294]), .Z(creg_next[294]) );
  AND U8035 ( .A(n3090), .B(n7011), .Z(n7010) );
  XNOR U8036 ( .A(c[294]), .B(n7012), .Z(n7011) );
  IV U8037 ( .A(o[294]), .Z(n7012) );
  XNOR U8038 ( .A(n7013), .B(n7014), .Z(o[294]) );
  XOR U8039 ( .A(n7015), .B(o[293]), .Z(creg_next[293]) );
  AND U8040 ( .A(n3090), .B(n7016), .Z(n7015) );
  XNOR U8041 ( .A(c[293]), .B(n7017), .Z(n7016) );
  IV U8042 ( .A(o[293]), .Z(n7017) );
  XNOR U8043 ( .A(n7018), .B(n7019), .Z(o[293]) );
  XOR U8044 ( .A(n7020), .B(o[292]), .Z(creg_next[292]) );
  AND U8045 ( .A(n3090), .B(n7021), .Z(n7020) );
  XNOR U8046 ( .A(c[292]), .B(n7022), .Z(n7021) );
  IV U8047 ( .A(o[292]), .Z(n7022) );
  XNOR U8048 ( .A(n7023), .B(n7024), .Z(o[292]) );
  XOR U8049 ( .A(n7025), .B(o[291]), .Z(creg_next[291]) );
  AND U8050 ( .A(n3090), .B(n7026), .Z(n7025) );
  XNOR U8051 ( .A(c[291]), .B(n7027), .Z(n7026) );
  IV U8052 ( .A(o[291]), .Z(n7027) );
  XNOR U8053 ( .A(n7028), .B(n7029), .Z(o[291]) );
  XOR U8054 ( .A(n7030), .B(o[290]), .Z(creg_next[290]) );
  AND U8055 ( .A(n3090), .B(n7031), .Z(n7030) );
  XNOR U8056 ( .A(c[290]), .B(n7032), .Z(n7031) );
  IV U8057 ( .A(o[290]), .Z(n7032) );
  XNOR U8058 ( .A(n7033), .B(n7034), .Z(o[290]) );
  XOR U8059 ( .A(n7035), .B(o[28]), .Z(creg_next[28]) );
  AND U8060 ( .A(n3090), .B(n7036), .Z(n7035) );
  XNOR U8061 ( .A(c[28]), .B(n7037), .Z(n7036) );
  IV U8062 ( .A(o[28]), .Z(n7037) );
  XNOR U8063 ( .A(n7038), .B(n7039), .Z(o[28]) );
  XOR U8064 ( .A(n7040), .B(o[289]), .Z(creg_next[289]) );
  AND U8065 ( .A(n3090), .B(n7041), .Z(n7040) );
  XNOR U8066 ( .A(c[289]), .B(n7042), .Z(n7041) );
  IV U8067 ( .A(o[289]), .Z(n7042) );
  XNOR U8068 ( .A(n7043), .B(n7044), .Z(o[289]) );
  XOR U8069 ( .A(n7045), .B(o[288]), .Z(creg_next[288]) );
  AND U8070 ( .A(n3090), .B(n7046), .Z(n7045) );
  XNOR U8071 ( .A(c[288]), .B(n7047), .Z(n7046) );
  IV U8072 ( .A(o[288]), .Z(n7047) );
  XNOR U8073 ( .A(n7048), .B(n7049), .Z(o[288]) );
  XOR U8074 ( .A(n7050), .B(o[287]), .Z(creg_next[287]) );
  AND U8075 ( .A(n3090), .B(n7051), .Z(n7050) );
  XNOR U8076 ( .A(c[287]), .B(n7052), .Z(n7051) );
  IV U8077 ( .A(o[287]), .Z(n7052) );
  XNOR U8078 ( .A(n7053), .B(n7054), .Z(o[287]) );
  XOR U8079 ( .A(n7055), .B(o[286]), .Z(creg_next[286]) );
  AND U8080 ( .A(n3090), .B(n7056), .Z(n7055) );
  XNOR U8081 ( .A(c[286]), .B(n7057), .Z(n7056) );
  IV U8082 ( .A(o[286]), .Z(n7057) );
  XNOR U8083 ( .A(n7058), .B(n7059), .Z(o[286]) );
  XOR U8084 ( .A(n7060), .B(o[285]), .Z(creg_next[285]) );
  AND U8085 ( .A(n3090), .B(n7061), .Z(n7060) );
  XNOR U8086 ( .A(c[285]), .B(n7062), .Z(n7061) );
  IV U8087 ( .A(o[285]), .Z(n7062) );
  XNOR U8088 ( .A(n7063), .B(n7064), .Z(o[285]) );
  XOR U8089 ( .A(n7065), .B(o[284]), .Z(creg_next[284]) );
  AND U8090 ( .A(n3090), .B(n7066), .Z(n7065) );
  XNOR U8091 ( .A(c[284]), .B(n7067), .Z(n7066) );
  IV U8092 ( .A(o[284]), .Z(n7067) );
  XNOR U8093 ( .A(n7068), .B(n7069), .Z(o[284]) );
  XOR U8094 ( .A(n7070), .B(o[283]), .Z(creg_next[283]) );
  AND U8095 ( .A(n3090), .B(n7071), .Z(n7070) );
  XNOR U8096 ( .A(c[283]), .B(n7072), .Z(n7071) );
  IV U8097 ( .A(o[283]), .Z(n7072) );
  XNOR U8098 ( .A(n7073), .B(n7074), .Z(o[283]) );
  XOR U8099 ( .A(n7075), .B(o[282]), .Z(creg_next[282]) );
  AND U8100 ( .A(n3090), .B(n7076), .Z(n7075) );
  XNOR U8101 ( .A(c[282]), .B(n7077), .Z(n7076) );
  IV U8102 ( .A(o[282]), .Z(n7077) );
  XNOR U8103 ( .A(n7078), .B(n7079), .Z(o[282]) );
  XOR U8104 ( .A(n7080), .B(o[281]), .Z(creg_next[281]) );
  AND U8105 ( .A(n3090), .B(n7081), .Z(n7080) );
  XNOR U8106 ( .A(c[281]), .B(n7082), .Z(n7081) );
  IV U8107 ( .A(o[281]), .Z(n7082) );
  XNOR U8108 ( .A(n7083), .B(n7084), .Z(o[281]) );
  XOR U8109 ( .A(n7085), .B(o[280]), .Z(creg_next[280]) );
  AND U8110 ( .A(n3090), .B(n7086), .Z(n7085) );
  XNOR U8111 ( .A(c[280]), .B(n7087), .Z(n7086) );
  IV U8112 ( .A(o[280]), .Z(n7087) );
  XNOR U8113 ( .A(n7088), .B(n7089), .Z(o[280]) );
  XOR U8114 ( .A(n7090), .B(o[27]), .Z(creg_next[27]) );
  AND U8115 ( .A(n3090), .B(n7091), .Z(n7090) );
  XNOR U8116 ( .A(c[27]), .B(n7092), .Z(n7091) );
  IV U8117 ( .A(o[27]), .Z(n7092) );
  XNOR U8118 ( .A(n7093), .B(n7094), .Z(o[27]) );
  XOR U8119 ( .A(n7095), .B(o[279]), .Z(creg_next[279]) );
  AND U8120 ( .A(n3090), .B(n7096), .Z(n7095) );
  XNOR U8121 ( .A(c[279]), .B(n7097), .Z(n7096) );
  IV U8122 ( .A(o[279]), .Z(n7097) );
  XNOR U8123 ( .A(n7098), .B(n7099), .Z(o[279]) );
  XOR U8124 ( .A(n7100), .B(o[278]), .Z(creg_next[278]) );
  AND U8125 ( .A(n3090), .B(n7101), .Z(n7100) );
  XNOR U8126 ( .A(c[278]), .B(n7102), .Z(n7101) );
  IV U8127 ( .A(o[278]), .Z(n7102) );
  XNOR U8128 ( .A(n7103), .B(n7104), .Z(o[278]) );
  XOR U8129 ( .A(n7105), .B(o[277]), .Z(creg_next[277]) );
  AND U8130 ( .A(n3090), .B(n7106), .Z(n7105) );
  XNOR U8131 ( .A(c[277]), .B(n7107), .Z(n7106) );
  IV U8132 ( .A(o[277]), .Z(n7107) );
  XNOR U8133 ( .A(n7108), .B(n7109), .Z(o[277]) );
  XOR U8134 ( .A(n7110), .B(o[276]), .Z(creg_next[276]) );
  AND U8135 ( .A(n3090), .B(n7111), .Z(n7110) );
  XNOR U8136 ( .A(c[276]), .B(n7112), .Z(n7111) );
  IV U8137 ( .A(o[276]), .Z(n7112) );
  XNOR U8138 ( .A(n7113), .B(n7114), .Z(o[276]) );
  XOR U8139 ( .A(n7115), .B(o[275]), .Z(creg_next[275]) );
  AND U8140 ( .A(n3090), .B(n7116), .Z(n7115) );
  XNOR U8141 ( .A(c[275]), .B(n7117), .Z(n7116) );
  IV U8142 ( .A(o[275]), .Z(n7117) );
  XNOR U8143 ( .A(n7118), .B(n7119), .Z(o[275]) );
  XOR U8144 ( .A(n7120), .B(o[274]), .Z(creg_next[274]) );
  AND U8145 ( .A(n3090), .B(n7121), .Z(n7120) );
  XNOR U8146 ( .A(c[274]), .B(n7122), .Z(n7121) );
  IV U8147 ( .A(o[274]), .Z(n7122) );
  XNOR U8148 ( .A(n7123), .B(n7124), .Z(o[274]) );
  XOR U8149 ( .A(n7125), .B(o[273]), .Z(creg_next[273]) );
  AND U8150 ( .A(n3090), .B(n7126), .Z(n7125) );
  XNOR U8151 ( .A(c[273]), .B(n7127), .Z(n7126) );
  IV U8152 ( .A(o[273]), .Z(n7127) );
  XNOR U8153 ( .A(n7128), .B(n7129), .Z(o[273]) );
  XOR U8154 ( .A(n7130), .B(o[272]), .Z(creg_next[272]) );
  AND U8155 ( .A(n3090), .B(n7131), .Z(n7130) );
  XNOR U8156 ( .A(c[272]), .B(n7132), .Z(n7131) );
  IV U8157 ( .A(o[272]), .Z(n7132) );
  XNOR U8158 ( .A(n7133), .B(n7134), .Z(o[272]) );
  XOR U8159 ( .A(n7135), .B(o[271]), .Z(creg_next[271]) );
  AND U8160 ( .A(n3090), .B(n7136), .Z(n7135) );
  XNOR U8161 ( .A(c[271]), .B(n7137), .Z(n7136) );
  IV U8162 ( .A(o[271]), .Z(n7137) );
  XNOR U8163 ( .A(n7138), .B(n7139), .Z(o[271]) );
  XOR U8164 ( .A(n7140), .B(o[270]), .Z(creg_next[270]) );
  AND U8165 ( .A(n3090), .B(n7141), .Z(n7140) );
  XNOR U8166 ( .A(c[270]), .B(n7142), .Z(n7141) );
  IV U8167 ( .A(o[270]), .Z(n7142) );
  XNOR U8168 ( .A(n7143), .B(n7144), .Z(o[270]) );
  XOR U8169 ( .A(n7145), .B(o[26]), .Z(creg_next[26]) );
  AND U8170 ( .A(n3090), .B(n7146), .Z(n7145) );
  XNOR U8171 ( .A(c[26]), .B(n7147), .Z(n7146) );
  IV U8172 ( .A(o[26]), .Z(n7147) );
  XNOR U8173 ( .A(n7148), .B(n7149), .Z(o[26]) );
  XOR U8174 ( .A(n7150), .B(o[269]), .Z(creg_next[269]) );
  AND U8175 ( .A(n3090), .B(n7151), .Z(n7150) );
  XNOR U8176 ( .A(c[269]), .B(n7152), .Z(n7151) );
  IV U8177 ( .A(o[269]), .Z(n7152) );
  XNOR U8178 ( .A(n7153), .B(n7154), .Z(o[269]) );
  XOR U8179 ( .A(n7155), .B(o[268]), .Z(creg_next[268]) );
  AND U8180 ( .A(n3090), .B(n7156), .Z(n7155) );
  XNOR U8181 ( .A(c[268]), .B(n7157), .Z(n7156) );
  IV U8182 ( .A(o[268]), .Z(n7157) );
  XNOR U8183 ( .A(n7158), .B(n7159), .Z(o[268]) );
  XOR U8184 ( .A(n7160), .B(o[267]), .Z(creg_next[267]) );
  AND U8185 ( .A(n3090), .B(n7161), .Z(n7160) );
  XNOR U8186 ( .A(c[267]), .B(n7162), .Z(n7161) );
  IV U8187 ( .A(o[267]), .Z(n7162) );
  XNOR U8188 ( .A(n7163), .B(n7164), .Z(o[267]) );
  XOR U8189 ( .A(n7165), .B(o[266]), .Z(creg_next[266]) );
  AND U8190 ( .A(n3090), .B(n7166), .Z(n7165) );
  XNOR U8191 ( .A(c[266]), .B(n7167), .Z(n7166) );
  IV U8192 ( .A(o[266]), .Z(n7167) );
  XNOR U8193 ( .A(n7168), .B(n7169), .Z(o[266]) );
  XOR U8194 ( .A(n7170), .B(o[265]), .Z(creg_next[265]) );
  AND U8195 ( .A(n3090), .B(n7171), .Z(n7170) );
  XNOR U8196 ( .A(c[265]), .B(n7172), .Z(n7171) );
  IV U8197 ( .A(o[265]), .Z(n7172) );
  XNOR U8198 ( .A(n7173), .B(n7174), .Z(o[265]) );
  XOR U8199 ( .A(n7175), .B(o[264]), .Z(creg_next[264]) );
  AND U8200 ( .A(n3090), .B(n7176), .Z(n7175) );
  XNOR U8201 ( .A(c[264]), .B(n7177), .Z(n7176) );
  IV U8202 ( .A(o[264]), .Z(n7177) );
  XNOR U8203 ( .A(n7178), .B(n7179), .Z(o[264]) );
  XOR U8204 ( .A(n7180), .B(o[263]), .Z(creg_next[263]) );
  AND U8205 ( .A(n3090), .B(n7181), .Z(n7180) );
  XNOR U8206 ( .A(c[263]), .B(n7182), .Z(n7181) );
  IV U8207 ( .A(o[263]), .Z(n7182) );
  XNOR U8208 ( .A(n7183), .B(n7184), .Z(o[263]) );
  XOR U8209 ( .A(n7185), .B(o[262]), .Z(creg_next[262]) );
  AND U8210 ( .A(n3090), .B(n7186), .Z(n7185) );
  XNOR U8211 ( .A(c[262]), .B(n7187), .Z(n7186) );
  IV U8212 ( .A(o[262]), .Z(n7187) );
  XNOR U8213 ( .A(n7188), .B(n7189), .Z(o[262]) );
  XOR U8214 ( .A(n7190), .B(o[261]), .Z(creg_next[261]) );
  AND U8215 ( .A(n3090), .B(n7191), .Z(n7190) );
  XNOR U8216 ( .A(c[261]), .B(n7192), .Z(n7191) );
  IV U8217 ( .A(o[261]), .Z(n7192) );
  XNOR U8218 ( .A(n7193), .B(n7194), .Z(o[261]) );
  XOR U8219 ( .A(n7195), .B(o[260]), .Z(creg_next[260]) );
  AND U8220 ( .A(n3090), .B(n7196), .Z(n7195) );
  XNOR U8221 ( .A(c[260]), .B(n7197), .Z(n7196) );
  IV U8222 ( .A(o[260]), .Z(n7197) );
  XNOR U8223 ( .A(n7198), .B(n7199), .Z(o[260]) );
  XOR U8224 ( .A(n7200), .B(o[25]), .Z(creg_next[25]) );
  AND U8225 ( .A(n3090), .B(n7201), .Z(n7200) );
  XNOR U8226 ( .A(c[25]), .B(n7202), .Z(n7201) );
  IV U8227 ( .A(o[25]), .Z(n7202) );
  XNOR U8228 ( .A(n7203), .B(n7204), .Z(o[25]) );
  XOR U8229 ( .A(n7205), .B(o[259]), .Z(creg_next[259]) );
  AND U8230 ( .A(n3090), .B(n7206), .Z(n7205) );
  XNOR U8231 ( .A(c[259]), .B(n7207), .Z(n7206) );
  IV U8232 ( .A(o[259]), .Z(n7207) );
  XNOR U8233 ( .A(n7208), .B(n7209), .Z(o[259]) );
  XOR U8234 ( .A(n7210), .B(o[258]), .Z(creg_next[258]) );
  AND U8235 ( .A(n3090), .B(n7211), .Z(n7210) );
  XNOR U8236 ( .A(c[258]), .B(n7212), .Z(n7211) );
  IV U8237 ( .A(o[258]), .Z(n7212) );
  XNOR U8238 ( .A(n7213), .B(n7214), .Z(o[258]) );
  XOR U8239 ( .A(n7215), .B(o[257]), .Z(creg_next[257]) );
  AND U8240 ( .A(n3090), .B(n7216), .Z(n7215) );
  XNOR U8241 ( .A(c[257]), .B(n7217), .Z(n7216) );
  IV U8242 ( .A(o[257]), .Z(n7217) );
  XNOR U8243 ( .A(n7218), .B(n7219), .Z(o[257]) );
  XOR U8244 ( .A(n7220), .B(o[256]), .Z(creg_next[256]) );
  AND U8245 ( .A(n3090), .B(n7221), .Z(n7220) );
  XNOR U8246 ( .A(c[256]), .B(n7222), .Z(n7221) );
  IV U8247 ( .A(o[256]), .Z(n7222) );
  XNOR U8248 ( .A(n7223), .B(n7224), .Z(o[256]) );
  XOR U8249 ( .A(n7225), .B(o[255]), .Z(creg_next[255]) );
  AND U8250 ( .A(n3090), .B(n7226), .Z(n7225) );
  XNOR U8251 ( .A(c[255]), .B(n7227), .Z(n7226) );
  IV U8252 ( .A(o[255]), .Z(n7227) );
  XNOR U8253 ( .A(n7228), .B(n7229), .Z(o[255]) );
  XOR U8254 ( .A(n7230), .B(o[254]), .Z(creg_next[254]) );
  AND U8255 ( .A(n3090), .B(n7231), .Z(n7230) );
  XNOR U8256 ( .A(c[254]), .B(n7232), .Z(n7231) );
  IV U8257 ( .A(o[254]), .Z(n7232) );
  XNOR U8258 ( .A(n7233), .B(n7234), .Z(o[254]) );
  XOR U8259 ( .A(n7235), .B(o[253]), .Z(creg_next[253]) );
  AND U8260 ( .A(n3090), .B(n7236), .Z(n7235) );
  XNOR U8261 ( .A(c[253]), .B(n7237), .Z(n7236) );
  IV U8262 ( .A(o[253]), .Z(n7237) );
  XNOR U8263 ( .A(n7238), .B(n7239), .Z(o[253]) );
  XOR U8264 ( .A(n7240), .B(o[252]), .Z(creg_next[252]) );
  AND U8265 ( .A(n3090), .B(n7241), .Z(n7240) );
  XNOR U8266 ( .A(c[252]), .B(n7242), .Z(n7241) );
  IV U8267 ( .A(o[252]), .Z(n7242) );
  XNOR U8268 ( .A(n7243), .B(n7244), .Z(o[252]) );
  XOR U8269 ( .A(n7245), .B(o[251]), .Z(creg_next[251]) );
  AND U8270 ( .A(n3090), .B(n7246), .Z(n7245) );
  XNOR U8271 ( .A(c[251]), .B(n7247), .Z(n7246) );
  IV U8272 ( .A(o[251]), .Z(n7247) );
  XNOR U8273 ( .A(n7248), .B(n7249), .Z(o[251]) );
  XOR U8274 ( .A(n7250), .B(o[250]), .Z(creg_next[250]) );
  AND U8275 ( .A(n3090), .B(n7251), .Z(n7250) );
  XNOR U8276 ( .A(c[250]), .B(n7252), .Z(n7251) );
  IV U8277 ( .A(o[250]), .Z(n7252) );
  XNOR U8278 ( .A(n7253), .B(n7254), .Z(o[250]) );
  XOR U8279 ( .A(n7255), .B(o[24]), .Z(creg_next[24]) );
  AND U8280 ( .A(n3090), .B(n7256), .Z(n7255) );
  XNOR U8281 ( .A(c[24]), .B(n7257), .Z(n7256) );
  IV U8282 ( .A(o[24]), .Z(n7257) );
  XNOR U8283 ( .A(n7258), .B(n7259), .Z(o[24]) );
  XOR U8284 ( .A(n7260), .B(o[249]), .Z(creg_next[249]) );
  AND U8285 ( .A(n3090), .B(n7261), .Z(n7260) );
  XNOR U8286 ( .A(c[249]), .B(n7262), .Z(n7261) );
  IV U8287 ( .A(o[249]), .Z(n7262) );
  XNOR U8288 ( .A(n7263), .B(n7264), .Z(o[249]) );
  XOR U8289 ( .A(n7265), .B(o[248]), .Z(creg_next[248]) );
  AND U8290 ( .A(n3090), .B(n7266), .Z(n7265) );
  XNOR U8291 ( .A(c[248]), .B(n7267), .Z(n7266) );
  IV U8292 ( .A(o[248]), .Z(n7267) );
  XNOR U8293 ( .A(n7268), .B(n7269), .Z(o[248]) );
  XOR U8294 ( .A(n7270), .B(o[247]), .Z(creg_next[247]) );
  AND U8295 ( .A(n3090), .B(n7271), .Z(n7270) );
  XNOR U8296 ( .A(c[247]), .B(n7272), .Z(n7271) );
  IV U8297 ( .A(o[247]), .Z(n7272) );
  XNOR U8298 ( .A(n7273), .B(n7274), .Z(o[247]) );
  XOR U8299 ( .A(n7275), .B(o[246]), .Z(creg_next[246]) );
  AND U8300 ( .A(n3090), .B(n7276), .Z(n7275) );
  XNOR U8301 ( .A(c[246]), .B(n7277), .Z(n7276) );
  IV U8302 ( .A(o[246]), .Z(n7277) );
  XNOR U8303 ( .A(n7278), .B(n7279), .Z(o[246]) );
  XOR U8304 ( .A(n7280), .B(o[245]), .Z(creg_next[245]) );
  AND U8305 ( .A(n3090), .B(n7281), .Z(n7280) );
  XNOR U8306 ( .A(c[245]), .B(n7282), .Z(n7281) );
  IV U8307 ( .A(o[245]), .Z(n7282) );
  XNOR U8308 ( .A(n7283), .B(n7284), .Z(o[245]) );
  XOR U8309 ( .A(n7285), .B(o[244]), .Z(creg_next[244]) );
  AND U8310 ( .A(n3090), .B(n7286), .Z(n7285) );
  XNOR U8311 ( .A(c[244]), .B(n7287), .Z(n7286) );
  IV U8312 ( .A(o[244]), .Z(n7287) );
  XNOR U8313 ( .A(n7288), .B(n7289), .Z(o[244]) );
  XOR U8314 ( .A(n7290), .B(o[243]), .Z(creg_next[243]) );
  AND U8315 ( .A(n3090), .B(n7291), .Z(n7290) );
  XNOR U8316 ( .A(c[243]), .B(n7292), .Z(n7291) );
  IV U8317 ( .A(o[243]), .Z(n7292) );
  XNOR U8318 ( .A(n7293), .B(n7294), .Z(o[243]) );
  XOR U8319 ( .A(n7295), .B(o[242]), .Z(creg_next[242]) );
  AND U8320 ( .A(n3090), .B(n7296), .Z(n7295) );
  XNOR U8321 ( .A(c[242]), .B(n7297), .Z(n7296) );
  IV U8322 ( .A(o[242]), .Z(n7297) );
  XNOR U8323 ( .A(n7298), .B(n7299), .Z(o[242]) );
  XOR U8324 ( .A(n7300), .B(o[241]), .Z(creg_next[241]) );
  AND U8325 ( .A(n3090), .B(n7301), .Z(n7300) );
  XNOR U8326 ( .A(c[241]), .B(n7302), .Z(n7301) );
  IV U8327 ( .A(o[241]), .Z(n7302) );
  XNOR U8328 ( .A(n7303), .B(n7304), .Z(o[241]) );
  XOR U8329 ( .A(n7305), .B(o[240]), .Z(creg_next[240]) );
  AND U8330 ( .A(n3090), .B(n7306), .Z(n7305) );
  XNOR U8331 ( .A(c[240]), .B(n7307), .Z(n7306) );
  IV U8332 ( .A(o[240]), .Z(n7307) );
  XNOR U8333 ( .A(n7308), .B(n7309), .Z(o[240]) );
  XOR U8334 ( .A(n7310), .B(o[23]), .Z(creg_next[23]) );
  AND U8335 ( .A(n3090), .B(n7311), .Z(n7310) );
  XNOR U8336 ( .A(c[23]), .B(n7312), .Z(n7311) );
  IV U8337 ( .A(o[23]), .Z(n7312) );
  XNOR U8338 ( .A(n7313), .B(n7314), .Z(o[23]) );
  XOR U8339 ( .A(n7315), .B(o[239]), .Z(creg_next[239]) );
  AND U8340 ( .A(n3090), .B(n7316), .Z(n7315) );
  XNOR U8341 ( .A(c[239]), .B(n7317), .Z(n7316) );
  IV U8342 ( .A(o[239]), .Z(n7317) );
  XNOR U8343 ( .A(n7318), .B(n7319), .Z(o[239]) );
  XOR U8344 ( .A(n7320), .B(o[238]), .Z(creg_next[238]) );
  AND U8345 ( .A(n3090), .B(n7321), .Z(n7320) );
  XNOR U8346 ( .A(c[238]), .B(n7322), .Z(n7321) );
  IV U8347 ( .A(o[238]), .Z(n7322) );
  XNOR U8348 ( .A(n7323), .B(n7324), .Z(o[238]) );
  XOR U8349 ( .A(n7325), .B(o[237]), .Z(creg_next[237]) );
  AND U8350 ( .A(n3090), .B(n7326), .Z(n7325) );
  XNOR U8351 ( .A(c[237]), .B(n7327), .Z(n7326) );
  IV U8352 ( .A(o[237]), .Z(n7327) );
  XNOR U8353 ( .A(n7328), .B(n7329), .Z(o[237]) );
  XOR U8354 ( .A(n7330), .B(o[236]), .Z(creg_next[236]) );
  AND U8355 ( .A(n3090), .B(n7331), .Z(n7330) );
  XNOR U8356 ( .A(c[236]), .B(n7332), .Z(n7331) );
  IV U8357 ( .A(o[236]), .Z(n7332) );
  XNOR U8358 ( .A(n7333), .B(n7334), .Z(o[236]) );
  XOR U8359 ( .A(n7335), .B(o[235]), .Z(creg_next[235]) );
  AND U8360 ( .A(n3090), .B(n7336), .Z(n7335) );
  XNOR U8361 ( .A(c[235]), .B(n7337), .Z(n7336) );
  IV U8362 ( .A(o[235]), .Z(n7337) );
  XNOR U8363 ( .A(n7338), .B(n7339), .Z(o[235]) );
  XOR U8364 ( .A(n7340), .B(o[234]), .Z(creg_next[234]) );
  AND U8365 ( .A(n3090), .B(n7341), .Z(n7340) );
  XNOR U8366 ( .A(c[234]), .B(n7342), .Z(n7341) );
  IV U8367 ( .A(o[234]), .Z(n7342) );
  XNOR U8368 ( .A(n7343), .B(n7344), .Z(o[234]) );
  XOR U8369 ( .A(n7345), .B(o[233]), .Z(creg_next[233]) );
  AND U8370 ( .A(n3090), .B(n7346), .Z(n7345) );
  XNOR U8371 ( .A(c[233]), .B(n7347), .Z(n7346) );
  IV U8372 ( .A(o[233]), .Z(n7347) );
  XNOR U8373 ( .A(n7348), .B(n7349), .Z(o[233]) );
  XOR U8374 ( .A(n7350), .B(o[232]), .Z(creg_next[232]) );
  AND U8375 ( .A(n3090), .B(n7351), .Z(n7350) );
  XNOR U8376 ( .A(c[232]), .B(n7352), .Z(n7351) );
  IV U8377 ( .A(o[232]), .Z(n7352) );
  XNOR U8378 ( .A(n7353), .B(n7354), .Z(o[232]) );
  XOR U8379 ( .A(n7355), .B(o[231]), .Z(creg_next[231]) );
  AND U8380 ( .A(n3090), .B(n7356), .Z(n7355) );
  XNOR U8381 ( .A(c[231]), .B(n7357), .Z(n7356) );
  IV U8382 ( .A(o[231]), .Z(n7357) );
  XNOR U8383 ( .A(n7358), .B(n7359), .Z(o[231]) );
  XOR U8384 ( .A(n7360), .B(o[230]), .Z(creg_next[230]) );
  AND U8385 ( .A(n3090), .B(n7361), .Z(n7360) );
  XNOR U8386 ( .A(c[230]), .B(n7362), .Z(n7361) );
  IV U8387 ( .A(o[230]), .Z(n7362) );
  XNOR U8388 ( .A(n7363), .B(n7364), .Z(o[230]) );
  XOR U8389 ( .A(n7365), .B(o[22]), .Z(creg_next[22]) );
  AND U8390 ( .A(n3090), .B(n7366), .Z(n7365) );
  XNOR U8391 ( .A(c[22]), .B(n7367), .Z(n7366) );
  IV U8392 ( .A(o[22]), .Z(n7367) );
  XNOR U8393 ( .A(n7368), .B(n7369), .Z(o[22]) );
  XOR U8394 ( .A(n7370), .B(o[229]), .Z(creg_next[229]) );
  AND U8395 ( .A(n3090), .B(n7371), .Z(n7370) );
  XNOR U8396 ( .A(c[229]), .B(n7372), .Z(n7371) );
  IV U8397 ( .A(o[229]), .Z(n7372) );
  XNOR U8398 ( .A(n7373), .B(n7374), .Z(o[229]) );
  XOR U8399 ( .A(n7375), .B(o[228]), .Z(creg_next[228]) );
  AND U8400 ( .A(n3090), .B(n7376), .Z(n7375) );
  XNOR U8401 ( .A(c[228]), .B(n7377), .Z(n7376) );
  IV U8402 ( .A(o[228]), .Z(n7377) );
  XNOR U8403 ( .A(n7378), .B(n7379), .Z(o[228]) );
  XOR U8404 ( .A(n7380), .B(o[227]), .Z(creg_next[227]) );
  AND U8405 ( .A(n3090), .B(n7381), .Z(n7380) );
  XNOR U8406 ( .A(c[227]), .B(n7382), .Z(n7381) );
  IV U8407 ( .A(o[227]), .Z(n7382) );
  XNOR U8408 ( .A(n7383), .B(n7384), .Z(o[227]) );
  XOR U8409 ( .A(n7385), .B(o[226]), .Z(creg_next[226]) );
  AND U8410 ( .A(n3090), .B(n7386), .Z(n7385) );
  XNOR U8411 ( .A(c[226]), .B(n7387), .Z(n7386) );
  IV U8412 ( .A(o[226]), .Z(n7387) );
  XNOR U8413 ( .A(n7388), .B(n7389), .Z(o[226]) );
  XOR U8414 ( .A(n7390), .B(o[225]), .Z(creg_next[225]) );
  AND U8415 ( .A(n3090), .B(n7391), .Z(n7390) );
  XNOR U8416 ( .A(c[225]), .B(n7392), .Z(n7391) );
  IV U8417 ( .A(o[225]), .Z(n7392) );
  XNOR U8418 ( .A(n7393), .B(n7394), .Z(o[225]) );
  XOR U8419 ( .A(n7395), .B(o[224]), .Z(creg_next[224]) );
  AND U8420 ( .A(n3090), .B(n7396), .Z(n7395) );
  XNOR U8421 ( .A(c[224]), .B(n7397), .Z(n7396) );
  IV U8422 ( .A(o[224]), .Z(n7397) );
  XNOR U8423 ( .A(n7398), .B(n7399), .Z(o[224]) );
  XOR U8424 ( .A(n7400), .B(o[223]), .Z(creg_next[223]) );
  AND U8425 ( .A(n3090), .B(n7401), .Z(n7400) );
  XNOR U8426 ( .A(c[223]), .B(n7402), .Z(n7401) );
  IV U8427 ( .A(o[223]), .Z(n7402) );
  XNOR U8428 ( .A(n7403), .B(n7404), .Z(o[223]) );
  XOR U8429 ( .A(n7405), .B(o[222]), .Z(creg_next[222]) );
  AND U8430 ( .A(n3090), .B(n7406), .Z(n7405) );
  XNOR U8431 ( .A(c[222]), .B(n7407), .Z(n7406) );
  IV U8432 ( .A(o[222]), .Z(n7407) );
  XNOR U8433 ( .A(n7408), .B(n7409), .Z(o[222]) );
  XOR U8434 ( .A(n7410), .B(o[221]), .Z(creg_next[221]) );
  AND U8435 ( .A(n3090), .B(n7411), .Z(n7410) );
  XNOR U8436 ( .A(c[221]), .B(n7412), .Z(n7411) );
  IV U8437 ( .A(o[221]), .Z(n7412) );
  XNOR U8438 ( .A(n7413), .B(n7414), .Z(o[221]) );
  XOR U8439 ( .A(n7415), .B(o[220]), .Z(creg_next[220]) );
  AND U8440 ( .A(n3090), .B(n7416), .Z(n7415) );
  XNOR U8441 ( .A(c[220]), .B(n7417), .Z(n7416) );
  IV U8442 ( .A(o[220]), .Z(n7417) );
  XNOR U8443 ( .A(n7418), .B(n7419), .Z(o[220]) );
  XOR U8444 ( .A(n7420), .B(o[21]), .Z(creg_next[21]) );
  AND U8445 ( .A(n3090), .B(n7421), .Z(n7420) );
  XNOR U8446 ( .A(c[21]), .B(n7422), .Z(n7421) );
  IV U8447 ( .A(o[21]), .Z(n7422) );
  XNOR U8448 ( .A(n7423), .B(n7424), .Z(o[21]) );
  XOR U8449 ( .A(n7425), .B(o[219]), .Z(creg_next[219]) );
  AND U8450 ( .A(n3090), .B(n7426), .Z(n7425) );
  XNOR U8451 ( .A(c[219]), .B(n7427), .Z(n7426) );
  IV U8452 ( .A(o[219]), .Z(n7427) );
  XNOR U8453 ( .A(n7428), .B(n7429), .Z(o[219]) );
  XOR U8454 ( .A(n7430), .B(o[218]), .Z(creg_next[218]) );
  AND U8455 ( .A(n3090), .B(n7431), .Z(n7430) );
  XNOR U8456 ( .A(c[218]), .B(n7432), .Z(n7431) );
  IV U8457 ( .A(o[218]), .Z(n7432) );
  XNOR U8458 ( .A(n7433), .B(n7434), .Z(o[218]) );
  XOR U8459 ( .A(n7435), .B(o[217]), .Z(creg_next[217]) );
  AND U8460 ( .A(n3090), .B(n7436), .Z(n7435) );
  XNOR U8461 ( .A(c[217]), .B(n7437), .Z(n7436) );
  IV U8462 ( .A(o[217]), .Z(n7437) );
  XNOR U8463 ( .A(n7438), .B(n7439), .Z(o[217]) );
  XOR U8464 ( .A(n7440), .B(o[216]), .Z(creg_next[216]) );
  AND U8465 ( .A(n3090), .B(n7441), .Z(n7440) );
  XNOR U8466 ( .A(c[216]), .B(n7442), .Z(n7441) );
  IV U8467 ( .A(o[216]), .Z(n7442) );
  XNOR U8468 ( .A(n7443), .B(n7444), .Z(o[216]) );
  XOR U8469 ( .A(n7445), .B(o[215]), .Z(creg_next[215]) );
  AND U8470 ( .A(n3090), .B(n7446), .Z(n7445) );
  XNOR U8471 ( .A(c[215]), .B(n7447), .Z(n7446) );
  IV U8472 ( .A(o[215]), .Z(n7447) );
  XNOR U8473 ( .A(n7448), .B(n7449), .Z(o[215]) );
  XOR U8474 ( .A(n7450), .B(o[214]), .Z(creg_next[214]) );
  AND U8475 ( .A(n3090), .B(n7451), .Z(n7450) );
  XNOR U8476 ( .A(c[214]), .B(n7452), .Z(n7451) );
  IV U8477 ( .A(o[214]), .Z(n7452) );
  XNOR U8478 ( .A(n7453), .B(n7454), .Z(o[214]) );
  XOR U8479 ( .A(n7455), .B(o[213]), .Z(creg_next[213]) );
  AND U8480 ( .A(n3090), .B(n7456), .Z(n7455) );
  XNOR U8481 ( .A(c[213]), .B(n7457), .Z(n7456) );
  IV U8482 ( .A(o[213]), .Z(n7457) );
  XNOR U8483 ( .A(n7458), .B(n7459), .Z(o[213]) );
  XOR U8484 ( .A(n7460), .B(o[212]), .Z(creg_next[212]) );
  AND U8485 ( .A(n3090), .B(n7461), .Z(n7460) );
  XNOR U8486 ( .A(c[212]), .B(n7462), .Z(n7461) );
  IV U8487 ( .A(o[212]), .Z(n7462) );
  XNOR U8488 ( .A(n7463), .B(n7464), .Z(o[212]) );
  XOR U8489 ( .A(n7465), .B(o[211]), .Z(creg_next[211]) );
  AND U8490 ( .A(n3090), .B(n7466), .Z(n7465) );
  XNOR U8491 ( .A(c[211]), .B(n7467), .Z(n7466) );
  IV U8492 ( .A(o[211]), .Z(n7467) );
  XNOR U8493 ( .A(n7468), .B(n7469), .Z(o[211]) );
  XOR U8494 ( .A(n7470), .B(o[210]), .Z(creg_next[210]) );
  AND U8495 ( .A(n3090), .B(n7471), .Z(n7470) );
  XNOR U8496 ( .A(c[210]), .B(n7472), .Z(n7471) );
  IV U8497 ( .A(o[210]), .Z(n7472) );
  XNOR U8498 ( .A(n7473), .B(n7474), .Z(o[210]) );
  XOR U8499 ( .A(n7475), .B(o[20]), .Z(creg_next[20]) );
  AND U8500 ( .A(n3090), .B(n7476), .Z(n7475) );
  XNOR U8501 ( .A(c[20]), .B(n7477), .Z(n7476) );
  IV U8502 ( .A(o[20]), .Z(n7477) );
  XNOR U8503 ( .A(n7478), .B(n7479), .Z(o[20]) );
  XOR U8504 ( .A(n7480), .B(o[209]), .Z(creg_next[209]) );
  AND U8505 ( .A(n3090), .B(n7481), .Z(n7480) );
  XNOR U8506 ( .A(c[209]), .B(n7482), .Z(n7481) );
  IV U8507 ( .A(o[209]), .Z(n7482) );
  XNOR U8508 ( .A(n7483), .B(n7484), .Z(o[209]) );
  XOR U8509 ( .A(n7485), .B(o[208]), .Z(creg_next[208]) );
  AND U8510 ( .A(n3090), .B(n7486), .Z(n7485) );
  XNOR U8511 ( .A(c[208]), .B(n7487), .Z(n7486) );
  IV U8512 ( .A(o[208]), .Z(n7487) );
  XNOR U8513 ( .A(n7488), .B(n7489), .Z(o[208]) );
  XOR U8514 ( .A(n7490), .B(o[207]), .Z(creg_next[207]) );
  AND U8515 ( .A(n3090), .B(n7491), .Z(n7490) );
  XNOR U8516 ( .A(c[207]), .B(n7492), .Z(n7491) );
  IV U8517 ( .A(o[207]), .Z(n7492) );
  XNOR U8518 ( .A(n7493), .B(n7494), .Z(o[207]) );
  XOR U8519 ( .A(n7495), .B(o[206]), .Z(creg_next[206]) );
  AND U8520 ( .A(n3090), .B(n7496), .Z(n7495) );
  XNOR U8521 ( .A(c[206]), .B(n7497), .Z(n7496) );
  IV U8522 ( .A(o[206]), .Z(n7497) );
  XNOR U8523 ( .A(n7498), .B(n7499), .Z(o[206]) );
  XOR U8524 ( .A(n7500), .B(o[205]), .Z(creg_next[205]) );
  AND U8525 ( .A(n3090), .B(n7501), .Z(n7500) );
  XNOR U8526 ( .A(c[205]), .B(n7502), .Z(n7501) );
  IV U8527 ( .A(o[205]), .Z(n7502) );
  XNOR U8528 ( .A(n7503), .B(n7504), .Z(o[205]) );
  XOR U8529 ( .A(n7505), .B(o[204]), .Z(creg_next[204]) );
  AND U8530 ( .A(n3090), .B(n7506), .Z(n7505) );
  XNOR U8531 ( .A(c[204]), .B(n7507), .Z(n7506) );
  IV U8532 ( .A(o[204]), .Z(n7507) );
  XNOR U8533 ( .A(n7508), .B(n7509), .Z(o[204]) );
  XOR U8534 ( .A(n7510), .B(o[203]), .Z(creg_next[203]) );
  AND U8535 ( .A(n3090), .B(n7511), .Z(n7510) );
  XNOR U8536 ( .A(c[203]), .B(n7512), .Z(n7511) );
  IV U8537 ( .A(o[203]), .Z(n7512) );
  XNOR U8538 ( .A(n7513), .B(n7514), .Z(o[203]) );
  XOR U8539 ( .A(n7515), .B(o[202]), .Z(creg_next[202]) );
  AND U8540 ( .A(n3090), .B(n7516), .Z(n7515) );
  XNOR U8541 ( .A(c[202]), .B(n7517), .Z(n7516) );
  IV U8542 ( .A(o[202]), .Z(n7517) );
  XNOR U8543 ( .A(n7518), .B(n7519), .Z(o[202]) );
  XOR U8544 ( .A(n7520), .B(o[201]), .Z(creg_next[201]) );
  AND U8545 ( .A(n3090), .B(n7521), .Z(n7520) );
  XNOR U8546 ( .A(c[201]), .B(n7522), .Z(n7521) );
  IV U8547 ( .A(o[201]), .Z(n7522) );
  XNOR U8548 ( .A(n7523), .B(n7524), .Z(o[201]) );
  XOR U8549 ( .A(n7525), .B(o[200]), .Z(creg_next[200]) );
  AND U8550 ( .A(n3090), .B(n7526), .Z(n7525) );
  XNOR U8551 ( .A(c[200]), .B(n7527), .Z(n7526) );
  IV U8552 ( .A(o[200]), .Z(n7527) );
  XNOR U8553 ( .A(n7528), .B(n7529), .Z(o[200]) );
  XOR U8554 ( .A(n7530), .B(o[1]), .Z(creg_next[1]) );
  AND U8555 ( .A(n3090), .B(n7531), .Z(n7530) );
  XNOR U8556 ( .A(c[1]), .B(n7532), .Z(n7531) );
  IV U8557 ( .A(o[1]), .Z(n7532) );
  XNOR U8558 ( .A(n7533), .B(n7534), .Z(o[1]) );
  XOR U8559 ( .A(n7535), .B(o[19]), .Z(creg_next[19]) );
  AND U8560 ( .A(n3090), .B(n7536), .Z(n7535) );
  XNOR U8561 ( .A(c[19]), .B(n7537), .Z(n7536) );
  IV U8562 ( .A(o[19]), .Z(n7537) );
  XNOR U8563 ( .A(n7538), .B(n7539), .Z(o[19]) );
  XOR U8564 ( .A(n7540), .B(o[199]), .Z(creg_next[199]) );
  AND U8565 ( .A(n3090), .B(n7541), .Z(n7540) );
  XNOR U8566 ( .A(c[199]), .B(n7542), .Z(n7541) );
  IV U8567 ( .A(o[199]), .Z(n7542) );
  XNOR U8568 ( .A(n7543), .B(n7544), .Z(o[199]) );
  XOR U8569 ( .A(n7545), .B(o[198]), .Z(creg_next[198]) );
  AND U8570 ( .A(n3090), .B(n7546), .Z(n7545) );
  XNOR U8571 ( .A(c[198]), .B(n7547), .Z(n7546) );
  IV U8572 ( .A(o[198]), .Z(n7547) );
  XNOR U8573 ( .A(n7548), .B(n7549), .Z(o[198]) );
  XOR U8574 ( .A(n7550), .B(o[197]), .Z(creg_next[197]) );
  AND U8575 ( .A(n3090), .B(n7551), .Z(n7550) );
  XNOR U8576 ( .A(c[197]), .B(n7552), .Z(n7551) );
  IV U8577 ( .A(o[197]), .Z(n7552) );
  XNOR U8578 ( .A(n7553), .B(n7554), .Z(o[197]) );
  XOR U8579 ( .A(n7555), .B(o[196]), .Z(creg_next[196]) );
  AND U8580 ( .A(n3090), .B(n7556), .Z(n7555) );
  XNOR U8581 ( .A(c[196]), .B(n7557), .Z(n7556) );
  IV U8582 ( .A(o[196]), .Z(n7557) );
  XNOR U8583 ( .A(n7558), .B(n7559), .Z(o[196]) );
  XOR U8584 ( .A(n7560), .B(o[195]), .Z(creg_next[195]) );
  AND U8585 ( .A(n3090), .B(n7561), .Z(n7560) );
  XNOR U8586 ( .A(c[195]), .B(n7562), .Z(n7561) );
  IV U8587 ( .A(o[195]), .Z(n7562) );
  XNOR U8588 ( .A(n7563), .B(n7564), .Z(o[195]) );
  XOR U8589 ( .A(n7565), .B(o[194]), .Z(creg_next[194]) );
  AND U8590 ( .A(n3090), .B(n7566), .Z(n7565) );
  XNOR U8591 ( .A(c[194]), .B(n7567), .Z(n7566) );
  IV U8592 ( .A(o[194]), .Z(n7567) );
  XNOR U8593 ( .A(n7568), .B(n7569), .Z(o[194]) );
  XOR U8594 ( .A(n7570), .B(o[193]), .Z(creg_next[193]) );
  AND U8595 ( .A(n3090), .B(n7571), .Z(n7570) );
  XNOR U8596 ( .A(c[193]), .B(n7572), .Z(n7571) );
  IV U8597 ( .A(o[193]), .Z(n7572) );
  XNOR U8598 ( .A(n7573), .B(n7574), .Z(o[193]) );
  XOR U8599 ( .A(n7575), .B(o[192]), .Z(creg_next[192]) );
  AND U8600 ( .A(n3090), .B(n7576), .Z(n7575) );
  XNOR U8601 ( .A(c[192]), .B(n7577), .Z(n7576) );
  IV U8602 ( .A(o[192]), .Z(n7577) );
  XNOR U8603 ( .A(n7578), .B(n7579), .Z(o[192]) );
  XOR U8604 ( .A(n7580), .B(o[191]), .Z(creg_next[191]) );
  AND U8605 ( .A(n3090), .B(n7581), .Z(n7580) );
  XNOR U8606 ( .A(c[191]), .B(n7582), .Z(n7581) );
  IV U8607 ( .A(o[191]), .Z(n7582) );
  XNOR U8608 ( .A(n7583), .B(n7584), .Z(o[191]) );
  XOR U8609 ( .A(n7585), .B(o[190]), .Z(creg_next[190]) );
  AND U8610 ( .A(n3090), .B(n7586), .Z(n7585) );
  XNOR U8611 ( .A(c[190]), .B(n7587), .Z(n7586) );
  IV U8612 ( .A(o[190]), .Z(n7587) );
  XNOR U8613 ( .A(n7588), .B(n7589), .Z(o[190]) );
  XOR U8614 ( .A(n7590), .B(o[18]), .Z(creg_next[18]) );
  AND U8615 ( .A(n3090), .B(n7591), .Z(n7590) );
  XNOR U8616 ( .A(c[18]), .B(n7592), .Z(n7591) );
  IV U8617 ( .A(o[18]), .Z(n7592) );
  XNOR U8618 ( .A(n7593), .B(n7594), .Z(o[18]) );
  XOR U8619 ( .A(n7595), .B(o[189]), .Z(creg_next[189]) );
  AND U8620 ( .A(n3090), .B(n7596), .Z(n7595) );
  XNOR U8621 ( .A(c[189]), .B(n7597), .Z(n7596) );
  IV U8622 ( .A(o[189]), .Z(n7597) );
  XNOR U8623 ( .A(n7598), .B(n7599), .Z(o[189]) );
  XOR U8624 ( .A(n7600), .B(o[188]), .Z(creg_next[188]) );
  AND U8625 ( .A(n3090), .B(n7601), .Z(n7600) );
  XNOR U8626 ( .A(c[188]), .B(n7602), .Z(n7601) );
  IV U8627 ( .A(o[188]), .Z(n7602) );
  XNOR U8628 ( .A(n7603), .B(n7604), .Z(o[188]) );
  XOR U8629 ( .A(n7605), .B(o[187]), .Z(creg_next[187]) );
  AND U8630 ( .A(n3090), .B(n7606), .Z(n7605) );
  XNOR U8631 ( .A(c[187]), .B(n7607), .Z(n7606) );
  IV U8632 ( .A(o[187]), .Z(n7607) );
  XNOR U8633 ( .A(n7608), .B(n7609), .Z(o[187]) );
  XOR U8634 ( .A(n7610), .B(o[186]), .Z(creg_next[186]) );
  AND U8635 ( .A(n3090), .B(n7611), .Z(n7610) );
  XNOR U8636 ( .A(c[186]), .B(n7612), .Z(n7611) );
  IV U8637 ( .A(o[186]), .Z(n7612) );
  XNOR U8638 ( .A(n7613), .B(n7614), .Z(o[186]) );
  XOR U8639 ( .A(n7615), .B(o[185]), .Z(creg_next[185]) );
  AND U8640 ( .A(n3090), .B(n7616), .Z(n7615) );
  XNOR U8641 ( .A(c[185]), .B(n7617), .Z(n7616) );
  IV U8642 ( .A(o[185]), .Z(n7617) );
  XNOR U8643 ( .A(n7618), .B(n7619), .Z(o[185]) );
  XOR U8644 ( .A(n7620), .B(o[184]), .Z(creg_next[184]) );
  AND U8645 ( .A(n3090), .B(n7621), .Z(n7620) );
  XNOR U8646 ( .A(c[184]), .B(n7622), .Z(n7621) );
  IV U8647 ( .A(o[184]), .Z(n7622) );
  XNOR U8648 ( .A(n7623), .B(n7624), .Z(o[184]) );
  XOR U8649 ( .A(n7625), .B(o[183]), .Z(creg_next[183]) );
  AND U8650 ( .A(n3090), .B(n7626), .Z(n7625) );
  XNOR U8651 ( .A(c[183]), .B(n7627), .Z(n7626) );
  IV U8652 ( .A(o[183]), .Z(n7627) );
  XNOR U8653 ( .A(n7628), .B(n7629), .Z(o[183]) );
  XOR U8654 ( .A(n7630), .B(o[182]), .Z(creg_next[182]) );
  AND U8655 ( .A(n3090), .B(n7631), .Z(n7630) );
  XNOR U8656 ( .A(c[182]), .B(n7632), .Z(n7631) );
  IV U8657 ( .A(o[182]), .Z(n7632) );
  XNOR U8658 ( .A(n7633), .B(n7634), .Z(o[182]) );
  XOR U8659 ( .A(n7635), .B(o[181]), .Z(creg_next[181]) );
  AND U8660 ( .A(n3090), .B(n7636), .Z(n7635) );
  XNOR U8661 ( .A(c[181]), .B(n7637), .Z(n7636) );
  IV U8662 ( .A(o[181]), .Z(n7637) );
  XNOR U8663 ( .A(n7638), .B(n7639), .Z(o[181]) );
  XOR U8664 ( .A(n7640), .B(o[180]), .Z(creg_next[180]) );
  AND U8665 ( .A(n3090), .B(n7641), .Z(n7640) );
  XNOR U8666 ( .A(c[180]), .B(n7642), .Z(n7641) );
  IV U8667 ( .A(o[180]), .Z(n7642) );
  XNOR U8668 ( .A(n7643), .B(n7644), .Z(o[180]) );
  XOR U8669 ( .A(n7645), .B(o[17]), .Z(creg_next[17]) );
  AND U8670 ( .A(n3090), .B(n7646), .Z(n7645) );
  XNOR U8671 ( .A(c[17]), .B(n7647), .Z(n7646) );
  IV U8672 ( .A(o[17]), .Z(n7647) );
  XNOR U8673 ( .A(n7648), .B(n7649), .Z(o[17]) );
  XOR U8674 ( .A(n7650), .B(o[179]), .Z(creg_next[179]) );
  AND U8675 ( .A(n3090), .B(n7651), .Z(n7650) );
  XNOR U8676 ( .A(c[179]), .B(n7652), .Z(n7651) );
  IV U8677 ( .A(o[179]), .Z(n7652) );
  XNOR U8678 ( .A(n7653), .B(n7654), .Z(o[179]) );
  XOR U8679 ( .A(n7655), .B(o[178]), .Z(creg_next[178]) );
  AND U8680 ( .A(n3090), .B(n7656), .Z(n7655) );
  XNOR U8681 ( .A(c[178]), .B(n7657), .Z(n7656) );
  IV U8682 ( .A(o[178]), .Z(n7657) );
  XNOR U8683 ( .A(n7658), .B(n7659), .Z(o[178]) );
  XOR U8684 ( .A(n7660), .B(o[177]), .Z(creg_next[177]) );
  AND U8685 ( .A(n3090), .B(n7661), .Z(n7660) );
  XNOR U8686 ( .A(c[177]), .B(n7662), .Z(n7661) );
  IV U8687 ( .A(o[177]), .Z(n7662) );
  XNOR U8688 ( .A(n7663), .B(n7664), .Z(o[177]) );
  XOR U8689 ( .A(n7665), .B(o[176]), .Z(creg_next[176]) );
  AND U8690 ( .A(n3090), .B(n7666), .Z(n7665) );
  XNOR U8691 ( .A(c[176]), .B(n7667), .Z(n7666) );
  IV U8692 ( .A(o[176]), .Z(n7667) );
  XNOR U8693 ( .A(n7668), .B(n7669), .Z(o[176]) );
  XOR U8694 ( .A(n7670), .B(o[175]), .Z(creg_next[175]) );
  AND U8695 ( .A(n3090), .B(n7671), .Z(n7670) );
  XNOR U8696 ( .A(c[175]), .B(n7672), .Z(n7671) );
  IV U8697 ( .A(o[175]), .Z(n7672) );
  XNOR U8698 ( .A(n7673), .B(n7674), .Z(o[175]) );
  XOR U8699 ( .A(n7675), .B(o[174]), .Z(creg_next[174]) );
  AND U8700 ( .A(n3090), .B(n7676), .Z(n7675) );
  XNOR U8701 ( .A(c[174]), .B(n7677), .Z(n7676) );
  IV U8702 ( .A(o[174]), .Z(n7677) );
  XNOR U8703 ( .A(n7678), .B(n7679), .Z(o[174]) );
  XOR U8704 ( .A(n7680), .B(o[173]), .Z(creg_next[173]) );
  AND U8705 ( .A(n3090), .B(n7681), .Z(n7680) );
  XNOR U8706 ( .A(c[173]), .B(n7682), .Z(n7681) );
  IV U8707 ( .A(o[173]), .Z(n7682) );
  XNOR U8708 ( .A(n7683), .B(n7684), .Z(o[173]) );
  XOR U8709 ( .A(n7685), .B(o[172]), .Z(creg_next[172]) );
  AND U8710 ( .A(n3090), .B(n7686), .Z(n7685) );
  XNOR U8711 ( .A(c[172]), .B(n7687), .Z(n7686) );
  IV U8712 ( .A(o[172]), .Z(n7687) );
  XNOR U8713 ( .A(n7688), .B(n7689), .Z(o[172]) );
  XOR U8714 ( .A(n7690), .B(o[171]), .Z(creg_next[171]) );
  AND U8715 ( .A(n3090), .B(n7691), .Z(n7690) );
  XNOR U8716 ( .A(c[171]), .B(n7692), .Z(n7691) );
  IV U8717 ( .A(o[171]), .Z(n7692) );
  XNOR U8718 ( .A(n7693), .B(n7694), .Z(o[171]) );
  XOR U8719 ( .A(n7695), .B(o[170]), .Z(creg_next[170]) );
  AND U8720 ( .A(n3090), .B(n7696), .Z(n7695) );
  XNOR U8721 ( .A(c[170]), .B(n7697), .Z(n7696) );
  IV U8722 ( .A(o[170]), .Z(n7697) );
  XNOR U8723 ( .A(n7698), .B(n7699), .Z(o[170]) );
  XOR U8724 ( .A(n7700), .B(o[16]), .Z(creg_next[16]) );
  AND U8725 ( .A(n3090), .B(n7701), .Z(n7700) );
  XNOR U8726 ( .A(c[16]), .B(n7702), .Z(n7701) );
  IV U8727 ( .A(o[16]), .Z(n7702) );
  XNOR U8728 ( .A(n7703), .B(n7704), .Z(o[16]) );
  XOR U8729 ( .A(n7705), .B(o[169]), .Z(creg_next[169]) );
  AND U8730 ( .A(n3090), .B(n7706), .Z(n7705) );
  XNOR U8731 ( .A(c[169]), .B(n7707), .Z(n7706) );
  IV U8732 ( .A(o[169]), .Z(n7707) );
  XNOR U8733 ( .A(n7708), .B(n7709), .Z(o[169]) );
  XOR U8734 ( .A(n7710), .B(o[168]), .Z(creg_next[168]) );
  AND U8735 ( .A(n3090), .B(n7711), .Z(n7710) );
  XNOR U8736 ( .A(c[168]), .B(n7712), .Z(n7711) );
  IV U8737 ( .A(o[168]), .Z(n7712) );
  XNOR U8738 ( .A(n7713), .B(n7714), .Z(o[168]) );
  XOR U8739 ( .A(n7715), .B(o[167]), .Z(creg_next[167]) );
  AND U8740 ( .A(n3090), .B(n7716), .Z(n7715) );
  XNOR U8741 ( .A(c[167]), .B(n7717), .Z(n7716) );
  IV U8742 ( .A(o[167]), .Z(n7717) );
  XNOR U8743 ( .A(n7718), .B(n7719), .Z(o[167]) );
  XOR U8744 ( .A(n7720), .B(o[166]), .Z(creg_next[166]) );
  AND U8745 ( .A(n3090), .B(n7721), .Z(n7720) );
  XNOR U8746 ( .A(c[166]), .B(n7722), .Z(n7721) );
  IV U8747 ( .A(o[166]), .Z(n7722) );
  XNOR U8748 ( .A(n7723), .B(n7724), .Z(o[166]) );
  XOR U8749 ( .A(n7725), .B(o[165]), .Z(creg_next[165]) );
  AND U8750 ( .A(n3090), .B(n7726), .Z(n7725) );
  XNOR U8751 ( .A(c[165]), .B(n7727), .Z(n7726) );
  IV U8752 ( .A(o[165]), .Z(n7727) );
  XNOR U8753 ( .A(n7728), .B(n7729), .Z(o[165]) );
  XOR U8754 ( .A(n7730), .B(o[164]), .Z(creg_next[164]) );
  AND U8755 ( .A(n3090), .B(n7731), .Z(n7730) );
  XNOR U8756 ( .A(c[164]), .B(n7732), .Z(n7731) );
  IV U8757 ( .A(o[164]), .Z(n7732) );
  XNOR U8758 ( .A(n7733), .B(n7734), .Z(o[164]) );
  XOR U8759 ( .A(n7735), .B(o[163]), .Z(creg_next[163]) );
  AND U8760 ( .A(n3090), .B(n7736), .Z(n7735) );
  XNOR U8761 ( .A(c[163]), .B(n7737), .Z(n7736) );
  IV U8762 ( .A(o[163]), .Z(n7737) );
  XNOR U8763 ( .A(n7738), .B(n7739), .Z(o[163]) );
  XOR U8764 ( .A(n7740), .B(o[162]), .Z(creg_next[162]) );
  AND U8765 ( .A(n3090), .B(n7741), .Z(n7740) );
  XNOR U8766 ( .A(c[162]), .B(n7742), .Z(n7741) );
  IV U8767 ( .A(o[162]), .Z(n7742) );
  XNOR U8768 ( .A(n7743), .B(n7744), .Z(o[162]) );
  XOR U8769 ( .A(n7745), .B(o[161]), .Z(creg_next[161]) );
  AND U8770 ( .A(n3090), .B(n7746), .Z(n7745) );
  XNOR U8771 ( .A(c[161]), .B(n7747), .Z(n7746) );
  IV U8772 ( .A(o[161]), .Z(n7747) );
  XNOR U8773 ( .A(n7748), .B(n7749), .Z(o[161]) );
  XOR U8774 ( .A(n7750), .B(o[160]), .Z(creg_next[160]) );
  AND U8775 ( .A(n3090), .B(n7751), .Z(n7750) );
  XNOR U8776 ( .A(c[160]), .B(n7752), .Z(n7751) );
  IV U8777 ( .A(o[160]), .Z(n7752) );
  XNOR U8778 ( .A(n7753), .B(n7754), .Z(o[160]) );
  XOR U8779 ( .A(n7755), .B(o[15]), .Z(creg_next[15]) );
  AND U8780 ( .A(n3090), .B(n7756), .Z(n7755) );
  XNOR U8781 ( .A(c[15]), .B(n7757), .Z(n7756) );
  IV U8782 ( .A(o[15]), .Z(n7757) );
  XNOR U8783 ( .A(n7758), .B(n7759), .Z(o[15]) );
  XOR U8784 ( .A(n7760), .B(o[159]), .Z(creg_next[159]) );
  AND U8785 ( .A(n3090), .B(n7761), .Z(n7760) );
  XNOR U8786 ( .A(c[159]), .B(n7762), .Z(n7761) );
  IV U8787 ( .A(o[159]), .Z(n7762) );
  XNOR U8788 ( .A(n7763), .B(n7764), .Z(o[159]) );
  XOR U8789 ( .A(n7765), .B(o[158]), .Z(creg_next[158]) );
  AND U8790 ( .A(n3090), .B(n7766), .Z(n7765) );
  XNOR U8791 ( .A(c[158]), .B(n7767), .Z(n7766) );
  IV U8792 ( .A(o[158]), .Z(n7767) );
  XNOR U8793 ( .A(n7768), .B(n7769), .Z(o[158]) );
  XOR U8794 ( .A(n7770), .B(o[157]), .Z(creg_next[157]) );
  AND U8795 ( .A(n3090), .B(n7771), .Z(n7770) );
  XNOR U8796 ( .A(c[157]), .B(n7772), .Z(n7771) );
  IV U8797 ( .A(o[157]), .Z(n7772) );
  XNOR U8798 ( .A(n7773), .B(n7774), .Z(o[157]) );
  XOR U8799 ( .A(n7775), .B(o[156]), .Z(creg_next[156]) );
  AND U8800 ( .A(n3090), .B(n7776), .Z(n7775) );
  XNOR U8801 ( .A(c[156]), .B(n7777), .Z(n7776) );
  IV U8802 ( .A(o[156]), .Z(n7777) );
  XNOR U8803 ( .A(n7778), .B(n7779), .Z(o[156]) );
  XOR U8804 ( .A(n7780), .B(o[155]), .Z(creg_next[155]) );
  AND U8805 ( .A(n3090), .B(n7781), .Z(n7780) );
  XNOR U8806 ( .A(c[155]), .B(n7782), .Z(n7781) );
  IV U8807 ( .A(o[155]), .Z(n7782) );
  XNOR U8808 ( .A(n7783), .B(n7784), .Z(o[155]) );
  XOR U8809 ( .A(n7785), .B(o[154]), .Z(creg_next[154]) );
  AND U8810 ( .A(n3090), .B(n7786), .Z(n7785) );
  XNOR U8811 ( .A(c[154]), .B(n7787), .Z(n7786) );
  IV U8812 ( .A(o[154]), .Z(n7787) );
  XNOR U8813 ( .A(n7788), .B(n7789), .Z(o[154]) );
  XOR U8814 ( .A(n7790), .B(o[153]), .Z(creg_next[153]) );
  AND U8815 ( .A(n3090), .B(n7791), .Z(n7790) );
  XNOR U8816 ( .A(c[153]), .B(n7792), .Z(n7791) );
  IV U8817 ( .A(o[153]), .Z(n7792) );
  XNOR U8818 ( .A(n7793), .B(n7794), .Z(o[153]) );
  XOR U8819 ( .A(n7795), .B(o[152]), .Z(creg_next[152]) );
  AND U8820 ( .A(n3090), .B(n7796), .Z(n7795) );
  XNOR U8821 ( .A(c[152]), .B(n7797), .Z(n7796) );
  IV U8822 ( .A(o[152]), .Z(n7797) );
  XNOR U8823 ( .A(n7798), .B(n7799), .Z(o[152]) );
  XOR U8824 ( .A(n7800), .B(o[151]), .Z(creg_next[151]) );
  AND U8825 ( .A(n3090), .B(n7801), .Z(n7800) );
  XNOR U8826 ( .A(c[151]), .B(n7802), .Z(n7801) );
  IV U8827 ( .A(o[151]), .Z(n7802) );
  XNOR U8828 ( .A(n7803), .B(n7804), .Z(o[151]) );
  XOR U8829 ( .A(n7805), .B(o[150]), .Z(creg_next[150]) );
  AND U8830 ( .A(n3090), .B(n7806), .Z(n7805) );
  XNOR U8831 ( .A(c[150]), .B(n7807), .Z(n7806) );
  IV U8832 ( .A(o[150]), .Z(n7807) );
  XNOR U8833 ( .A(n7808), .B(n7809), .Z(o[150]) );
  XOR U8834 ( .A(n7810), .B(o[14]), .Z(creg_next[14]) );
  AND U8835 ( .A(n3090), .B(n7811), .Z(n7810) );
  XNOR U8836 ( .A(c[14]), .B(n7812), .Z(n7811) );
  IV U8837 ( .A(o[14]), .Z(n7812) );
  XNOR U8838 ( .A(n7813), .B(n7814), .Z(o[14]) );
  XOR U8839 ( .A(n7815), .B(o[149]), .Z(creg_next[149]) );
  AND U8840 ( .A(n3090), .B(n7816), .Z(n7815) );
  XNOR U8841 ( .A(c[149]), .B(n7817), .Z(n7816) );
  IV U8842 ( .A(o[149]), .Z(n7817) );
  XNOR U8843 ( .A(n7818), .B(n7819), .Z(o[149]) );
  XOR U8844 ( .A(n7820), .B(o[148]), .Z(creg_next[148]) );
  AND U8845 ( .A(n3090), .B(n7821), .Z(n7820) );
  XNOR U8846 ( .A(c[148]), .B(n7822), .Z(n7821) );
  IV U8847 ( .A(o[148]), .Z(n7822) );
  XNOR U8848 ( .A(n7823), .B(n7824), .Z(o[148]) );
  XOR U8849 ( .A(n7825), .B(o[147]), .Z(creg_next[147]) );
  AND U8850 ( .A(n3090), .B(n7826), .Z(n7825) );
  XNOR U8851 ( .A(c[147]), .B(n7827), .Z(n7826) );
  IV U8852 ( .A(o[147]), .Z(n7827) );
  XNOR U8853 ( .A(n7828), .B(n7829), .Z(o[147]) );
  XOR U8854 ( .A(n7830), .B(o[146]), .Z(creg_next[146]) );
  AND U8855 ( .A(n3090), .B(n7831), .Z(n7830) );
  XNOR U8856 ( .A(c[146]), .B(n7832), .Z(n7831) );
  IV U8857 ( .A(o[146]), .Z(n7832) );
  XNOR U8858 ( .A(n7833), .B(n7834), .Z(o[146]) );
  XOR U8859 ( .A(n7835), .B(o[145]), .Z(creg_next[145]) );
  AND U8860 ( .A(n3090), .B(n7836), .Z(n7835) );
  XNOR U8861 ( .A(c[145]), .B(n7837), .Z(n7836) );
  IV U8862 ( .A(o[145]), .Z(n7837) );
  XNOR U8863 ( .A(n7838), .B(n7839), .Z(o[145]) );
  XOR U8864 ( .A(n7840), .B(o[144]), .Z(creg_next[144]) );
  AND U8865 ( .A(n3090), .B(n7841), .Z(n7840) );
  XNOR U8866 ( .A(c[144]), .B(n7842), .Z(n7841) );
  IV U8867 ( .A(o[144]), .Z(n7842) );
  XNOR U8868 ( .A(n7843), .B(n7844), .Z(o[144]) );
  XOR U8869 ( .A(n7845), .B(o[143]), .Z(creg_next[143]) );
  AND U8870 ( .A(n3090), .B(n7846), .Z(n7845) );
  XNOR U8871 ( .A(c[143]), .B(n7847), .Z(n7846) );
  IV U8872 ( .A(o[143]), .Z(n7847) );
  XNOR U8873 ( .A(n7848), .B(n7849), .Z(o[143]) );
  XOR U8874 ( .A(n7850), .B(o[142]), .Z(creg_next[142]) );
  AND U8875 ( .A(n3090), .B(n7851), .Z(n7850) );
  XNOR U8876 ( .A(c[142]), .B(n7852), .Z(n7851) );
  IV U8877 ( .A(o[142]), .Z(n7852) );
  XNOR U8878 ( .A(n7853), .B(n7854), .Z(o[142]) );
  XOR U8879 ( .A(n7855), .B(o[141]), .Z(creg_next[141]) );
  AND U8880 ( .A(n3090), .B(n7856), .Z(n7855) );
  XNOR U8881 ( .A(c[141]), .B(n7857), .Z(n7856) );
  IV U8882 ( .A(o[141]), .Z(n7857) );
  XNOR U8883 ( .A(n7858), .B(n7859), .Z(o[141]) );
  XOR U8884 ( .A(n7860), .B(o[140]), .Z(creg_next[140]) );
  AND U8885 ( .A(n3090), .B(n7861), .Z(n7860) );
  XNOR U8886 ( .A(c[140]), .B(n7862), .Z(n7861) );
  IV U8887 ( .A(o[140]), .Z(n7862) );
  XNOR U8888 ( .A(n7863), .B(n7864), .Z(o[140]) );
  XOR U8889 ( .A(n7865), .B(o[13]), .Z(creg_next[13]) );
  AND U8890 ( .A(n3090), .B(n7866), .Z(n7865) );
  XNOR U8891 ( .A(c[13]), .B(n7867), .Z(n7866) );
  IV U8892 ( .A(o[13]), .Z(n7867) );
  XNOR U8893 ( .A(n7868), .B(n7869), .Z(o[13]) );
  XOR U8894 ( .A(n7870), .B(o[139]), .Z(creg_next[139]) );
  AND U8895 ( .A(n3090), .B(n7871), .Z(n7870) );
  XNOR U8896 ( .A(c[139]), .B(n7872), .Z(n7871) );
  IV U8897 ( .A(o[139]), .Z(n7872) );
  XNOR U8898 ( .A(n7873), .B(n7874), .Z(o[139]) );
  XOR U8899 ( .A(n7875), .B(o[138]), .Z(creg_next[138]) );
  AND U8900 ( .A(n3090), .B(n7876), .Z(n7875) );
  XNOR U8901 ( .A(c[138]), .B(n7877), .Z(n7876) );
  IV U8902 ( .A(o[138]), .Z(n7877) );
  XNOR U8903 ( .A(n7878), .B(n7879), .Z(o[138]) );
  XOR U8904 ( .A(n7880), .B(o[137]), .Z(creg_next[137]) );
  AND U8905 ( .A(n3090), .B(n7881), .Z(n7880) );
  XNOR U8906 ( .A(c[137]), .B(n7882), .Z(n7881) );
  IV U8907 ( .A(o[137]), .Z(n7882) );
  XNOR U8908 ( .A(n7883), .B(n7884), .Z(o[137]) );
  XOR U8909 ( .A(n7885), .B(o[136]), .Z(creg_next[136]) );
  AND U8910 ( .A(n3090), .B(n7886), .Z(n7885) );
  XNOR U8911 ( .A(c[136]), .B(n7887), .Z(n7886) );
  IV U8912 ( .A(o[136]), .Z(n7887) );
  XNOR U8913 ( .A(n7888), .B(n7889), .Z(o[136]) );
  XOR U8914 ( .A(n7890), .B(o[135]), .Z(creg_next[135]) );
  AND U8915 ( .A(n3090), .B(n7891), .Z(n7890) );
  XNOR U8916 ( .A(c[135]), .B(n7892), .Z(n7891) );
  IV U8917 ( .A(o[135]), .Z(n7892) );
  XNOR U8918 ( .A(n7893), .B(n7894), .Z(o[135]) );
  XOR U8919 ( .A(n7895), .B(o[134]), .Z(creg_next[134]) );
  AND U8920 ( .A(n3090), .B(n7896), .Z(n7895) );
  XNOR U8921 ( .A(c[134]), .B(n7897), .Z(n7896) );
  IV U8922 ( .A(o[134]), .Z(n7897) );
  XNOR U8923 ( .A(n7898), .B(n7899), .Z(o[134]) );
  XOR U8924 ( .A(n7900), .B(o[133]), .Z(creg_next[133]) );
  AND U8925 ( .A(n3090), .B(n7901), .Z(n7900) );
  XNOR U8926 ( .A(c[133]), .B(n7902), .Z(n7901) );
  IV U8927 ( .A(o[133]), .Z(n7902) );
  XNOR U8928 ( .A(n7903), .B(n7904), .Z(o[133]) );
  XOR U8929 ( .A(n7905), .B(o[132]), .Z(creg_next[132]) );
  AND U8930 ( .A(n3090), .B(n7906), .Z(n7905) );
  XNOR U8931 ( .A(c[132]), .B(n7907), .Z(n7906) );
  IV U8932 ( .A(o[132]), .Z(n7907) );
  XNOR U8933 ( .A(n7908), .B(n7909), .Z(o[132]) );
  XOR U8934 ( .A(n7910), .B(o[131]), .Z(creg_next[131]) );
  AND U8935 ( .A(n3090), .B(n7911), .Z(n7910) );
  XNOR U8936 ( .A(c[131]), .B(n7912), .Z(n7911) );
  IV U8937 ( .A(o[131]), .Z(n7912) );
  XNOR U8938 ( .A(n7913), .B(n7914), .Z(o[131]) );
  XOR U8939 ( .A(n7915), .B(o[130]), .Z(creg_next[130]) );
  AND U8940 ( .A(n3090), .B(n7916), .Z(n7915) );
  XNOR U8941 ( .A(c[130]), .B(n7917), .Z(n7916) );
  IV U8942 ( .A(o[130]), .Z(n7917) );
  XNOR U8943 ( .A(n7918), .B(n7919), .Z(o[130]) );
  XOR U8944 ( .A(n7920), .B(o[12]), .Z(creg_next[12]) );
  AND U8945 ( .A(n3090), .B(n7921), .Z(n7920) );
  XNOR U8946 ( .A(c[12]), .B(n7922), .Z(n7921) );
  IV U8947 ( .A(o[12]), .Z(n7922) );
  XNOR U8948 ( .A(n7923), .B(n7924), .Z(o[12]) );
  XOR U8949 ( .A(n7925), .B(o[129]), .Z(creg_next[129]) );
  AND U8950 ( .A(n3090), .B(n7926), .Z(n7925) );
  XNOR U8951 ( .A(c[129]), .B(n7927), .Z(n7926) );
  IV U8952 ( .A(o[129]), .Z(n7927) );
  XNOR U8953 ( .A(n7928), .B(n7929), .Z(o[129]) );
  XOR U8954 ( .A(n7930), .B(o[128]), .Z(creg_next[128]) );
  AND U8955 ( .A(n3090), .B(n7931), .Z(n7930) );
  XNOR U8956 ( .A(c[128]), .B(n7932), .Z(n7931) );
  IV U8957 ( .A(o[128]), .Z(n7932) );
  XNOR U8958 ( .A(n7933), .B(n7934), .Z(o[128]) );
  XOR U8959 ( .A(n7935), .B(o[127]), .Z(creg_next[127]) );
  AND U8960 ( .A(n3090), .B(n7936), .Z(n7935) );
  XNOR U8961 ( .A(c[127]), .B(n7937), .Z(n7936) );
  IV U8962 ( .A(o[127]), .Z(n7937) );
  XNOR U8963 ( .A(n7938), .B(n7939), .Z(o[127]) );
  XOR U8964 ( .A(n7940), .B(o[126]), .Z(creg_next[126]) );
  AND U8965 ( .A(n3090), .B(n7941), .Z(n7940) );
  XNOR U8966 ( .A(c[126]), .B(n7942), .Z(n7941) );
  IV U8967 ( .A(o[126]), .Z(n7942) );
  XNOR U8968 ( .A(n7943), .B(n7944), .Z(o[126]) );
  XOR U8969 ( .A(n7945), .B(o[125]), .Z(creg_next[125]) );
  AND U8970 ( .A(n3090), .B(n7946), .Z(n7945) );
  XNOR U8971 ( .A(c[125]), .B(n7947), .Z(n7946) );
  IV U8972 ( .A(o[125]), .Z(n7947) );
  XNOR U8973 ( .A(n7948), .B(n7949), .Z(o[125]) );
  XOR U8974 ( .A(n7950), .B(o[124]), .Z(creg_next[124]) );
  AND U8975 ( .A(n3090), .B(n7951), .Z(n7950) );
  XNOR U8976 ( .A(c[124]), .B(n7952), .Z(n7951) );
  IV U8977 ( .A(o[124]), .Z(n7952) );
  XNOR U8978 ( .A(n7953), .B(n7954), .Z(o[124]) );
  XOR U8979 ( .A(n7955), .B(o[123]), .Z(creg_next[123]) );
  AND U8980 ( .A(n3090), .B(n7956), .Z(n7955) );
  XNOR U8981 ( .A(c[123]), .B(n7957), .Z(n7956) );
  IV U8982 ( .A(o[123]), .Z(n7957) );
  XNOR U8983 ( .A(n7958), .B(n7959), .Z(o[123]) );
  XOR U8984 ( .A(n7960), .B(o[122]), .Z(creg_next[122]) );
  AND U8985 ( .A(n3090), .B(n7961), .Z(n7960) );
  XNOR U8986 ( .A(c[122]), .B(n7962), .Z(n7961) );
  IV U8987 ( .A(o[122]), .Z(n7962) );
  XNOR U8988 ( .A(n7963), .B(n7964), .Z(o[122]) );
  XOR U8989 ( .A(n7965), .B(o[121]), .Z(creg_next[121]) );
  AND U8990 ( .A(n3090), .B(n7966), .Z(n7965) );
  XNOR U8991 ( .A(c[121]), .B(n7967), .Z(n7966) );
  IV U8992 ( .A(o[121]), .Z(n7967) );
  XNOR U8993 ( .A(n7968), .B(n7969), .Z(o[121]) );
  XOR U8994 ( .A(n7970), .B(o[120]), .Z(creg_next[120]) );
  AND U8995 ( .A(n3090), .B(n7971), .Z(n7970) );
  XNOR U8996 ( .A(c[120]), .B(n7972), .Z(n7971) );
  IV U8997 ( .A(o[120]), .Z(n7972) );
  XNOR U8998 ( .A(n7973), .B(n7974), .Z(o[120]) );
  XOR U8999 ( .A(n7975), .B(o[11]), .Z(creg_next[11]) );
  AND U9000 ( .A(n3090), .B(n7976), .Z(n7975) );
  XNOR U9001 ( .A(c[11]), .B(n7977), .Z(n7976) );
  IV U9002 ( .A(o[11]), .Z(n7977) );
  XNOR U9003 ( .A(n7978), .B(n7979), .Z(o[11]) );
  XOR U9004 ( .A(n7980), .B(o[119]), .Z(creg_next[119]) );
  AND U9005 ( .A(n3090), .B(n7981), .Z(n7980) );
  XNOR U9006 ( .A(c[119]), .B(n7982), .Z(n7981) );
  IV U9007 ( .A(o[119]), .Z(n7982) );
  XNOR U9008 ( .A(n7983), .B(n7984), .Z(o[119]) );
  XOR U9009 ( .A(n7985), .B(o[118]), .Z(creg_next[118]) );
  AND U9010 ( .A(n3090), .B(n7986), .Z(n7985) );
  XNOR U9011 ( .A(c[118]), .B(n7987), .Z(n7986) );
  IV U9012 ( .A(o[118]), .Z(n7987) );
  XNOR U9013 ( .A(n7988), .B(n7989), .Z(o[118]) );
  XOR U9014 ( .A(n7990), .B(o[117]), .Z(creg_next[117]) );
  AND U9015 ( .A(n3090), .B(n7991), .Z(n7990) );
  XNOR U9016 ( .A(c[117]), .B(n7992), .Z(n7991) );
  IV U9017 ( .A(o[117]), .Z(n7992) );
  XNOR U9018 ( .A(n7993), .B(n7994), .Z(o[117]) );
  XOR U9019 ( .A(n7995), .B(o[116]), .Z(creg_next[116]) );
  AND U9020 ( .A(n3090), .B(n7996), .Z(n7995) );
  XNOR U9021 ( .A(c[116]), .B(n7997), .Z(n7996) );
  IV U9022 ( .A(o[116]), .Z(n7997) );
  XNOR U9023 ( .A(n7998), .B(n7999), .Z(o[116]) );
  XOR U9024 ( .A(n8000), .B(o[115]), .Z(creg_next[115]) );
  AND U9025 ( .A(n3090), .B(n8001), .Z(n8000) );
  XNOR U9026 ( .A(c[115]), .B(n8002), .Z(n8001) );
  IV U9027 ( .A(o[115]), .Z(n8002) );
  XNOR U9028 ( .A(n8003), .B(n8004), .Z(o[115]) );
  XOR U9029 ( .A(n8005), .B(o[114]), .Z(creg_next[114]) );
  AND U9030 ( .A(n3090), .B(n8006), .Z(n8005) );
  XNOR U9031 ( .A(c[114]), .B(n8007), .Z(n8006) );
  IV U9032 ( .A(o[114]), .Z(n8007) );
  XNOR U9033 ( .A(n8008), .B(n8009), .Z(o[114]) );
  XOR U9034 ( .A(n8010), .B(o[113]), .Z(creg_next[113]) );
  AND U9035 ( .A(n3090), .B(n8011), .Z(n8010) );
  XNOR U9036 ( .A(c[113]), .B(n8012), .Z(n8011) );
  IV U9037 ( .A(o[113]), .Z(n8012) );
  XNOR U9038 ( .A(n8013), .B(n8014), .Z(o[113]) );
  XOR U9039 ( .A(n8015), .B(o[112]), .Z(creg_next[112]) );
  AND U9040 ( .A(n3090), .B(n8016), .Z(n8015) );
  XNOR U9041 ( .A(c[112]), .B(n8017), .Z(n8016) );
  IV U9042 ( .A(o[112]), .Z(n8017) );
  XNOR U9043 ( .A(n8018), .B(n8019), .Z(o[112]) );
  XOR U9044 ( .A(n8020), .B(o[111]), .Z(creg_next[111]) );
  AND U9045 ( .A(n3090), .B(n8021), .Z(n8020) );
  XNOR U9046 ( .A(c[111]), .B(n8022), .Z(n8021) );
  IV U9047 ( .A(o[111]), .Z(n8022) );
  XNOR U9048 ( .A(n8023), .B(n8024), .Z(o[111]) );
  XOR U9049 ( .A(n8025), .B(o[110]), .Z(creg_next[110]) );
  AND U9050 ( .A(n3090), .B(n8026), .Z(n8025) );
  XNOR U9051 ( .A(c[110]), .B(n8027), .Z(n8026) );
  IV U9052 ( .A(o[110]), .Z(n8027) );
  XNOR U9053 ( .A(n8028), .B(n8029), .Z(o[110]) );
  XOR U9054 ( .A(n8030), .B(o[10]), .Z(creg_next[10]) );
  AND U9055 ( .A(n3090), .B(n8031), .Z(n8030) );
  XNOR U9056 ( .A(c[10]), .B(n8032), .Z(n8031) );
  IV U9057 ( .A(o[10]), .Z(n8032) );
  XNOR U9058 ( .A(n8033), .B(n8034), .Z(o[10]) );
  XOR U9059 ( .A(n8035), .B(o[109]), .Z(creg_next[109]) );
  AND U9060 ( .A(n3090), .B(n8036), .Z(n8035) );
  XNOR U9061 ( .A(c[109]), .B(n8037), .Z(n8036) );
  IV U9062 ( .A(o[109]), .Z(n8037) );
  XNOR U9063 ( .A(n8038), .B(n8039), .Z(o[109]) );
  XOR U9064 ( .A(n8040), .B(o[108]), .Z(creg_next[108]) );
  AND U9065 ( .A(n3090), .B(n8041), .Z(n8040) );
  XNOR U9066 ( .A(c[108]), .B(n8042), .Z(n8041) );
  IV U9067 ( .A(o[108]), .Z(n8042) );
  XNOR U9068 ( .A(n8043), .B(n8044), .Z(o[108]) );
  XOR U9069 ( .A(n8045), .B(o[107]), .Z(creg_next[107]) );
  AND U9070 ( .A(n3090), .B(n8046), .Z(n8045) );
  XNOR U9071 ( .A(c[107]), .B(n8047), .Z(n8046) );
  IV U9072 ( .A(o[107]), .Z(n8047) );
  XNOR U9073 ( .A(n8048), .B(n8049), .Z(o[107]) );
  XOR U9074 ( .A(n8050), .B(o[106]), .Z(creg_next[106]) );
  AND U9075 ( .A(n3090), .B(n8051), .Z(n8050) );
  XNOR U9076 ( .A(c[106]), .B(n8052), .Z(n8051) );
  IV U9077 ( .A(o[106]), .Z(n8052) );
  XNOR U9078 ( .A(n8053), .B(n8054), .Z(o[106]) );
  XOR U9079 ( .A(n8055), .B(o[105]), .Z(creg_next[105]) );
  AND U9080 ( .A(n3090), .B(n8056), .Z(n8055) );
  XNOR U9081 ( .A(c[105]), .B(n8057), .Z(n8056) );
  IV U9082 ( .A(o[105]), .Z(n8057) );
  XNOR U9083 ( .A(n8058), .B(n8059), .Z(o[105]) );
  XOR U9084 ( .A(n8060), .B(o[104]), .Z(creg_next[104]) );
  AND U9085 ( .A(n3090), .B(n8061), .Z(n8060) );
  XNOR U9086 ( .A(c[104]), .B(n8062), .Z(n8061) );
  IV U9087 ( .A(o[104]), .Z(n8062) );
  XNOR U9088 ( .A(n8063), .B(n8064), .Z(o[104]) );
  XOR U9089 ( .A(n8065), .B(o[103]), .Z(creg_next[103]) );
  AND U9090 ( .A(n3090), .B(n8066), .Z(n8065) );
  XNOR U9091 ( .A(c[103]), .B(n8067), .Z(n8066) );
  IV U9092 ( .A(o[103]), .Z(n8067) );
  XNOR U9093 ( .A(n8068), .B(n8069), .Z(o[103]) );
  XOR U9094 ( .A(n8070), .B(o[102]), .Z(creg_next[102]) );
  AND U9095 ( .A(n3090), .B(n8071), .Z(n8070) );
  XNOR U9096 ( .A(c[102]), .B(n8072), .Z(n8071) );
  IV U9097 ( .A(o[102]), .Z(n8072) );
  XNOR U9098 ( .A(n8073), .B(n8074), .Z(o[102]) );
  XOR U9099 ( .A(n8075), .B(o[1023]), .Z(creg_next[1023]) );
  AND U9100 ( .A(n3090), .B(n8076), .Z(n8075) );
  XNOR U9101 ( .A(c[1023]), .B(n8077), .Z(n8076) );
  IV U9102 ( .A(o[1023]), .Z(n8077) );
  XNOR U9103 ( .A(n1041), .B(n1040), .Z(o[1023]) );
  XNOR U9104 ( .A(n8078), .B(n1035), .Z(n1040) );
  IV U9105 ( .A(n1042), .Z(n1035) );
  XOR U9106 ( .A(n8079), .B(n8080), .Z(n1042) );
  ANDN U9107 ( .B(n8081), .A(n8082), .Z(n8079) );
  XOR U9108 ( .A(n8083), .B(n8080), .Z(n8081) );
  NAND U9109 ( .A(n8084), .B(n[1023]), .Z(n1041) );
  NAND U9110 ( .A(n8085), .B(n[1023]), .Z(n8084) );
  XOR U9111 ( .A(n8086), .B(o[1022]), .Z(creg_next[1022]) );
  AND U9112 ( .A(n3090), .B(n8087), .Z(n8086) );
  XNOR U9113 ( .A(c[1022]), .B(n8088), .Z(n8087) );
  IV U9114 ( .A(o[1022]), .Z(n8088) );
  XNOR U9115 ( .A(n8083), .B(n8082), .Z(o[1022]) );
  XNOR U9116 ( .A(n8089), .B(n8090), .Z(n8082) );
  IV U9117 ( .A(n8080), .Z(n8090) );
  XOR U9118 ( .A(n8091), .B(n8092), .Z(n8080) );
  ANDN U9119 ( .B(n8093), .A(n8094), .Z(n8091) );
  XOR U9120 ( .A(n8095), .B(n8092), .Z(n8093) );
  NAND U9121 ( .A(n8096), .B(n[1022]), .Z(n8083) );
  NAND U9122 ( .A(n8085), .B(n[1022]), .Z(n8096) );
  XOR U9123 ( .A(n8097), .B(o[1021]), .Z(creg_next[1021]) );
  AND U9124 ( .A(n3090), .B(n8098), .Z(n8097) );
  XNOR U9125 ( .A(c[1021]), .B(n8099), .Z(n8098) );
  IV U9126 ( .A(o[1021]), .Z(n8099) );
  XNOR U9127 ( .A(n8095), .B(n8094), .Z(o[1021]) );
  XNOR U9128 ( .A(n8100), .B(n8101), .Z(n8094) );
  IV U9129 ( .A(n8092), .Z(n8101) );
  XOR U9130 ( .A(n8102), .B(n8103), .Z(n8092) );
  ANDN U9131 ( .B(n8104), .A(n8105), .Z(n8102) );
  XOR U9132 ( .A(n8106), .B(n8103), .Z(n8104) );
  NAND U9133 ( .A(n8107), .B(n[1021]), .Z(n8095) );
  NAND U9134 ( .A(n8085), .B(n[1021]), .Z(n8107) );
  XOR U9135 ( .A(n8108), .B(o[1020]), .Z(creg_next[1020]) );
  AND U9136 ( .A(n3090), .B(n8109), .Z(n8108) );
  XNOR U9137 ( .A(c[1020]), .B(n8110), .Z(n8109) );
  IV U9138 ( .A(o[1020]), .Z(n8110) );
  XNOR U9139 ( .A(n8106), .B(n8105), .Z(o[1020]) );
  XNOR U9140 ( .A(n8111), .B(n8112), .Z(n8105) );
  IV U9141 ( .A(n8103), .Z(n8112) );
  XOR U9142 ( .A(n8113), .B(n8114), .Z(n8103) );
  ANDN U9143 ( .B(n8115), .A(n8116), .Z(n8113) );
  XOR U9144 ( .A(n8117), .B(n8114), .Z(n8115) );
  NAND U9145 ( .A(n8118), .B(n[1020]), .Z(n8106) );
  NAND U9146 ( .A(n8085), .B(n[1020]), .Z(n8118) );
  XOR U9147 ( .A(n8119), .B(o[101]), .Z(creg_next[101]) );
  AND U9148 ( .A(n3090), .B(n8120), .Z(n8119) );
  XNOR U9149 ( .A(c[101]), .B(n8121), .Z(n8120) );
  IV U9150 ( .A(o[101]), .Z(n8121) );
  XNOR U9151 ( .A(n8122), .B(n8123), .Z(o[101]) );
  XOR U9152 ( .A(n8124), .B(o[1019]), .Z(creg_next[1019]) );
  AND U9153 ( .A(n3090), .B(n8125), .Z(n8124) );
  XNOR U9154 ( .A(c[1019]), .B(n8126), .Z(n8125) );
  IV U9155 ( .A(o[1019]), .Z(n8126) );
  XNOR U9156 ( .A(n8117), .B(n8116), .Z(o[1019]) );
  XNOR U9157 ( .A(n8127), .B(n8128), .Z(n8116) );
  IV U9158 ( .A(n8114), .Z(n8128) );
  XOR U9159 ( .A(n8129), .B(n8130), .Z(n8114) );
  ANDN U9160 ( .B(n8131), .A(n8132), .Z(n8129) );
  XOR U9161 ( .A(n8133), .B(n8130), .Z(n8131) );
  NAND U9162 ( .A(n8134), .B(n[1019]), .Z(n8117) );
  NAND U9163 ( .A(n8085), .B(n[1019]), .Z(n8134) );
  XOR U9164 ( .A(n8135), .B(o[1018]), .Z(creg_next[1018]) );
  AND U9165 ( .A(n3090), .B(n8136), .Z(n8135) );
  XNOR U9166 ( .A(c[1018]), .B(n8137), .Z(n8136) );
  IV U9167 ( .A(o[1018]), .Z(n8137) );
  XNOR U9168 ( .A(n8133), .B(n8132), .Z(o[1018]) );
  XNOR U9169 ( .A(n8138), .B(n8139), .Z(n8132) );
  IV U9170 ( .A(n8130), .Z(n8139) );
  XOR U9171 ( .A(n8140), .B(n8141), .Z(n8130) );
  ANDN U9172 ( .B(n8142), .A(n8143), .Z(n8140) );
  XOR U9173 ( .A(n8144), .B(n8141), .Z(n8142) );
  NAND U9174 ( .A(n8145), .B(n[1018]), .Z(n8133) );
  NAND U9175 ( .A(n8085), .B(n[1018]), .Z(n8145) );
  XOR U9176 ( .A(n8146), .B(o[1017]), .Z(creg_next[1017]) );
  AND U9177 ( .A(n3090), .B(n8147), .Z(n8146) );
  XNOR U9178 ( .A(c[1017]), .B(n8148), .Z(n8147) );
  IV U9179 ( .A(o[1017]), .Z(n8148) );
  XNOR U9180 ( .A(n8144), .B(n8143), .Z(o[1017]) );
  XNOR U9181 ( .A(n8149), .B(n8150), .Z(n8143) );
  IV U9182 ( .A(n8141), .Z(n8150) );
  XOR U9183 ( .A(n8151), .B(n8152), .Z(n8141) );
  ANDN U9184 ( .B(n8153), .A(n8154), .Z(n8151) );
  XOR U9185 ( .A(n8155), .B(n8152), .Z(n8153) );
  NAND U9186 ( .A(n8156), .B(n[1017]), .Z(n8144) );
  NAND U9187 ( .A(n8085), .B(n[1017]), .Z(n8156) );
  XOR U9188 ( .A(n8157), .B(o[1016]), .Z(creg_next[1016]) );
  AND U9189 ( .A(n3090), .B(n8158), .Z(n8157) );
  XNOR U9190 ( .A(c[1016]), .B(n8159), .Z(n8158) );
  IV U9191 ( .A(o[1016]), .Z(n8159) );
  XNOR U9192 ( .A(n8155), .B(n8154), .Z(o[1016]) );
  XNOR U9193 ( .A(n8160), .B(n8161), .Z(n8154) );
  IV U9194 ( .A(n8152), .Z(n8161) );
  XOR U9195 ( .A(n8162), .B(n8163), .Z(n8152) );
  ANDN U9196 ( .B(n8164), .A(n8165), .Z(n8162) );
  XOR U9197 ( .A(n8166), .B(n8163), .Z(n8164) );
  NAND U9198 ( .A(n8167), .B(n[1016]), .Z(n8155) );
  NAND U9199 ( .A(n8085), .B(n[1016]), .Z(n8167) );
  XOR U9200 ( .A(n8168), .B(o[1015]), .Z(creg_next[1015]) );
  AND U9201 ( .A(n3090), .B(n8169), .Z(n8168) );
  XNOR U9202 ( .A(c[1015]), .B(n8170), .Z(n8169) );
  IV U9203 ( .A(o[1015]), .Z(n8170) );
  XNOR U9204 ( .A(n8166), .B(n8165), .Z(o[1015]) );
  XNOR U9205 ( .A(n8171), .B(n8172), .Z(n8165) );
  IV U9206 ( .A(n8163), .Z(n8172) );
  XOR U9207 ( .A(n8173), .B(n8174), .Z(n8163) );
  ANDN U9208 ( .B(n8175), .A(n8176), .Z(n8173) );
  XOR U9209 ( .A(n8177), .B(n8174), .Z(n8175) );
  NAND U9210 ( .A(n8178), .B(n[1015]), .Z(n8166) );
  NAND U9211 ( .A(n8085), .B(n[1015]), .Z(n8178) );
  XOR U9212 ( .A(n8179), .B(o[1014]), .Z(creg_next[1014]) );
  AND U9213 ( .A(n3090), .B(n8180), .Z(n8179) );
  XNOR U9214 ( .A(c[1014]), .B(n8181), .Z(n8180) );
  IV U9215 ( .A(o[1014]), .Z(n8181) );
  XNOR U9216 ( .A(n8177), .B(n8176), .Z(o[1014]) );
  XNOR U9217 ( .A(n8182), .B(n8183), .Z(n8176) );
  IV U9218 ( .A(n8174), .Z(n8183) );
  XOR U9219 ( .A(n8184), .B(n8185), .Z(n8174) );
  ANDN U9220 ( .B(n8186), .A(n8187), .Z(n8184) );
  XOR U9221 ( .A(n8188), .B(n8185), .Z(n8186) );
  NAND U9222 ( .A(n8189), .B(n[1014]), .Z(n8177) );
  NAND U9223 ( .A(n8085), .B(n[1014]), .Z(n8189) );
  XOR U9224 ( .A(n8190), .B(o[1013]), .Z(creg_next[1013]) );
  AND U9225 ( .A(n3090), .B(n8191), .Z(n8190) );
  XNOR U9226 ( .A(c[1013]), .B(n8192), .Z(n8191) );
  IV U9227 ( .A(o[1013]), .Z(n8192) );
  XNOR U9228 ( .A(n8188), .B(n8187), .Z(o[1013]) );
  XNOR U9229 ( .A(n8193), .B(n8194), .Z(n8187) );
  IV U9230 ( .A(n8185), .Z(n8194) );
  XOR U9231 ( .A(n8195), .B(n8196), .Z(n8185) );
  ANDN U9232 ( .B(n8197), .A(n8198), .Z(n8195) );
  XOR U9233 ( .A(n8199), .B(n8196), .Z(n8197) );
  NAND U9234 ( .A(n8200), .B(n[1013]), .Z(n8188) );
  NAND U9235 ( .A(n8085), .B(n[1013]), .Z(n8200) );
  XOR U9236 ( .A(n8201), .B(o[1012]), .Z(creg_next[1012]) );
  AND U9237 ( .A(n3090), .B(n8202), .Z(n8201) );
  XNOR U9238 ( .A(c[1012]), .B(n8203), .Z(n8202) );
  IV U9239 ( .A(o[1012]), .Z(n8203) );
  XNOR U9240 ( .A(n8199), .B(n8198), .Z(o[1012]) );
  XNOR U9241 ( .A(n8204), .B(n8205), .Z(n8198) );
  IV U9242 ( .A(n8196), .Z(n8205) );
  XOR U9243 ( .A(n8206), .B(n8207), .Z(n8196) );
  ANDN U9244 ( .B(n8208), .A(n8209), .Z(n8206) );
  XOR U9245 ( .A(n8210), .B(n8207), .Z(n8208) );
  NAND U9246 ( .A(n8211), .B(n[1012]), .Z(n8199) );
  NAND U9247 ( .A(n8085), .B(n[1012]), .Z(n8211) );
  XOR U9248 ( .A(n8212), .B(o[1011]), .Z(creg_next[1011]) );
  AND U9249 ( .A(n3090), .B(n8213), .Z(n8212) );
  XNOR U9250 ( .A(c[1011]), .B(n8214), .Z(n8213) );
  IV U9251 ( .A(o[1011]), .Z(n8214) );
  XNOR U9252 ( .A(n8210), .B(n8209), .Z(o[1011]) );
  XNOR U9253 ( .A(n8215), .B(n8216), .Z(n8209) );
  IV U9254 ( .A(n8207), .Z(n8216) );
  XOR U9255 ( .A(n8217), .B(n8218), .Z(n8207) );
  ANDN U9256 ( .B(n8219), .A(n8220), .Z(n8217) );
  XOR U9257 ( .A(n8221), .B(n8218), .Z(n8219) );
  NAND U9258 ( .A(n8222), .B(n[1011]), .Z(n8210) );
  NAND U9259 ( .A(n8085), .B(n[1011]), .Z(n8222) );
  XOR U9260 ( .A(n8223), .B(o[1010]), .Z(creg_next[1010]) );
  AND U9261 ( .A(n3090), .B(n8224), .Z(n8223) );
  XNOR U9262 ( .A(c[1010]), .B(n8225), .Z(n8224) );
  IV U9263 ( .A(o[1010]), .Z(n8225) );
  XNOR U9264 ( .A(n8221), .B(n8220), .Z(o[1010]) );
  XNOR U9265 ( .A(n8226), .B(n8227), .Z(n8220) );
  IV U9266 ( .A(n8218), .Z(n8227) );
  XOR U9267 ( .A(n8228), .B(n8229), .Z(n8218) );
  ANDN U9268 ( .B(n8230), .A(n8231), .Z(n8228) );
  XOR U9269 ( .A(n8232), .B(n8229), .Z(n8230) );
  NAND U9270 ( .A(n8233), .B(n[1010]), .Z(n8221) );
  NAND U9271 ( .A(n8085), .B(n[1010]), .Z(n8233) );
  XOR U9272 ( .A(n8234), .B(o[100]), .Z(creg_next[100]) );
  AND U9273 ( .A(n3090), .B(n8235), .Z(n8234) );
  XNOR U9274 ( .A(c[100]), .B(n8236), .Z(n8235) );
  IV U9275 ( .A(o[100]), .Z(n8236) );
  XNOR U9276 ( .A(n8237), .B(n8238), .Z(o[100]) );
  XOR U9277 ( .A(n8239), .B(o[1009]), .Z(creg_next[1009]) );
  AND U9278 ( .A(n3090), .B(n8240), .Z(n8239) );
  XNOR U9279 ( .A(c[1009]), .B(n8241), .Z(n8240) );
  IV U9280 ( .A(o[1009]), .Z(n8241) );
  XNOR U9281 ( .A(n8232), .B(n8231), .Z(o[1009]) );
  XNOR U9282 ( .A(n8242), .B(n8243), .Z(n8231) );
  IV U9283 ( .A(n8229), .Z(n8243) );
  XOR U9284 ( .A(n8244), .B(n8245), .Z(n8229) );
  ANDN U9285 ( .B(n8246), .A(n8247), .Z(n8244) );
  XOR U9286 ( .A(n8248), .B(n8245), .Z(n8246) );
  NAND U9287 ( .A(n8249), .B(n[1009]), .Z(n8232) );
  NAND U9288 ( .A(n8085), .B(n[1009]), .Z(n8249) );
  XOR U9289 ( .A(n8250), .B(o[1008]), .Z(creg_next[1008]) );
  AND U9290 ( .A(n3090), .B(n8251), .Z(n8250) );
  XNOR U9291 ( .A(c[1008]), .B(n8252), .Z(n8251) );
  IV U9292 ( .A(o[1008]), .Z(n8252) );
  XNOR U9293 ( .A(n8248), .B(n8247), .Z(o[1008]) );
  XNOR U9294 ( .A(n8253), .B(n8254), .Z(n8247) );
  IV U9295 ( .A(n8245), .Z(n8254) );
  XOR U9296 ( .A(n8255), .B(n8256), .Z(n8245) );
  ANDN U9297 ( .B(n8257), .A(n8258), .Z(n8255) );
  XOR U9298 ( .A(n8259), .B(n8256), .Z(n8257) );
  NAND U9299 ( .A(n8260), .B(n[1008]), .Z(n8248) );
  NAND U9300 ( .A(n8085), .B(n[1008]), .Z(n8260) );
  XOR U9301 ( .A(n8261), .B(o[1007]), .Z(creg_next[1007]) );
  AND U9302 ( .A(n3090), .B(n8262), .Z(n8261) );
  XNOR U9303 ( .A(c[1007]), .B(n8263), .Z(n8262) );
  IV U9304 ( .A(o[1007]), .Z(n8263) );
  XNOR U9305 ( .A(n8259), .B(n8258), .Z(o[1007]) );
  XNOR U9306 ( .A(n8264), .B(n8265), .Z(n8258) );
  IV U9307 ( .A(n8256), .Z(n8265) );
  XOR U9308 ( .A(n8266), .B(n8267), .Z(n8256) );
  ANDN U9309 ( .B(n8268), .A(n8269), .Z(n8266) );
  XOR U9310 ( .A(n8270), .B(n8267), .Z(n8268) );
  NAND U9311 ( .A(n8271), .B(n[1007]), .Z(n8259) );
  NAND U9312 ( .A(n8085), .B(n[1007]), .Z(n8271) );
  XOR U9313 ( .A(n8272), .B(o[1006]), .Z(creg_next[1006]) );
  AND U9314 ( .A(n3090), .B(n8273), .Z(n8272) );
  XNOR U9315 ( .A(c[1006]), .B(n8274), .Z(n8273) );
  IV U9316 ( .A(o[1006]), .Z(n8274) );
  XNOR U9317 ( .A(n8270), .B(n8269), .Z(o[1006]) );
  XNOR U9318 ( .A(n8275), .B(n8276), .Z(n8269) );
  IV U9319 ( .A(n8267), .Z(n8276) );
  XOR U9320 ( .A(n8277), .B(n8278), .Z(n8267) );
  ANDN U9321 ( .B(n8279), .A(n8280), .Z(n8277) );
  XOR U9322 ( .A(n8281), .B(n8278), .Z(n8279) );
  NAND U9323 ( .A(n8282), .B(n[1006]), .Z(n8270) );
  NAND U9324 ( .A(n8085), .B(n[1006]), .Z(n8282) );
  XOR U9325 ( .A(n8283), .B(o[1005]), .Z(creg_next[1005]) );
  AND U9326 ( .A(n3090), .B(n8284), .Z(n8283) );
  XNOR U9327 ( .A(c[1005]), .B(n8285), .Z(n8284) );
  IV U9328 ( .A(o[1005]), .Z(n8285) );
  XNOR U9329 ( .A(n8281), .B(n8280), .Z(o[1005]) );
  XNOR U9330 ( .A(n8286), .B(n8287), .Z(n8280) );
  IV U9331 ( .A(n8278), .Z(n8287) );
  XOR U9332 ( .A(n8288), .B(n8289), .Z(n8278) );
  ANDN U9333 ( .B(n8290), .A(n8291), .Z(n8288) );
  XOR U9334 ( .A(n8292), .B(n8289), .Z(n8290) );
  NAND U9335 ( .A(n8293), .B(n[1005]), .Z(n8281) );
  NAND U9336 ( .A(n8085), .B(n[1005]), .Z(n8293) );
  XOR U9337 ( .A(n8294), .B(o[1004]), .Z(creg_next[1004]) );
  AND U9338 ( .A(n3090), .B(n8295), .Z(n8294) );
  XNOR U9339 ( .A(c[1004]), .B(n8296), .Z(n8295) );
  IV U9340 ( .A(o[1004]), .Z(n8296) );
  XNOR U9341 ( .A(n8292), .B(n8291), .Z(o[1004]) );
  XNOR U9342 ( .A(n8297), .B(n8298), .Z(n8291) );
  IV U9343 ( .A(n8289), .Z(n8298) );
  XOR U9344 ( .A(n8299), .B(n8300), .Z(n8289) );
  ANDN U9345 ( .B(n8301), .A(n8302), .Z(n8299) );
  XOR U9346 ( .A(n8303), .B(n8300), .Z(n8301) );
  NAND U9347 ( .A(n8304), .B(n[1004]), .Z(n8292) );
  NAND U9348 ( .A(n8085), .B(n[1004]), .Z(n8304) );
  XOR U9349 ( .A(n8305), .B(o[1003]), .Z(creg_next[1003]) );
  AND U9350 ( .A(n3090), .B(n8306), .Z(n8305) );
  XNOR U9351 ( .A(c[1003]), .B(n8307), .Z(n8306) );
  IV U9352 ( .A(o[1003]), .Z(n8307) );
  XNOR U9353 ( .A(n8303), .B(n8302), .Z(o[1003]) );
  XNOR U9354 ( .A(n8308), .B(n8309), .Z(n8302) );
  IV U9355 ( .A(n8300), .Z(n8309) );
  XOR U9356 ( .A(n8310), .B(n8311), .Z(n8300) );
  ANDN U9357 ( .B(n8312), .A(n8313), .Z(n8310) );
  XOR U9358 ( .A(n8314), .B(n8311), .Z(n8312) );
  NAND U9359 ( .A(n8315), .B(n[1003]), .Z(n8303) );
  NAND U9360 ( .A(n8085), .B(n[1003]), .Z(n8315) );
  XOR U9361 ( .A(n8316), .B(o[1002]), .Z(creg_next[1002]) );
  AND U9362 ( .A(n3090), .B(n8317), .Z(n8316) );
  XNOR U9363 ( .A(c[1002]), .B(n8318), .Z(n8317) );
  IV U9364 ( .A(o[1002]), .Z(n8318) );
  XNOR U9365 ( .A(n8314), .B(n8313), .Z(o[1002]) );
  XNOR U9366 ( .A(n8319), .B(n8320), .Z(n8313) );
  IV U9367 ( .A(n8311), .Z(n8320) );
  XOR U9368 ( .A(n8321), .B(n8322), .Z(n8311) );
  ANDN U9369 ( .B(n8323), .A(n8324), .Z(n8321) );
  XOR U9370 ( .A(n8325), .B(n8322), .Z(n8323) );
  NAND U9371 ( .A(n8326), .B(n[1002]), .Z(n8314) );
  NAND U9372 ( .A(n8085), .B(n[1002]), .Z(n8326) );
  XOR U9373 ( .A(n8327), .B(o[1001]), .Z(creg_next[1001]) );
  AND U9374 ( .A(n3090), .B(n8328), .Z(n8327) );
  XNOR U9375 ( .A(c[1001]), .B(n8329), .Z(n8328) );
  IV U9376 ( .A(o[1001]), .Z(n8329) );
  XNOR U9377 ( .A(n8325), .B(n8324), .Z(o[1001]) );
  XNOR U9378 ( .A(n8330), .B(n8331), .Z(n8324) );
  IV U9379 ( .A(n8322), .Z(n8331) );
  XOR U9380 ( .A(n8332), .B(n8333), .Z(n8322) );
  ANDN U9381 ( .B(n8334), .A(n8335), .Z(n8332) );
  XOR U9382 ( .A(n8336), .B(n8333), .Z(n8334) );
  NAND U9383 ( .A(n8337), .B(n[1001]), .Z(n8325) );
  NAND U9384 ( .A(n8085), .B(n[1001]), .Z(n8337) );
  XOR U9385 ( .A(n8338), .B(o[1000]), .Z(creg_next[1000]) );
  AND U9386 ( .A(n3090), .B(n8339), .Z(n8338) );
  XNOR U9387 ( .A(c[1000]), .B(n8340), .Z(n8339) );
  IV U9388 ( .A(o[1000]), .Z(n8340) );
  XNOR U9389 ( .A(n8336), .B(n8335), .Z(o[1000]) );
  XNOR U9390 ( .A(n8341), .B(n8342), .Z(n8335) );
  IV U9391 ( .A(n8333), .Z(n8342) );
  XOR U9392 ( .A(n8343), .B(n8344), .Z(n8333) );
  ANDN U9393 ( .B(n8345), .A(n3104), .Z(n8343) );
  XNOR U9394 ( .A(n8346), .B(n8347), .Z(n3104) );
  IV U9395 ( .A(n8344), .Z(n8347) );
  XOR U9396 ( .A(n3103), .B(n8344), .Z(n8345) );
  XOR U9397 ( .A(n8348), .B(n8349), .Z(n8344) );
  ANDN U9398 ( .B(n8350), .A(n3109), .Z(n8348) );
  XNOR U9399 ( .A(n8351), .B(n8352), .Z(n3109) );
  IV U9400 ( .A(n8349), .Z(n8352) );
  XOR U9401 ( .A(n3108), .B(n8349), .Z(n8350) );
  XOR U9402 ( .A(n8353), .B(n8354), .Z(n8349) );
  ANDN U9403 ( .B(n8355), .A(n3114), .Z(n8353) );
  XNOR U9404 ( .A(n8356), .B(n8357), .Z(n3114) );
  IV U9405 ( .A(n8354), .Z(n8357) );
  XOR U9406 ( .A(n3113), .B(n8354), .Z(n8355) );
  XOR U9407 ( .A(n8358), .B(n8359), .Z(n8354) );
  ANDN U9408 ( .B(n8360), .A(n3119), .Z(n8358) );
  XNOR U9409 ( .A(n8361), .B(n8362), .Z(n3119) );
  IV U9410 ( .A(n8359), .Z(n8362) );
  XOR U9411 ( .A(n3118), .B(n8359), .Z(n8360) );
  XOR U9412 ( .A(n8363), .B(n8364), .Z(n8359) );
  ANDN U9413 ( .B(n8365), .A(n3124), .Z(n8363) );
  XNOR U9414 ( .A(n8366), .B(n8367), .Z(n3124) );
  IV U9415 ( .A(n8364), .Z(n8367) );
  XOR U9416 ( .A(n3123), .B(n8364), .Z(n8365) );
  XOR U9417 ( .A(n8368), .B(n8369), .Z(n8364) );
  ANDN U9418 ( .B(n8370), .A(n3129), .Z(n8368) );
  XNOR U9419 ( .A(n8371), .B(n8372), .Z(n3129) );
  IV U9420 ( .A(n8369), .Z(n8372) );
  XOR U9421 ( .A(n3128), .B(n8369), .Z(n8370) );
  XOR U9422 ( .A(n8373), .B(n8374), .Z(n8369) );
  ANDN U9423 ( .B(n8375), .A(n3134), .Z(n8373) );
  XNOR U9424 ( .A(n8376), .B(n8377), .Z(n3134) );
  IV U9425 ( .A(n8374), .Z(n8377) );
  XOR U9426 ( .A(n3133), .B(n8374), .Z(n8375) );
  XOR U9427 ( .A(n8378), .B(n8379), .Z(n8374) );
  ANDN U9428 ( .B(n8380), .A(n3139), .Z(n8378) );
  XNOR U9429 ( .A(n8381), .B(n8382), .Z(n3139) );
  IV U9430 ( .A(n8379), .Z(n8382) );
  XOR U9431 ( .A(n3138), .B(n8379), .Z(n8380) );
  XOR U9432 ( .A(n8383), .B(n8384), .Z(n8379) );
  ANDN U9433 ( .B(n8385), .A(n3144), .Z(n8383) );
  XNOR U9434 ( .A(n8386), .B(n8387), .Z(n3144) );
  IV U9435 ( .A(n8384), .Z(n8387) );
  XOR U9436 ( .A(n3143), .B(n8384), .Z(n8385) );
  XOR U9437 ( .A(n8388), .B(n8389), .Z(n8384) );
  ANDN U9438 ( .B(n8390), .A(n3149), .Z(n8388) );
  XNOR U9439 ( .A(n8391), .B(n8392), .Z(n3149) );
  IV U9440 ( .A(n8389), .Z(n8392) );
  XOR U9441 ( .A(n3148), .B(n8389), .Z(n8390) );
  XOR U9442 ( .A(n8393), .B(n8394), .Z(n8389) );
  ANDN U9443 ( .B(n8395), .A(n3159), .Z(n8393) );
  XNOR U9444 ( .A(n8396), .B(n8397), .Z(n3159) );
  IV U9445 ( .A(n8394), .Z(n8397) );
  XOR U9446 ( .A(n3158), .B(n8394), .Z(n8395) );
  XOR U9447 ( .A(n8398), .B(n8399), .Z(n8394) );
  ANDN U9448 ( .B(n8400), .A(n3164), .Z(n8398) );
  XNOR U9449 ( .A(n8401), .B(n8402), .Z(n3164) );
  IV U9450 ( .A(n8399), .Z(n8402) );
  XOR U9451 ( .A(n3163), .B(n8399), .Z(n8400) );
  XOR U9452 ( .A(n8403), .B(n8404), .Z(n8399) );
  ANDN U9453 ( .B(n8405), .A(n3169), .Z(n8403) );
  XNOR U9454 ( .A(n8406), .B(n8407), .Z(n3169) );
  IV U9455 ( .A(n8404), .Z(n8407) );
  XOR U9456 ( .A(n3168), .B(n8404), .Z(n8405) );
  XOR U9457 ( .A(n8408), .B(n8409), .Z(n8404) );
  ANDN U9458 ( .B(n8410), .A(n3174), .Z(n8408) );
  XNOR U9459 ( .A(n8411), .B(n8412), .Z(n3174) );
  IV U9460 ( .A(n8409), .Z(n8412) );
  XOR U9461 ( .A(n3173), .B(n8409), .Z(n8410) );
  XOR U9462 ( .A(n8413), .B(n8414), .Z(n8409) );
  ANDN U9463 ( .B(n8415), .A(n3179), .Z(n8413) );
  XNOR U9464 ( .A(n8416), .B(n8417), .Z(n3179) );
  IV U9465 ( .A(n8414), .Z(n8417) );
  XOR U9466 ( .A(n3178), .B(n8414), .Z(n8415) );
  XOR U9467 ( .A(n8418), .B(n8419), .Z(n8414) );
  ANDN U9468 ( .B(n8420), .A(n3184), .Z(n8418) );
  XNOR U9469 ( .A(n8421), .B(n8422), .Z(n3184) );
  IV U9470 ( .A(n8419), .Z(n8422) );
  XOR U9471 ( .A(n3183), .B(n8419), .Z(n8420) );
  XOR U9472 ( .A(n8423), .B(n8424), .Z(n8419) );
  ANDN U9473 ( .B(n8425), .A(n3189), .Z(n8423) );
  XNOR U9474 ( .A(n8426), .B(n8427), .Z(n3189) );
  IV U9475 ( .A(n8424), .Z(n8427) );
  XOR U9476 ( .A(n3188), .B(n8424), .Z(n8425) );
  XOR U9477 ( .A(n8428), .B(n8429), .Z(n8424) );
  ANDN U9478 ( .B(n8430), .A(n3194), .Z(n8428) );
  XNOR U9479 ( .A(n8431), .B(n8432), .Z(n3194) );
  IV U9480 ( .A(n8429), .Z(n8432) );
  XOR U9481 ( .A(n3193), .B(n8429), .Z(n8430) );
  XOR U9482 ( .A(n8433), .B(n8434), .Z(n8429) );
  ANDN U9483 ( .B(n8435), .A(n3199), .Z(n8433) );
  XNOR U9484 ( .A(n8436), .B(n8437), .Z(n3199) );
  IV U9485 ( .A(n8434), .Z(n8437) );
  XOR U9486 ( .A(n3198), .B(n8434), .Z(n8435) );
  XOR U9487 ( .A(n8438), .B(n8439), .Z(n8434) );
  ANDN U9488 ( .B(n8440), .A(n3204), .Z(n8438) );
  XNOR U9489 ( .A(n8441), .B(n8442), .Z(n3204) );
  IV U9490 ( .A(n8439), .Z(n8442) );
  XOR U9491 ( .A(n3203), .B(n8439), .Z(n8440) );
  XOR U9492 ( .A(n8443), .B(n8444), .Z(n8439) );
  ANDN U9493 ( .B(n8445), .A(n3214), .Z(n8443) );
  XNOR U9494 ( .A(n8446), .B(n8447), .Z(n3214) );
  IV U9495 ( .A(n8444), .Z(n8447) );
  XOR U9496 ( .A(n3213), .B(n8444), .Z(n8445) );
  XOR U9497 ( .A(n8448), .B(n8449), .Z(n8444) );
  ANDN U9498 ( .B(n8450), .A(n3219), .Z(n8448) );
  XNOR U9499 ( .A(n8451), .B(n8452), .Z(n3219) );
  IV U9500 ( .A(n8449), .Z(n8452) );
  XOR U9501 ( .A(n3218), .B(n8449), .Z(n8450) );
  XOR U9502 ( .A(n8453), .B(n8454), .Z(n8449) );
  ANDN U9503 ( .B(n8455), .A(n3224), .Z(n8453) );
  XNOR U9504 ( .A(n8456), .B(n8457), .Z(n3224) );
  IV U9505 ( .A(n8454), .Z(n8457) );
  XOR U9506 ( .A(n3223), .B(n8454), .Z(n8455) );
  XOR U9507 ( .A(n8458), .B(n8459), .Z(n8454) );
  ANDN U9508 ( .B(n8460), .A(n3229), .Z(n8458) );
  XNOR U9509 ( .A(n8461), .B(n8462), .Z(n3229) );
  IV U9510 ( .A(n8459), .Z(n8462) );
  XOR U9511 ( .A(n3228), .B(n8459), .Z(n8460) );
  XOR U9512 ( .A(n8463), .B(n8464), .Z(n8459) );
  ANDN U9513 ( .B(n8465), .A(n3234), .Z(n8463) );
  XNOR U9514 ( .A(n8466), .B(n8467), .Z(n3234) );
  IV U9515 ( .A(n8464), .Z(n8467) );
  XOR U9516 ( .A(n3233), .B(n8464), .Z(n8465) );
  XOR U9517 ( .A(n8468), .B(n8469), .Z(n8464) );
  ANDN U9518 ( .B(n8470), .A(n3239), .Z(n8468) );
  XNOR U9519 ( .A(n8471), .B(n8472), .Z(n3239) );
  IV U9520 ( .A(n8469), .Z(n8472) );
  XOR U9521 ( .A(n3238), .B(n8469), .Z(n8470) );
  XOR U9522 ( .A(n8473), .B(n8474), .Z(n8469) );
  ANDN U9523 ( .B(n8475), .A(n3244), .Z(n8473) );
  XNOR U9524 ( .A(n8476), .B(n8477), .Z(n3244) );
  IV U9525 ( .A(n8474), .Z(n8477) );
  XOR U9526 ( .A(n3243), .B(n8474), .Z(n8475) );
  XOR U9527 ( .A(n8478), .B(n8479), .Z(n8474) );
  ANDN U9528 ( .B(n8480), .A(n3249), .Z(n8478) );
  XNOR U9529 ( .A(n8481), .B(n8482), .Z(n3249) );
  IV U9530 ( .A(n8479), .Z(n8482) );
  XOR U9531 ( .A(n3248), .B(n8479), .Z(n8480) );
  XOR U9532 ( .A(n8483), .B(n8484), .Z(n8479) );
  ANDN U9533 ( .B(n8485), .A(n3254), .Z(n8483) );
  XNOR U9534 ( .A(n8486), .B(n8487), .Z(n3254) );
  IV U9535 ( .A(n8484), .Z(n8487) );
  XOR U9536 ( .A(n3253), .B(n8484), .Z(n8485) );
  XOR U9537 ( .A(n8488), .B(n8489), .Z(n8484) );
  ANDN U9538 ( .B(n8490), .A(n3259), .Z(n8488) );
  XNOR U9539 ( .A(n8491), .B(n8492), .Z(n3259) );
  IV U9540 ( .A(n8489), .Z(n8492) );
  XOR U9541 ( .A(n3258), .B(n8489), .Z(n8490) );
  XOR U9542 ( .A(n8493), .B(n8494), .Z(n8489) );
  ANDN U9543 ( .B(n8495), .A(n3269), .Z(n8493) );
  XNOR U9544 ( .A(n8496), .B(n8497), .Z(n3269) );
  IV U9545 ( .A(n8494), .Z(n8497) );
  XOR U9546 ( .A(n3268), .B(n8494), .Z(n8495) );
  XOR U9547 ( .A(n8498), .B(n8499), .Z(n8494) );
  ANDN U9548 ( .B(n8500), .A(n3274), .Z(n8498) );
  XNOR U9549 ( .A(n8501), .B(n8502), .Z(n3274) );
  IV U9550 ( .A(n8499), .Z(n8502) );
  XOR U9551 ( .A(n3273), .B(n8499), .Z(n8500) );
  XOR U9552 ( .A(n8503), .B(n8504), .Z(n8499) );
  ANDN U9553 ( .B(n8505), .A(n3279), .Z(n8503) );
  XNOR U9554 ( .A(n8506), .B(n8507), .Z(n3279) );
  IV U9555 ( .A(n8504), .Z(n8507) );
  XOR U9556 ( .A(n3278), .B(n8504), .Z(n8505) );
  XOR U9557 ( .A(n8508), .B(n8509), .Z(n8504) );
  ANDN U9558 ( .B(n8510), .A(n3284), .Z(n8508) );
  XNOR U9559 ( .A(n8511), .B(n8512), .Z(n3284) );
  IV U9560 ( .A(n8509), .Z(n8512) );
  XOR U9561 ( .A(n3283), .B(n8509), .Z(n8510) );
  XOR U9562 ( .A(n8513), .B(n8514), .Z(n8509) );
  ANDN U9563 ( .B(n8515), .A(n3289), .Z(n8513) );
  XNOR U9564 ( .A(n8516), .B(n8517), .Z(n3289) );
  IV U9565 ( .A(n8514), .Z(n8517) );
  XOR U9566 ( .A(n3288), .B(n8514), .Z(n8515) );
  XOR U9567 ( .A(n8518), .B(n8519), .Z(n8514) );
  ANDN U9568 ( .B(n8520), .A(n3294), .Z(n8518) );
  XNOR U9569 ( .A(n8521), .B(n8522), .Z(n3294) );
  IV U9570 ( .A(n8519), .Z(n8522) );
  XOR U9571 ( .A(n3293), .B(n8519), .Z(n8520) );
  XOR U9572 ( .A(n8523), .B(n8524), .Z(n8519) );
  ANDN U9573 ( .B(n8525), .A(n3299), .Z(n8523) );
  XNOR U9574 ( .A(n8526), .B(n8527), .Z(n3299) );
  IV U9575 ( .A(n8524), .Z(n8527) );
  XOR U9576 ( .A(n3298), .B(n8524), .Z(n8525) );
  XOR U9577 ( .A(n8528), .B(n8529), .Z(n8524) );
  ANDN U9578 ( .B(n8530), .A(n3304), .Z(n8528) );
  XNOR U9579 ( .A(n8531), .B(n8532), .Z(n3304) );
  IV U9580 ( .A(n8529), .Z(n8532) );
  XOR U9581 ( .A(n3303), .B(n8529), .Z(n8530) );
  XOR U9582 ( .A(n8533), .B(n8534), .Z(n8529) );
  ANDN U9583 ( .B(n8535), .A(n3309), .Z(n8533) );
  XNOR U9584 ( .A(n8536), .B(n8537), .Z(n3309) );
  IV U9585 ( .A(n8534), .Z(n8537) );
  XOR U9586 ( .A(n3308), .B(n8534), .Z(n8535) );
  XOR U9587 ( .A(n8538), .B(n8539), .Z(n8534) );
  ANDN U9588 ( .B(n8540), .A(n3314), .Z(n8538) );
  XNOR U9589 ( .A(n8541), .B(n8542), .Z(n3314) );
  IV U9590 ( .A(n8539), .Z(n8542) );
  XOR U9591 ( .A(n3313), .B(n8539), .Z(n8540) );
  XOR U9592 ( .A(n8543), .B(n8544), .Z(n8539) );
  ANDN U9593 ( .B(n8545), .A(n3324), .Z(n8543) );
  XNOR U9594 ( .A(n8546), .B(n8547), .Z(n3324) );
  IV U9595 ( .A(n8544), .Z(n8547) );
  XOR U9596 ( .A(n3323), .B(n8544), .Z(n8545) );
  XOR U9597 ( .A(n8548), .B(n8549), .Z(n8544) );
  ANDN U9598 ( .B(n8550), .A(n3329), .Z(n8548) );
  XNOR U9599 ( .A(n8551), .B(n8552), .Z(n3329) );
  IV U9600 ( .A(n8549), .Z(n8552) );
  XOR U9601 ( .A(n3328), .B(n8549), .Z(n8550) );
  XOR U9602 ( .A(n8553), .B(n8554), .Z(n8549) );
  ANDN U9603 ( .B(n8555), .A(n3334), .Z(n8553) );
  XNOR U9604 ( .A(n8556), .B(n8557), .Z(n3334) );
  IV U9605 ( .A(n8554), .Z(n8557) );
  XOR U9606 ( .A(n3333), .B(n8554), .Z(n8555) );
  XOR U9607 ( .A(n8558), .B(n8559), .Z(n8554) );
  ANDN U9608 ( .B(n8560), .A(n3339), .Z(n8558) );
  XNOR U9609 ( .A(n8561), .B(n8562), .Z(n3339) );
  IV U9610 ( .A(n8559), .Z(n8562) );
  XOR U9611 ( .A(n3338), .B(n8559), .Z(n8560) );
  XOR U9612 ( .A(n8563), .B(n8564), .Z(n8559) );
  ANDN U9613 ( .B(n8565), .A(n3344), .Z(n8563) );
  XNOR U9614 ( .A(n8566), .B(n8567), .Z(n3344) );
  IV U9615 ( .A(n8564), .Z(n8567) );
  XOR U9616 ( .A(n3343), .B(n8564), .Z(n8565) );
  XOR U9617 ( .A(n8568), .B(n8569), .Z(n8564) );
  ANDN U9618 ( .B(n8570), .A(n3349), .Z(n8568) );
  XNOR U9619 ( .A(n8571), .B(n8572), .Z(n3349) );
  IV U9620 ( .A(n8569), .Z(n8572) );
  XOR U9621 ( .A(n3348), .B(n8569), .Z(n8570) );
  XOR U9622 ( .A(n8573), .B(n8574), .Z(n8569) );
  ANDN U9623 ( .B(n8575), .A(n3354), .Z(n8573) );
  XNOR U9624 ( .A(n8576), .B(n8577), .Z(n3354) );
  IV U9625 ( .A(n8574), .Z(n8577) );
  XOR U9626 ( .A(n3353), .B(n8574), .Z(n8575) );
  XOR U9627 ( .A(n8578), .B(n8579), .Z(n8574) );
  ANDN U9628 ( .B(n8580), .A(n3359), .Z(n8578) );
  XNOR U9629 ( .A(n8581), .B(n8582), .Z(n3359) );
  IV U9630 ( .A(n8579), .Z(n8582) );
  XOR U9631 ( .A(n3358), .B(n8579), .Z(n8580) );
  XOR U9632 ( .A(n8583), .B(n8584), .Z(n8579) );
  ANDN U9633 ( .B(n8585), .A(n3364), .Z(n8583) );
  XNOR U9634 ( .A(n8586), .B(n8587), .Z(n3364) );
  IV U9635 ( .A(n8584), .Z(n8587) );
  XOR U9636 ( .A(n3363), .B(n8584), .Z(n8585) );
  XOR U9637 ( .A(n8588), .B(n8589), .Z(n8584) );
  ANDN U9638 ( .B(n8590), .A(n3369), .Z(n8588) );
  XNOR U9639 ( .A(n8591), .B(n8592), .Z(n3369) );
  IV U9640 ( .A(n8589), .Z(n8592) );
  XOR U9641 ( .A(n3368), .B(n8589), .Z(n8590) );
  XOR U9642 ( .A(n8593), .B(n8594), .Z(n8589) );
  ANDN U9643 ( .B(n8595), .A(n3379), .Z(n8593) );
  XNOR U9644 ( .A(n8596), .B(n8597), .Z(n3379) );
  IV U9645 ( .A(n8594), .Z(n8597) );
  XOR U9646 ( .A(n3378), .B(n8594), .Z(n8595) );
  XOR U9647 ( .A(n8598), .B(n8599), .Z(n8594) );
  ANDN U9648 ( .B(n8600), .A(n3384), .Z(n8598) );
  XNOR U9649 ( .A(n8601), .B(n8602), .Z(n3384) );
  IV U9650 ( .A(n8599), .Z(n8602) );
  XOR U9651 ( .A(n3383), .B(n8599), .Z(n8600) );
  XOR U9652 ( .A(n8603), .B(n8604), .Z(n8599) );
  ANDN U9653 ( .B(n8605), .A(n3389), .Z(n8603) );
  XNOR U9654 ( .A(n8606), .B(n8607), .Z(n3389) );
  IV U9655 ( .A(n8604), .Z(n8607) );
  XOR U9656 ( .A(n3388), .B(n8604), .Z(n8605) );
  XOR U9657 ( .A(n8608), .B(n8609), .Z(n8604) );
  ANDN U9658 ( .B(n8610), .A(n3394), .Z(n8608) );
  XNOR U9659 ( .A(n8611), .B(n8612), .Z(n3394) );
  IV U9660 ( .A(n8609), .Z(n8612) );
  XOR U9661 ( .A(n3393), .B(n8609), .Z(n8610) );
  XOR U9662 ( .A(n8613), .B(n8614), .Z(n8609) );
  ANDN U9663 ( .B(n8615), .A(n3399), .Z(n8613) );
  XNOR U9664 ( .A(n8616), .B(n8617), .Z(n3399) );
  IV U9665 ( .A(n8614), .Z(n8617) );
  XOR U9666 ( .A(n3398), .B(n8614), .Z(n8615) );
  XOR U9667 ( .A(n8618), .B(n8619), .Z(n8614) );
  ANDN U9668 ( .B(n8620), .A(n3404), .Z(n8618) );
  XNOR U9669 ( .A(n8621), .B(n8622), .Z(n3404) );
  IV U9670 ( .A(n8619), .Z(n8622) );
  XOR U9671 ( .A(n3403), .B(n8619), .Z(n8620) );
  XOR U9672 ( .A(n8623), .B(n8624), .Z(n8619) );
  ANDN U9673 ( .B(n8625), .A(n3409), .Z(n8623) );
  XNOR U9674 ( .A(n8626), .B(n8627), .Z(n3409) );
  IV U9675 ( .A(n8624), .Z(n8627) );
  XOR U9676 ( .A(n3408), .B(n8624), .Z(n8625) );
  XOR U9677 ( .A(n8628), .B(n8629), .Z(n8624) );
  ANDN U9678 ( .B(n8630), .A(n3414), .Z(n8628) );
  XNOR U9679 ( .A(n8631), .B(n8632), .Z(n3414) );
  IV U9680 ( .A(n8629), .Z(n8632) );
  XOR U9681 ( .A(n3413), .B(n8629), .Z(n8630) );
  XOR U9682 ( .A(n8633), .B(n8634), .Z(n8629) );
  ANDN U9683 ( .B(n8635), .A(n3419), .Z(n8633) );
  XNOR U9684 ( .A(n8636), .B(n8637), .Z(n3419) );
  IV U9685 ( .A(n8634), .Z(n8637) );
  XOR U9686 ( .A(n3418), .B(n8634), .Z(n8635) );
  XOR U9687 ( .A(n8638), .B(n8639), .Z(n8634) );
  ANDN U9688 ( .B(n8640), .A(n3424), .Z(n8638) );
  XNOR U9689 ( .A(n8641), .B(n8642), .Z(n3424) );
  IV U9690 ( .A(n8639), .Z(n8642) );
  XOR U9691 ( .A(n3423), .B(n8639), .Z(n8640) );
  XOR U9692 ( .A(n8643), .B(n8644), .Z(n8639) );
  ANDN U9693 ( .B(n8645), .A(n3434), .Z(n8643) );
  XNOR U9694 ( .A(n8646), .B(n8647), .Z(n3434) );
  IV U9695 ( .A(n8644), .Z(n8647) );
  XOR U9696 ( .A(n3433), .B(n8644), .Z(n8645) );
  XOR U9697 ( .A(n8648), .B(n8649), .Z(n8644) );
  ANDN U9698 ( .B(n8650), .A(n3439), .Z(n8648) );
  XNOR U9699 ( .A(n8651), .B(n8652), .Z(n3439) );
  IV U9700 ( .A(n8649), .Z(n8652) );
  XOR U9701 ( .A(n3438), .B(n8649), .Z(n8650) );
  XOR U9702 ( .A(n8653), .B(n8654), .Z(n8649) );
  ANDN U9703 ( .B(n8655), .A(n3444), .Z(n8653) );
  XNOR U9704 ( .A(n8656), .B(n8657), .Z(n3444) );
  IV U9705 ( .A(n8654), .Z(n8657) );
  XOR U9706 ( .A(n3443), .B(n8654), .Z(n8655) );
  XOR U9707 ( .A(n8658), .B(n8659), .Z(n8654) );
  ANDN U9708 ( .B(n8660), .A(n3449), .Z(n8658) );
  XNOR U9709 ( .A(n8661), .B(n8662), .Z(n3449) );
  IV U9710 ( .A(n8659), .Z(n8662) );
  XOR U9711 ( .A(n3448), .B(n8659), .Z(n8660) );
  XOR U9712 ( .A(n8663), .B(n8664), .Z(n8659) );
  ANDN U9713 ( .B(n8665), .A(n3454), .Z(n8663) );
  XNOR U9714 ( .A(n8666), .B(n8667), .Z(n3454) );
  IV U9715 ( .A(n8664), .Z(n8667) );
  XOR U9716 ( .A(n3453), .B(n8664), .Z(n8665) );
  XOR U9717 ( .A(n8668), .B(n8669), .Z(n8664) );
  ANDN U9718 ( .B(n8670), .A(n3459), .Z(n8668) );
  XNOR U9719 ( .A(n8671), .B(n8672), .Z(n3459) );
  IV U9720 ( .A(n8669), .Z(n8672) );
  XOR U9721 ( .A(n3458), .B(n8669), .Z(n8670) );
  XOR U9722 ( .A(n8673), .B(n8674), .Z(n8669) );
  ANDN U9723 ( .B(n8675), .A(n3464), .Z(n8673) );
  XNOR U9724 ( .A(n8676), .B(n8677), .Z(n3464) );
  IV U9725 ( .A(n8674), .Z(n8677) );
  XOR U9726 ( .A(n3463), .B(n8674), .Z(n8675) );
  XOR U9727 ( .A(n8678), .B(n8679), .Z(n8674) );
  ANDN U9728 ( .B(n8680), .A(n3469), .Z(n8678) );
  XNOR U9729 ( .A(n8681), .B(n8682), .Z(n3469) );
  IV U9730 ( .A(n8679), .Z(n8682) );
  XOR U9731 ( .A(n3468), .B(n8679), .Z(n8680) );
  XOR U9732 ( .A(n8683), .B(n8684), .Z(n8679) );
  ANDN U9733 ( .B(n8685), .A(n3474), .Z(n8683) );
  XNOR U9734 ( .A(n8686), .B(n8687), .Z(n3474) );
  IV U9735 ( .A(n8684), .Z(n8687) );
  XOR U9736 ( .A(n3473), .B(n8684), .Z(n8685) );
  XOR U9737 ( .A(n8688), .B(n8689), .Z(n8684) );
  ANDN U9738 ( .B(n8690), .A(n3479), .Z(n8688) );
  XNOR U9739 ( .A(n8691), .B(n8692), .Z(n3479) );
  IV U9740 ( .A(n8689), .Z(n8692) );
  XOR U9741 ( .A(n3478), .B(n8689), .Z(n8690) );
  XOR U9742 ( .A(n8693), .B(n8694), .Z(n8689) );
  ANDN U9743 ( .B(n8695), .A(n3489), .Z(n8693) );
  XNOR U9744 ( .A(n8696), .B(n8697), .Z(n3489) );
  IV U9745 ( .A(n8694), .Z(n8697) );
  XOR U9746 ( .A(n3488), .B(n8694), .Z(n8695) );
  XOR U9747 ( .A(n8698), .B(n8699), .Z(n8694) );
  ANDN U9748 ( .B(n8700), .A(n3494), .Z(n8698) );
  XNOR U9749 ( .A(n8701), .B(n8702), .Z(n3494) );
  IV U9750 ( .A(n8699), .Z(n8702) );
  XOR U9751 ( .A(n3493), .B(n8699), .Z(n8700) );
  XOR U9752 ( .A(n8703), .B(n8704), .Z(n8699) );
  ANDN U9753 ( .B(n8705), .A(n3499), .Z(n8703) );
  XNOR U9754 ( .A(n8706), .B(n8707), .Z(n3499) );
  IV U9755 ( .A(n8704), .Z(n8707) );
  XOR U9756 ( .A(n3498), .B(n8704), .Z(n8705) );
  XOR U9757 ( .A(n8708), .B(n8709), .Z(n8704) );
  ANDN U9758 ( .B(n8710), .A(n3504), .Z(n8708) );
  XNOR U9759 ( .A(n8711), .B(n8712), .Z(n3504) );
  IV U9760 ( .A(n8709), .Z(n8712) );
  XOR U9761 ( .A(n3503), .B(n8709), .Z(n8710) );
  XOR U9762 ( .A(n8713), .B(n8714), .Z(n8709) );
  ANDN U9763 ( .B(n8715), .A(n3509), .Z(n8713) );
  XNOR U9764 ( .A(n8716), .B(n8717), .Z(n3509) );
  IV U9765 ( .A(n8714), .Z(n8717) );
  XOR U9766 ( .A(n3508), .B(n8714), .Z(n8715) );
  XOR U9767 ( .A(n8718), .B(n8719), .Z(n8714) );
  ANDN U9768 ( .B(n8720), .A(n3514), .Z(n8718) );
  XNOR U9769 ( .A(n8721), .B(n8722), .Z(n3514) );
  IV U9770 ( .A(n8719), .Z(n8722) );
  XOR U9771 ( .A(n3513), .B(n8719), .Z(n8720) );
  XOR U9772 ( .A(n8723), .B(n8724), .Z(n8719) );
  ANDN U9773 ( .B(n8725), .A(n3519), .Z(n8723) );
  XNOR U9774 ( .A(n8726), .B(n8727), .Z(n3519) );
  IV U9775 ( .A(n8724), .Z(n8727) );
  XOR U9776 ( .A(n3518), .B(n8724), .Z(n8725) );
  XOR U9777 ( .A(n8728), .B(n8729), .Z(n8724) );
  ANDN U9778 ( .B(n8730), .A(n3524), .Z(n8728) );
  XNOR U9779 ( .A(n8731), .B(n8732), .Z(n3524) );
  IV U9780 ( .A(n8729), .Z(n8732) );
  XOR U9781 ( .A(n3523), .B(n8729), .Z(n8730) );
  XOR U9782 ( .A(n8733), .B(n8734), .Z(n8729) );
  ANDN U9783 ( .B(n8735), .A(n3529), .Z(n8733) );
  XNOR U9784 ( .A(n8736), .B(n8737), .Z(n3529) );
  IV U9785 ( .A(n8734), .Z(n8737) );
  XOR U9786 ( .A(n3528), .B(n8734), .Z(n8735) );
  XOR U9787 ( .A(n8738), .B(n8739), .Z(n8734) );
  ANDN U9788 ( .B(n8740), .A(n3534), .Z(n8738) );
  XNOR U9789 ( .A(n8741), .B(n8742), .Z(n3534) );
  IV U9790 ( .A(n8739), .Z(n8742) );
  XOR U9791 ( .A(n3533), .B(n8739), .Z(n8740) );
  XOR U9792 ( .A(n8743), .B(n8744), .Z(n8739) );
  ANDN U9793 ( .B(n8745), .A(n3544), .Z(n8743) );
  XNOR U9794 ( .A(n8746), .B(n8747), .Z(n3544) );
  IV U9795 ( .A(n8744), .Z(n8747) );
  XOR U9796 ( .A(n3543), .B(n8744), .Z(n8745) );
  XOR U9797 ( .A(n8748), .B(n8749), .Z(n8744) );
  ANDN U9798 ( .B(n8750), .A(n3549), .Z(n8748) );
  XNOR U9799 ( .A(n8751), .B(n8752), .Z(n3549) );
  IV U9800 ( .A(n8749), .Z(n8752) );
  XOR U9801 ( .A(n3548), .B(n8749), .Z(n8750) );
  XOR U9802 ( .A(n8753), .B(n8754), .Z(n8749) );
  ANDN U9803 ( .B(n8755), .A(n3554), .Z(n8753) );
  XNOR U9804 ( .A(n8756), .B(n8757), .Z(n3554) );
  IV U9805 ( .A(n8754), .Z(n8757) );
  XOR U9806 ( .A(n3553), .B(n8754), .Z(n8755) );
  XOR U9807 ( .A(n8758), .B(n8759), .Z(n8754) );
  ANDN U9808 ( .B(n8760), .A(n3559), .Z(n8758) );
  XNOR U9809 ( .A(n8761), .B(n8762), .Z(n3559) );
  IV U9810 ( .A(n8759), .Z(n8762) );
  XOR U9811 ( .A(n3558), .B(n8759), .Z(n8760) );
  XOR U9812 ( .A(n8763), .B(n8764), .Z(n8759) );
  ANDN U9813 ( .B(n8765), .A(n3564), .Z(n8763) );
  XNOR U9814 ( .A(n8766), .B(n8767), .Z(n3564) );
  IV U9815 ( .A(n8764), .Z(n8767) );
  XOR U9816 ( .A(n3563), .B(n8764), .Z(n8765) );
  XOR U9817 ( .A(n8768), .B(n8769), .Z(n8764) );
  ANDN U9818 ( .B(n8770), .A(n3569), .Z(n8768) );
  XNOR U9819 ( .A(n8771), .B(n8772), .Z(n3569) );
  IV U9820 ( .A(n8769), .Z(n8772) );
  XOR U9821 ( .A(n3568), .B(n8769), .Z(n8770) );
  XOR U9822 ( .A(n8773), .B(n8774), .Z(n8769) );
  ANDN U9823 ( .B(n8775), .A(n3574), .Z(n8773) );
  XNOR U9824 ( .A(n8776), .B(n8777), .Z(n3574) );
  IV U9825 ( .A(n8774), .Z(n8777) );
  XOR U9826 ( .A(n3573), .B(n8774), .Z(n8775) );
  XOR U9827 ( .A(n8778), .B(n8779), .Z(n8774) );
  ANDN U9828 ( .B(n8780), .A(n3579), .Z(n8778) );
  XNOR U9829 ( .A(n8781), .B(n8782), .Z(n3579) );
  IV U9830 ( .A(n8779), .Z(n8782) );
  XOR U9831 ( .A(n3578), .B(n8779), .Z(n8780) );
  XOR U9832 ( .A(n8783), .B(n8784), .Z(n8779) );
  ANDN U9833 ( .B(n8785), .A(n3584), .Z(n8783) );
  XNOR U9834 ( .A(n8786), .B(n8787), .Z(n3584) );
  IV U9835 ( .A(n8784), .Z(n8787) );
  XOR U9836 ( .A(n3583), .B(n8784), .Z(n8785) );
  XOR U9837 ( .A(n8788), .B(n8789), .Z(n8784) );
  ANDN U9838 ( .B(n8790), .A(n3589), .Z(n8788) );
  XNOR U9839 ( .A(n8791), .B(n8792), .Z(n3589) );
  IV U9840 ( .A(n8789), .Z(n8792) );
  XOR U9841 ( .A(n3588), .B(n8789), .Z(n8790) );
  XOR U9842 ( .A(n8793), .B(n8794), .Z(n8789) );
  ANDN U9843 ( .B(n8795), .A(n3599), .Z(n8793) );
  XNOR U9844 ( .A(n8796), .B(n8797), .Z(n3599) );
  IV U9845 ( .A(n8794), .Z(n8797) );
  XOR U9846 ( .A(n3598), .B(n8794), .Z(n8795) );
  XOR U9847 ( .A(n8798), .B(n8799), .Z(n8794) );
  ANDN U9848 ( .B(n8800), .A(n3604), .Z(n8798) );
  XNOR U9849 ( .A(n8801), .B(n8802), .Z(n3604) );
  IV U9850 ( .A(n8799), .Z(n8802) );
  XOR U9851 ( .A(n3603), .B(n8799), .Z(n8800) );
  XOR U9852 ( .A(n8803), .B(n8804), .Z(n8799) );
  ANDN U9853 ( .B(n8805), .A(n3609), .Z(n8803) );
  XNOR U9854 ( .A(n8806), .B(n8807), .Z(n3609) );
  IV U9855 ( .A(n8804), .Z(n8807) );
  XOR U9856 ( .A(n3608), .B(n8804), .Z(n8805) );
  XOR U9857 ( .A(n8808), .B(n8809), .Z(n8804) );
  ANDN U9858 ( .B(n8810), .A(n3614), .Z(n8808) );
  XNOR U9859 ( .A(n8811), .B(n8812), .Z(n3614) );
  IV U9860 ( .A(n8809), .Z(n8812) );
  XOR U9861 ( .A(n3613), .B(n8809), .Z(n8810) );
  XOR U9862 ( .A(n8813), .B(n8814), .Z(n8809) );
  ANDN U9863 ( .B(n8815), .A(n3619), .Z(n8813) );
  XNOR U9864 ( .A(n8816), .B(n8817), .Z(n3619) );
  IV U9865 ( .A(n8814), .Z(n8817) );
  XOR U9866 ( .A(n3618), .B(n8814), .Z(n8815) );
  XOR U9867 ( .A(n8818), .B(n8819), .Z(n8814) );
  ANDN U9868 ( .B(n8820), .A(n3624), .Z(n8818) );
  XNOR U9869 ( .A(n8821), .B(n8822), .Z(n3624) );
  IV U9870 ( .A(n8819), .Z(n8822) );
  XOR U9871 ( .A(n3623), .B(n8819), .Z(n8820) );
  XOR U9872 ( .A(n8823), .B(n8824), .Z(n8819) );
  ANDN U9873 ( .B(n8825), .A(n3629), .Z(n8823) );
  XNOR U9874 ( .A(n8826), .B(n8827), .Z(n3629) );
  IV U9875 ( .A(n8824), .Z(n8827) );
  XOR U9876 ( .A(n3628), .B(n8824), .Z(n8825) );
  XOR U9877 ( .A(n8828), .B(n8829), .Z(n8824) );
  ANDN U9878 ( .B(n8830), .A(n3634), .Z(n8828) );
  XNOR U9879 ( .A(n8831), .B(n8832), .Z(n3634) );
  IV U9880 ( .A(n8829), .Z(n8832) );
  XOR U9881 ( .A(n3633), .B(n8829), .Z(n8830) );
  XOR U9882 ( .A(n8833), .B(n8834), .Z(n8829) );
  ANDN U9883 ( .B(n8835), .A(n3639), .Z(n8833) );
  XNOR U9884 ( .A(n8836), .B(n8837), .Z(n3639) );
  IV U9885 ( .A(n8834), .Z(n8837) );
  XOR U9886 ( .A(n3638), .B(n8834), .Z(n8835) );
  XOR U9887 ( .A(n8838), .B(n8839), .Z(n8834) );
  ANDN U9888 ( .B(n8840), .A(n3644), .Z(n8838) );
  XNOR U9889 ( .A(n8841), .B(n8842), .Z(n3644) );
  IV U9890 ( .A(n8839), .Z(n8842) );
  XOR U9891 ( .A(n3643), .B(n8839), .Z(n8840) );
  XOR U9892 ( .A(n8843), .B(n8844), .Z(n8839) );
  ANDN U9893 ( .B(n8845), .A(n3659), .Z(n8843) );
  XNOR U9894 ( .A(n8846), .B(n8847), .Z(n3659) );
  IV U9895 ( .A(n8844), .Z(n8847) );
  XOR U9896 ( .A(n3658), .B(n8844), .Z(n8845) );
  XOR U9897 ( .A(n8848), .B(n8849), .Z(n8844) );
  ANDN U9898 ( .B(n8850), .A(n3664), .Z(n8848) );
  XNOR U9899 ( .A(n8851), .B(n8852), .Z(n3664) );
  IV U9900 ( .A(n8849), .Z(n8852) );
  XOR U9901 ( .A(n3663), .B(n8849), .Z(n8850) );
  XOR U9902 ( .A(n8853), .B(n8854), .Z(n8849) );
  ANDN U9903 ( .B(n8855), .A(n3669), .Z(n8853) );
  XNOR U9904 ( .A(n8856), .B(n8857), .Z(n3669) );
  IV U9905 ( .A(n8854), .Z(n8857) );
  XOR U9906 ( .A(n3668), .B(n8854), .Z(n8855) );
  XOR U9907 ( .A(n8858), .B(n8859), .Z(n8854) );
  ANDN U9908 ( .B(n8860), .A(n3674), .Z(n8858) );
  XNOR U9909 ( .A(n8861), .B(n8862), .Z(n3674) );
  IV U9910 ( .A(n8859), .Z(n8862) );
  XOR U9911 ( .A(n3673), .B(n8859), .Z(n8860) );
  XOR U9912 ( .A(n8863), .B(n8864), .Z(n8859) );
  ANDN U9913 ( .B(n8865), .A(n3679), .Z(n8863) );
  XNOR U9914 ( .A(n8866), .B(n8867), .Z(n3679) );
  IV U9915 ( .A(n8864), .Z(n8867) );
  XOR U9916 ( .A(n3678), .B(n8864), .Z(n8865) );
  XOR U9917 ( .A(n8868), .B(n8869), .Z(n8864) );
  ANDN U9918 ( .B(n8870), .A(n3684), .Z(n8868) );
  XNOR U9919 ( .A(n8871), .B(n8872), .Z(n3684) );
  IV U9920 ( .A(n8869), .Z(n8872) );
  XOR U9921 ( .A(n3683), .B(n8869), .Z(n8870) );
  XOR U9922 ( .A(n8873), .B(n8874), .Z(n8869) );
  ANDN U9923 ( .B(n8875), .A(n3689), .Z(n8873) );
  XNOR U9924 ( .A(n8876), .B(n8877), .Z(n3689) );
  IV U9925 ( .A(n8874), .Z(n8877) );
  XOR U9926 ( .A(n3688), .B(n8874), .Z(n8875) );
  XOR U9927 ( .A(n8878), .B(n8879), .Z(n8874) );
  ANDN U9928 ( .B(n8880), .A(n3694), .Z(n8878) );
  XNOR U9929 ( .A(n8881), .B(n8882), .Z(n3694) );
  IV U9930 ( .A(n8879), .Z(n8882) );
  XOR U9931 ( .A(n3693), .B(n8879), .Z(n8880) );
  XOR U9932 ( .A(n8883), .B(n8884), .Z(n8879) );
  ANDN U9933 ( .B(n8885), .A(n3699), .Z(n8883) );
  XNOR U9934 ( .A(n8886), .B(n8887), .Z(n3699) );
  IV U9935 ( .A(n8884), .Z(n8887) );
  XOR U9936 ( .A(n3698), .B(n8884), .Z(n8885) );
  XOR U9937 ( .A(n8888), .B(n8889), .Z(n8884) );
  ANDN U9938 ( .B(n8890), .A(n3704), .Z(n8888) );
  XNOR U9939 ( .A(n8891), .B(n8892), .Z(n3704) );
  IV U9940 ( .A(n8889), .Z(n8892) );
  XOR U9941 ( .A(n3703), .B(n8889), .Z(n8890) );
  XOR U9942 ( .A(n8893), .B(n8894), .Z(n8889) );
  ANDN U9943 ( .B(n8895), .A(n3714), .Z(n8893) );
  XNOR U9944 ( .A(n8896), .B(n8897), .Z(n3714) );
  IV U9945 ( .A(n8894), .Z(n8897) );
  XOR U9946 ( .A(n3713), .B(n8894), .Z(n8895) );
  XOR U9947 ( .A(n8898), .B(n8899), .Z(n8894) );
  ANDN U9948 ( .B(n8900), .A(n3719), .Z(n8898) );
  XNOR U9949 ( .A(n8901), .B(n8902), .Z(n3719) );
  IV U9950 ( .A(n8899), .Z(n8902) );
  XOR U9951 ( .A(n3718), .B(n8899), .Z(n8900) );
  XOR U9952 ( .A(n8903), .B(n8904), .Z(n8899) );
  ANDN U9953 ( .B(n8905), .A(n3724), .Z(n8903) );
  XNOR U9954 ( .A(n8906), .B(n8907), .Z(n3724) );
  IV U9955 ( .A(n8904), .Z(n8907) );
  XOR U9956 ( .A(n3723), .B(n8904), .Z(n8905) );
  XOR U9957 ( .A(n8908), .B(n8909), .Z(n8904) );
  ANDN U9958 ( .B(n8910), .A(n3729), .Z(n8908) );
  XNOR U9959 ( .A(n8911), .B(n8912), .Z(n3729) );
  IV U9960 ( .A(n8909), .Z(n8912) );
  XOR U9961 ( .A(n3728), .B(n8909), .Z(n8910) );
  XOR U9962 ( .A(n8913), .B(n8914), .Z(n8909) );
  ANDN U9963 ( .B(n8915), .A(n3734), .Z(n8913) );
  XNOR U9964 ( .A(n8916), .B(n8917), .Z(n3734) );
  IV U9965 ( .A(n8914), .Z(n8917) );
  XOR U9966 ( .A(n3733), .B(n8914), .Z(n8915) );
  XOR U9967 ( .A(n8918), .B(n8919), .Z(n8914) );
  ANDN U9968 ( .B(n8920), .A(n3739), .Z(n8918) );
  XNOR U9969 ( .A(n8921), .B(n8922), .Z(n3739) );
  IV U9970 ( .A(n8919), .Z(n8922) );
  XOR U9971 ( .A(n3738), .B(n8919), .Z(n8920) );
  XOR U9972 ( .A(n8923), .B(n8924), .Z(n8919) );
  ANDN U9973 ( .B(n8925), .A(n3744), .Z(n8923) );
  XNOR U9974 ( .A(n8926), .B(n8927), .Z(n3744) );
  IV U9975 ( .A(n8924), .Z(n8927) );
  XOR U9976 ( .A(n3743), .B(n8924), .Z(n8925) );
  XOR U9977 ( .A(n8928), .B(n8929), .Z(n8924) );
  ANDN U9978 ( .B(n8930), .A(n3749), .Z(n8928) );
  XNOR U9979 ( .A(n8931), .B(n8932), .Z(n3749) );
  IV U9980 ( .A(n8929), .Z(n8932) );
  XOR U9981 ( .A(n3748), .B(n8929), .Z(n8930) );
  XOR U9982 ( .A(n8933), .B(n8934), .Z(n8929) );
  ANDN U9983 ( .B(n8935), .A(n3754), .Z(n8933) );
  XNOR U9984 ( .A(n8936), .B(n8937), .Z(n3754) );
  IV U9985 ( .A(n8934), .Z(n8937) );
  XOR U9986 ( .A(n3753), .B(n8934), .Z(n8935) );
  XOR U9987 ( .A(n8938), .B(n8939), .Z(n8934) );
  ANDN U9988 ( .B(n8940), .A(n3759), .Z(n8938) );
  XNOR U9989 ( .A(n8941), .B(n8942), .Z(n3759) );
  IV U9990 ( .A(n8939), .Z(n8942) );
  XOR U9991 ( .A(n3758), .B(n8939), .Z(n8940) );
  XOR U9992 ( .A(n8943), .B(n8944), .Z(n8939) );
  ANDN U9993 ( .B(n8945), .A(n3769), .Z(n8943) );
  XNOR U9994 ( .A(n8946), .B(n8947), .Z(n3769) );
  IV U9995 ( .A(n8944), .Z(n8947) );
  XOR U9996 ( .A(n3768), .B(n8944), .Z(n8945) );
  XOR U9997 ( .A(n8948), .B(n8949), .Z(n8944) );
  ANDN U9998 ( .B(n8950), .A(n3774), .Z(n8948) );
  XNOR U9999 ( .A(n8951), .B(n8952), .Z(n3774) );
  IV U10000 ( .A(n8949), .Z(n8952) );
  XOR U10001 ( .A(n3773), .B(n8949), .Z(n8950) );
  XOR U10002 ( .A(n8953), .B(n8954), .Z(n8949) );
  ANDN U10003 ( .B(n8955), .A(n3779), .Z(n8953) );
  XNOR U10004 ( .A(n8956), .B(n8957), .Z(n3779) );
  IV U10005 ( .A(n8954), .Z(n8957) );
  XOR U10006 ( .A(n3778), .B(n8954), .Z(n8955) );
  XOR U10007 ( .A(n8958), .B(n8959), .Z(n8954) );
  ANDN U10008 ( .B(n8960), .A(n3784), .Z(n8958) );
  XNOR U10009 ( .A(n8961), .B(n8962), .Z(n3784) );
  IV U10010 ( .A(n8959), .Z(n8962) );
  XOR U10011 ( .A(n3783), .B(n8959), .Z(n8960) );
  XOR U10012 ( .A(n8963), .B(n8964), .Z(n8959) );
  ANDN U10013 ( .B(n8965), .A(n3789), .Z(n8963) );
  XNOR U10014 ( .A(n8966), .B(n8967), .Z(n3789) );
  IV U10015 ( .A(n8964), .Z(n8967) );
  XOR U10016 ( .A(n3788), .B(n8964), .Z(n8965) );
  XOR U10017 ( .A(n8968), .B(n8969), .Z(n8964) );
  ANDN U10018 ( .B(n8970), .A(n3794), .Z(n8968) );
  XNOR U10019 ( .A(n8971), .B(n8972), .Z(n3794) );
  IV U10020 ( .A(n8969), .Z(n8972) );
  XOR U10021 ( .A(n3793), .B(n8969), .Z(n8970) );
  XOR U10022 ( .A(n8973), .B(n8974), .Z(n8969) );
  ANDN U10023 ( .B(n8975), .A(n3799), .Z(n8973) );
  XNOR U10024 ( .A(n8976), .B(n8977), .Z(n3799) );
  IV U10025 ( .A(n8974), .Z(n8977) );
  XOR U10026 ( .A(n3798), .B(n8974), .Z(n8975) );
  XOR U10027 ( .A(n8978), .B(n8979), .Z(n8974) );
  ANDN U10028 ( .B(n8980), .A(n3804), .Z(n8978) );
  XNOR U10029 ( .A(n8981), .B(n8982), .Z(n3804) );
  IV U10030 ( .A(n8979), .Z(n8982) );
  XOR U10031 ( .A(n3803), .B(n8979), .Z(n8980) );
  XOR U10032 ( .A(n8983), .B(n8984), .Z(n8979) );
  ANDN U10033 ( .B(n8985), .A(n3809), .Z(n8983) );
  XNOR U10034 ( .A(n8986), .B(n8987), .Z(n3809) );
  IV U10035 ( .A(n8984), .Z(n8987) );
  XOR U10036 ( .A(n3808), .B(n8984), .Z(n8985) );
  XOR U10037 ( .A(n8988), .B(n8989), .Z(n8984) );
  ANDN U10038 ( .B(n8990), .A(n3814), .Z(n8988) );
  XNOR U10039 ( .A(n8991), .B(n8992), .Z(n3814) );
  IV U10040 ( .A(n8989), .Z(n8992) );
  XOR U10041 ( .A(n3813), .B(n8989), .Z(n8990) );
  XOR U10042 ( .A(n8993), .B(n8994), .Z(n8989) );
  ANDN U10043 ( .B(n8995), .A(n3824), .Z(n8993) );
  XNOR U10044 ( .A(n8996), .B(n8997), .Z(n3824) );
  IV U10045 ( .A(n8994), .Z(n8997) );
  XOR U10046 ( .A(n3823), .B(n8994), .Z(n8995) );
  XOR U10047 ( .A(n8998), .B(n8999), .Z(n8994) );
  ANDN U10048 ( .B(n9000), .A(n3829), .Z(n8998) );
  XNOR U10049 ( .A(n9001), .B(n9002), .Z(n3829) );
  IV U10050 ( .A(n8999), .Z(n9002) );
  XOR U10051 ( .A(n3828), .B(n8999), .Z(n9000) );
  XOR U10052 ( .A(n9003), .B(n9004), .Z(n8999) );
  ANDN U10053 ( .B(n9005), .A(n3834), .Z(n9003) );
  XNOR U10054 ( .A(n9006), .B(n9007), .Z(n3834) );
  IV U10055 ( .A(n9004), .Z(n9007) );
  XOR U10056 ( .A(n3833), .B(n9004), .Z(n9005) );
  XOR U10057 ( .A(n9008), .B(n9009), .Z(n9004) );
  ANDN U10058 ( .B(n9010), .A(n3839), .Z(n9008) );
  XNOR U10059 ( .A(n9011), .B(n9012), .Z(n3839) );
  IV U10060 ( .A(n9009), .Z(n9012) );
  XOR U10061 ( .A(n3838), .B(n9009), .Z(n9010) );
  XOR U10062 ( .A(n9013), .B(n9014), .Z(n9009) );
  ANDN U10063 ( .B(n9015), .A(n3844), .Z(n9013) );
  XNOR U10064 ( .A(n9016), .B(n9017), .Z(n3844) );
  IV U10065 ( .A(n9014), .Z(n9017) );
  XOR U10066 ( .A(n3843), .B(n9014), .Z(n9015) );
  XOR U10067 ( .A(n9018), .B(n9019), .Z(n9014) );
  ANDN U10068 ( .B(n9020), .A(n3849), .Z(n9018) );
  XNOR U10069 ( .A(n9021), .B(n9022), .Z(n3849) );
  IV U10070 ( .A(n9019), .Z(n9022) );
  XOR U10071 ( .A(n3848), .B(n9019), .Z(n9020) );
  XOR U10072 ( .A(n9023), .B(n9024), .Z(n9019) );
  ANDN U10073 ( .B(n9025), .A(n3854), .Z(n9023) );
  XNOR U10074 ( .A(n9026), .B(n9027), .Z(n3854) );
  IV U10075 ( .A(n9024), .Z(n9027) );
  XOR U10076 ( .A(n3853), .B(n9024), .Z(n9025) );
  XOR U10077 ( .A(n9028), .B(n9029), .Z(n9024) );
  ANDN U10078 ( .B(n9030), .A(n3859), .Z(n9028) );
  XNOR U10079 ( .A(n9031), .B(n9032), .Z(n3859) );
  IV U10080 ( .A(n9029), .Z(n9032) );
  XOR U10081 ( .A(n3858), .B(n9029), .Z(n9030) );
  XOR U10082 ( .A(n9033), .B(n9034), .Z(n9029) );
  ANDN U10083 ( .B(n9035), .A(n3864), .Z(n9033) );
  XNOR U10084 ( .A(n9036), .B(n9037), .Z(n3864) );
  IV U10085 ( .A(n9034), .Z(n9037) );
  XOR U10086 ( .A(n3863), .B(n9034), .Z(n9035) );
  XOR U10087 ( .A(n9038), .B(n9039), .Z(n9034) );
  ANDN U10088 ( .B(n9040), .A(n3869), .Z(n9038) );
  XNOR U10089 ( .A(n9041), .B(n9042), .Z(n3869) );
  IV U10090 ( .A(n9039), .Z(n9042) );
  XOR U10091 ( .A(n3868), .B(n9039), .Z(n9040) );
  XOR U10092 ( .A(n9043), .B(n9044), .Z(n9039) );
  ANDN U10093 ( .B(n9045), .A(n3879), .Z(n9043) );
  XNOR U10094 ( .A(n9046), .B(n9047), .Z(n3879) );
  IV U10095 ( .A(n9044), .Z(n9047) );
  XOR U10096 ( .A(n3878), .B(n9044), .Z(n9045) );
  XOR U10097 ( .A(n9048), .B(n9049), .Z(n9044) );
  ANDN U10098 ( .B(n9050), .A(n3884), .Z(n9048) );
  XNOR U10099 ( .A(n9051), .B(n9052), .Z(n3884) );
  IV U10100 ( .A(n9049), .Z(n9052) );
  XOR U10101 ( .A(n3883), .B(n9049), .Z(n9050) );
  XOR U10102 ( .A(n9053), .B(n9054), .Z(n9049) );
  ANDN U10103 ( .B(n9055), .A(n3889), .Z(n9053) );
  XNOR U10104 ( .A(n9056), .B(n9057), .Z(n3889) );
  IV U10105 ( .A(n9054), .Z(n9057) );
  XOR U10106 ( .A(n3888), .B(n9054), .Z(n9055) );
  XOR U10107 ( .A(n9058), .B(n9059), .Z(n9054) );
  ANDN U10108 ( .B(n9060), .A(n3894), .Z(n9058) );
  XNOR U10109 ( .A(n9061), .B(n9062), .Z(n3894) );
  IV U10110 ( .A(n9059), .Z(n9062) );
  XOR U10111 ( .A(n3893), .B(n9059), .Z(n9060) );
  XOR U10112 ( .A(n9063), .B(n9064), .Z(n9059) );
  ANDN U10113 ( .B(n9065), .A(n3899), .Z(n9063) );
  XNOR U10114 ( .A(n9066), .B(n9067), .Z(n3899) );
  IV U10115 ( .A(n9064), .Z(n9067) );
  XOR U10116 ( .A(n3898), .B(n9064), .Z(n9065) );
  XOR U10117 ( .A(n9068), .B(n9069), .Z(n9064) );
  ANDN U10118 ( .B(n9070), .A(n3904), .Z(n9068) );
  XNOR U10119 ( .A(n9071), .B(n9072), .Z(n3904) );
  IV U10120 ( .A(n9069), .Z(n9072) );
  XOR U10121 ( .A(n3903), .B(n9069), .Z(n9070) );
  XOR U10122 ( .A(n9073), .B(n9074), .Z(n9069) );
  ANDN U10123 ( .B(n9075), .A(n3909), .Z(n9073) );
  XNOR U10124 ( .A(n9076), .B(n9077), .Z(n3909) );
  IV U10125 ( .A(n9074), .Z(n9077) );
  XOR U10126 ( .A(n3908), .B(n9074), .Z(n9075) );
  XOR U10127 ( .A(n9078), .B(n9079), .Z(n9074) );
  ANDN U10128 ( .B(n9080), .A(n3914), .Z(n9078) );
  XNOR U10129 ( .A(n9081), .B(n9082), .Z(n3914) );
  IV U10130 ( .A(n9079), .Z(n9082) );
  XOR U10131 ( .A(n3913), .B(n9079), .Z(n9080) );
  XOR U10132 ( .A(n9083), .B(n9084), .Z(n9079) );
  ANDN U10133 ( .B(n9085), .A(n3919), .Z(n9083) );
  XNOR U10134 ( .A(n9086), .B(n9087), .Z(n3919) );
  IV U10135 ( .A(n9084), .Z(n9087) );
  XOR U10136 ( .A(n3918), .B(n9084), .Z(n9085) );
  XOR U10137 ( .A(n9088), .B(n9089), .Z(n9084) );
  ANDN U10138 ( .B(n9090), .A(n3924), .Z(n9088) );
  XNOR U10139 ( .A(n9091), .B(n9092), .Z(n3924) );
  IV U10140 ( .A(n9089), .Z(n9092) );
  XOR U10141 ( .A(n3923), .B(n9089), .Z(n9090) );
  XOR U10142 ( .A(n9093), .B(n9094), .Z(n9089) );
  ANDN U10143 ( .B(n9095), .A(n3934), .Z(n9093) );
  XNOR U10144 ( .A(n9096), .B(n9097), .Z(n3934) );
  IV U10145 ( .A(n9094), .Z(n9097) );
  XOR U10146 ( .A(n3933), .B(n9094), .Z(n9095) );
  XOR U10147 ( .A(n9098), .B(n9099), .Z(n9094) );
  ANDN U10148 ( .B(n9100), .A(n3939), .Z(n9098) );
  XNOR U10149 ( .A(n9101), .B(n9102), .Z(n3939) );
  IV U10150 ( .A(n9099), .Z(n9102) );
  XOR U10151 ( .A(n3938), .B(n9099), .Z(n9100) );
  XOR U10152 ( .A(n9103), .B(n9104), .Z(n9099) );
  ANDN U10153 ( .B(n9105), .A(n3944), .Z(n9103) );
  XNOR U10154 ( .A(n9106), .B(n9107), .Z(n3944) );
  IV U10155 ( .A(n9104), .Z(n9107) );
  XOR U10156 ( .A(n3943), .B(n9104), .Z(n9105) );
  XOR U10157 ( .A(n9108), .B(n9109), .Z(n9104) );
  ANDN U10158 ( .B(n9110), .A(n3949), .Z(n9108) );
  XNOR U10159 ( .A(n9111), .B(n9112), .Z(n3949) );
  IV U10160 ( .A(n9109), .Z(n9112) );
  XOR U10161 ( .A(n3948), .B(n9109), .Z(n9110) );
  XOR U10162 ( .A(n9113), .B(n9114), .Z(n9109) );
  ANDN U10163 ( .B(n9115), .A(n3954), .Z(n9113) );
  XNOR U10164 ( .A(n9116), .B(n9117), .Z(n3954) );
  IV U10165 ( .A(n9114), .Z(n9117) );
  XOR U10166 ( .A(n3953), .B(n9114), .Z(n9115) );
  XOR U10167 ( .A(n9118), .B(n9119), .Z(n9114) );
  ANDN U10168 ( .B(n9120), .A(n3959), .Z(n9118) );
  XNOR U10169 ( .A(n9121), .B(n9122), .Z(n3959) );
  IV U10170 ( .A(n9119), .Z(n9122) );
  XOR U10171 ( .A(n3958), .B(n9119), .Z(n9120) );
  XOR U10172 ( .A(n9123), .B(n9124), .Z(n9119) );
  ANDN U10173 ( .B(n9125), .A(n3964), .Z(n9123) );
  XNOR U10174 ( .A(n9126), .B(n9127), .Z(n3964) );
  IV U10175 ( .A(n9124), .Z(n9127) );
  XOR U10176 ( .A(n3963), .B(n9124), .Z(n9125) );
  XOR U10177 ( .A(n9128), .B(n9129), .Z(n9124) );
  ANDN U10178 ( .B(n9130), .A(n3969), .Z(n9128) );
  XNOR U10179 ( .A(n9131), .B(n9132), .Z(n3969) );
  IV U10180 ( .A(n9129), .Z(n9132) );
  XOR U10181 ( .A(n3968), .B(n9129), .Z(n9130) );
  XOR U10182 ( .A(n9133), .B(n9134), .Z(n9129) );
  ANDN U10183 ( .B(n9135), .A(n3974), .Z(n9133) );
  XNOR U10184 ( .A(n9136), .B(n9137), .Z(n3974) );
  IV U10185 ( .A(n9134), .Z(n9137) );
  XOR U10186 ( .A(n3973), .B(n9134), .Z(n9135) );
  XOR U10187 ( .A(n9138), .B(n9139), .Z(n9134) );
  ANDN U10188 ( .B(n9140), .A(n3979), .Z(n9138) );
  XNOR U10189 ( .A(n9141), .B(n9142), .Z(n3979) );
  IV U10190 ( .A(n9139), .Z(n9142) );
  XOR U10191 ( .A(n3978), .B(n9139), .Z(n9140) );
  XOR U10192 ( .A(n9143), .B(n9144), .Z(n9139) );
  ANDN U10193 ( .B(n9145), .A(n3989), .Z(n9143) );
  XNOR U10194 ( .A(n9146), .B(n9147), .Z(n3989) );
  IV U10195 ( .A(n9144), .Z(n9147) );
  XOR U10196 ( .A(n3988), .B(n9144), .Z(n9145) );
  XOR U10197 ( .A(n9148), .B(n9149), .Z(n9144) );
  ANDN U10198 ( .B(n9150), .A(n3994), .Z(n9148) );
  XNOR U10199 ( .A(n9151), .B(n9152), .Z(n3994) );
  IV U10200 ( .A(n9149), .Z(n9152) );
  XOR U10201 ( .A(n3993), .B(n9149), .Z(n9150) );
  XOR U10202 ( .A(n9153), .B(n9154), .Z(n9149) );
  ANDN U10203 ( .B(n9155), .A(n3999), .Z(n9153) );
  XNOR U10204 ( .A(n9156), .B(n9157), .Z(n3999) );
  IV U10205 ( .A(n9154), .Z(n9157) );
  XOR U10206 ( .A(n3998), .B(n9154), .Z(n9155) );
  XOR U10207 ( .A(n9158), .B(n9159), .Z(n9154) );
  ANDN U10208 ( .B(n9160), .A(n4004), .Z(n9158) );
  XNOR U10209 ( .A(n9161), .B(n9162), .Z(n4004) );
  IV U10210 ( .A(n9159), .Z(n9162) );
  XOR U10211 ( .A(n4003), .B(n9159), .Z(n9160) );
  XOR U10212 ( .A(n9163), .B(n9164), .Z(n9159) );
  ANDN U10213 ( .B(n9165), .A(n4009), .Z(n9163) );
  XNOR U10214 ( .A(n9166), .B(n9167), .Z(n4009) );
  IV U10215 ( .A(n9164), .Z(n9167) );
  XOR U10216 ( .A(n4008), .B(n9164), .Z(n9165) );
  XOR U10217 ( .A(n9168), .B(n9169), .Z(n9164) );
  ANDN U10218 ( .B(n9170), .A(n4014), .Z(n9168) );
  XNOR U10219 ( .A(n9171), .B(n9172), .Z(n4014) );
  IV U10220 ( .A(n9169), .Z(n9172) );
  XOR U10221 ( .A(n4013), .B(n9169), .Z(n9170) );
  XOR U10222 ( .A(n9173), .B(n9174), .Z(n9169) );
  ANDN U10223 ( .B(n9175), .A(n4019), .Z(n9173) );
  XNOR U10224 ( .A(n9176), .B(n9177), .Z(n4019) );
  IV U10225 ( .A(n9174), .Z(n9177) );
  XOR U10226 ( .A(n4018), .B(n9174), .Z(n9175) );
  XOR U10227 ( .A(n9178), .B(n9179), .Z(n9174) );
  ANDN U10228 ( .B(n9180), .A(n4024), .Z(n9178) );
  XNOR U10229 ( .A(n9181), .B(n9182), .Z(n4024) );
  IV U10230 ( .A(n9179), .Z(n9182) );
  XOR U10231 ( .A(n4023), .B(n9179), .Z(n9180) );
  XOR U10232 ( .A(n9183), .B(n9184), .Z(n9179) );
  ANDN U10233 ( .B(n9185), .A(n4029), .Z(n9183) );
  XNOR U10234 ( .A(n9186), .B(n9187), .Z(n4029) );
  IV U10235 ( .A(n9184), .Z(n9187) );
  XOR U10236 ( .A(n4028), .B(n9184), .Z(n9185) );
  XOR U10237 ( .A(n9188), .B(n9189), .Z(n9184) );
  ANDN U10238 ( .B(n9190), .A(n4034), .Z(n9188) );
  XNOR U10239 ( .A(n9191), .B(n9192), .Z(n4034) );
  IV U10240 ( .A(n9189), .Z(n9192) );
  XOR U10241 ( .A(n4033), .B(n9189), .Z(n9190) );
  XOR U10242 ( .A(n9193), .B(n9194), .Z(n9189) );
  ANDN U10243 ( .B(n9195), .A(n4044), .Z(n9193) );
  XNOR U10244 ( .A(n9196), .B(n9197), .Z(n4044) );
  IV U10245 ( .A(n9194), .Z(n9197) );
  XOR U10246 ( .A(n4043), .B(n9194), .Z(n9195) );
  XOR U10247 ( .A(n9198), .B(n9199), .Z(n9194) );
  ANDN U10248 ( .B(n9200), .A(n4049), .Z(n9198) );
  XNOR U10249 ( .A(n9201), .B(n9202), .Z(n4049) );
  IV U10250 ( .A(n9199), .Z(n9202) );
  XOR U10251 ( .A(n4048), .B(n9199), .Z(n9200) );
  XOR U10252 ( .A(n9203), .B(n9204), .Z(n9199) );
  ANDN U10253 ( .B(n9205), .A(n4054), .Z(n9203) );
  XNOR U10254 ( .A(n9206), .B(n9207), .Z(n4054) );
  IV U10255 ( .A(n9204), .Z(n9207) );
  XOR U10256 ( .A(n4053), .B(n9204), .Z(n9205) );
  XOR U10257 ( .A(n9208), .B(n9209), .Z(n9204) );
  ANDN U10258 ( .B(n9210), .A(n4059), .Z(n9208) );
  XNOR U10259 ( .A(n9211), .B(n9212), .Z(n4059) );
  IV U10260 ( .A(n9209), .Z(n9212) );
  XOR U10261 ( .A(n4058), .B(n9209), .Z(n9210) );
  XOR U10262 ( .A(n9213), .B(n9214), .Z(n9209) );
  ANDN U10263 ( .B(n9215), .A(n4064), .Z(n9213) );
  XNOR U10264 ( .A(n9216), .B(n9217), .Z(n4064) );
  IV U10265 ( .A(n9214), .Z(n9217) );
  XOR U10266 ( .A(n4063), .B(n9214), .Z(n9215) );
  XOR U10267 ( .A(n9218), .B(n9219), .Z(n9214) );
  ANDN U10268 ( .B(n9220), .A(n4069), .Z(n9218) );
  XNOR U10269 ( .A(n9221), .B(n9222), .Z(n4069) );
  IV U10270 ( .A(n9219), .Z(n9222) );
  XOR U10271 ( .A(n4068), .B(n9219), .Z(n9220) );
  XOR U10272 ( .A(n9223), .B(n9224), .Z(n9219) );
  ANDN U10273 ( .B(n9225), .A(n4074), .Z(n9223) );
  XNOR U10274 ( .A(n9226), .B(n9227), .Z(n4074) );
  IV U10275 ( .A(n9224), .Z(n9227) );
  XOR U10276 ( .A(n4073), .B(n9224), .Z(n9225) );
  XOR U10277 ( .A(n9228), .B(n9229), .Z(n9224) );
  ANDN U10278 ( .B(n9230), .A(n4079), .Z(n9228) );
  XNOR U10279 ( .A(n9231), .B(n9232), .Z(n4079) );
  IV U10280 ( .A(n9229), .Z(n9232) );
  XOR U10281 ( .A(n4078), .B(n9229), .Z(n9230) );
  XOR U10282 ( .A(n9233), .B(n9234), .Z(n9229) );
  ANDN U10283 ( .B(n9235), .A(n4084), .Z(n9233) );
  XNOR U10284 ( .A(n9236), .B(n9237), .Z(n4084) );
  IV U10285 ( .A(n9234), .Z(n9237) );
  XOR U10286 ( .A(n4083), .B(n9234), .Z(n9235) );
  XOR U10287 ( .A(n9238), .B(n9239), .Z(n9234) );
  ANDN U10288 ( .B(n9240), .A(n4089), .Z(n9238) );
  XNOR U10289 ( .A(n9241), .B(n9242), .Z(n4089) );
  IV U10290 ( .A(n9239), .Z(n9242) );
  XOR U10291 ( .A(n4088), .B(n9239), .Z(n9240) );
  XOR U10292 ( .A(n9243), .B(n9244), .Z(n9239) );
  ANDN U10293 ( .B(n9245), .A(n4099), .Z(n9243) );
  XNOR U10294 ( .A(n9246), .B(n9247), .Z(n4099) );
  IV U10295 ( .A(n9244), .Z(n9247) );
  XOR U10296 ( .A(n4098), .B(n9244), .Z(n9245) );
  XOR U10297 ( .A(n9248), .B(n9249), .Z(n9244) );
  ANDN U10298 ( .B(n9250), .A(n4104), .Z(n9248) );
  XNOR U10299 ( .A(n9251), .B(n9252), .Z(n4104) );
  IV U10300 ( .A(n9249), .Z(n9252) );
  XOR U10301 ( .A(n4103), .B(n9249), .Z(n9250) );
  XOR U10302 ( .A(n9253), .B(n9254), .Z(n9249) );
  ANDN U10303 ( .B(n9255), .A(n4109), .Z(n9253) );
  XNOR U10304 ( .A(n9256), .B(n9257), .Z(n4109) );
  IV U10305 ( .A(n9254), .Z(n9257) );
  XOR U10306 ( .A(n4108), .B(n9254), .Z(n9255) );
  XOR U10307 ( .A(n9258), .B(n9259), .Z(n9254) );
  ANDN U10308 ( .B(n9260), .A(n4114), .Z(n9258) );
  XNOR U10309 ( .A(n9261), .B(n9262), .Z(n4114) );
  IV U10310 ( .A(n9259), .Z(n9262) );
  XOR U10311 ( .A(n4113), .B(n9259), .Z(n9260) );
  XOR U10312 ( .A(n9263), .B(n9264), .Z(n9259) );
  ANDN U10313 ( .B(n9265), .A(n4119), .Z(n9263) );
  XNOR U10314 ( .A(n9266), .B(n9267), .Z(n4119) );
  IV U10315 ( .A(n9264), .Z(n9267) );
  XOR U10316 ( .A(n4118), .B(n9264), .Z(n9265) );
  XOR U10317 ( .A(n9268), .B(n9269), .Z(n9264) );
  ANDN U10318 ( .B(n9270), .A(n4124), .Z(n9268) );
  XNOR U10319 ( .A(n9271), .B(n9272), .Z(n4124) );
  IV U10320 ( .A(n9269), .Z(n9272) );
  XOR U10321 ( .A(n4123), .B(n9269), .Z(n9270) );
  XOR U10322 ( .A(n9273), .B(n9274), .Z(n9269) );
  ANDN U10323 ( .B(n9275), .A(n4129), .Z(n9273) );
  XNOR U10324 ( .A(n9276), .B(n9277), .Z(n4129) );
  IV U10325 ( .A(n9274), .Z(n9277) );
  XOR U10326 ( .A(n4128), .B(n9274), .Z(n9275) );
  XOR U10327 ( .A(n9278), .B(n9279), .Z(n9274) );
  ANDN U10328 ( .B(n9280), .A(n4134), .Z(n9278) );
  XNOR U10329 ( .A(n9281), .B(n9282), .Z(n4134) );
  IV U10330 ( .A(n9279), .Z(n9282) );
  XOR U10331 ( .A(n4133), .B(n9279), .Z(n9280) );
  XOR U10332 ( .A(n9283), .B(n9284), .Z(n9279) );
  ANDN U10333 ( .B(n9285), .A(n4139), .Z(n9283) );
  XNOR U10334 ( .A(n9286), .B(n9287), .Z(n4139) );
  IV U10335 ( .A(n9284), .Z(n9287) );
  XOR U10336 ( .A(n4138), .B(n9284), .Z(n9285) );
  XOR U10337 ( .A(n9288), .B(n9289), .Z(n9284) );
  ANDN U10338 ( .B(n9290), .A(n4144), .Z(n9288) );
  XNOR U10339 ( .A(n9291), .B(n9292), .Z(n4144) );
  IV U10340 ( .A(n9289), .Z(n9292) );
  XOR U10341 ( .A(n4143), .B(n9289), .Z(n9290) );
  XOR U10342 ( .A(n9293), .B(n9294), .Z(n9289) );
  ANDN U10343 ( .B(n9295), .A(n4154), .Z(n9293) );
  XNOR U10344 ( .A(n9296), .B(n9297), .Z(n4154) );
  IV U10345 ( .A(n9294), .Z(n9297) );
  XOR U10346 ( .A(n4153), .B(n9294), .Z(n9295) );
  XOR U10347 ( .A(n9298), .B(n9299), .Z(n9294) );
  ANDN U10348 ( .B(n9300), .A(n4159), .Z(n9298) );
  XNOR U10349 ( .A(n9301), .B(n9302), .Z(n4159) );
  IV U10350 ( .A(n9299), .Z(n9302) );
  XOR U10351 ( .A(n4158), .B(n9299), .Z(n9300) );
  XOR U10352 ( .A(n9303), .B(n9304), .Z(n9299) );
  ANDN U10353 ( .B(n9305), .A(n4164), .Z(n9303) );
  XNOR U10354 ( .A(n9306), .B(n9307), .Z(n4164) );
  IV U10355 ( .A(n9304), .Z(n9307) );
  XOR U10356 ( .A(n4163), .B(n9304), .Z(n9305) );
  XOR U10357 ( .A(n9308), .B(n9309), .Z(n9304) );
  ANDN U10358 ( .B(n9310), .A(n4169), .Z(n9308) );
  XNOR U10359 ( .A(n9311), .B(n9312), .Z(n4169) );
  IV U10360 ( .A(n9309), .Z(n9312) );
  XOR U10361 ( .A(n4168), .B(n9309), .Z(n9310) );
  XOR U10362 ( .A(n9313), .B(n9314), .Z(n9309) );
  ANDN U10363 ( .B(n9315), .A(n4174), .Z(n9313) );
  XNOR U10364 ( .A(n9316), .B(n9317), .Z(n4174) );
  IV U10365 ( .A(n9314), .Z(n9317) );
  XOR U10366 ( .A(n4173), .B(n9314), .Z(n9315) );
  XOR U10367 ( .A(n9318), .B(n9319), .Z(n9314) );
  ANDN U10368 ( .B(n9320), .A(n4179), .Z(n9318) );
  XNOR U10369 ( .A(n9321), .B(n9322), .Z(n4179) );
  IV U10370 ( .A(n9319), .Z(n9322) );
  XOR U10371 ( .A(n4178), .B(n9319), .Z(n9320) );
  XOR U10372 ( .A(n9323), .B(n9324), .Z(n9319) );
  ANDN U10373 ( .B(n9325), .A(n4184), .Z(n9323) );
  XNOR U10374 ( .A(n9326), .B(n9327), .Z(n4184) );
  IV U10375 ( .A(n9324), .Z(n9327) );
  XOR U10376 ( .A(n4183), .B(n9324), .Z(n9325) );
  XOR U10377 ( .A(n9328), .B(n9329), .Z(n9324) );
  ANDN U10378 ( .B(n9330), .A(n4189), .Z(n9328) );
  XNOR U10379 ( .A(n9331), .B(n9332), .Z(n4189) );
  IV U10380 ( .A(n9329), .Z(n9332) );
  XOR U10381 ( .A(n4188), .B(n9329), .Z(n9330) );
  XOR U10382 ( .A(n9333), .B(n9334), .Z(n9329) );
  ANDN U10383 ( .B(n9335), .A(n4194), .Z(n9333) );
  XNOR U10384 ( .A(n9336), .B(n9337), .Z(n4194) );
  IV U10385 ( .A(n9334), .Z(n9337) );
  XOR U10386 ( .A(n4193), .B(n9334), .Z(n9335) );
  XOR U10387 ( .A(n9338), .B(n9339), .Z(n9334) );
  ANDN U10388 ( .B(n9340), .A(n4199), .Z(n9338) );
  XNOR U10389 ( .A(n9341), .B(n9342), .Z(n4199) );
  IV U10390 ( .A(n9339), .Z(n9342) );
  XOR U10391 ( .A(n4198), .B(n9339), .Z(n9340) );
  XOR U10392 ( .A(n9343), .B(n9344), .Z(n9339) );
  ANDN U10393 ( .B(n9345), .A(n4214), .Z(n9343) );
  XNOR U10394 ( .A(n9346), .B(n9347), .Z(n4214) );
  IV U10395 ( .A(n9344), .Z(n9347) );
  XOR U10396 ( .A(n4213), .B(n9344), .Z(n9345) );
  XOR U10397 ( .A(n9348), .B(n9349), .Z(n9344) );
  ANDN U10398 ( .B(n9350), .A(n4219), .Z(n9348) );
  XNOR U10399 ( .A(n9351), .B(n9352), .Z(n4219) );
  IV U10400 ( .A(n9349), .Z(n9352) );
  XOR U10401 ( .A(n4218), .B(n9349), .Z(n9350) );
  XOR U10402 ( .A(n9353), .B(n9354), .Z(n9349) );
  ANDN U10403 ( .B(n9355), .A(n4224), .Z(n9353) );
  XNOR U10404 ( .A(n9356), .B(n9357), .Z(n4224) );
  IV U10405 ( .A(n9354), .Z(n9357) );
  XOR U10406 ( .A(n4223), .B(n9354), .Z(n9355) );
  XOR U10407 ( .A(n9358), .B(n9359), .Z(n9354) );
  ANDN U10408 ( .B(n9360), .A(n4229), .Z(n9358) );
  XNOR U10409 ( .A(n9361), .B(n9362), .Z(n4229) );
  IV U10410 ( .A(n9359), .Z(n9362) );
  XOR U10411 ( .A(n4228), .B(n9359), .Z(n9360) );
  XOR U10412 ( .A(n9363), .B(n9364), .Z(n9359) );
  ANDN U10413 ( .B(n9365), .A(n4234), .Z(n9363) );
  XNOR U10414 ( .A(n9366), .B(n9367), .Z(n4234) );
  IV U10415 ( .A(n9364), .Z(n9367) );
  XOR U10416 ( .A(n4233), .B(n9364), .Z(n9365) );
  XOR U10417 ( .A(n9368), .B(n9369), .Z(n9364) );
  ANDN U10418 ( .B(n9370), .A(n4239), .Z(n9368) );
  XNOR U10419 ( .A(n9371), .B(n9372), .Z(n4239) );
  IV U10420 ( .A(n9369), .Z(n9372) );
  XOR U10421 ( .A(n4238), .B(n9369), .Z(n9370) );
  XOR U10422 ( .A(n9373), .B(n9374), .Z(n9369) );
  ANDN U10423 ( .B(n9375), .A(n4244), .Z(n9373) );
  XNOR U10424 ( .A(n9376), .B(n9377), .Z(n4244) );
  IV U10425 ( .A(n9374), .Z(n9377) );
  XOR U10426 ( .A(n4243), .B(n9374), .Z(n9375) );
  XOR U10427 ( .A(n9378), .B(n9379), .Z(n9374) );
  ANDN U10428 ( .B(n9380), .A(n4249), .Z(n9378) );
  XNOR U10429 ( .A(n9381), .B(n9382), .Z(n4249) );
  IV U10430 ( .A(n9379), .Z(n9382) );
  XOR U10431 ( .A(n4248), .B(n9379), .Z(n9380) );
  XOR U10432 ( .A(n9383), .B(n9384), .Z(n9379) );
  ANDN U10433 ( .B(n9385), .A(n4254), .Z(n9383) );
  XNOR U10434 ( .A(n9386), .B(n9387), .Z(n4254) );
  IV U10435 ( .A(n9384), .Z(n9387) );
  XOR U10436 ( .A(n4253), .B(n9384), .Z(n9385) );
  XOR U10437 ( .A(n9388), .B(n9389), .Z(n9384) );
  ANDN U10438 ( .B(n9390), .A(n4259), .Z(n9388) );
  XNOR U10439 ( .A(n9391), .B(n9392), .Z(n4259) );
  IV U10440 ( .A(n9389), .Z(n9392) );
  XOR U10441 ( .A(n4258), .B(n9389), .Z(n9390) );
  XOR U10442 ( .A(n9393), .B(n9394), .Z(n9389) );
  ANDN U10443 ( .B(n9395), .A(n4269), .Z(n9393) );
  XNOR U10444 ( .A(n9396), .B(n9397), .Z(n4269) );
  IV U10445 ( .A(n9394), .Z(n9397) );
  XOR U10446 ( .A(n4268), .B(n9394), .Z(n9395) );
  XOR U10447 ( .A(n9398), .B(n9399), .Z(n9394) );
  ANDN U10448 ( .B(n9400), .A(n4274), .Z(n9398) );
  XNOR U10449 ( .A(n9401), .B(n9402), .Z(n4274) );
  IV U10450 ( .A(n9399), .Z(n9402) );
  XOR U10451 ( .A(n4273), .B(n9399), .Z(n9400) );
  XOR U10452 ( .A(n9403), .B(n9404), .Z(n9399) );
  ANDN U10453 ( .B(n9405), .A(n4279), .Z(n9403) );
  XNOR U10454 ( .A(n9406), .B(n9407), .Z(n4279) );
  IV U10455 ( .A(n9404), .Z(n9407) );
  XOR U10456 ( .A(n4278), .B(n9404), .Z(n9405) );
  XOR U10457 ( .A(n9408), .B(n9409), .Z(n9404) );
  ANDN U10458 ( .B(n9410), .A(n4284), .Z(n9408) );
  XNOR U10459 ( .A(n9411), .B(n9412), .Z(n4284) );
  IV U10460 ( .A(n9409), .Z(n9412) );
  XOR U10461 ( .A(n4283), .B(n9409), .Z(n9410) );
  XOR U10462 ( .A(n9413), .B(n9414), .Z(n9409) );
  ANDN U10463 ( .B(n9415), .A(n4289), .Z(n9413) );
  XNOR U10464 ( .A(n9416), .B(n9417), .Z(n4289) );
  IV U10465 ( .A(n9414), .Z(n9417) );
  XOR U10466 ( .A(n4288), .B(n9414), .Z(n9415) );
  XOR U10467 ( .A(n9418), .B(n9419), .Z(n9414) );
  ANDN U10468 ( .B(n9420), .A(n4294), .Z(n9418) );
  XNOR U10469 ( .A(n9421), .B(n9422), .Z(n4294) );
  IV U10470 ( .A(n9419), .Z(n9422) );
  XOR U10471 ( .A(n4293), .B(n9419), .Z(n9420) );
  XOR U10472 ( .A(n9423), .B(n9424), .Z(n9419) );
  ANDN U10473 ( .B(n9425), .A(n4299), .Z(n9423) );
  XNOR U10474 ( .A(n9426), .B(n9427), .Z(n4299) );
  IV U10475 ( .A(n9424), .Z(n9427) );
  XOR U10476 ( .A(n4298), .B(n9424), .Z(n9425) );
  XOR U10477 ( .A(n9428), .B(n9429), .Z(n9424) );
  ANDN U10478 ( .B(n9430), .A(n4304), .Z(n9428) );
  XNOR U10479 ( .A(n9431), .B(n9432), .Z(n4304) );
  IV U10480 ( .A(n9429), .Z(n9432) );
  XOR U10481 ( .A(n4303), .B(n9429), .Z(n9430) );
  XOR U10482 ( .A(n9433), .B(n9434), .Z(n9429) );
  ANDN U10483 ( .B(n9435), .A(n4309), .Z(n9433) );
  XNOR U10484 ( .A(n9436), .B(n9437), .Z(n4309) );
  IV U10485 ( .A(n9434), .Z(n9437) );
  XOR U10486 ( .A(n4308), .B(n9434), .Z(n9435) );
  XOR U10487 ( .A(n9438), .B(n9439), .Z(n9434) );
  ANDN U10488 ( .B(n9440), .A(n4314), .Z(n9438) );
  XNOR U10489 ( .A(n9441), .B(n9442), .Z(n4314) );
  IV U10490 ( .A(n9439), .Z(n9442) );
  XOR U10491 ( .A(n4313), .B(n9439), .Z(n9440) );
  XOR U10492 ( .A(n9443), .B(n9444), .Z(n9439) );
  ANDN U10493 ( .B(n9445), .A(n4324), .Z(n9443) );
  XNOR U10494 ( .A(n9446), .B(n9447), .Z(n4324) );
  IV U10495 ( .A(n9444), .Z(n9447) );
  XOR U10496 ( .A(n4323), .B(n9444), .Z(n9445) );
  XOR U10497 ( .A(n9448), .B(n9449), .Z(n9444) );
  ANDN U10498 ( .B(n9450), .A(n4329), .Z(n9448) );
  XNOR U10499 ( .A(n9451), .B(n9452), .Z(n4329) );
  IV U10500 ( .A(n9449), .Z(n9452) );
  XOR U10501 ( .A(n4328), .B(n9449), .Z(n9450) );
  XOR U10502 ( .A(n9453), .B(n9454), .Z(n9449) );
  ANDN U10503 ( .B(n9455), .A(n4334), .Z(n9453) );
  XNOR U10504 ( .A(n9456), .B(n9457), .Z(n4334) );
  IV U10505 ( .A(n9454), .Z(n9457) );
  XOR U10506 ( .A(n4333), .B(n9454), .Z(n9455) );
  XOR U10507 ( .A(n9458), .B(n9459), .Z(n9454) );
  ANDN U10508 ( .B(n9460), .A(n4339), .Z(n9458) );
  XNOR U10509 ( .A(n9461), .B(n9462), .Z(n4339) );
  IV U10510 ( .A(n9459), .Z(n9462) );
  XOR U10511 ( .A(n4338), .B(n9459), .Z(n9460) );
  XOR U10512 ( .A(n9463), .B(n9464), .Z(n9459) );
  ANDN U10513 ( .B(n9465), .A(n4344), .Z(n9463) );
  XNOR U10514 ( .A(n9466), .B(n9467), .Z(n4344) );
  IV U10515 ( .A(n9464), .Z(n9467) );
  XOR U10516 ( .A(n4343), .B(n9464), .Z(n9465) );
  XOR U10517 ( .A(n9468), .B(n9469), .Z(n9464) );
  ANDN U10518 ( .B(n9470), .A(n4349), .Z(n9468) );
  XNOR U10519 ( .A(n9471), .B(n9472), .Z(n4349) );
  IV U10520 ( .A(n9469), .Z(n9472) );
  XOR U10521 ( .A(n4348), .B(n9469), .Z(n9470) );
  XOR U10522 ( .A(n9473), .B(n9474), .Z(n9469) );
  ANDN U10523 ( .B(n9475), .A(n4354), .Z(n9473) );
  XNOR U10524 ( .A(n9476), .B(n9477), .Z(n4354) );
  IV U10525 ( .A(n9474), .Z(n9477) );
  XOR U10526 ( .A(n4353), .B(n9474), .Z(n9475) );
  XOR U10527 ( .A(n9478), .B(n9479), .Z(n9474) );
  ANDN U10528 ( .B(n9480), .A(n4359), .Z(n9478) );
  XNOR U10529 ( .A(n9481), .B(n9482), .Z(n4359) );
  IV U10530 ( .A(n9479), .Z(n9482) );
  XOR U10531 ( .A(n4358), .B(n9479), .Z(n9480) );
  XOR U10532 ( .A(n9483), .B(n9484), .Z(n9479) );
  ANDN U10533 ( .B(n9485), .A(n4364), .Z(n9483) );
  XNOR U10534 ( .A(n9486), .B(n9487), .Z(n4364) );
  IV U10535 ( .A(n9484), .Z(n9487) );
  XOR U10536 ( .A(n4363), .B(n9484), .Z(n9485) );
  XOR U10537 ( .A(n9488), .B(n9489), .Z(n9484) );
  ANDN U10538 ( .B(n9490), .A(n4369), .Z(n9488) );
  XNOR U10539 ( .A(n9491), .B(n9492), .Z(n4369) );
  IV U10540 ( .A(n9489), .Z(n9492) );
  XOR U10541 ( .A(n4368), .B(n9489), .Z(n9490) );
  XOR U10542 ( .A(n9493), .B(n9494), .Z(n9489) );
  ANDN U10543 ( .B(n9495), .A(n4379), .Z(n9493) );
  XNOR U10544 ( .A(n9496), .B(n9497), .Z(n4379) );
  IV U10545 ( .A(n9494), .Z(n9497) );
  XOR U10546 ( .A(n4378), .B(n9494), .Z(n9495) );
  XOR U10547 ( .A(n9498), .B(n9499), .Z(n9494) );
  ANDN U10548 ( .B(n9500), .A(n4384), .Z(n9498) );
  XNOR U10549 ( .A(n9501), .B(n9502), .Z(n4384) );
  IV U10550 ( .A(n9499), .Z(n9502) );
  XOR U10551 ( .A(n4383), .B(n9499), .Z(n9500) );
  XOR U10552 ( .A(n9503), .B(n9504), .Z(n9499) );
  ANDN U10553 ( .B(n9505), .A(n4389), .Z(n9503) );
  XNOR U10554 ( .A(n9506), .B(n9507), .Z(n4389) );
  IV U10555 ( .A(n9504), .Z(n9507) );
  XOR U10556 ( .A(n4388), .B(n9504), .Z(n9505) );
  XOR U10557 ( .A(n9508), .B(n9509), .Z(n9504) );
  ANDN U10558 ( .B(n9510), .A(n4394), .Z(n9508) );
  XNOR U10559 ( .A(n9511), .B(n9512), .Z(n4394) );
  IV U10560 ( .A(n9509), .Z(n9512) );
  XOR U10561 ( .A(n4393), .B(n9509), .Z(n9510) );
  XOR U10562 ( .A(n9513), .B(n9514), .Z(n9509) );
  ANDN U10563 ( .B(n9515), .A(n4399), .Z(n9513) );
  XNOR U10564 ( .A(n9516), .B(n9517), .Z(n4399) );
  IV U10565 ( .A(n9514), .Z(n9517) );
  XOR U10566 ( .A(n4398), .B(n9514), .Z(n9515) );
  XOR U10567 ( .A(n9518), .B(n9519), .Z(n9514) );
  ANDN U10568 ( .B(n9520), .A(n4404), .Z(n9518) );
  XNOR U10569 ( .A(n9521), .B(n9522), .Z(n4404) );
  IV U10570 ( .A(n9519), .Z(n9522) );
  XOR U10571 ( .A(n4403), .B(n9519), .Z(n9520) );
  XOR U10572 ( .A(n9523), .B(n9524), .Z(n9519) );
  ANDN U10573 ( .B(n9525), .A(n4409), .Z(n9523) );
  XNOR U10574 ( .A(n9526), .B(n9527), .Z(n4409) );
  IV U10575 ( .A(n9524), .Z(n9527) );
  XOR U10576 ( .A(n4408), .B(n9524), .Z(n9525) );
  XOR U10577 ( .A(n9528), .B(n9529), .Z(n9524) );
  ANDN U10578 ( .B(n9530), .A(n4414), .Z(n9528) );
  XNOR U10579 ( .A(n9531), .B(n9532), .Z(n4414) );
  IV U10580 ( .A(n9529), .Z(n9532) );
  XOR U10581 ( .A(n4413), .B(n9529), .Z(n9530) );
  XOR U10582 ( .A(n9533), .B(n9534), .Z(n9529) );
  ANDN U10583 ( .B(n9535), .A(n4419), .Z(n9533) );
  XNOR U10584 ( .A(n9536), .B(n9537), .Z(n4419) );
  IV U10585 ( .A(n9534), .Z(n9537) );
  XOR U10586 ( .A(n4418), .B(n9534), .Z(n9535) );
  XOR U10587 ( .A(n9538), .B(n9539), .Z(n9534) );
  ANDN U10588 ( .B(n9540), .A(n4424), .Z(n9538) );
  XNOR U10589 ( .A(n9541), .B(n9542), .Z(n4424) );
  IV U10590 ( .A(n9539), .Z(n9542) );
  XOR U10591 ( .A(n4423), .B(n9539), .Z(n9540) );
  XOR U10592 ( .A(n9543), .B(n9544), .Z(n9539) );
  ANDN U10593 ( .B(n9545), .A(n4434), .Z(n9543) );
  XNOR U10594 ( .A(n9546), .B(n9547), .Z(n4434) );
  IV U10595 ( .A(n9544), .Z(n9547) );
  XOR U10596 ( .A(n4433), .B(n9544), .Z(n9545) );
  XOR U10597 ( .A(n9548), .B(n9549), .Z(n9544) );
  ANDN U10598 ( .B(n9550), .A(n4439), .Z(n9548) );
  XNOR U10599 ( .A(n9551), .B(n9552), .Z(n4439) );
  IV U10600 ( .A(n9549), .Z(n9552) );
  XOR U10601 ( .A(n4438), .B(n9549), .Z(n9550) );
  XOR U10602 ( .A(n9553), .B(n9554), .Z(n9549) );
  ANDN U10603 ( .B(n9555), .A(n4444), .Z(n9553) );
  XNOR U10604 ( .A(n9556), .B(n9557), .Z(n4444) );
  IV U10605 ( .A(n9554), .Z(n9557) );
  XOR U10606 ( .A(n4443), .B(n9554), .Z(n9555) );
  XOR U10607 ( .A(n9558), .B(n9559), .Z(n9554) );
  ANDN U10608 ( .B(n9560), .A(n4449), .Z(n9558) );
  XNOR U10609 ( .A(n9561), .B(n9562), .Z(n4449) );
  IV U10610 ( .A(n9559), .Z(n9562) );
  XOR U10611 ( .A(n4448), .B(n9559), .Z(n9560) );
  XOR U10612 ( .A(n9563), .B(n9564), .Z(n9559) );
  ANDN U10613 ( .B(n9565), .A(n4454), .Z(n9563) );
  XNOR U10614 ( .A(n9566), .B(n9567), .Z(n4454) );
  IV U10615 ( .A(n9564), .Z(n9567) );
  XOR U10616 ( .A(n4453), .B(n9564), .Z(n9565) );
  XOR U10617 ( .A(n9568), .B(n9569), .Z(n9564) );
  ANDN U10618 ( .B(n9570), .A(n4459), .Z(n9568) );
  XNOR U10619 ( .A(n9571), .B(n9572), .Z(n4459) );
  IV U10620 ( .A(n9569), .Z(n9572) );
  XOR U10621 ( .A(n4458), .B(n9569), .Z(n9570) );
  XOR U10622 ( .A(n9573), .B(n9574), .Z(n9569) );
  ANDN U10623 ( .B(n9575), .A(n4464), .Z(n9573) );
  XNOR U10624 ( .A(n9576), .B(n9577), .Z(n4464) );
  IV U10625 ( .A(n9574), .Z(n9577) );
  XOR U10626 ( .A(n4463), .B(n9574), .Z(n9575) );
  XOR U10627 ( .A(n9578), .B(n9579), .Z(n9574) );
  ANDN U10628 ( .B(n9580), .A(n4469), .Z(n9578) );
  XNOR U10629 ( .A(n9581), .B(n9582), .Z(n4469) );
  IV U10630 ( .A(n9579), .Z(n9582) );
  XOR U10631 ( .A(n4468), .B(n9579), .Z(n9580) );
  XOR U10632 ( .A(n9583), .B(n9584), .Z(n9579) );
  ANDN U10633 ( .B(n9585), .A(n4474), .Z(n9583) );
  XNOR U10634 ( .A(n9586), .B(n9587), .Z(n4474) );
  IV U10635 ( .A(n9584), .Z(n9587) );
  XOR U10636 ( .A(n4473), .B(n9584), .Z(n9585) );
  XOR U10637 ( .A(n9588), .B(n9589), .Z(n9584) );
  ANDN U10638 ( .B(n9590), .A(n4479), .Z(n9588) );
  XNOR U10639 ( .A(n9591), .B(n9592), .Z(n4479) );
  IV U10640 ( .A(n9589), .Z(n9592) );
  XOR U10641 ( .A(n4478), .B(n9589), .Z(n9590) );
  XOR U10642 ( .A(n9593), .B(n9594), .Z(n9589) );
  ANDN U10643 ( .B(n9595), .A(n4489), .Z(n9593) );
  XNOR U10644 ( .A(n9596), .B(n9597), .Z(n4489) );
  IV U10645 ( .A(n9594), .Z(n9597) );
  XOR U10646 ( .A(n4488), .B(n9594), .Z(n9595) );
  XOR U10647 ( .A(n9598), .B(n9599), .Z(n9594) );
  ANDN U10648 ( .B(n9600), .A(n4494), .Z(n9598) );
  XNOR U10649 ( .A(n9601), .B(n9602), .Z(n4494) );
  IV U10650 ( .A(n9599), .Z(n9602) );
  XOR U10651 ( .A(n4493), .B(n9599), .Z(n9600) );
  XOR U10652 ( .A(n9603), .B(n9604), .Z(n9599) );
  ANDN U10653 ( .B(n9605), .A(n4499), .Z(n9603) );
  XNOR U10654 ( .A(n9606), .B(n9607), .Z(n4499) );
  IV U10655 ( .A(n9604), .Z(n9607) );
  XOR U10656 ( .A(n4498), .B(n9604), .Z(n9605) );
  XOR U10657 ( .A(n9608), .B(n9609), .Z(n9604) );
  ANDN U10658 ( .B(n9610), .A(n4504), .Z(n9608) );
  XNOR U10659 ( .A(n9611), .B(n9612), .Z(n4504) );
  IV U10660 ( .A(n9609), .Z(n9612) );
  XOR U10661 ( .A(n4503), .B(n9609), .Z(n9610) );
  XOR U10662 ( .A(n9613), .B(n9614), .Z(n9609) );
  ANDN U10663 ( .B(n9615), .A(n4509), .Z(n9613) );
  XNOR U10664 ( .A(n9616), .B(n9617), .Z(n4509) );
  IV U10665 ( .A(n9614), .Z(n9617) );
  XOR U10666 ( .A(n4508), .B(n9614), .Z(n9615) );
  XOR U10667 ( .A(n9618), .B(n9619), .Z(n9614) );
  ANDN U10668 ( .B(n9620), .A(n4514), .Z(n9618) );
  XNOR U10669 ( .A(n9621), .B(n9622), .Z(n4514) );
  IV U10670 ( .A(n9619), .Z(n9622) );
  XOR U10671 ( .A(n4513), .B(n9619), .Z(n9620) );
  XOR U10672 ( .A(n9623), .B(n9624), .Z(n9619) );
  ANDN U10673 ( .B(n9625), .A(n4519), .Z(n9623) );
  XNOR U10674 ( .A(n9626), .B(n9627), .Z(n4519) );
  IV U10675 ( .A(n9624), .Z(n9627) );
  XOR U10676 ( .A(n4518), .B(n9624), .Z(n9625) );
  XOR U10677 ( .A(n9628), .B(n9629), .Z(n9624) );
  ANDN U10678 ( .B(n9630), .A(n4524), .Z(n9628) );
  XNOR U10679 ( .A(n9631), .B(n9632), .Z(n4524) );
  IV U10680 ( .A(n9629), .Z(n9632) );
  XOR U10681 ( .A(n4523), .B(n9629), .Z(n9630) );
  XOR U10682 ( .A(n9633), .B(n9634), .Z(n9629) );
  ANDN U10683 ( .B(n9635), .A(n4529), .Z(n9633) );
  XNOR U10684 ( .A(n9636), .B(n9637), .Z(n4529) );
  IV U10685 ( .A(n9634), .Z(n9637) );
  XOR U10686 ( .A(n4528), .B(n9634), .Z(n9635) );
  XOR U10687 ( .A(n9638), .B(n9639), .Z(n9634) );
  ANDN U10688 ( .B(n9640), .A(n4534), .Z(n9638) );
  XNOR U10689 ( .A(n9641), .B(n9642), .Z(n4534) );
  IV U10690 ( .A(n9639), .Z(n9642) );
  XOR U10691 ( .A(n4533), .B(n9639), .Z(n9640) );
  XOR U10692 ( .A(n9643), .B(n9644), .Z(n9639) );
  ANDN U10693 ( .B(n9645), .A(n4544), .Z(n9643) );
  XNOR U10694 ( .A(n9646), .B(n9647), .Z(n4544) );
  IV U10695 ( .A(n9644), .Z(n9647) );
  XOR U10696 ( .A(n4543), .B(n9644), .Z(n9645) );
  XOR U10697 ( .A(n9648), .B(n9649), .Z(n9644) );
  ANDN U10698 ( .B(n9650), .A(n4549), .Z(n9648) );
  XNOR U10699 ( .A(n9651), .B(n9652), .Z(n4549) );
  IV U10700 ( .A(n9649), .Z(n9652) );
  XOR U10701 ( .A(n4548), .B(n9649), .Z(n9650) );
  XOR U10702 ( .A(n9653), .B(n9654), .Z(n9649) );
  ANDN U10703 ( .B(n9655), .A(n4554), .Z(n9653) );
  XNOR U10704 ( .A(n9656), .B(n9657), .Z(n4554) );
  IV U10705 ( .A(n9654), .Z(n9657) );
  XOR U10706 ( .A(n4553), .B(n9654), .Z(n9655) );
  XOR U10707 ( .A(n9658), .B(n9659), .Z(n9654) );
  ANDN U10708 ( .B(n9660), .A(n4559), .Z(n9658) );
  XNOR U10709 ( .A(n9661), .B(n9662), .Z(n4559) );
  IV U10710 ( .A(n9659), .Z(n9662) );
  XOR U10711 ( .A(n4558), .B(n9659), .Z(n9660) );
  XOR U10712 ( .A(n9663), .B(n9664), .Z(n9659) );
  ANDN U10713 ( .B(n9665), .A(n4564), .Z(n9663) );
  XNOR U10714 ( .A(n9666), .B(n9667), .Z(n4564) );
  IV U10715 ( .A(n9664), .Z(n9667) );
  XOR U10716 ( .A(n4563), .B(n9664), .Z(n9665) );
  XOR U10717 ( .A(n9668), .B(n9669), .Z(n9664) );
  ANDN U10718 ( .B(n9670), .A(n4569), .Z(n9668) );
  XNOR U10719 ( .A(n9671), .B(n9672), .Z(n4569) );
  IV U10720 ( .A(n9669), .Z(n9672) );
  XOR U10721 ( .A(n4568), .B(n9669), .Z(n9670) );
  XOR U10722 ( .A(n9673), .B(n9674), .Z(n9669) );
  ANDN U10723 ( .B(n9675), .A(n4574), .Z(n9673) );
  XNOR U10724 ( .A(n9676), .B(n9677), .Z(n4574) );
  IV U10725 ( .A(n9674), .Z(n9677) );
  XOR U10726 ( .A(n4573), .B(n9674), .Z(n9675) );
  XOR U10727 ( .A(n9678), .B(n9679), .Z(n9674) );
  ANDN U10728 ( .B(n9680), .A(n4579), .Z(n9678) );
  XNOR U10729 ( .A(n9681), .B(n9682), .Z(n4579) );
  IV U10730 ( .A(n9679), .Z(n9682) );
  XOR U10731 ( .A(n4578), .B(n9679), .Z(n9680) );
  XOR U10732 ( .A(n9683), .B(n9684), .Z(n9679) );
  ANDN U10733 ( .B(n9685), .A(n4584), .Z(n9683) );
  XNOR U10734 ( .A(n9686), .B(n9687), .Z(n4584) );
  IV U10735 ( .A(n9684), .Z(n9687) );
  XOR U10736 ( .A(n4583), .B(n9684), .Z(n9685) );
  XOR U10737 ( .A(n9688), .B(n9689), .Z(n9684) );
  ANDN U10738 ( .B(n9690), .A(n4589), .Z(n9688) );
  XNOR U10739 ( .A(n9691), .B(n9692), .Z(n4589) );
  IV U10740 ( .A(n9689), .Z(n9692) );
  XOR U10741 ( .A(n4588), .B(n9689), .Z(n9690) );
  XOR U10742 ( .A(n9693), .B(n9694), .Z(n9689) );
  ANDN U10743 ( .B(n9695), .A(n4599), .Z(n9693) );
  XNOR U10744 ( .A(n9696), .B(n9697), .Z(n4599) );
  IV U10745 ( .A(n9694), .Z(n9697) );
  XOR U10746 ( .A(n4598), .B(n9694), .Z(n9695) );
  XOR U10747 ( .A(n9698), .B(n9699), .Z(n9694) );
  ANDN U10748 ( .B(n9700), .A(n4604), .Z(n9698) );
  XNOR U10749 ( .A(n9701), .B(n9702), .Z(n4604) );
  IV U10750 ( .A(n9699), .Z(n9702) );
  XOR U10751 ( .A(n4603), .B(n9699), .Z(n9700) );
  XOR U10752 ( .A(n9703), .B(n9704), .Z(n9699) );
  ANDN U10753 ( .B(n9705), .A(n4609), .Z(n9703) );
  XNOR U10754 ( .A(n9706), .B(n9707), .Z(n4609) );
  IV U10755 ( .A(n9704), .Z(n9707) );
  XOR U10756 ( .A(n4608), .B(n9704), .Z(n9705) );
  XOR U10757 ( .A(n9708), .B(n9709), .Z(n9704) );
  ANDN U10758 ( .B(n9710), .A(n4614), .Z(n9708) );
  XNOR U10759 ( .A(n9711), .B(n9712), .Z(n4614) );
  IV U10760 ( .A(n9709), .Z(n9712) );
  XOR U10761 ( .A(n4613), .B(n9709), .Z(n9710) );
  XOR U10762 ( .A(n9713), .B(n9714), .Z(n9709) );
  ANDN U10763 ( .B(n9715), .A(n4619), .Z(n9713) );
  XNOR U10764 ( .A(n9716), .B(n9717), .Z(n4619) );
  IV U10765 ( .A(n9714), .Z(n9717) );
  XOR U10766 ( .A(n4618), .B(n9714), .Z(n9715) );
  XOR U10767 ( .A(n9718), .B(n9719), .Z(n9714) );
  ANDN U10768 ( .B(n9720), .A(n4624), .Z(n9718) );
  XNOR U10769 ( .A(n9721), .B(n9722), .Z(n4624) );
  IV U10770 ( .A(n9719), .Z(n9722) );
  XOR U10771 ( .A(n4623), .B(n9719), .Z(n9720) );
  XOR U10772 ( .A(n9723), .B(n9724), .Z(n9719) );
  ANDN U10773 ( .B(n9725), .A(n4629), .Z(n9723) );
  XNOR U10774 ( .A(n9726), .B(n9727), .Z(n4629) );
  IV U10775 ( .A(n9724), .Z(n9727) );
  XOR U10776 ( .A(n4628), .B(n9724), .Z(n9725) );
  XOR U10777 ( .A(n9728), .B(n9729), .Z(n9724) );
  ANDN U10778 ( .B(n9730), .A(n4634), .Z(n9728) );
  XNOR U10779 ( .A(n9731), .B(n9732), .Z(n4634) );
  IV U10780 ( .A(n9729), .Z(n9732) );
  XOR U10781 ( .A(n4633), .B(n9729), .Z(n9730) );
  XOR U10782 ( .A(n9733), .B(n9734), .Z(n9729) );
  ANDN U10783 ( .B(n9735), .A(n4639), .Z(n9733) );
  XNOR U10784 ( .A(n9736), .B(n9737), .Z(n4639) );
  IV U10785 ( .A(n9734), .Z(n9737) );
  XOR U10786 ( .A(n4638), .B(n9734), .Z(n9735) );
  XOR U10787 ( .A(n9738), .B(n9739), .Z(n9734) );
  ANDN U10788 ( .B(n9740), .A(n4644), .Z(n9738) );
  XNOR U10789 ( .A(n9741), .B(n9742), .Z(n4644) );
  IV U10790 ( .A(n9739), .Z(n9742) );
  XOR U10791 ( .A(n4643), .B(n9739), .Z(n9740) );
  XOR U10792 ( .A(n9743), .B(n9744), .Z(n9739) );
  ANDN U10793 ( .B(n9745), .A(n4654), .Z(n9743) );
  XNOR U10794 ( .A(n9746), .B(n9747), .Z(n4654) );
  IV U10795 ( .A(n9744), .Z(n9747) );
  XOR U10796 ( .A(n4653), .B(n9744), .Z(n9745) );
  XOR U10797 ( .A(n9748), .B(n9749), .Z(n9744) );
  ANDN U10798 ( .B(n9750), .A(n4659), .Z(n9748) );
  XNOR U10799 ( .A(n9751), .B(n9752), .Z(n4659) );
  IV U10800 ( .A(n9749), .Z(n9752) );
  XOR U10801 ( .A(n4658), .B(n9749), .Z(n9750) );
  XOR U10802 ( .A(n9753), .B(n9754), .Z(n9749) );
  ANDN U10803 ( .B(n9755), .A(n4664), .Z(n9753) );
  XNOR U10804 ( .A(n9756), .B(n9757), .Z(n4664) );
  IV U10805 ( .A(n9754), .Z(n9757) );
  XOR U10806 ( .A(n4663), .B(n9754), .Z(n9755) );
  XOR U10807 ( .A(n9758), .B(n9759), .Z(n9754) );
  ANDN U10808 ( .B(n9760), .A(n4669), .Z(n9758) );
  XNOR U10809 ( .A(n9761), .B(n9762), .Z(n4669) );
  IV U10810 ( .A(n9759), .Z(n9762) );
  XOR U10811 ( .A(n4668), .B(n9759), .Z(n9760) );
  XOR U10812 ( .A(n9763), .B(n9764), .Z(n9759) );
  ANDN U10813 ( .B(n9765), .A(n4674), .Z(n9763) );
  XNOR U10814 ( .A(n9766), .B(n9767), .Z(n4674) );
  IV U10815 ( .A(n9764), .Z(n9767) );
  XOR U10816 ( .A(n4673), .B(n9764), .Z(n9765) );
  XOR U10817 ( .A(n9768), .B(n9769), .Z(n9764) );
  ANDN U10818 ( .B(n9770), .A(n4679), .Z(n9768) );
  XNOR U10819 ( .A(n9771), .B(n9772), .Z(n4679) );
  IV U10820 ( .A(n9769), .Z(n9772) );
  XOR U10821 ( .A(n4678), .B(n9769), .Z(n9770) );
  XOR U10822 ( .A(n9773), .B(n9774), .Z(n9769) );
  ANDN U10823 ( .B(n9775), .A(n4684), .Z(n9773) );
  XNOR U10824 ( .A(n9776), .B(n9777), .Z(n4684) );
  IV U10825 ( .A(n9774), .Z(n9777) );
  XOR U10826 ( .A(n4683), .B(n9774), .Z(n9775) );
  XOR U10827 ( .A(n9778), .B(n9779), .Z(n9774) );
  ANDN U10828 ( .B(n9780), .A(n4689), .Z(n9778) );
  XNOR U10829 ( .A(n9781), .B(n9782), .Z(n4689) );
  IV U10830 ( .A(n9779), .Z(n9782) );
  XOR U10831 ( .A(n4688), .B(n9779), .Z(n9780) );
  XOR U10832 ( .A(n9783), .B(n9784), .Z(n9779) );
  ANDN U10833 ( .B(n9785), .A(n4694), .Z(n9783) );
  XNOR U10834 ( .A(n9786), .B(n9787), .Z(n4694) );
  IV U10835 ( .A(n9784), .Z(n9787) );
  XOR U10836 ( .A(n4693), .B(n9784), .Z(n9785) );
  XOR U10837 ( .A(n9788), .B(n9789), .Z(n9784) );
  ANDN U10838 ( .B(n9790), .A(n4699), .Z(n9788) );
  XNOR U10839 ( .A(n9791), .B(n9792), .Z(n4699) );
  IV U10840 ( .A(n9789), .Z(n9792) );
  XOR U10841 ( .A(n4698), .B(n9789), .Z(n9790) );
  XOR U10842 ( .A(n9793), .B(n9794), .Z(n9789) );
  ANDN U10843 ( .B(n9795), .A(n4709), .Z(n9793) );
  XNOR U10844 ( .A(n9796), .B(n9797), .Z(n4709) );
  IV U10845 ( .A(n9794), .Z(n9797) );
  XOR U10846 ( .A(n4708), .B(n9794), .Z(n9795) );
  XOR U10847 ( .A(n9798), .B(n9799), .Z(n9794) );
  ANDN U10848 ( .B(n9800), .A(n4714), .Z(n9798) );
  XNOR U10849 ( .A(n9801), .B(n9802), .Z(n4714) );
  IV U10850 ( .A(n9799), .Z(n9802) );
  XOR U10851 ( .A(n4713), .B(n9799), .Z(n9800) );
  XOR U10852 ( .A(n9803), .B(n9804), .Z(n9799) );
  ANDN U10853 ( .B(n9805), .A(n4719), .Z(n9803) );
  XNOR U10854 ( .A(n9806), .B(n9807), .Z(n4719) );
  IV U10855 ( .A(n9804), .Z(n9807) );
  XOR U10856 ( .A(n4718), .B(n9804), .Z(n9805) );
  XOR U10857 ( .A(n9808), .B(n9809), .Z(n9804) );
  ANDN U10858 ( .B(n9810), .A(n4724), .Z(n9808) );
  XNOR U10859 ( .A(n9811), .B(n9812), .Z(n4724) );
  IV U10860 ( .A(n9809), .Z(n9812) );
  XOR U10861 ( .A(n4723), .B(n9809), .Z(n9810) );
  XOR U10862 ( .A(n9813), .B(n9814), .Z(n9809) );
  ANDN U10863 ( .B(n9815), .A(n4729), .Z(n9813) );
  XNOR U10864 ( .A(n9816), .B(n9817), .Z(n4729) );
  IV U10865 ( .A(n9814), .Z(n9817) );
  XOR U10866 ( .A(n4728), .B(n9814), .Z(n9815) );
  XOR U10867 ( .A(n9818), .B(n9819), .Z(n9814) );
  ANDN U10868 ( .B(n9820), .A(n4734), .Z(n9818) );
  XNOR U10869 ( .A(n9821), .B(n9822), .Z(n4734) );
  IV U10870 ( .A(n9819), .Z(n9822) );
  XOR U10871 ( .A(n4733), .B(n9819), .Z(n9820) );
  XOR U10872 ( .A(n9823), .B(n9824), .Z(n9819) );
  ANDN U10873 ( .B(n9825), .A(n4739), .Z(n9823) );
  XNOR U10874 ( .A(n9826), .B(n9827), .Z(n4739) );
  IV U10875 ( .A(n9824), .Z(n9827) );
  XOR U10876 ( .A(n4738), .B(n9824), .Z(n9825) );
  XOR U10877 ( .A(n9828), .B(n9829), .Z(n9824) );
  ANDN U10878 ( .B(n9830), .A(n4744), .Z(n9828) );
  XNOR U10879 ( .A(n9831), .B(n9832), .Z(n4744) );
  IV U10880 ( .A(n9829), .Z(n9832) );
  XOR U10881 ( .A(n4743), .B(n9829), .Z(n9830) );
  XOR U10882 ( .A(n9833), .B(n9834), .Z(n9829) );
  ANDN U10883 ( .B(n9835), .A(n4749), .Z(n9833) );
  XNOR U10884 ( .A(n9836), .B(n9837), .Z(n4749) );
  IV U10885 ( .A(n9834), .Z(n9837) );
  XOR U10886 ( .A(n4748), .B(n9834), .Z(n9835) );
  XOR U10887 ( .A(n9838), .B(n9839), .Z(n9834) );
  ANDN U10888 ( .B(n9840), .A(n4754), .Z(n9838) );
  XNOR U10889 ( .A(n9841), .B(n9842), .Z(n4754) );
  IV U10890 ( .A(n9839), .Z(n9842) );
  XOR U10891 ( .A(n4753), .B(n9839), .Z(n9840) );
  XOR U10892 ( .A(n9843), .B(n9844), .Z(n9839) );
  ANDN U10893 ( .B(n9845), .A(n4769), .Z(n9843) );
  XNOR U10894 ( .A(n9846), .B(n9847), .Z(n4769) );
  IV U10895 ( .A(n9844), .Z(n9847) );
  XOR U10896 ( .A(n4768), .B(n9844), .Z(n9845) );
  XOR U10897 ( .A(n9848), .B(n9849), .Z(n9844) );
  ANDN U10898 ( .B(n9850), .A(n4774), .Z(n9848) );
  XNOR U10899 ( .A(n9851), .B(n9852), .Z(n4774) );
  IV U10900 ( .A(n9849), .Z(n9852) );
  XOR U10901 ( .A(n4773), .B(n9849), .Z(n9850) );
  XOR U10902 ( .A(n9853), .B(n9854), .Z(n9849) );
  ANDN U10903 ( .B(n9855), .A(n4779), .Z(n9853) );
  XNOR U10904 ( .A(n9856), .B(n9857), .Z(n4779) );
  IV U10905 ( .A(n9854), .Z(n9857) );
  XOR U10906 ( .A(n4778), .B(n9854), .Z(n9855) );
  XOR U10907 ( .A(n9858), .B(n9859), .Z(n9854) );
  ANDN U10908 ( .B(n9860), .A(n4784), .Z(n9858) );
  XNOR U10909 ( .A(n9861), .B(n9862), .Z(n4784) );
  IV U10910 ( .A(n9859), .Z(n9862) );
  XOR U10911 ( .A(n4783), .B(n9859), .Z(n9860) );
  XOR U10912 ( .A(n9863), .B(n9864), .Z(n9859) );
  ANDN U10913 ( .B(n9865), .A(n4789), .Z(n9863) );
  XNOR U10914 ( .A(n9866), .B(n9867), .Z(n4789) );
  IV U10915 ( .A(n9864), .Z(n9867) );
  XOR U10916 ( .A(n4788), .B(n9864), .Z(n9865) );
  XOR U10917 ( .A(n9868), .B(n9869), .Z(n9864) );
  ANDN U10918 ( .B(n9870), .A(n4794), .Z(n9868) );
  XNOR U10919 ( .A(n9871), .B(n9872), .Z(n4794) );
  IV U10920 ( .A(n9869), .Z(n9872) );
  XOR U10921 ( .A(n4793), .B(n9869), .Z(n9870) );
  XOR U10922 ( .A(n9873), .B(n9874), .Z(n9869) );
  ANDN U10923 ( .B(n9875), .A(n4799), .Z(n9873) );
  XNOR U10924 ( .A(n9876), .B(n9877), .Z(n4799) );
  IV U10925 ( .A(n9874), .Z(n9877) );
  XOR U10926 ( .A(n4798), .B(n9874), .Z(n9875) );
  XOR U10927 ( .A(n9878), .B(n9879), .Z(n9874) );
  ANDN U10928 ( .B(n9880), .A(n4804), .Z(n9878) );
  XNOR U10929 ( .A(n9881), .B(n9882), .Z(n4804) );
  IV U10930 ( .A(n9879), .Z(n9882) );
  XOR U10931 ( .A(n4803), .B(n9879), .Z(n9880) );
  XOR U10932 ( .A(n9883), .B(n9884), .Z(n9879) );
  ANDN U10933 ( .B(n9885), .A(n4809), .Z(n9883) );
  XNOR U10934 ( .A(n9886), .B(n9887), .Z(n4809) );
  IV U10935 ( .A(n9884), .Z(n9887) );
  XOR U10936 ( .A(n4808), .B(n9884), .Z(n9885) );
  XOR U10937 ( .A(n9888), .B(n9889), .Z(n9884) );
  ANDN U10938 ( .B(n9890), .A(n4814), .Z(n9888) );
  XNOR U10939 ( .A(n9891), .B(n9892), .Z(n4814) );
  IV U10940 ( .A(n9889), .Z(n9892) );
  XOR U10941 ( .A(n4813), .B(n9889), .Z(n9890) );
  XOR U10942 ( .A(n9893), .B(n9894), .Z(n9889) );
  ANDN U10943 ( .B(n9895), .A(n4824), .Z(n9893) );
  XNOR U10944 ( .A(n9896), .B(n9897), .Z(n4824) );
  IV U10945 ( .A(n9894), .Z(n9897) );
  XOR U10946 ( .A(n4823), .B(n9894), .Z(n9895) );
  XOR U10947 ( .A(n9898), .B(n9899), .Z(n9894) );
  ANDN U10948 ( .B(n9900), .A(n4829), .Z(n9898) );
  XNOR U10949 ( .A(n9901), .B(n9902), .Z(n4829) );
  IV U10950 ( .A(n9899), .Z(n9902) );
  XOR U10951 ( .A(n4828), .B(n9899), .Z(n9900) );
  XOR U10952 ( .A(n9903), .B(n9904), .Z(n9899) );
  ANDN U10953 ( .B(n9905), .A(n4834), .Z(n9903) );
  XNOR U10954 ( .A(n9906), .B(n9907), .Z(n4834) );
  IV U10955 ( .A(n9904), .Z(n9907) );
  XOR U10956 ( .A(n4833), .B(n9904), .Z(n9905) );
  XOR U10957 ( .A(n9908), .B(n9909), .Z(n9904) );
  ANDN U10958 ( .B(n9910), .A(n4839), .Z(n9908) );
  XNOR U10959 ( .A(n9911), .B(n9912), .Z(n4839) );
  IV U10960 ( .A(n9909), .Z(n9912) );
  XOR U10961 ( .A(n4838), .B(n9909), .Z(n9910) );
  XOR U10962 ( .A(n9913), .B(n9914), .Z(n9909) );
  ANDN U10963 ( .B(n9915), .A(n4844), .Z(n9913) );
  XNOR U10964 ( .A(n9916), .B(n9917), .Z(n4844) );
  IV U10965 ( .A(n9914), .Z(n9917) );
  XOR U10966 ( .A(n4843), .B(n9914), .Z(n9915) );
  XOR U10967 ( .A(n9918), .B(n9919), .Z(n9914) );
  ANDN U10968 ( .B(n9920), .A(n4849), .Z(n9918) );
  XNOR U10969 ( .A(n9921), .B(n9922), .Z(n4849) );
  IV U10970 ( .A(n9919), .Z(n9922) );
  XOR U10971 ( .A(n4848), .B(n9919), .Z(n9920) );
  XOR U10972 ( .A(n9923), .B(n9924), .Z(n9919) );
  ANDN U10973 ( .B(n9925), .A(n4854), .Z(n9923) );
  XNOR U10974 ( .A(n9926), .B(n9927), .Z(n4854) );
  IV U10975 ( .A(n9924), .Z(n9927) );
  XOR U10976 ( .A(n4853), .B(n9924), .Z(n9925) );
  XOR U10977 ( .A(n9928), .B(n9929), .Z(n9924) );
  ANDN U10978 ( .B(n9930), .A(n4859), .Z(n9928) );
  XNOR U10979 ( .A(n9931), .B(n9932), .Z(n4859) );
  IV U10980 ( .A(n9929), .Z(n9932) );
  XOR U10981 ( .A(n4858), .B(n9929), .Z(n9930) );
  XOR U10982 ( .A(n9933), .B(n9934), .Z(n9929) );
  ANDN U10983 ( .B(n9935), .A(n4864), .Z(n9933) );
  XNOR U10984 ( .A(n9936), .B(n9937), .Z(n4864) );
  IV U10985 ( .A(n9934), .Z(n9937) );
  XOR U10986 ( .A(n4863), .B(n9934), .Z(n9935) );
  XOR U10987 ( .A(n9938), .B(n9939), .Z(n9934) );
  ANDN U10988 ( .B(n9940), .A(n4869), .Z(n9938) );
  XNOR U10989 ( .A(n9941), .B(n9942), .Z(n4869) );
  IV U10990 ( .A(n9939), .Z(n9942) );
  XOR U10991 ( .A(n4868), .B(n9939), .Z(n9940) );
  XOR U10992 ( .A(n9943), .B(n9944), .Z(n9939) );
  ANDN U10993 ( .B(n9945), .A(n4879), .Z(n9943) );
  XNOR U10994 ( .A(n9946), .B(n9947), .Z(n4879) );
  IV U10995 ( .A(n9944), .Z(n9947) );
  XOR U10996 ( .A(n4878), .B(n9944), .Z(n9945) );
  XOR U10997 ( .A(n9948), .B(n9949), .Z(n9944) );
  ANDN U10998 ( .B(n9950), .A(n4884), .Z(n9948) );
  XNOR U10999 ( .A(n9951), .B(n9952), .Z(n4884) );
  IV U11000 ( .A(n9949), .Z(n9952) );
  XOR U11001 ( .A(n4883), .B(n9949), .Z(n9950) );
  XOR U11002 ( .A(n9953), .B(n9954), .Z(n9949) );
  ANDN U11003 ( .B(n9955), .A(n4889), .Z(n9953) );
  XNOR U11004 ( .A(n9956), .B(n9957), .Z(n4889) );
  IV U11005 ( .A(n9954), .Z(n9957) );
  XOR U11006 ( .A(n4888), .B(n9954), .Z(n9955) );
  XOR U11007 ( .A(n9958), .B(n9959), .Z(n9954) );
  ANDN U11008 ( .B(n9960), .A(n4894), .Z(n9958) );
  XNOR U11009 ( .A(n9961), .B(n9962), .Z(n4894) );
  IV U11010 ( .A(n9959), .Z(n9962) );
  XOR U11011 ( .A(n4893), .B(n9959), .Z(n9960) );
  XOR U11012 ( .A(n9963), .B(n9964), .Z(n9959) );
  ANDN U11013 ( .B(n9965), .A(n4899), .Z(n9963) );
  XNOR U11014 ( .A(n9966), .B(n9967), .Z(n4899) );
  IV U11015 ( .A(n9964), .Z(n9967) );
  XOR U11016 ( .A(n4898), .B(n9964), .Z(n9965) );
  XOR U11017 ( .A(n9968), .B(n9969), .Z(n9964) );
  ANDN U11018 ( .B(n9970), .A(n4904), .Z(n9968) );
  XNOR U11019 ( .A(n9971), .B(n9972), .Z(n4904) );
  IV U11020 ( .A(n9969), .Z(n9972) );
  XOR U11021 ( .A(n4903), .B(n9969), .Z(n9970) );
  XOR U11022 ( .A(n9973), .B(n9974), .Z(n9969) );
  ANDN U11023 ( .B(n9975), .A(n4909), .Z(n9973) );
  XNOR U11024 ( .A(n9976), .B(n9977), .Z(n4909) );
  IV U11025 ( .A(n9974), .Z(n9977) );
  XOR U11026 ( .A(n4908), .B(n9974), .Z(n9975) );
  XOR U11027 ( .A(n9978), .B(n9979), .Z(n9974) );
  ANDN U11028 ( .B(n9980), .A(n4914), .Z(n9978) );
  XNOR U11029 ( .A(n9981), .B(n9982), .Z(n4914) );
  IV U11030 ( .A(n9979), .Z(n9982) );
  XOR U11031 ( .A(n4913), .B(n9979), .Z(n9980) );
  XOR U11032 ( .A(n9983), .B(n9984), .Z(n9979) );
  ANDN U11033 ( .B(n9985), .A(n4919), .Z(n9983) );
  XNOR U11034 ( .A(n9986), .B(n9987), .Z(n4919) );
  IV U11035 ( .A(n9984), .Z(n9987) );
  XOR U11036 ( .A(n4918), .B(n9984), .Z(n9985) );
  XOR U11037 ( .A(n9988), .B(n9989), .Z(n9984) );
  ANDN U11038 ( .B(n9990), .A(n4924), .Z(n9988) );
  XNOR U11039 ( .A(n9991), .B(n9992), .Z(n4924) );
  IV U11040 ( .A(n9989), .Z(n9992) );
  XOR U11041 ( .A(n4923), .B(n9989), .Z(n9990) );
  XOR U11042 ( .A(n9993), .B(n9994), .Z(n9989) );
  ANDN U11043 ( .B(n9995), .A(n4934), .Z(n9993) );
  XNOR U11044 ( .A(n9996), .B(n9997), .Z(n4934) );
  IV U11045 ( .A(n9994), .Z(n9997) );
  XOR U11046 ( .A(n4933), .B(n9994), .Z(n9995) );
  XOR U11047 ( .A(n9998), .B(n9999), .Z(n9994) );
  ANDN U11048 ( .B(n10000), .A(n4939), .Z(n9998) );
  XNOR U11049 ( .A(n10001), .B(n10002), .Z(n4939) );
  IV U11050 ( .A(n9999), .Z(n10002) );
  XOR U11051 ( .A(n4938), .B(n9999), .Z(n10000) );
  XOR U11052 ( .A(n10003), .B(n10004), .Z(n9999) );
  ANDN U11053 ( .B(n10005), .A(n4944), .Z(n10003) );
  XNOR U11054 ( .A(n10006), .B(n10007), .Z(n4944) );
  IV U11055 ( .A(n10004), .Z(n10007) );
  XOR U11056 ( .A(n4943), .B(n10004), .Z(n10005) );
  XOR U11057 ( .A(n10008), .B(n10009), .Z(n10004) );
  ANDN U11058 ( .B(n10010), .A(n4949), .Z(n10008) );
  XNOR U11059 ( .A(n10011), .B(n10012), .Z(n4949) );
  IV U11060 ( .A(n10009), .Z(n10012) );
  XOR U11061 ( .A(n4948), .B(n10009), .Z(n10010) );
  XOR U11062 ( .A(n10013), .B(n10014), .Z(n10009) );
  ANDN U11063 ( .B(n10015), .A(n4954), .Z(n10013) );
  XNOR U11064 ( .A(n10016), .B(n10017), .Z(n4954) );
  IV U11065 ( .A(n10014), .Z(n10017) );
  XOR U11066 ( .A(n4953), .B(n10014), .Z(n10015) );
  XOR U11067 ( .A(n10018), .B(n10019), .Z(n10014) );
  ANDN U11068 ( .B(n10020), .A(n4959), .Z(n10018) );
  XNOR U11069 ( .A(n10021), .B(n10022), .Z(n4959) );
  IV U11070 ( .A(n10019), .Z(n10022) );
  XOR U11071 ( .A(n4958), .B(n10019), .Z(n10020) );
  XOR U11072 ( .A(n10023), .B(n10024), .Z(n10019) );
  ANDN U11073 ( .B(n10025), .A(n4964), .Z(n10023) );
  XNOR U11074 ( .A(n10026), .B(n10027), .Z(n4964) );
  IV U11075 ( .A(n10024), .Z(n10027) );
  XOR U11076 ( .A(n4963), .B(n10024), .Z(n10025) );
  XOR U11077 ( .A(n10028), .B(n10029), .Z(n10024) );
  ANDN U11078 ( .B(n10030), .A(n4969), .Z(n10028) );
  XNOR U11079 ( .A(n10031), .B(n10032), .Z(n4969) );
  IV U11080 ( .A(n10029), .Z(n10032) );
  XOR U11081 ( .A(n4968), .B(n10029), .Z(n10030) );
  XOR U11082 ( .A(n10033), .B(n10034), .Z(n10029) );
  ANDN U11083 ( .B(n10035), .A(n4974), .Z(n10033) );
  XNOR U11084 ( .A(n10036), .B(n10037), .Z(n4974) );
  IV U11085 ( .A(n10034), .Z(n10037) );
  XOR U11086 ( .A(n4973), .B(n10034), .Z(n10035) );
  XOR U11087 ( .A(n10038), .B(n10039), .Z(n10034) );
  ANDN U11088 ( .B(n10040), .A(n4979), .Z(n10038) );
  XNOR U11089 ( .A(n10041), .B(n10042), .Z(n4979) );
  IV U11090 ( .A(n10039), .Z(n10042) );
  XOR U11091 ( .A(n4978), .B(n10039), .Z(n10040) );
  XOR U11092 ( .A(n10043), .B(n10044), .Z(n10039) );
  ANDN U11093 ( .B(n10045), .A(n4989), .Z(n10043) );
  XNOR U11094 ( .A(n10046), .B(n10047), .Z(n4989) );
  IV U11095 ( .A(n10044), .Z(n10047) );
  XOR U11096 ( .A(n4988), .B(n10044), .Z(n10045) );
  XOR U11097 ( .A(n10048), .B(n10049), .Z(n10044) );
  ANDN U11098 ( .B(n10050), .A(n4994), .Z(n10048) );
  XNOR U11099 ( .A(n10051), .B(n10052), .Z(n4994) );
  IV U11100 ( .A(n10049), .Z(n10052) );
  XOR U11101 ( .A(n4993), .B(n10049), .Z(n10050) );
  XOR U11102 ( .A(n10053), .B(n10054), .Z(n10049) );
  ANDN U11103 ( .B(n10055), .A(n4999), .Z(n10053) );
  XNOR U11104 ( .A(n10056), .B(n10057), .Z(n4999) );
  IV U11105 ( .A(n10054), .Z(n10057) );
  XOR U11106 ( .A(n4998), .B(n10054), .Z(n10055) );
  XOR U11107 ( .A(n10058), .B(n10059), .Z(n10054) );
  ANDN U11108 ( .B(n10060), .A(n5004), .Z(n10058) );
  XNOR U11109 ( .A(n10061), .B(n10062), .Z(n5004) );
  IV U11110 ( .A(n10059), .Z(n10062) );
  XOR U11111 ( .A(n5003), .B(n10059), .Z(n10060) );
  XOR U11112 ( .A(n10063), .B(n10064), .Z(n10059) );
  ANDN U11113 ( .B(n10065), .A(n5009), .Z(n10063) );
  XNOR U11114 ( .A(n10066), .B(n10067), .Z(n5009) );
  IV U11115 ( .A(n10064), .Z(n10067) );
  XOR U11116 ( .A(n5008), .B(n10064), .Z(n10065) );
  XOR U11117 ( .A(n10068), .B(n10069), .Z(n10064) );
  ANDN U11118 ( .B(n10070), .A(n5014), .Z(n10068) );
  XNOR U11119 ( .A(n10071), .B(n10072), .Z(n5014) );
  IV U11120 ( .A(n10069), .Z(n10072) );
  XOR U11121 ( .A(n5013), .B(n10069), .Z(n10070) );
  XOR U11122 ( .A(n10073), .B(n10074), .Z(n10069) );
  ANDN U11123 ( .B(n10075), .A(n5019), .Z(n10073) );
  XNOR U11124 ( .A(n10076), .B(n10077), .Z(n5019) );
  IV U11125 ( .A(n10074), .Z(n10077) );
  XOR U11126 ( .A(n5018), .B(n10074), .Z(n10075) );
  XOR U11127 ( .A(n10078), .B(n10079), .Z(n10074) );
  ANDN U11128 ( .B(n10080), .A(n5024), .Z(n10078) );
  XNOR U11129 ( .A(n10081), .B(n10082), .Z(n5024) );
  IV U11130 ( .A(n10079), .Z(n10082) );
  XOR U11131 ( .A(n5023), .B(n10079), .Z(n10080) );
  XOR U11132 ( .A(n10083), .B(n10084), .Z(n10079) );
  ANDN U11133 ( .B(n10085), .A(n5029), .Z(n10083) );
  XNOR U11134 ( .A(n10086), .B(n10087), .Z(n5029) );
  IV U11135 ( .A(n10084), .Z(n10087) );
  XOR U11136 ( .A(n5028), .B(n10084), .Z(n10085) );
  XOR U11137 ( .A(n10088), .B(n10089), .Z(n10084) );
  ANDN U11138 ( .B(n10090), .A(n5034), .Z(n10088) );
  XNOR U11139 ( .A(n10091), .B(n10092), .Z(n5034) );
  IV U11140 ( .A(n10089), .Z(n10092) );
  XOR U11141 ( .A(n5033), .B(n10089), .Z(n10090) );
  XOR U11142 ( .A(n10093), .B(n10094), .Z(n10089) );
  ANDN U11143 ( .B(n10095), .A(n5044), .Z(n10093) );
  XNOR U11144 ( .A(n10096), .B(n10097), .Z(n5044) );
  IV U11145 ( .A(n10094), .Z(n10097) );
  XOR U11146 ( .A(n5043), .B(n10094), .Z(n10095) );
  XOR U11147 ( .A(n10098), .B(n10099), .Z(n10094) );
  ANDN U11148 ( .B(n10100), .A(n5049), .Z(n10098) );
  XNOR U11149 ( .A(n10101), .B(n10102), .Z(n5049) );
  IV U11150 ( .A(n10099), .Z(n10102) );
  XOR U11151 ( .A(n5048), .B(n10099), .Z(n10100) );
  XOR U11152 ( .A(n10103), .B(n10104), .Z(n10099) );
  ANDN U11153 ( .B(n10105), .A(n5054), .Z(n10103) );
  XNOR U11154 ( .A(n10106), .B(n10107), .Z(n5054) );
  IV U11155 ( .A(n10104), .Z(n10107) );
  XOR U11156 ( .A(n5053), .B(n10104), .Z(n10105) );
  XOR U11157 ( .A(n10108), .B(n10109), .Z(n10104) );
  ANDN U11158 ( .B(n10110), .A(n5059), .Z(n10108) );
  XNOR U11159 ( .A(n10111), .B(n10112), .Z(n5059) );
  IV U11160 ( .A(n10109), .Z(n10112) );
  XOR U11161 ( .A(n5058), .B(n10109), .Z(n10110) );
  XOR U11162 ( .A(n10113), .B(n10114), .Z(n10109) );
  ANDN U11163 ( .B(n10115), .A(n5064), .Z(n10113) );
  XNOR U11164 ( .A(n10116), .B(n10117), .Z(n5064) );
  IV U11165 ( .A(n10114), .Z(n10117) );
  XOR U11166 ( .A(n5063), .B(n10114), .Z(n10115) );
  XOR U11167 ( .A(n10118), .B(n10119), .Z(n10114) );
  ANDN U11168 ( .B(n10120), .A(n5069), .Z(n10118) );
  XNOR U11169 ( .A(n10121), .B(n10122), .Z(n5069) );
  IV U11170 ( .A(n10119), .Z(n10122) );
  XOR U11171 ( .A(n5068), .B(n10119), .Z(n10120) );
  XOR U11172 ( .A(n10123), .B(n10124), .Z(n10119) );
  ANDN U11173 ( .B(n10125), .A(n5074), .Z(n10123) );
  XNOR U11174 ( .A(n10126), .B(n10127), .Z(n5074) );
  IV U11175 ( .A(n10124), .Z(n10127) );
  XOR U11176 ( .A(n5073), .B(n10124), .Z(n10125) );
  XOR U11177 ( .A(n10128), .B(n10129), .Z(n10124) );
  ANDN U11178 ( .B(n10130), .A(n5079), .Z(n10128) );
  XNOR U11179 ( .A(n10131), .B(n10132), .Z(n5079) );
  IV U11180 ( .A(n10129), .Z(n10132) );
  XOR U11181 ( .A(n5078), .B(n10129), .Z(n10130) );
  XOR U11182 ( .A(n10133), .B(n10134), .Z(n10129) );
  ANDN U11183 ( .B(n10135), .A(n5084), .Z(n10133) );
  XNOR U11184 ( .A(n10136), .B(n10137), .Z(n5084) );
  IV U11185 ( .A(n10134), .Z(n10137) );
  XOR U11186 ( .A(n5083), .B(n10134), .Z(n10135) );
  XOR U11187 ( .A(n10138), .B(n10139), .Z(n10134) );
  ANDN U11188 ( .B(n10140), .A(n5089), .Z(n10138) );
  XNOR U11189 ( .A(n10141), .B(n10142), .Z(n5089) );
  IV U11190 ( .A(n10139), .Z(n10142) );
  XOR U11191 ( .A(n5088), .B(n10139), .Z(n10140) );
  XOR U11192 ( .A(n10143), .B(n10144), .Z(n10139) );
  ANDN U11193 ( .B(n10145), .A(n5099), .Z(n10143) );
  XNOR U11194 ( .A(n10146), .B(n10147), .Z(n5099) );
  IV U11195 ( .A(n10144), .Z(n10147) );
  XOR U11196 ( .A(n5098), .B(n10144), .Z(n10145) );
  XOR U11197 ( .A(n10148), .B(n10149), .Z(n10144) );
  ANDN U11198 ( .B(n10150), .A(n5104), .Z(n10148) );
  XNOR U11199 ( .A(n10151), .B(n10152), .Z(n5104) );
  IV U11200 ( .A(n10149), .Z(n10152) );
  XOR U11201 ( .A(n5103), .B(n10149), .Z(n10150) );
  XOR U11202 ( .A(n10153), .B(n10154), .Z(n10149) );
  ANDN U11203 ( .B(n10155), .A(n5109), .Z(n10153) );
  XNOR U11204 ( .A(n10156), .B(n10157), .Z(n5109) );
  IV U11205 ( .A(n10154), .Z(n10157) );
  XOR U11206 ( .A(n5108), .B(n10154), .Z(n10155) );
  XOR U11207 ( .A(n10158), .B(n10159), .Z(n10154) );
  ANDN U11208 ( .B(n10160), .A(n5114), .Z(n10158) );
  XNOR U11209 ( .A(n10161), .B(n10162), .Z(n5114) );
  IV U11210 ( .A(n10159), .Z(n10162) );
  XOR U11211 ( .A(n5113), .B(n10159), .Z(n10160) );
  XOR U11212 ( .A(n10163), .B(n10164), .Z(n10159) );
  ANDN U11213 ( .B(n10165), .A(n5119), .Z(n10163) );
  XNOR U11214 ( .A(n10166), .B(n10167), .Z(n5119) );
  IV U11215 ( .A(n10164), .Z(n10167) );
  XOR U11216 ( .A(n5118), .B(n10164), .Z(n10165) );
  XOR U11217 ( .A(n10168), .B(n10169), .Z(n10164) );
  ANDN U11218 ( .B(n10170), .A(n5124), .Z(n10168) );
  XNOR U11219 ( .A(n10171), .B(n10172), .Z(n5124) );
  IV U11220 ( .A(n10169), .Z(n10172) );
  XOR U11221 ( .A(n5123), .B(n10169), .Z(n10170) );
  XOR U11222 ( .A(n10173), .B(n10174), .Z(n10169) );
  ANDN U11223 ( .B(n10175), .A(n5129), .Z(n10173) );
  XNOR U11224 ( .A(n10176), .B(n10177), .Z(n5129) );
  IV U11225 ( .A(n10174), .Z(n10177) );
  XOR U11226 ( .A(n5128), .B(n10174), .Z(n10175) );
  XOR U11227 ( .A(n10178), .B(n10179), .Z(n10174) );
  ANDN U11228 ( .B(n10180), .A(n5134), .Z(n10178) );
  XNOR U11229 ( .A(n10181), .B(n10182), .Z(n5134) );
  IV U11230 ( .A(n10179), .Z(n10182) );
  XOR U11231 ( .A(n5133), .B(n10179), .Z(n10180) );
  XOR U11232 ( .A(n10183), .B(n10184), .Z(n10179) );
  ANDN U11233 ( .B(n10185), .A(n5139), .Z(n10183) );
  XNOR U11234 ( .A(n10186), .B(n10187), .Z(n5139) );
  IV U11235 ( .A(n10184), .Z(n10187) );
  XOR U11236 ( .A(n5138), .B(n10184), .Z(n10185) );
  XOR U11237 ( .A(n10188), .B(n10189), .Z(n10184) );
  ANDN U11238 ( .B(n10190), .A(n5144), .Z(n10188) );
  XNOR U11239 ( .A(n10191), .B(n10192), .Z(n5144) );
  IV U11240 ( .A(n10189), .Z(n10192) );
  XOR U11241 ( .A(n5143), .B(n10189), .Z(n10190) );
  XOR U11242 ( .A(n10193), .B(n10194), .Z(n10189) );
  ANDN U11243 ( .B(n10195), .A(n5154), .Z(n10193) );
  XNOR U11244 ( .A(n10196), .B(n10197), .Z(n5154) );
  IV U11245 ( .A(n10194), .Z(n10197) );
  XOR U11246 ( .A(n5153), .B(n10194), .Z(n10195) );
  XOR U11247 ( .A(n10198), .B(n10199), .Z(n10194) );
  ANDN U11248 ( .B(n10200), .A(n5159), .Z(n10198) );
  XNOR U11249 ( .A(n10201), .B(n10202), .Z(n5159) );
  IV U11250 ( .A(n10199), .Z(n10202) );
  XOR U11251 ( .A(n5158), .B(n10199), .Z(n10200) );
  XOR U11252 ( .A(n10203), .B(n10204), .Z(n10199) );
  ANDN U11253 ( .B(n10205), .A(n5164), .Z(n10203) );
  XNOR U11254 ( .A(n10206), .B(n10207), .Z(n5164) );
  IV U11255 ( .A(n10204), .Z(n10207) );
  XOR U11256 ( .A(n5163), .B(n10204), .Z(n10205) );
  XOR U11257 ( .A(n10208), .B(n10209), .Z(n10204) );
  ANDN U11258 ( .B(n10210), .A(n5169), .Z(n10208) );
  XNOR U11259 ( .A(n10211), .B(n10212), .Z(n5169) );
  IV U11260 ( .A(n10209), .Z(n10212) );
  XOR U11261 ( .A(n5168), .B(n10209), .Z(n10210) );
  XOR U11262 ( .A(n10213), .B(n10214), .Z(n10209) );
  ANDN U11263 ( .B(n10215), .A(n5174), .Z(n10213) );
  XNOR U11264 ( .A(n10216), .B(n10217), .Z(n5174) );
  IV U11265 ( .A(n10214), .Z(n10217) );
  XOR U11266 ( .A(n5173), .B(n10214), .Z(n10215) );
  XOR U11267 ( .A(n10218), .B(n10219), .Z(n10214) );
  ANDN U11268 ( .B(n10220), .A(n5179), .Z(n10218) );
  XNOR U11269 ( .A(n10221), .B(n10222), .Z(n5179) );
  IV U11270 ( .A(n10219), .Z(n10222) );
  XOR U11271 ( .A(n5178), .B(n10219), .Z(n10220) );
  XOR U11272 ( .A(n10223), .B(n10224), .Z(n10219) );
  ANDN U11273 ( .B(n10225), .A(n5184), .Z(n10223) );
  XNOR U11274 ( .A(n10226), .B(n10227), .Z(n5184) );
  IV U11275 ( .A(n10224), .Z(n10227) );
  XOR U11276 ( .A(n5183), .B(n10224), .Z(n10225) );
  XOR U11277 ( .A(n10228), .B(n10229), .Z(n10224) );
  ANDN U11278 ( .B(n10230), .A(n5189), .Z(n10228) );
  XNOR U11279 ( .A(n10231), .B(n10232), .Z(n5189) );
  IV U11280 ( .A(n10229), .Z(n10232) );
  XOR U11281 ( .A(n5188), .B(n10229), .Z(n10230) );
  XOR U11282 ( .A(n10233), .B(n10234), .Z(n10229) );
  ANDN U11283 ( .B(n10235), .A(n5194), .Z(n10233) );
  XNOR U11284 ( .A(n10236), .B(n10237), .Z(n5194) );
  IV U11285 ( .A(n10234), .Z(n10237) );
  XOR U11286 ( .A(n5193), .B(n10234), .Z(n10235) );
  XOR U11287 ( .A(n10238), .B(n10239), .Z(n10234) );
  ANDN U11288 ( .B(n10240), .A(n5199), .Z(n10238) );
  XNOR U11289 ( .A(n10241), .B(n10242), .Z(n5199) );
  IV U11290 ( .A(n10239), .Z(n10242) );
  XOR U11291 ( .A(n5198), .B(n10239), .Z(n10240) );
  XOR U11292 ( .A(n10243), .B(n10244), .Z(n10239) );
  ANDN U11293 ( .B(n10245), .A(n5209), .Z(n10243) );
  XNOR U11294 ( .A(n10246), .B(n10247), .Z(n5209) );
  IV U11295 ( .A(n10244), .Z(n10247) );
  XOR U11296 ( .A(n5208), .B(n10244), .Z(n10245) );
  XOR U11297 ( .A(n10248), .B(n10249), .Z(n10244) );
  ANDN U11298 ( .B(n10250), .A(n5214), .Z(n10248) );
  XNOR U11299 ( .A(n10251), .B(n10252), .Z(n5214) );
  IV U11300 ( .A(n10249), .Z(n10252) );
  XOR U11301 ( .A(n5213), .B(n10249), .Z(n10250) );
  XOR U11302 ( .A(n10253), .B(n10254), .Z(n10249) );
  ANDN U11303 ( .B(n10255), .A(n5219), .Z(n10253) );
  XNOR U11304 ( .A(n10256), .B(n10257), .Z(n5219) );
  IV U11305 ( .A(n10254), .Z(n10257) );
  XOR U11306 ( .A(n5218), .B(n10254), .Z(n10255) );
  XOR U11307 ( .A(n10258), .B(n10259), .Z(n10254) );
  ANDN U11308 ( .B(n10260), .A(n5224), .Z(n10258) );
  XNOR U11309 ( .A(n10261), .B(n10262), .Z(n5224) );
  IV U11310 ( .A(n10259), .Z(n10262) );
  XOR U11311 ( .A(n5223), .B(n10259), .Z(n10260) );
  XOR U11312 ( .A(n10263), .B(n10264), .Z(n10259) );
  ANDN U11313 ( .B(n10265), .A(n5229), .Z(n10263) );
  XNOR U11314 ( .A(n10266), .B(n10267), .Z(n5229) );
  IV U11315 ( .A(n10264), .Z(n10267) );
  XOR U11316 ( .A(n5228), .B(n10264), .Z(n10265) );
  XOR U11317 ( .A(n10268), .B(n10269), .Z(n10264) );
  ANDN U11318 ( .B(n10270), .A(n5234), .Z(n10268) );
  XNOR U11319 ( .A(n10271), .B(n10272), .Z(n5234) );
  IV U11320 ( .A(n10269), .Z(n10272) );
  XOR U11321 ( .A(n5233), .B(n10269), .Z(n10270) );
  XOR U11322 ( .A(n10273), .B(n10274), .Z(n10269) );
  ANDN U11323 ( .B(n10275), .A(n5239), .Z(n10273) );
  XNOR U11324 ( .A(n10276), .B(n10277), .Z(n5239) );
  IV U11325 ( .A(n10274), .Z(n10277) );
  XOR U11326 ( .A(n5238), .B(n10274), .Z(n10275) );
  XOR U11327 ( .A(n10278), .B(n10279), .Z(n10274) );
  ANDN U11328 ( .B(n10280), .A(n5244), .Z(n10278) );
  XNOR U11329 ( .A(n10281), .B(n10282), .Z(n5244) );
  IV U11330 ( .A(n10279), .Z(n10282) );
  XOR U11331 ( .A(n5243), .B(n10279), .Z(n10280) );
  XOR U11332 ( .A(n10283), .B(n10284), .Z(n10279) );
  ANDN U11333 ( .B(n10285), .A(n5249), .Z(n10283) );
  XNOR U11334 ( .A(n10286), .B(n10287), .Z(n5249) );
  IV U11335 ( .A(n10284), .Z(n10287) );
  XOR U11336 ( .A(n5248), .B(n10284), .Z(n10285) );
  XOR U11337 ( .A(n10288), .B(n10289), .Z(n10284) );
  ANDN U11338 ( .B(n10290), .A(n5254), .Z(n10288) );
  XNOR U11339 ( .A(n10291), .B(n10292), .Z(n5254) );
  IV U11340 ( .A(n10289), .Z(n10292) );
  XOR U11341 ( .A(n5253), .B(n10289), .Z(n10290) );
  XOR U11342 ( .A(n10293), .B(n10294), .Z(n10289) );
  ANDN U11343 ( .B(n10295), .A(n5264), .Z(n10293) );
  XNOR U11344 ( .A(n10296), .B(n10297), .Z(n5264) );
  IV U11345 ( .A(n10294), .Z(n10297) );
  XOR U11346 ( .A(n5263), .B(n10294), .Z(n10295) );
  XOR U11347 ( .A(n10298), .B(n10299), .Z(n10294) );
  ANDN U11348 ( .B(n10300), .A(n5269), .Z(n10298) );
  XNOR U11349 ( .A(n10301), .B(n10302), .Z(n5269) );
  IV U11350 ( .A(n10299), .Z(n10302) );
  XOR U11351 ( .A(n5268), .B(n10299), .Z(n10300) );
  XOR U11352 ( .A(n10303), .B(n10304), .Z(n10299) );
  ANDN U11353 ( .B(n10305), .A(n5274), .Z(n10303) );
  XNOR U11354 ( .A(n10306), .B(n10307), .Z(n5274) );
  IV U11355 ( .A(n10304), .Z(n10307) );
  XOR U11356 ( .A(n5273), .B(n10304), .Z(n10305) );
  XOR U11357 ( .A(n10308), .B(n10309), .Z(n10304) );
  ANDN U11358 ( .B(n10310), .A(n5279), .Z(n10308) );
  XNOR U11359 ( .A(n10311), .B(n10312), .Z(n5279) );
  IV U11360 ( .A(n10309), .Z(n10312) );
  XOR U11361 ( .A(n5278), .B(n10309), .Z(n10310) );
  XOR U11362 ( .A(n10313), .B(n10314), .Z(n10309) );
  ANDN U11363 ( .B(n10315), .A(n5284), .Z(n10313) );
  XNOR U11364 ( .A(n10316), .B(n10317), .Z(n5284) );
  IV U11365 ( .A(n10314), .Z(n10317) );
  XOR U11366 ( .A(n5283), .B(n10314), .Z(n10315) );
  XOR U11367 ( .A(n10318), .B(n10319), .Z(n10314) );
  ANDN U11368 ( .B(n10320), .A(n5289), .Z(n10318) );
  XNOR U11369 ( .A(n10321), .B(n10322), .Z(n5289) );
  IV U11370 ( .A(n10319), .Z(n10322) );
  XOR U11371 ( .A(n5288), .B(n10319), .Z(n10320) );
  XOR U11372 ( .A(n10323), .B(n10324), .Z(n10319) );
  ANDN U11373 ( .B(n10325), .A(n5294), .Z(n10323) );
  XNOR U11374 ( .A(n10326), .B(n10327), .Z(n5294) );
  IV U11375 ( .A(n10324), .Z(n10327) );
  XOR U11376 ( .A(n5293), .B(n10324), .Z(n10325) );
  XOR U11377 ( .A(n10328), .B(n10329), .Z(n10324) );
  ANDN U11378 ( .B(n10330), .A(n5299), .Z(n10328) );
  XNOR U11379 ( .A(n10331), .B(n10332), .Z(n5299) );
  IV U11380 ( .A(n10329), .Z(n10332) );
  XOR U11381 ( .A(n5298), .B(n10329), .Z(n10330) );
  XOR U11382 ( .A(n10333), .B(n10334), .Z(n10329) );
  ANDN U11383 ( .B(n10335), .A(n5304), .Z(n10333) );
  XNOR U11384 ( .A(n10336), .B(n10337), .Z(n5304) );
  IV U11385 ( .A(n10334), .Z(n10337) );
  XOR U11386 ( .A(n5303), .B(n10334), .Z(n10335) );
  XOR U11387 ( .A(n10338), .B(n10339), .Z(n10334) );
  ANDN U11388 ( .B(n10340), .A(n5309), .Z(n10338) );
  XNOR U11389 ( .A(n10341), .B(n10342), .Z(n5309) );
  IV U11390 ( .A(n10339), .Z(n10342) );
  XOR U11391 ( .A(n5308), .B(n10339), .Z(n10340) );
  XOR U11392 ( .A(n10343), .B(n10344), .Z(n10339) );
  ANDN U11393 ( .B(n10345), .A(n5324), .Z(n10343) );
  XNOR U11394 ( .A(n10346), .B(n10347), .Z(n5324) );
  IV U11395 ( .A(n10344), .Z(n10347) );
  XOR U11396 ( .A(n5323), .B(n10344), .Z(n10345) );
  XOR U11397 ( .A(n10348), .B(n10349), .Z(n10344) );
  ANDN U11398 ( .B(n10350), .A(n5329), .Z(n10348) );
  XNOR U11399 ( .A(n10351), .B(n10352), .Z(n5329) );
  IV U11400 ( .A(n10349), .Z(n10352) );
  XOR U11401 ( .A(n5328), .B(n10349), .Z(n10350) );
  XOR U11402 ( .A(n10353), .B(n10354), .Z(n10349) );
  ANDN U11403 ( .B(n10355), .A(n5334), .Z(n10353) );
  XNOR U11404 ( .A(n10356), .B(n10357), .Z(n5334) );
  IV U11405 ( .A(n10354), .Z(n10357) );
  XOR U11406 ( .A(n5333), .B(n10354), .Z(n10355) );
  XOR U11407 ( .A(n10358), .B(n10359), .Z(n10354) );
  ANDN U11408 ( .B(n10360), .A(n5339), .Z(n10358) );
  XNOR U11409 ( .A(n10361), .B(n10362), .Z(n5339) );
  IV U11410 ( .A(n10359), .Z(n10362) );
  XOR U11411 ( .A(n5338), .B(n10359), .Z(n10360) );
  XOR U11412 ( .A(n10363), .B(n10364), .Z(n10359) );
  ANDN U11413 ( .B(n10365), .A(n5344), .Z(n10363) );
  XNOR U11414 ( .A(n10366), .B(n10367), .Z(n5344) );
  IV U11415 ( .A(n10364), .Z(n10367) );
  XOR U11416 ( .A(n5343), .B(n10364), .Z(n10365) );
  XOR U11417 ( .A(n10368), .B(n10369), .Z(n10364) );
  ANDN U11418 ( .B(n10370), .A(n5349), .Z(n10368) );
  XNOR U11419 ( .A(n10371), .B(n10372), .Z(n5349) );
  IV U11420 ( .A(n10369), .Z(n10372) );
  XOR U11421 ( .A(n5348), .B(n10369), .Z(n10370) );
  XOR U11422 ( .A(n10373), .B(n10374), .Z(n10369) );
  ANDN U11423 ( .B(n10375), .A(n5354), .Z(n10373) );
  XNOR U11424 ( .A(n10376), .B(n10377), .Z(n5354) );
  IV U11425 ( .A(n10374), .Z(n10377) );
  XOR U11426 ( .A(n5353), .B(n10374), .Z(n10375) );
  XOR U11427 ( .A(n10378), .B(n10379), .Z(n10374) );
  ANDN U11428 ( .B(n10380), .A(n5359), .Z(n10378) );
  XNOR U11429 ( .A(n10381), .B(n10382), .Z(n5359) );
  IV U11430 ( .A(n10379), .Z(n10382) );
  XOR U11431 ( .A(n5358), .B(n10379), .Z(n10380) );
  XOR U11432 ( .A(n10383), .B(n10384), .Z(n10379) );
  ANDN U11433 ( .B(n10385), .A(n5364), .Z(n10383) );
  XNOR U11434 ( .A(n10386), .B(n10387), .Z(n5364) );
  IV U11435 ( .A(n10384), .Z(n10387) );
  XOR U11436 ( .A(n5363), .B(n10384), .Z(n10385) );
  XOR U11437 ( .A(n10388), .B(n10389), .Z(n10384) );
  ANDN U11438 ( .B(n10390), .A(n5369), .Z(n10388) );
  XNOR U11439 ( .A(n10391), .B(n10392), .Z(n5369) );
  IV U11440 ( .A(n10389), .Z(n10392) );
  XOR U11441 ( .A(n5368), .B(n10389), .Z(n10390) );
  XOR U11442 ( .A(n10393), .B(n10394), .Z(n10389) );
  ANDN U11443 ( .B(n10395), .A(n5379), .Z(n10393) );
  XNOR U11444 ( .A(n10396), .B(n10397), .Z(n5379) );
  IV U11445 ( .A(n10394), .Z(n10397) );
  XOR U11446 ( .A(n5378), .B(n10394), .Z(n10395) );
  XOR U11447 ( .A(n10398), .B(n10399), .Z(n10394) );
  ANDN U11448 ( .B(n10400), .A(n5384), .Z(n10398) );
  XNOR U11449 ( .A(n10401), .B(n10402), .Z(n5384) );
  IV U11450 ( .A(n10399), .Z(n10402) );
  XOR U11451 ( .A(n5383), .B(n10399), .Z(n10400) );
  XOR U11452 ( .A(n10403), .B(n10404), .Z(n10399) );
  ANDN U11453 ( .B(n10405), .A(n5389), .Z(n10403) );
  XNOR U11454 ( .A(n10406), .B(n10407), .Z(n5389) );
  IV U11455 ( .A(n10404), .Z(n10407) );
  XOR U11456 ( .A(n5388), .B(n10404), .Z(n10405) );
  XOR U11457 ( .A(n10408), .B(n10409), .Z(n10404) );
  ANDN U11458 ( .B(n10410), .A(n5394), .Z(n10408) );
  XNOR U11459 ( .A(n10411), .B(n10412), .Z(n5394) );
  IV U11460 ( .A(n10409), .Z(n10412) );
  XOR U11461 ( .A(n5393), .B(n10409), .Z(n10410) );
  XOR U11462 ( .A(n10413), .B(n10414), .Z(n10409) );
  ANDN U11463 ( .B(n10415), .A(n5399), .Z(n10413) );
  XNOR U11464 ( .A(n10416), .B(n10417), .Z(n5399) );
  IV U11465 ( .A(n10414), .Z(n10417) );
  XOR U11466 ( .A(n5398), .B(n10414), .Z(n10415) );
  XOR U11467 ( .A(n10418), .B(n10419), .Z(n10414) );
  ANDN U11468 ( .B(n10420), .A(n5404), .Z(n10418) );
  XNOR U11469 ( .A(n10421), .B(n10422), .Z(n5404) );
  IV U11470 ( .A(n10419), .Z(n10422) );
  XOR U11471 ( .A(n5403), .B(n10419), .Z(n10420) );
  XOR U11472 ( .A(n10423), .B(n10424), .Z(n10419) );
  ANDN U11473 ( .B(n10425), .A(n5409), .Z(n10423) );
  XNOR U11474 ( .A(n10426), .B(n10427), .Z(n5409) );
  IV U11475 ( .A(n10424), .Z(n10427) );
  XOR U11476 ( .A(n5408), .B(n10424), .Z(n10425) );
  XOR U11477 ( .A(n10428), .B(n10429), .Z(n10424) );
  ANDN U11478 ( .B(n10430), .A(n5414), .Z(n10428) );
  XNOR U11479 ( .A(n10431), .B(n10432), .Z(n5414) );
  IV U11480 ( .A(n10429), .Z(n10432) );
  XOR U11481 ( .A(n5413), .B(n10429), .Z(n10430) );
  XOR U11482 ( .A(n10433), .B(n10434), .Z(n10429) );
  ANDN U11483 ( .B(n10435), .A(n5419), .Z(n10433) );
  XNOR U11484 ( .A(n10436), .B(n10437), .Z(n5419) );
  IV U11485 ( .A(n10434), .Z(n10437) );
  XOR U11486 ( .A(n5418), .B(n10434), .Z(n10435) );
  XOR U11487 ( .A(n10438), .B(n10439), .Z(n10434) );
  ANDN U11488 ( .B(n10440), .A(n5424), .Z(n10438) );
  XNOR U11489 ( .A(n10441), .B(n10442), .Z(n5424) );
  IV U11490 ( .A(n10439), .Z(n10442) );
  XOR U11491 ( .A(n5423), .B(n10439), .Z(n10440) );
  XOR U11492 ( .A(n10443), .B(n10444), .Z(n10439) );
  ANDN U11493 ( .B(n10445), .A(n5434), .Z(n10443) );
  XNOR U11494 ( .A(n10446), .B(n10447), .Z(n5434) );
  IV U11495 ( .A(n10444), .Z(n10447) );
  XOR U11496 ( .A(n5433), .B(n10444), .Z(n10445) );
  XOR U11497 ( .A(n10448), .B(n10449), .Z(n10444) );
  ANDN U11498 ( .B(n10450), .A(n5439), .Z(n10448) );
  XNOR U11499 ( .A(n10451), .B(n10452), .Z(n5439) );
  IV U11500 ( .A(n10449), .Z(n10452) );
  XOR U11501 ( .A(n5438), .B(n10449), .Z(n10450) );
  XOR U11502 ( .A(n10453), .B(n10454), .Z(n10449) );
  ANDN U11503 ( .B(n10455), .A(n5444), .Z(n10453) );
  XNOR U11504 ( .A(n10456), .B(n10457), .Z(n5444) );
  IV U11505 ( .A(n10454), .Z(n10457) );
  XOR U11506 ( .A(n5443), .B(n10454), .Z(n10455) );
  XOR U11507 ( .A(n10458), .B(n10459), .Z(n10454) );
  ANDN U11508 ( .B(n10460), .A(n5449), .Z(n10458) );
  XNOR U11509 ( .A(n10461), .B(n10462), .Z(n5449) );
  IV U11510 ( .A(n10459), .Z(n10462) );
  XOR U11511 ( .A(n5448), .B(n10459), .Z(n10460) );
  XOR U11512 ( .A(n10463), .B(n10464), .Z(n10459) );
  ANDN U11513 ( .B(n10465), .A(n5454), .Z(n10463) );
  XNOR U11514 ( .A(n10466), .B(n10467), .Z(n5454) );
  IV U11515 ( .A(n10464), .Z(n10467) );
  XOR U11516 ( .A(n5453), .B(n10464), .Z(n10465) );
  XOR U11517 ( .A(n10468), .B(n10469), .Z(n10464) );
  ANDN U11518 ( .B(n10470), .A(n5459), .Z(n10468) );
  XNOR U11519 ( .A(n10471), .B(n10472), .Z(n5459) );
  IV U11520 ( .A(n10469), .Z(n10472) );
  XOR U11521 ( .A(n5458), .B(n10469), .Z(n10470) );
  XOR U11522 ( .A(n10473), .B(n10474), .Z(n10469) );
  ANDN U11523 ( .B(n10475), .A(n5464), .Z(n10473) );
  XNOR U11524 ( .A(n10476), .B(n10477), .Z(n5464) );
  IV U11525 ( .A(n10474), .Z(n10477) );
  XOR U11526 ( .A(n5463), .B(n10474), .Z(n10475) );
  XOR U11527 ( .A(n10478), .B(n10479), .Z(n10474) );
  ANDN U11528 ( .B(n10480), .A(n5469), .Z(n10478) );
  XNOR U11529 ( .A(n10481), .B(n10482), .Z(n5469) );
  IV U11530 ( .A(n10479), .Z(n10482) );
  XOR U11531 ( .A(n5468), .B(n10479), .Z(n10480) );
  XOR U11532 ( .A(n10483), .B(n10484), .Z(n10479) );
  ANDN U11533 ( .B(n10485), .A(n5474), .Z(n10483) );
  XNOR U11534 ( .A(n10486), .B(n10487), .Z(n5474) );
  IV U11535 ( .A(n10484), .Z(n10487) );
  XOR U11536 ( .A(n5473), .B(n10484), .Z(n10485) );
  XOR U11537 ( .A(n10488), .B(n10489), .Z(n10484) );
  ANDN U11538 ( .B(n10490), .A(n5479), .Z(n10488) );
  XNOR U11539 ( .A(n10491), .B(n10492), .Z(n5479) );
  IV U11540 ( .A(n10489), .Z(n10492) );
  XOR U11541 ( .A(n5478), .B(n10489), .Z(n10490) );
  XOR U11542 ( .A(n10493), .B(n10494), .Z(n10489) );
  ANDN U11543 ( .B(n10495), .A(n5489), .Z(n10493) );
  XNOR U11544 ( .A(n10496), .B(n10497), .Z(n5489) );
  IV U11545 ( .A(n10494), .Z(n10497) );
  XOR U11546 ( .A(n5488), .B(n10494), .Z(n10495) );
  XOR U11547 ( .A(n10498), .B(n10499), .Z(n10494) );
  ANDN U11548 ( .B(n10500), .A(n5494), .Z(n10498) );
  XNOR U11549 ( .A(n10501), .B(n10502), .Z(n5494) );
  IV U11550 ( .A(n10499), .Z(n10502) );
  XOR U11551 ( .A(n5493), .B(n10499), .Z(n10500) );
  XOR U11552 ( .A(n10503), .B(n10504), .Z(n10499) );
  ANDN U11553 ( .B(n10505), .A(n5499), .Z(n10503) );
  XNOR U11554 ( .A(n10506), .B(n10507), .Z(n5499) );
  IV U11555 ( .A(n10504), .Z(n10507) );
  XOR U11556 ( .A(n5498), .B(n10504), .Z(n10505) );
  XOR U11557 ( .A(n10508), .B(n10509), .Z(n10504) );
  ANDN U11558 ( .B(n10510), .A(n5504), .Z(n10508) );
  XNOR U11559 ( .A(n10511), .B(n10512), .Z(n5504) );
  IV U11560 ( .A(n10509), .Z(n10512) );
  XOR U11561 ( .A(n5503), .B(n10509), .Z(n10510) );
  XOR U11562 ( .A(n10513), .B(n10514), .Z(n10509) );
  ANDN U11563 ( .B(n10515), .A(n5509), .Z(n10513) );
  XNOR U11564 ( .A(n10516), .B(n10517), .Z(n5509) );
  IV U11565 ( .A(n10514), .Z(n10517) );
  XOR U11566 ( .A(n5508), .B(n10514), .Z(n10515) );
  XOR U11567 ( .A(n10518), .B(n10519), .Z(n10514) );
  ANDN U11568 ( .B(n10520), .A(n5514), .Z(n10518) );
  XNOR U11569 ( .A(n10521), .B(n10522), .Z(n5514) );
  IV U11570 ( .A(n10519), .Z(n10522) );
  XOR U11571 ( .A(n5513), .B(n10519), .Z(n10520) );
  XOR U11572 ( .A(n10523), .B(n10524), .Z(n10519) );
  ANDN U11573 ( .B(n10525), .A(n5519), .Z(n10523) );
  XNOR U11574 ( .A(n10526), .B(n10527), .Z(n5519) );
  IV U11575 ( .A(n10524), .Z(n10527) );
  XOR U11576 ( .A(n5518), .B(n10524), .Z(n10525) );
  XOR U11577 ( .A(n10528), .B(n10529), .Z(n10524) );
  ANDN U11578 ( .B(n10530), .A(n5524), .Z(n10528) );
  XNOR U11579 ( .A(n10531), .B(n10532), .Z(n5524) );
  IV U11580 ( .A(n10529), .Z(n10532) );
  XOR U11581 ( .A(n5523), .B(n10529), .Z(n10530) );
  XOR U11582 ( .A(n10533), .B(n10534), .Z(n10529) );
  ANDN U11583 ( .B(n10535), .A(n5529), .Z(n10533) );
  XNOR U11584 ( .A(n10536), .B(n10537), .Z(n5529) );
  IV U11585 ( .A(n10534), .Z(n10537) );
  XOR U11586 ( .A(n5528), .B(n10534), .Z(n10535) );
  XOR U11587 ( .A(n10538), .B(n10539), .Z(n10534) );
  ANDN U11588 ( .B(n10540), .A(n5534), .Z(n10538) );
  XNOR U11589 ( .A(n10541), .B(n10542), .Z(n5534) );
  IV U11590 ( .A(n10539), .Z(n10542) );
  XOR U11591 ( .A(n5533), .B(n10539), .Z(n10540) );
  XOR U11592 ( .A(n10543), .B(n10544), .Z(n10539) );
  ANDN U11593 ( .B(n10545), .A(n5544), .Z(n10543) );
  XNOR U11594 ( .A(n10546), .B(n10547), .Z(n5544) );
  IV U11595 ( .A(n10544), .Z(n10547) );
  XOR U11596 ( .A(n5543), .B(n10544), .Z(n10545) );
  XOR U11597 ( .A(n10548), .B(n10549), .Z(n10544) );
  ANDN U11598 ( .B(n10550), .A(n5549), .Z(n10548) );
  XNOR U11599 ( .A(n10551), .B(n10552), .Z(n5549) );
  IV U11600 ( .A(n10549), .Z(n10552) );
  XOR U11601 ( .A(n5548), .B(n10549), .Z(n10550) );
  XOR U11602 ( .A(n10553), .B(n10554), .Z(n10549) );
  ANDN U11603 ( .B(n10555), .A(n5554), .Z(n10553) );
  XNOR U11604 ( .A(n10556), .B(n10557), .Z(n5554) );
  IV U11605 ( .A(n10554), .Z(n10557) );
  XOR U11606 ( .A(n5553), .B(n10554), .Z(n10555) );
  XOR U11607 ( .A(n10558), .B(n10559), .Z(n10554) );
  ANDN U11608 ( .B(n10560), .A(n5559), .Z(n10558) );
  XNOR U11609 ( .A(n10561), .B(n10562), .Z(n5559) );
  IV U11610 ( .A(n10559), .Z(n10562) );
  XOR U11611 ( .A(n5558), .B(n10559), .Z(n10560) );
  XOR U11612 ( .A(n10563), .B(n10564), .Z(n10559) );
  ANDN U11613 ( .B(n10565), .A(n5564), .Z(n10563) );
  XNOR U11614 ( .A(n10566), .B(n10567), .Z(n5564) );
  IV U11615 ( .A(n10564), .Z(n10567) );
  XOR U11616 ( .A(n5563), .B(n10564), .Z(n10565) );
  XOR U11617 ( .A(n10568), .B(n10569), .Z(n10564) );
  ANDN U11618 ( .B(n10570), .A(n5569), .Z(n10568) );
  XNOR U11619 ( .A(n10571), .B(n10572), .Z(n5569) );
  IV U11620 ( .A(n10569), .Z(n10572) );
  XOR U11621 ( .A(n5568), .B(n10569), .Z(n10570) );
  XOR U11622 ( .A(n10573), .B(n10574), .Z(n10569) );
  ANDN U11623 ( .B(n10575), .A(n5574), .Z(n10573) );
  XNOR U11624 ( .A(n10576), .B(n10577), .Z(n5574) );
  IV U11625 ( .A(n10574), .Z(n10577) );
  XOR U11626 ( .A(n5573), .B(n10574), .Z(n10575) );
  XOR U11627 ( .A(n10578), .B(n10579), .Z(n10574) );
  ANDN U11628 ( .B(n10580), .A(n5579), .Z(n10578) );
  XNOR U11629 ( .A(n10581), .B(n10582), .Z(n5579) );
  IV U11630 ( .A(n10579), .Z(n10582) );
  XOR U11631 ( .A(n5578), .B(n10579), .Z(n10580) );
  XOR U11632 ( .A(n10583), .B(n10584), .Z(n10579) );
  ANDN U11633 ( .B(n10585), .A(n5584), .Z(n10583) );
  XNOR U11634 ( .A(n10586), .B(n10587), .Z(n5584) );
  IV U11635 ( .A(n10584), .Z(n10587) );
  XOR U11636 ( .A(n5583), .B(n10584), .Z(n10585) );
  XOR U11637 ( .A(n10588), .B(n10589), .Z(n10584) );
  ANDN U11638 ( .B(n10590), .A(n5589), .Z(n10588) );
  XNOR U11639 ( .A(n10591), .B(n10592), .Z(n5589) );
  IV U11640 ( .A(n10589), .Z(n10592) );
  XOR U11641 ( .A(n5588), .B(n10589), .Z(n10590) );
  XOR U11642 ( .A(n10593), .B(n10594), .Z(n10589) );
  ANDN U11643 ( .B(n10595), .A(n5599), .Z(n10593) );
  XNOR U11644 ( .A(n10596), .B(n10597), .Z(n5599) );
  IV U11645 ( .A(n10594), .Z(n10597) );
  XOR U11646 ( .A(n5598), .B(n10594), .Z(n10595) );
  XOR U11647 ( .A(n10598), .B(n10599), .Z(n10594) );
  ANDN U11648 ( .B(n10600), .A(n5604), .Z(n10598) );
  XNOR U11649 ( .A(n10601), .B(n10602), .Z(n5604) );
  IV U11650 ( .A(n10599), .Z(n10602) );
  XOR U11651 ( .A(n5603), .B(n10599), .Z(n10600) );
  XOR U11652 ( .A(n10603), .B(n10604), .Z(n10599) );
  ANDN U11653 ( .B(n10605), .A(n5609), .Z(n10603) );
  XNOR U11654 ( .A(n10606), .B(n10607), .Z(n5609) );
  IV U11655 ( .A(n10604), .Z(n10607) );
  XOR U11656 ( .A(n5608), .B(n10604), .Z(n10605) );
  XOR U11657 ( .A(n10608), .B(n10609), .Z(n10604) );
  ANDN U11658 ( .B(n10610), .A(n5614), .Z(n10608) );
  XNOR U11659 ( .A(n10611), .B(n10612), .Z(n5614) );
  IV U11660 ( .A(n10609), .Z(n10612) );
  XOR U11661 ( .A(n5613), .B(n10609), .Z(n10610) );
  XOR U11662 ( .A(n10613), .B(n10614), .Z(n10609) );
  ANDN U11663 ( .B(n10615), .A(n5619), .Z(n10613) );
  XNOR U11664 ( .A(n10616), .B(n10617), .Z(n5619) );
  IV U11665 ( .A(n10614), .Z(n10617) );
  XOR U11666 ( .A(n5618), .B(n10614), .Z(n10615) );
  XOR U11667 ( .A(n10618), .B(n10619), .Z(n10614) );
  ANDN U11668 ( .B(n10620), .A(n5624), .Z(n10618) );
  XNOR U11669 ( .A(n10621), .B(n10622), .Z(n5624) );
  IV U11670 ( .A(n10619), .Z(n10622) );
  XOR U11671 ( .A(n5623), .B(n10619), .Z(n10620) );
  XOR U11672 ( .A(n10623), .B(n10624), .Z(n10619) );
  ANDN U11673 ( .B(n10625), .A(n5629), .Z(n10623) );
  XNOR U11674 ( .A(n10626), .B(n10627), .Z(n5629) );
  IV U11675 ( .A(n10624), .Z(n10627) );
  XOR U11676 ( .A(n5628), .B(n10624), .Z(n10625) );
  XOR U11677 ( .A(n10628), .B(n10629), .Z(n10624) );
  ANDN U11678 ( .B(n10630), .A(n5634), .Z(n10628) );
  XNOR U11679 ( .A(n10631), .B(n10632), .Z(n5634) );
  IV U11680 ( .A(n10629), .Z(n10632) );
  XOR U11681 ( .A(n5633), .B(n10629), .Z(n10630) );
  XOR U11682 ( .A(n10633), .B(n10634), .Z(n10629) );
  ANDN U11683 ( .B(n10635), .A(n5639), .Z(n10633) );
  XNOR U11684 ( .A(n10636), .B(n10637), .Z(n5639) );
  IV U11685 ( .A(n10634), .Z(n10637) );
  XOR U11686 ( .A(n5638), .B(n10634), .Z(n10635) );
  XOR U11687 ( .A(n10638), .B(n10639), .Z(n10634) );
  ANDN U11688 ( .B(n10640), .A(n5644), .Z(n10638) );
  XNOR U11689 ( .A(n10641), .B(n10642), .Z(n5644) );
  IV U11690 ( .A(n10639), .Z(n10642) );
  XOR U11691 ( .A(n5643), .B(n10639), .Z(n10640) );
  XOR U11692 ( .A(n10643), .B(n10644), .Z(n10639) );
  ANDN U11693 ( .B(n10645), .A(n5654), .Z(n10643) );
  XNOR U11694 ( .A(n10646), .B(n10647), .Z(n5654) );
  IV U11695 ( .A(n10644), .Z(n10647) );
  XOR U11696 ( .A(n5653), .B(n10644), .Z(n10645) );
  XOR U11697 ( .A(n10648), .B(n10649), .Z(n10644) );
  ANDN U11698 ( .B(n10650), .A(n5659), .Z(n10648) );
  XNOR U11699 ( .A(n10651), .B(n10652), .Z(n5659) );
  IV U11700 ( .A(n10649), .Z(n10652) );
  XOR U11701 ( .A(n5658), .B(n10649), .Z(n10650) );
  XOR U11702 ( .A(n10653), .B(n10654), .Z(n10649) );
  ANDN U11703 ( .B(n10655), .A(n5664), .Z(n10653) );
  XNOR U11704 ( .A(n10656), .B(n10657), .Z(n5664) );
  IV U11705 ( .A(n10654), .Z(n10657) );
  XOR U11706 ( .A(n5663), .B(n10654), .Z(n10655) );
  XOR U11707 ( .A(n10658), .B(n10659), .Z(n10654) );
  ANDN U11708 ( .B(n10660), .A(n5669), .Z(n10658) );
  XNOR U11709 ( .A(n10661), .B(n10662), .Z(n5669) );
  IV U11710 ( .A(n10659), .Z(n10662) );
  XOR U11711 ( .A(n5668), .B(n10659), .Z(n10660) );
  XOR U11712 ( .A(n10663), .B(n10664), .Z(n10659) );
  ANDN U11713 ( .B(n10665), .A(n5674), .Z(n10663) );
  XNOR U11714 ( .A(n10666), .B(n10667), .Z(n5674) );
  IV U11715 ( .A(n10664), .Z(n10667) );
  XOR U11716 ( .A(n5673), .B(n10664), .Z(n10665) );
  XOR U11717 ( .A(n10668), .B(n10669), .Z(n10664) );
  ANDN U11718 ( .B(n10670), .A(n5679), .Z(n10668) );
  XNOR U11719 ( .A(n10671), .B(n10672), .Z(n5679) );
  IV U11720 ( .A(n10669), .Z(n10672) );
  XOR U11721 ( .A(n5678), .B(n10669), .Z(n10670) );
  XOR U11722 ( .A(n10673), .B(n10674), .Z(n10669) );
  ANDN U11723 ( .B(n10675), .A(n5684), .Z(n10673) );
  XNOR U11724 ( .A(n10676), .B(n10677), .Z(n5684) );
  IV U11725 ( .A(n10674), .Z(n10677) );
  XOR U11726 ( .A(n5683), .B(n10674), .Z(n10675) );
  XOR U11727 ( .A(n10678), .B(n10679), .Z(n10674) );
  ANDN U11728 ( .B(n10680), .A(n5689), .Z(n10678) );
  XNOR U11729 ( .A(n10681), .B(n10682), .Z(n5689) );
  IV U11730 ( .A(n10679), .Z(n10682) );
  XOR U11731 ( .A(n5688), .B(n10679), .Z(n10680) );
  XOR U11732 ( .A(n10683), .B(n10684), .Z(n10679) );
  ANDN U11733 ( .B(n10685), .A(n5694), .Z(n10683) );
  XNOR U11734 ( .A(n10686), .B(n10687), .Z(n5694) );
  IV U11735 ( .A(n10684), .Z(n10687) );
  XOR U11736 ( .A(n5693), .B(n10684), .Z(n10685) );
  XOR U11737 ( .A(n10688), .B(n10689), .Z(n10684) );
  ANDN U11738 ( .B(n10690), .A(n5699), .Z(n10688) );
  XNOR U11739 ( .A(n10691), .B(n10692), .Z(n5699) );
  IV U11740 ( .A(n10689), .Z(n10692) );
  XOR U11741 ( .A(n5698), .B(n10689), .Z(n10690) );
  XOR U11742 ( .A(n10693), .B(n10694), .Z(n10689) );
  ANDN U11743 ( .B(n10695), .A(n5709), .Z(n10693) );
  XNOR U11744 ( .A(n10696), .B(n10697), .Z(n5709) );
  IV U11745 ( .A(n10694), .Z(n10697) );
  XOR U11746 ( .A(n5708), .B(n10694), .Z(n10695) );
  XOR U11747 ( .A(n10698), .B(n10699), .Z(n10694) );
  ANDN U11748 ( .B(n10700), .A(n5714), .Z(n10698) );
  XNOR U11749 ( .A(n10701), .B(n10702), .Z(n5714) );
  IV U11750 ( .A(n10699), .Z(n10702) );
  XOR U11751 ( .A(n5713), .B(n10699), .Z(n10700) );
  XOR U11752 ( .A(n10703), .B(n10704), .Z(n10699) );
  ANDN U11753 ( .B(n10705), .A(n5719), .Z(n10703) );
  XNOR U11754 ( .A(n10706), .B(n10707), .Z(n5719) );
  IV U11755 ( .A(n10704), .Z(n10707) );
  XOR U11756 ( .A(n5718), .B(n10704), .Z(n10705) );
  XOR U11757 ( .A(n10708), .B(n10709), .Z(n10704) );
  ANDN U11758 ( .B(n10710), .A(n5724), .Z(n10708) );
  XNOR U11759 ( .A(n10711), .B(n10712), .Z(n5724) );
  IV U11760 ( .A(n10709), .Z(n10712) );
  XOR U11761 ( .A(n5723), .B(n10709), .Z(n10710) );
  XOR U11762 ( .A(n10713), .B(n10714), .Z(n10709) );
  ANDN U11763 ( .B(n10715), .A(n5729), .Z(n10713) );
  XNOR U11764 ( .A(n10716), .B(n10717), .Z(n5729) );
  IV U11765 ( .A(n10714), .Z(n10717) );
  XOR U11766 ( .A(n5728), .B(n10714), .Z(n10715) );
  XOR U11767 ( .A(n10718), .B(n10719), .Z(n10714) );
  ANDN U11768 ( .B(n10720), .A(n5734), .Z(n10718) );
  XNOR U11769 ( .A(n10721), .B(n10722), .Z(n5734) );
  IV U11770 ( .A(n10719), .Z(n10722) );
  XOR U11771 ( .A(n5733), .B(n10719), .Z(n10720) );
  XOR U11772 ( .A(n10723), .B(n10724), .Z(n10719) );
  ANDN U11773 ( .B(n10725), .A(n5739), .Z(n10723) );
  XNOR U11774 ( .A(n10726), .B(n10727), .Z(n5739) );
  IV U11775 ( .A(n10724), .Z(n10727) );
  XOR U11776 ( .A(n5738), .B(n10724), .Z(n10725) );
  XOR U11777 ( .A(n10728), .B(n10729), .Z(n10724) );
  ANDN U11778 ( .B(n10730), .A(n5744), .Z(n10728) );
  XNOR U11779 ( .A(n10731), .B(n10732), .Z(n5744) );
  IV U11780 ( .A(n10729), .Z(n10732) );
  XOR U11781 ( .A(n5743), .B(n10729), .Z(n10730) );
  XOR U11782 ( .A(n10733), .B(n10734), .Z(n10729) );
  ANDN U11783 ( .B(n10735), .A(n5749), .Z(n10733) );
  XNOR U11784 ( .A(n10736), .B(n10737), .Z(n5749) );
  IV U11785 ( .A(n10734), .Z(n10737) );
  XOR U11786 ( .A(n5748), .B(n10734), .Z(n10735) );
  XOR U11787 ( .A(n10738), .B(n10739), .Z(n10734) );
  ANDN U11788 ( .B(n10740), .A(n5754), .Z(n10738) );
  XNOR U11789 ( .A(n10741), .B(n10742), .Z(n5754) );
  IV U11790 ( .A(n10739), .Z(n10742) );
  XOR U11791 ( .A(n5753), .B(n10739), .Z(n10740) );
  XOR U11792 ( .A(n10743), .B(n10744), .Z(n10739) );
  ANDN U11793 ( .B(n10745), .A(n5764), .Z(n10743) );
  XNOR U11794 ( .A(n10746), .B(n10747), .Z(n5764) );
  IV U11795 ( .A(n10744), .Z(n10747) );
  XOR U11796 ( .A(n5763), .B(n10744), .Z(n10745) );
  XOR U11797 ( .A(n10748), .B(n10749), .Z(n10744) );
  ANDN U11798 ( .B(n10750), .A(n5769), .Z(n10748) );
  XNOR U11799 ( .A(n10751), .B(n10752), .Z(n5769) );
  IV U11800 ( .A(n10749), .Z(n10752) );
  XOR U11801 ( .A(n5768), .B(n10749), .Z(n10750) );
  XOR U11802 ( .A(n10753), .B(n10754), .Z(n10749) );
  ANDN U11803 ( .B(n10755), .A(n5774), .Z(n10753) );
  XNOR U11804 ( .A(n10756), .B(n10757), .Z(n5774) );
  IV U11805 ( .A(n10754), .Z(n10757) );
  XOR U11806 ( .A(n5773), .B(n10754), .Z(n10755) );
  XOR U11807 ( .A(n10758), .B(n10759), .Z(n10754) );
  ANDN U11808 ( .B(n10760), .A(n5779), .Z(n10758) );
  XNOR U11809 ( .A(n10761), .B(n10762), .Z(n5779) );
  IV U11810 ( .A(n10759), .Z(n10762) );
  XOR U11811 ( .A(n5778), .B(n10759), .Z(n10760) );
  XOR U11812 ( .A(n10763), .B(n10764), .Z(n10759) );
  ANDN U11813 ( .B(n10765), .A(n5784), .Z(n10763) );
  XNOR U11814 ( .A(n10766), .B(n10767), .Z(n5784) );
  IV U11815 ( .A(n10764), .Z(n10767) );
  XOR U11816 ( .A(n5783), .B(n10764), .Z(n10765) );
  XOR U11817 ( .A(n10768), .B(n10769), .Z(n10764) );
  ANDN U11818 ( .B(n10770), .A(n5789), .Z(n10768) );
  XNOR U11819 ( .A(n10771), .B(n10772), .Z(n5789) );
  IV U11820 ( .A(n10769), .Z(n10772) );
  XOR U11821 ( .A(n5788), .B(n10769), .Z(n10770) );
  XOR U11822 ( .A(n10773), .B(n10774), .Z(n10769) );
  ANDN U11823 ( .B(n10775), .A(n5794), .Z(n10773) );
  XNOR U11824 ( .A(n10776), .B(n10777), .Z(n5794) );
  IV U11825 ( .A(n10774), .Z(n10777) );
  XOR U11826 ( .A(n5793), .B(n10774), .Z(n10775) );
  XOR U11827 ( .A(n10778), .B(n10779), .Z(n10774) );
  ANDN U11828 ( .B(n10780), .A(n5799), .Z(n10778) );
  XNOR U11829 ( .A(n10781), .B(n10782), .Z(n5799) );
  IV U11830 ( .A(n10779), .Z(n10782) );
  XOR U11831 ( .A(n5798), .B(n10779), .Z(n10780) );
  XOR U11832 ( .A(n10783), .B(n10784), .Z(n10779) );
  ANDN U11833 ( .B(n10785), .A(n5804), .Z(n10783) );
  XNOR U11834 ( .A(n10786), .B(n10787), .Z(n5804) );
  IV U11835 ( .A(n10784), .Z(n10787) );
  XOR U11836 ( .A(n5803), .B(n10784), .Z(n10785) );
  XOR U11837 ( .A(n10788), .B(n10789), .Z(n10784) );
  ANDN U11838 ( .B(n10790), .A(n5809), .Z(n10788) );
  XNOR U11839 ( .A(n10791), .B(n10792), .Z(n5809) );
  IV U11840 ( .A(n10789), .Z(n10792) );
  XOR U11841 ( .A(n5808), .B(n10789), .Z(n10790) );
  XOR U11842 ( .A(n10793), .B(n10794), .Z(n10789) );
  ANDN U11843 ( .B(n10795), .A(n5819), .Z(n10793) );
  XNOR U11844 ( .A(n10796), .B(n10797), .Z(n5819) );
  IV U11845 ( .A(n10794), .Z(n10797) );
  XOR U11846 ( .A(n5818), .B(n10794), .Z(n10795) );
  XOR U11847 ( .A(n10798), .B(n10799), .Z(n10794) );
  ANDN U11848 ( .B(n10800), .A(n5824), .Z(n10798) );
  XNOR U11849 ( .A(n10801), .B(n10802), .Z(n5824) );
  IV U11850 ( .A(n10799), .Z(n10802) );
  XOR U11851 ( .A(n5823), .B(n10799), .Z(n10800) );
  XOR U11852 ( .A(n10803), .B(n10804), .Z(n10799) );
  ANDN U11853 ( .B(n10805), .A(n5829), .Z(n10803) );
  XNOR U11854 ( .A(n10806), .B(n10807), .Z(n5829) );
  IV U11855 ( .A(n10804), .Z(n10807) );
  XOR U11856 ( .A(n5828), .B(n10804), .Z(n10805) );
  XOR U11857 ( .A(n10808), .B(n10809), .Z(n10804) );
  ANDN U11858 ( .B(n10810), .A(n5834), .Z(n10808) );
  XNOR U11859 ( .A(n10811), .B(n10812), .Z(n5834) );
  IV U11860 ( .A(n10809), .Z(n10812) );
  XOR U11861 ( .A(n5833), .B(n10809), .Z(n10810) );
  XOR U11862 ( .A(n10813), .B(n10814), .Z(n10809) );
  ANDN U11863 ( .B(n10815), .A(n5839), .Z(n10813) );
  XNOR U11864 ( .A(n10816), .B(n10817), .Z(n5839) );
  IV U11865 ( .A(n10814), .Z(n10817) );
  XOR U11866 ( .A(n5838), .B(n10814), .Z(n10815) );
  XOR U11867 ( .A(n10818), .B(n10819), .Z(n10814) );
  ANDN U11868 ( .B(n10820), .A(n5844), .Z(n10818) );
  XNOR U11869 ( .A(n10821), .B(n10822), .Z(n5844) );
  IV U11870 ( .A(n10819), .Z(n10822) );
  XOR U11871 ( .A(n5843), .B(n10819), .Z(n10820) );
  XOR U11872 ( .A(n10823), .B(n10824), .Z(n10819) );
  ANDN U11873 ( .B(n10825), .A(n5849), .Z(n10823) );
  XNOR U11874 ( .A(n10826), .B(n10827), .Z(n5849) );
  IV U11875 ( .A(n10824), .Z(n10827) );
  XOR U11876 ( .A(n5848), .B(n10824), .Z(n10825) );
  XOR U11877 ( .A(n10828), .B(n10829), .Z(n10824) );
  ANDN U11878 ( .B(n10830), .A(n5854), .Z(n10828) );
  XNOR U11879 ( .A(n10831), .B(n10832), .Z(n5854) );
  IV U11880 ( .A(n10829), .Z(n10832) );
  XOR U11881 ( .A(n5853), .B(n10829), .Z(n10830) );
  XOR U11882 ( .A(n10833), .B(n10834), .Z(n10829) );
  ANDN U11883 ( .B(n10835), .A(n5859), .Z(n10833) );
  XNOR U11884 ( .A(n10836), .B(n10837), .Z(n5859) );
  IV U11885 ( .A(n10834), .Z(n10837) );
  XOR U11886 ( .A(n5858), .B(n10834), .Z(n10835) );
  XOR U11887 ( .A(n10838), .B(n10839), .Z(n10834) );
  ANDN U11888 ( .B(n10840), .A(n5864), .Z(n10838) );
  XNOR U11889 ( .A(n10841), .B(n10842), .Z(n5864) );
  IV U11890 ( .A(n10839), .Z(n10842) );
  XOR U11891 ( .A(n5863), .B(n10839), .Z(n10840) );
  XOR U11892 ( .A(n10843), .B(n10844), .Z(n10839) );
  ANDN U11893 ( .B(n10845), .A(n5879), .Z(n10843) );
  XNOR U11894 ( .A(n10846), .B(n10847), .Z(n5879) );
  IV U11895 ( .A(n10844), .Z(n10847) );
  XOR U11896 ( .A(n5878), .B(n10844), .Z(n10845) );
  XOR U11897 ( .A(n10848), .B(n10849), .Z(n10844) );
  ANDN U11898 ( .B(n10850), .A(n5884), .Z(n10848) );
  XNOR U11899 ( .A(n10851), .B(n10852), .Z(n5884) );
  IV U11900 ( .A(n10849), .Z(n10852) );
  XOR U11901 ( .A(n5883), .B(n10849), .Z(n10850) );
  XOR U11902 ( .A(n10853), .B(n10854), .Z(n10849) );
  ANDN U11903 ( .B(n10855), .A(n5889), .Z(n10853) );
  XNOR U11904 ( .A(n10856), .B(n10857), .Z(n5889) );
  IV U11905 ( .A(n10854), .Z(n10857) );
  XOR U11906 ( .A(n5888), .B(n10854), .Z(n10855) );
  XOR U11907 ( .A(n10858), .B(n10859), .Z(n10854) );
  ANDN U11908 ( .B(n10860), .A(n5894), .Z(n10858) );
  XNOR U11909 ( .A(n10861), .B(n10862), .Z(n5894) );
  IV U11910 ( .A(n10859), .Z(n10862) );
  XOR U11911 ( .A(n5893), .B(n10859), .Z(n10860) );
  XOR U11912 ( .A(n10863), .B(n10864), .Z(n10859) );
  ANDN U11913 ( .B(n10865), .A(n5899), .Z(n10863) );
  XNOR U11914 ( .A(n10866), .B(n10867), .Z(n5899) );
  IV U11915 ( .A(n10864), .Z(n10867) );
  XOR U11916 ( .A(n5898), .B(n10864), .Z(n10865) );
  XOR U11917 ( .A(n10868), .B(n10869), .Z(n10864) );
  ANDN U11918 ( .B(n10870), .A(n5904), .Z(n10868) );
  XNOR U11919 ( .A(n10871), .B(n10872), .Z(n5904) );
  IV U11920 ( .A(n10869), .Z(n10872) );
  XOR U11921 ( .A(n5903), .B(n10869), .Z(n10870) );
  XOR U11922 ( .A(n10873), .B(n10874), .Z(n10869) );
  ANDN U11923 ( .B(n10875), .A(n5909), .Z(n10873) );
  XNOR U11924 ( .A(n10876), .B(n10877), .Z(n5909) );
  IV U11925 ( .A(n10874), .Z(n10877) );
  XOR U11926 ( .A(n5908), .B(n10874), .Z(n10875) );
  XOR U11927 ( .A(n10878), .B(n10879), .Z(n10874) );
  ANDN U11928 ( .B(n10880), .A(n5914), .Z(n10878) );
  XNOR U11929 ( .A(n10881), .B(n10882), .Z(n5914) );
  IV U11930 ( .A(n10879), .Z(n10882) );
  XOR U11931 ( .A(n5913), .B(n10879), .Z(n10880) );
  XOR U11932 ( .A(n10883), .B(n10884), .Z(n10879) );
  ANDN U11933 ( .B(n10885), .A(n5919), .Z(n10883) );
  XNOR U11934 ( .A(n10886), .B(n10887), .Z(n5919) );
  IV U11935 ( .A(n10884), .Z(n10887) );
  XOR U11936 ( .A(n5918), .B(n10884), .Z(n10885) );
  XOR U11937 ( .A(n10888), .B(n10889), .Z(n10884) );
  ANDN U11938 ( .B(n10890), .A(n5924), .Z(n10888) );
  XNOR U11939 ( .A(n10891), .B(n10892), .Z(n5924) );
  IV U11940 ( .A(n10889), .Z(n10892) );
  XOR U11941 ( .A(n5923), .B(n10889), .Z(n10890) );
  XOR U11942 ( .A(n10893), .B(n10894), .Z(n10889) );
  ANDN U11943 ( .B(n10895), .A(n5934), .Z(n10893) );
  XNOR U11944 ( .A(n10896), .B(n10897), .Z(n5934) );
  IV U11945 ( .A(n10894), .Z(n10897) );
  XOR U11946 ( .A(n5933), .B(n10894), .Z(n10895) );
  XOR U11947 ( .A(n10898), .B(n10899), .Z(n10894) );
  ANDN U11948 ( .B(n10900), .A(n5939), .Z(n10898) );
  XNOR U11949 ( .A(n10901), .B(n10902), .Z(n5939) );
  IV U11950 ( .A(n10899), .Z(n10902) );
  XOR U11951 ( .A(n5938), .B(n10899), .Z(n10900) );
  XOR U11952 ( .A(n10903), .B(n10904), .Z(n10899) );
  ANDN U11953 ( .B(n10905), .A(n5944), .Z(n10903) );
  XNOR U11954 ( .A(n10906), .B(n10907), .Z(n5944) );
  IV U11955 ( .A(n10904), .Z(n10907) );
  XOR U11956 ( .A(n5943), .B(n10904), .Z(n10905) );
  XOR U11957 ( .A(n10908), .B(n10909), .Z(n10904) );
  ANDN U11958 ( .B(n10910), .A(n5949), .Z(n10908) );
  XNOR U11959 ( .A(n10911), .B(n10912), .Z(n5949) );
  IV U11960 ( .A(n10909), .Z(n10912) );
  XOR U11961 ( .A(n5948), .B(n10909), .Z(n10910) );
  XOR U11962 ( .A(n10913), .B(n10914), .Z(n10909) );
  ANDN U11963 ( .B(n10915), .A(n5954), .Z(n10913) );
  XNOR U11964 ( .A(n10916), .B(n10917), .Z(n5954) );
  IV U11965 ( .A(n10914), .Z(n10917) );
  XOR U11966 ( .A(n5953), .B(n10914), .Z(n10915) );
  XOR U11967 ( .A(n10918), .B(n10919), .Z(n10914) );
  ANDN U11968 ( .B(n10920), .A(n5959), .Z(n10918) );
  XNOR U11969 ( .A(n10921), .B(n10922), .Z(n5959) );
  IV U11970 ( .A(n10919), .Z(n10922) );
  XOR U11971 ( .A(n5958), .B(n10919), .Z(n10920) );
  XOR U11972 ( .A(n10923), .B(n10924), .Z(n10919) );
  ANDN U11973 ( .B(n10925), .A(n5964), .Z(n10923) );
  XNOR U11974 ( .A(n10926), .B(n10927), .Z(n5964) );
  IV U11975 ( .A(n10924), .Z(n10927) );
  XOR U11976 ( .A(n5963), .B(n10924), .Z(n10925) );
  XOR U11977 ( .A(n10928), .B(n10929), .Z(n10924) );
  ANDN U11978 ( .B(n10930), .A(n5969), .Z(n10928) );
  XNOR U11979 ( .A(n10931), .B(n10932), .Z(n5969) );
  IV U11980 ( .A(n10929), .Z(n10932) );
  XOR U11981 ( .A(n5968), .B(n10929), .Z(n10930) );
  XOR U11982 ( .A(n10933), .B(n10934), .Z(n10929) );
  ANDN U11983 ( .B(n10935), .A(n5974), .Z(n10933) );
  XNOR U11984 ( .A(n10936), .B(n10937), .Z(n5974) );
  IV U11985 ( .A(n10934), .Z(n10937) );
  XOR U11986 ( .A(n5973), .B(n10934), .Z(n10935) );
  XOR U11987 ( .A(n10938), .B(n10939), .Z(n10934) );
  ANDN U11988 ( .B(n10940), .A(n5979), .Z(n10938) );
  XNOR U11989 ( .A(n10941), .B(n10942), .Z(n5979) );
  IV U11990 ( .A(n10939), .Z(n10942) );
  XOR U11991 ( .A(n5978), .B(n10939), .Z(n10940) );
  XOR U11992 ( .A(n10943), .B(n10944), .Z(n10939) );
  ANDN U11993 ( .B(n10945), .A(n5989), .Z(n10943) );
  XNOR U11994 ( .A(n10946), .B(n10947), .Z(n5989) );
  IV U11995 ( .A(n10944), .Z(n10947) );
  XOR U11996 ( .A(n5988), .B(n10944), .Z(n10945) );
  XOR U11997 ( .A(n10948), .B(n10949), .Z(n10944) );
  ANDN U11998 ( .B(n10950), .A(n5994), .Z(n10948) );
  XNOR U11999 ( .A(n10951), .B(n10952), .Z(n5994) );
  IV U12000 ( .A(n10949), .Z(n10952) );
  XOR U12001 ( .A(n5993), .B(n10949), .Z(n10950) );
  XOR U12002 ( .A(n10953), .B(n10954), .Z(n10949) );
  ANDN U12003 ( .B(n10955), .A(n5999), .Z(n10953) );
  XNOR U12004 ( .A(n10956), .B(n10957), .Z(n5999) );
  IV U12005 ( .A(n10954), .Z(n10957) );
  XOR U12006 ( .A(n5998), .B(n10954), .Z(n10955) );
  XOR U12007 ( .A(n10958), .B(n10959), .Z(n10954) );
  ANDN U12008 ( .B(n10960), .A(n6004), .Z(n10958) );
  XNOR U12009 ( .A(n10961), .B(n10962), .Z(n6004) );
  IV U12010 ( .A(n10959), .Z(n10962) );
  XOR U12011 ( .A(n6003), .B(n10959), .Z(n10960) );
  XOR U12012 ( .A(n10963), .B(n10964), .Z(n10959) );
  ANDN U12013 ( .B(n10965), .A(n6009), .Z(n10963) );
  XNOR U12014 ( .A(n10966), .B(n10967), .Z(n6009) );
  IV U12015 ( .A(n10964), .Z(n10967) );
  XOR U12016 ( .A(n6008), .B(n10964), .Z(n10965) );
  XOR U12017 ( .A(n10968), .B(n10969), .Z(n10964) );
  ANDN U12018 ( .B(n10970), .A(n6014), .Z(n10968) );
  XNOR U12019 ( .A(n10971), .B(n10972), .Z(n6014) );
  IV U12020 ( .A(n10969), .Z(n10972) );
  XOR U12021 ( .A(n6013), .B(n10969), .Z(n10970) );
  XOR U12022 ( .A(n10973), .B(n10974), .Z(n10969) );
  ANDN U12023 ( .B(n10975), .A(n6019), .Z(n10973) );
  XNOR U12024 ( .A(n10976), .B(n10977), .Z(n6019) );
  IV U12025 ( .A(n10974), .Z(n10977) );
  XOR U12026 ( .A(n6018), .B(n10974), .Z(n10975) );
  XOR U12027 ( .A(n10978), .B(n10979), .Z(n10974) );
  ANDN U12028 ( .B(n10980), .A(n6024), .Z(n10978) );
  XNOR U12029 ( .A(n10981), .B(n10982), .Z(n6024) );
  IV U12030 ( .A(n10979), .Z(n10982) );
  XOR U12031 ( .A(n6023), .B(n10979), .Z(n10980) );
  XOR U12032 ( .A(n10983), .B(n10984), .Z(n10979) );
  ANDN U12033 ( .B(n10985), .A(n6029), .Z(n10983) );
  XNOR U12034 ( .A(n10986), .B(n10987), .Z(n6029) );
  IV U12035 ( .A(n10984), .Z(n10987) );
  XOR U12036 ( .A(n6028), .B(n10984), .Z(n10985) );
  XOR U12037 ( .A(n10988), .B(n10989), .Z(n10984) );
  ANDN U12038 ( .B(n10990), .A(n6034), .Z(n10988) );
  XNOR U12039 ( .A(n10991), .B(n10992), .Z(n6034) );
  IV U12040 ( .A(n10989), .Z(n10992) );
  XOR U12041 ( .A(n6033), .B(n10989), .Z(n10990) );
  XOR U12042 ( .A(n10993), .B(n10994), .Z(n10989) );
  ANDN U12043 ( .B(n10995), .A(n6044), .Z(n10993) );
  XNOR U12044 ( .A(n10996), .B(n10997), .Z(n6044) );
  IV U12045 ( .A(n10994), .Z(n10997) );
  XOR U12046 ( .A(n6043), .B(n10994), .Z(n10995) );
  XOR U12047 ( .A(n10998), .B(n10999), .Z(n10994) );
  ANDN U12048 ( .B(n11000), .A(n6049), .Z(n10998) );
  XNOR U12049 ( .A(n11001), .B(n11002), .Z(n6049) );
  IV U12050 ( .A(n10999), .Z(n11002) );
  XOR U12051 ( .A(n6048), .B(n10999), .Z(n11000) );
  XOR U12052 ( .A(n11003), .B(n11004), .Z(n10999) );
  ANDN U12053 ( .B(n11005), .A(n6054), .Z(n11003) );
  XNOR U12054 ( .A(n11006), .B(n11007), .Z(n6054) );
  IV U12055 ( .A(n11004), .Z(n11007) );
  XOR U12056 ( .A(n6053), .B(n11004), .Z(n11005) );
  XOR U12057 ( .A(n11008), .B(n11009), .Z(n11004) );
  ANDN U12058 ( .B(n11010), .A(n6059), .Z(n11008) );
  XNOR U12059 ( .A(n11011), .B(n11012), .Z(n6059) );
  IV U12060 ( .A(n11009), .Z(n11012) );
  XOR U12061 ( .A(n6058), .B(n11009), .Z(n11010) );
  XOR U12062 ( .A(n11013), .B(n11014), .Z(n11009) );
  ANDN U12063 ( .B(n11015), .A(n6064), .Z(n11013) );
  XNOR U12064 ( .A(n11016), .B(n11017), .Z(n6064) );
  IV U12065 ( .A(n11014), .Z(n11017) );
  XOR U12066 ( .A(n6063), .B(n11014), .Z(n11015) );
  XOR U12067 ( .A(n11018), .B(n11019), .Z(n11014) );
  ANDN U12068 ( .B(n11020), .A(n6069), .Z(n11018) );
  XNOR U12069 ( .A(n11021), .B(n11022), .Z(n6069) );
  IV U12070 ( .A(n11019), .Z(n11022) );
  XOR U12071 ( .A(n6068), .B(n11019), .Z(n11020) );
  XOR U12072 ( .A(n11023), .B(n11024), .Z(n11019) );
  ANDN U12073 ( .B(n11025), .A(n6074), .Z(n11023) );
  XNOR U12074 ( .A(n11026), .B(n11027), .Z(n6074) );
  IV U12075 ( .A(n11024), .Z(n11027) );
  XOR U12076 ( .A(n6073), .B(n11024), .Z(n11025) );
  XOR U12077 ( .A(n11028), .B(n11029), .Z(n11024) );
  ANDN U12078 ( .B(n11030), .A(n6079), .Z(n11028) );
  XNOR U12079 ( .A(n11031), .B(n11032), .Z(n6079) );
  IV U12080 ( .A(n11029), .Z(n11032) );
  XOR U12081 ( .A(n6078), .B(n11029), .Z(n11030) );
  XOR U12082 ( .A(n11033), .B(n11034), .Z(n11029) );
  ANDN U12083 ( .B(n11035), .A(n6084), .Z(n11033) );
  XNOR U12084 ( .A(n11036), .B(n11037), .Z(n6084) );
  IV U12085 ( .A(n11034), .Z(n11037) );
  XOR U12086 ( .A(n6083), .B(n11034), .Z(n11035) );
  XOR U12087 ( .A(n11038), .B(n11039), .Z(n11034) );
  ANDN U12088 ( .B(n11040), .A(n6089), .Z(n11038) );
  XNOR U12089 ( .A(n11041), .B(n11042), .Z(n6089) );
  IV U12090 ( .A(n11039), .Z(n11042) );
  XOR U12091 ( .A(n6088), .B(n11039), .Z(n11040) );
  XOR U12092 ( .A(n11043), .B(n11044), .Z(n11039) );
  ANDN U12093 ( .B(n11045), .A(n6099), .Z(n11043) );
  XNOR U12094 ( .A(n11046), .B(n11047), .Z(n6099) );
  IV U12095 ( .A(n11044), .Z(n11047) );
  XOR U12096 ( .A(n6098), .B(n11044), .Z(n11045) );
  XOR U12097 ( .A(n11048), .B(n11049), .Z(n11044) );
  ANDN U12098 ( .B(n11050), .A(n6104), .Z(n11048) );
  XNOR U12099 ( .A(n11051), .B(n11052), .Z(n6104) );
  IV U12100 ( .A(n11049), .Z(n11052) );
  XOR U12101 ( .A(n6103), .B(n11049), .Z(n11050) );
  XOR U12102 ( .A(n11053), .B(n11054), .Z(n11049) );
  ANDN U12103 ( .B(n11055), .A(n6109), .Z(n11053) );
  XNOR U12104 ( .A(n11056), .B(n11057), .Z(n6109) );
  IV U12105 ( .A(n11054), .Z(n11057) );
  XOR U12106 ( .A(n6108), .B(n11054), .Z(n11055) );
  XOR U12107 ( .A(n11058), .B(n11059), .Z(n11054) );
  ANDN U12108 ( .B(n11060), .A(n6114), .Z(n11058) );
  XNOR U12109 ( .A(n11061), .B(n11062), .Z(n6114) );
  IV U12110 ( .A(n11059), .Z(n11062) );
  XOR U12111 ( .A(n6113), .B(n11059), .Z(n11060) );
  XOR U12112 ( .A(n11063), .B(n11064), .Z(n11059) );
  ANDN U12113 ( .B(n11065), .A(n6119), .Z(n11063) );
  XNOR U12114 ( .A(n11066), .B(n11067), .Z(n6119) );
  IV U12115 ( .A(n11064), .Z(n11067) );
  XOR U12116 ( .A(n6118), .B(n11064), .Z(n11065) );
  XOR U12117 ( .A(n11068), .B(n11069), .Z(n11064) );
  ANDN U12118 ( .B(n11070), .A(n6124), .Z(n11068) );
  XNOR U12119 ( .A(n11071), .B(n11072), .Z(n6124) );
  IV U12120 ( .A(n11069), .Z(n11072) );
  XOR U12121 ( .A(n6123), .B(n11069), .Z(n11070) );
  XOR U12122 ( .A(n11073), .B(n11074), .Z(n11069) );
  ANDN U12123 ( .B(n11075), .A(n6129), .Z(n11073) );
  XNOR U12124 ( .A(n11076), .B(n11077), .Z(n6129) );
  IV U12125 ( .A(n11074), .Z(n11077) );
  XOR U12126 ( .A(n6128), .B(n11074), .Z(n11075) );
  XOR U12127 ( .A(n11078), .B(n11079), .Z(n11074) );
  ANDN U12128 ( .B(n11080), .A(n6134), .Z(n11078) );
  XNOR U12129 ( .A(n11081), .B(n11082), .Z(n6134) );
  IV U12130 ( .A(n11079), .Z(n11082) );
  XOR U12131 ( .A(n6133), .B(n11079), .Z(n11080) );
  XOR U12132 ( .A(n11083), .B(n11084), .Z(n11079) );
  ANDN U12133 ( .B(n11085), .A(n6139), .Z(n11083) );
  XNOR U12134 ( .A(n11086), .B(n11087), .Z(n6139) );
  IV U12135 ( .A(n11084), .Z(n11087) );
  XOR U12136 ( .A(n6138), .B(n11084), .Z(n11085) );
  XOR U12137 ( .A(n11088), .B(n11089), .Z(n11084) );
  ANDN U12138 ( .B(n11090), .A(n6144), .Z(n11088) );
  XNOR U12139 ( .A(n11091), .B(n11092), .Z(n6144) );
  IV U12140 ( .A(n11089), .Z(n11092) );
  XOR U12141 ( .A(n6143), .B(n11089), .Z(n11090) );
  XOR U12142 ( .A(n11093), .B(n11094), .Z(n11089) );
  ANDN U12143 ( .B(n11095), .A(n6154), .Z(n11093) );
  XNOR U12144 ( .A(n11096), .B(n11097), .Z(n6154) );
  IV U12145 ( .A(n11094), .Z(n11097) );
  XOR U12146 ( .A(n6153), .B(n11094), .Z(n11095) );
  XOR U12147 ( .A(n11098), .B(n11099), .Z(n11094) );
  ANDN U12148 ( .B(n11100), .A(n6159), .Z(n11098) );
  XNOR U12149 ( .A(n11101), .B(n11102), .Z(n6159) );
  IV U12150 ( .A(n11099), .Z(n11102) );
  XOR U12151 ( .A(n6158), .B(n11099), .Z(n11100) );
  XOR U12152 ( .A(n11103), .B(n11104), .Z(n11099) );
  ANDN U12153 ( .B(n11105), .A(n6164), .Z(n11103) );
  XNOR U12154 ( .A(n11106), .B(n11107), .Z(n6164) );
  IV U12155 ( .A(n11104), .Z(n11107) );
  XOR U12156 ( .A(n6163), .B(n11104), .Z(n11105) );
  XOR U12157 ( .A(n11108), .B(n11109), .Z(n11104) );
  ANDN U12158 ( .B(n11110), .A(n6169), .Z(n11108) );
  XNOR U12159 ( .A(n11111), .B(n11112), .Z(n6169) );
  IV U12160 ( .A(n11109), .Z(n11112) );
  XOR U12161 ( .A(n6168), .B(n11109), .Z(n11110) );
  XOR U12162 ( .A(n11113), .B(n11114), .Z(n11109) );
  ANDN U12163 ( .B(n11115), .A(n6174), .Z(n11113) );
  XNOR U12164 ( .A(n11116), .B(n11117), .Z(n6174) );
  IV U12165 ( .A(n11114), .Z(n11117) );
  XOR U12166 ( .A(n6173), .B(n11114), .Z(n11115) );
  XOR U12167 ( .A(n11118), .B(n11119), .Z(n11114) );
  ANDN U12168 ( .B(n11120), .A(n6179), .Z(n11118) );
  XNOR U12169 ( .A(n11121), .B(n11122), .Z(n6179) );
  IV U12170 ( .A(n11119), .Z(n11122) );
  XOR U12171 ( .A(n6178), .B(n11119), .Z(n11120) );
  XOR U12172 ( .A(n11123), .B(n11124), .Z(n11119) );
  ANDN U12173 ( .B(n11125), .A(n6184), .Z(n11123) );
  XNOR U12174 ( .A(n11126), .B(n11127), .Z(n6184) );
  IV U12175 ( .A(n11124), .Z(n11127) );
  XOR U12176 ( .A(n6183), .B(n11124), .Z(n11125) );
  XOR U12177 ( .A(n11128), .B(n11129), .Z(n11124) );
  ANDN U12178 ( .B(n11130), .A(n6189), .Z(n11128) );
  XNOR U12179 ( .A(n11131), .B(n11132), .Z(n6189) );
  IV U12180 ( .A(n11129), .Z(n11132) );
  XOR U12181 ( .A(n6188), .B(n11129), .Z(n11130) );
  XOR U12182 ( .A(n11133), .B(n11134), .Z(n11129) );
  ANDN U12183 ( .B(n11135), .A(n6194), .Z(n11133) );
  XNOR U12184 ( .A(n11136), .B(n11137), .Z(n6194) );
  IV U12185 ( .A(n11134), .Z(n11137) );
  XOR U12186 ( .A(n6193), .B(n11134), .Z(n11135) );
  XOR U12187 ( .A(n11138), .B(n11139), .Z(n11134) );
  ANDN U12188 ( .B(n11140), .A(n6199), .Z(n11138) );
  XNOR U12189 ( .A(n11141), .B(n11142), .Z(n6199) );
  IV U12190 ( .A(n11139), .Z(n11142) );
  XOR U12191 ( .A(n6198), .B(n11139), .Z(n11140) );
  XOR U12192 ( .A(n11143), .B(n11144), .Z(n11139) );
  ANDN U12193 ( .B(n11145), .A(n6209), .Z(n11143) );
  XNOR U12194 ( .A(n11146), .B(n11147), .Z(n6209) );
  IV U12195 ( .A(n11144), .Z(n11147) );
  XOR U12196 ( .A(n6208), .B(n11144), .Z(n11145) );
  XOR U12197 ( .A(n11148), .B(n11149), .Z(n11144) );
  ANDN U12198 ( .B(n11150), .A(n6214), .Z(n11148) );
  XNOR U12199 ( .A(n11151), .B(n11152), .Z(n6214) );
  IV U12200 ( .A(n11149), .Z(n11152) );
  XOR U12201 ( .A(n6213), .B(n11149), .Z(n11150) );
  XOR U12202 ( .A(n11153), .B(n11154), .Z(n11149) );
  ANDN U12203 ( .B(n11155), .A(n6219), .Z(n11153) );
  XNOR U12204 ( .A(n11156), .B(n11157), .Z(n6219) );
  IV U12205 ( .A(n11154), .Z(n11157) );
  XOR U12206 ( .A(n6218), .B(n11154), .Z(n11155) );
  XOR U12207 ( .A(n11158), .B(n11159), .Z(n11154) );
  ANDN U12208 ( .B(n11160), .A(n6224), .Z(n11158) );
  XNOR U12209 ( .A(n11161), .B(n11162), .Z(n6224) );
  IV U12210 ( .A(n11159), .Z(n11162) );
  XOR U12211 ( .A(n6223), .B(n11159), .Z(n11160) );
  XOR U12212 ( .A(n11163), .B(n11164), .Z(n11159) );
  ANDN U12213 ( .B(n11165), .A(n6229), .Z(n11163) );
  XNOR U12214 ( .A(n11166), .B(n11167), .Z(n6229) );
  IV U12215 ( .A(n11164), .Z(n11167) );
  XOR U12216 ( .A(n6228), .B(n11164), .Z(n11165) );
  XOR U12217 ( .A(n11168), .B(n11169), .Z(n11164) );
  ANDN U12218 ( .B(n11170), .A(n6234), .Z(n11168) );
  XNOR U12219 ( .A(n11171), .B(n11172), .Z(n6234) );
  IV U12220 ( .A(n11169), .Z(n11172) );
  XOR U12221 ( .A(n6233), .B(n11169), .Z(n11170) );
  XOR U12222 ( .A(n11173), .B(n11174), .Z(n11169) );
  ANDN U12223 ( .B(n11175), .A(n6239), .Z(n11173) );
  XNOR U12224 ( .A(n11176), .B(n11177), .Z(n6239) );
  IV U12225 ( .A(n11174), .Z(n11177) );
  XOR U12226 ( .A(n6238), .B(n11174), .Z(n11175) );
  XOR U12227 ( .A(n11178), .B(n11179), .Z(n11174) );
  ANDN U12228 ( .B(n11180), .A(n6244), .Z(n11178) );
  XNOR U12229 ( .A(n11181), .B(n11182), .Z(n6244) );
  IV U12230 ( .A(n11179), .Z(n11182) );
  XOR U12231 ( .A(n6243), .B(n11179), .Z(n11180) );
  XOR U12232 ( .A(n11183), .B(n11184), .Z(n11179) );
  ANDN U12233 ( .B(n11185), .A(n6249), .Z(n11183) );
  XNOR U12234 ( .A(n11186), .B(n11187), .Z(n6249) );
  IV U12235 ( .A(n11184), .Z(n11187) );
  XOR U12236 ( .A(n6248), .B(n11184), .Z(n11185) );
  XOR U12237 ( .A(n11188), .B(n11189), .Z(n11184) );
  ANDN U12238 ( .B(n11190), .A(n6254), .Z(n11188) );
  XNOR U12239 ( .A(n11191), .B(n11192), .Z(n6254) );
  IV U12240 ( .A(n11189), .Z(n11192) );
  XOR U12241 ( .A(n6253), .B(n11189), .Z(n11190) );
  XOR U12242 ( .A(n11193), .B(n11194), .Z(n11189) );
  ANDN U12243 ( .B(n11195), .A(n6264), .Z(n11193) );
  XNOR U12244 ( .A(n11196), .B(n11197), .Z(n6264) );
  IV U12245 ( .A(n11194), .Z(n11197) );
  XOR U12246 ( .A(n6263), .B(n11194), .Z(n11195) );
  XOR U12247 ( .A(n11198), .B(n11199), .Z(n11194) );
  ANDN U12248 ( .B(n11200), .A(n6269), .Z(n11198) );
  XNOR U12249 ( .A(n11201), .B(n11202), .Z(n6269) );
  IV U12250 ( .A(n11199), .Z(n11202) );
  XOR U12251 ( .A(n6268), .B(n11199), .Z(n11200) );
  XOR U12252 ( .A(n11203), .B(n11204), .Z(n11199) );
  ANDN U12253 ( .B(n11205), .A(n6274), .Z(n11203) );
  XNOR U12254 ( .A(n11206), .B(n11207), .Z(n6274) );
  IV U12255 ( .A(n11204), .Z(n11207) );
  XOR U12256 ( .A(n6273), .B(n11204), .Z(n11205) );
  XOR U12257 ( .A(n11208), .B(n11209), .Z(n11204) );
  ANDN U12258 ( .B(n11210), .A(n6279), .Z(n11208) );
  XNOR U12259 ( .A(n11211), .B(n11212), .Z(n6279) );
  IV U12260 ( .A(n11209), .Z(n11212) );
  XOR U12261 ( .A(n6278), .B(n11209), .Z(n11210) );
  XOR U12262 ( .A(n11213), .B(n11214), .Z(n11209) );
  ANDN U12263 ( .B(n11215), .A(n6284), .Z(n11213) );
  XNOR U12264 ( .A(n11216), .B(n11217), .Z(n6284) );
  IV U12265 ( .A(n11214), .Z(n11217) );
  XOR U12266 ( .A(n6283), .B(n11214), .Z(n11215) );
  XOR U12267 ( .A(n11218), .B(n11219), .Z(n11214) );
  ANDN U12268 ( .B(n11220), .A(n6289), .Z(n11218) );
  XNOR U12269 ( .A(n11221), .B(n11222), .Z(n6289) );
  IV U12270 ( .A(n11219), .Z(n11222) );
  XOR U12271 ( .A(n6288), .B(n11219), .Z(n11220) );
  XOR U12272 ( .A(n11223), .B(n11224), .Z(n11219) );
  ANDN U12273 ( .B(n11225), .A(n6294), .Z(n11223) );
  XNOR U12274 ( .A(n11226), .B(n11227), .Z(n6294) );
  IV U12275 ( .A(n11224), .Z(n11227) );
  XOR U12276 ( .A(n6293), .B(n11224), .Z(n11225) );
  XOR U12277 ( .A(n11228), .B(n11229), .Z(n11224) );
  ANDN U12278 ( .B(n11230), .A(n6299), .Z(n11228) );
  XNOR U12279 ( .A(n11231), .B(n11232), .Z(n6299) );
  IV U12280 ( .A(n11229), .Z(n11232) );
  XOR U12281 ( .A(n6298), .B(n11229), .Z(n11230) );
  XOR U12282 ( .A(n11233), .B(n11234), .Z(n11229) );
  ANDN U12283 ( .B(n11235), .A(n6304), .Z(n11233) );
  XNOR U12284 ( .A(n11236), .B(n11237), .Z(n6304) );
  IV U12285 ( .A(n11234), .Z(n11237) );
  XOR U12286 ( .A(n6303), .B(n11234), .Z(n11235) );
  XOR U12287 ( .A(n11238), .B(n11239), .Z(n11234) );
  ANDN U12288 ( .B(n11240), .A(n6309), .Z(n11238) );
  XNOR U12289 ( .A(n11241), .B(n11242), .Z(n6309) );
  IV U12290 ( .A(n11239), .Z(n11242) );
  XOR U12291 ( .A(n6308), .B(n11239), .Z(n11240) );
  XOR U12292 ( .A(n11243), .B(n11244), .Z(n11239) );
  ANDN U12293 ( .B(n11245), .A(n6319), .Z(n11243) );
  XNOR U12294 ( .A(n11246), .B(n11247), .Z(n6319) );
  IV U12295 ( .A(n11244), .Z(n11247) );
  XOR U12296 ( .A(n6318), .B(n11244), .Z(n11245) );
  XOR U12297 ( .A(n11248), .B(n11249), .Z(n11244) );
  ANDN U12298 ( .B(n11250), .A(n6324), .Z(n11248) );
  XNOR U12299 ( .A(n11251), .B(n11252), .Z(n6324) );
  IV U12300 ( .A(n11249), .Z(n11252) );
  XOR U12301 ( .A(n6323), .B(n11249), .Z(n11250) );
  XOR U12302 ( .A(n11253), .B(n11254), .Z(n11249) );
  ANDN U12303 ( .B(n11255), .A(n6329), .Z(n11253) );
  XNOR U12304 ( .A(n11256), .B(n11257), .Z(n6329) );
  IV U12305 ( .A(n11254), .Z(n11257) );
  XOR U12306 ( .A(n6328), .B(n11254), .Z(n11255) );
  XOR U12307 ( .A(n11258), .B(n11259), .Z(n11254) );
  ANDN U12308 ( .B(n11260), .A(n6334), .Z(n11258) );
  XNOR U12309 ( .A(n11261), .B(n11262), .Z(n6334) );
  IV U12310 ( .A(n11259), .Z(n11262) );
  XOR U12311 ( .A(n6333), .B(n11259), .Z(n11260) );
  XOR U12312 ( .A(n11263), .B(n11264), .Z(n11259) );
  ANDN U12313 ( .B(n11265), .A(n6339), .Z(n11263) );
  XNOR U12314 ( .A(n11266), .B(n11267), .Z(n6339) );
  IV U12315 ( .A(n11264), .Z(n11267) );
  XOR U12316 ( .A(n6338), .B(n11264), .Z(n11265) );
  XOR U12317 ( .A(n11268), .B(n11269), .Z(n11264) );
  ANDN U12318 ( .B(n11270), .A(n6344), .Z(n11268) );
  XNOR U12319 ( .A(n11271), .B(n11272), .Z(n6344) );
  IV U12320 ( .A(n11269), .Z(n11272) );
  XOR U12321 ( .A(n6343), .B(n11269), .Z(n11270) );
  XOR U12322 ( .A(n11273), .B(n11274), .Z(n11269) );
  ANDN U12323 ( .B(n11275), .A(n6349), .Z(n11273) );
  XNOR U12324 ( .A(n11276), .B(n11277), .Z(n6349) );
  IV U12325 ( .A(n11274), .Z(n11277) );
  XOR U12326 ( .A(n6348), .B(n11274), .Z(n11275) );
  XOR U12327 ( .A(n11278), .B(n11279), .Z(n11274) );
  ANDN U12328 ( .B(n11280), .A(n6354), .Z(n11278) );
  XNOR U12329 ( .A(n11281), .B(n11282), .Z(n6354) );
  IV U12330 ( .A(n11279), .Z(n11282) );
  XOR U12331 ( .A(n6353), .B(n11279), .Z(n11280) );
  XOR U12332 ( .A(n11283), .B(n11284), .Z(n11279) );
  ANDN U12333 ( .B(n11285), .A(n6359), .Z(n11283) );
  XNOR U12334 ( .A(n11286), .B(n11287), .Z(n6359) );
  IV U12335 ( .A(n11284), .Z(n11287) );
  XOR U12336 ( .A(n6358), .B(n11284), .Z(n11285) );
  XOR U12337 ( .A(n11288), .B(n11289), .Z(n11284) );
  ANDN U12338 ( .B(n11290), .A(n6364), .Z(n11288) );
  XNOR U12339 ( .A(n11291), .B(n11292), .Z(n6364) );
  IV U12340 ( .A(n11289), .Z(n11292) );
  XOR U12341 ( .A(n6363), .B(n11289), .Z(n11290) );
  XOR U12342 ( .A(n11293), .B(n11294), .Z(n11289) );
  ANDN U12343 ( .B(n11295), .A(n6374), .Z(n11293) );
  XNOR U12344 ( .A(n11296), .B(n11297), .Z(n6374) );
  IV U12345 ( .A(n11294), .Z(n11297) );
  XOR U12346 ( .A(n6373), .B(n11294), .Z(n11295) );
  XOR U12347 ( .A(n11298), .B(n11299), .Z(n11294) );
  ANDN U12348 ( .B(n11300), .A(n6379), .Z(n11298) );
  XNOR U12349 ( .A(n11301), .B(n11302), .Z(n6379) );
  IV U12350 ( .A(n11299), .Z(n11302) );
  XOR U12351 ( .A(n6378), .B(n11299), .Z(n11300) );
  XOR U12352 ( .A(n11303), .B(n11304), .Z(n11299) );
  ANDN U12353 ( .B(n11305), .A(n6384), .Z(n11303) );
  XNOR U12354 ( .A(n11306), .B(n11307), .Z(n6384) );
  IV U12355 ( .A(n11304), .Z(n11307) );
  XOR U12356 ( .A(n6383), .B(n11304), .Z(n11305) );
  XOR U12357 ( .A(n11308), .B(n11309), .Z(n11304) );
  ANDN U12358 ( .B(n11310), .A(n6389), .Z(n11308) );
  XNOR U12359 ( .A(n11311), .B(n11312), .Z(n6389) );
  IV U12360 ( .A(n11309), .Z(n11312) );
  XOR U12361 ( .A(n6388), .B(n11309), .Z(n11310) );
  XOR U12362 ( .A(n11313), .B(n11314), .Z(n11309) );
  ANDN U12363 ( .B(n11315), .A(n6394), .Z(n11313) );
  XNOR U12364 ( .A(n11316), .B(n11317), .Z(n6394) );
  IV U12365 ( .A(n11314), .Z(n11317) );
  XOR U12366 ( .A(n6393), .B(n11314), .Z(n11315) );
  XOR U12367 ( .A(n11318), .B(n11319), .Z(n11314) );
  ANDN U12368 ( .B(n11320), .A(n6399), .Z(n11318) );
  XNOR U12369 ( .A(n11321), .B(n11322), .Z(n6399) );
  IV U12370 ( .A(n11319), .Z(n11322) );
  XOR U12371 ( .A(n6398), .B(n11319), .Z(n11320) );
  XOR U12372 ( .A(n11323), .B(n11324), .Z(n11319) );
  ANDN U12373 ( .B(n11325), .A(n6404), .Z(n11323) );
  XNOR U12374 ( .A(n11326), .B(n11327), .Z(n6404) );
  IV U12375 ( .A(n11324), .Z(n11327) );
  XOR U12376 ( .A(n6403), .B(n11324), .Z(n11325) );
  XOR U12377 ( .A(n11328), .B(n11329), .Z(n11324) );
  ANDN U12378 ( .B(n11330), .A(n6409), .Z(n11328) );
  XNOR U12379 ( .A(n11331), .B(n11332), .Z(n6409) );
  IV U12380 ( .A(n11329), .Z(n11332) );
  XOR U12381 ( .A(n6408), .B(n11329), .Z(n11330) );
  XOR U12382 ( .A(n11333), .B(n11334), .Z(n11329) );
  ANDN U12383 ( .B(n11335), .A(n6414), .Z(n11333) );
  XNOR U12384 ( .A(n11336), .B(n11337), .Z(n6414) );
  IV U12385 ( .A(n11334), .Z(n11337) );
  XOR U12386 ( .A(n6413), .B(n11334), .Z(n11335) );
  XOR U12387 ( .A(n11338), .B(n11339), .Z(n11334) );
  ANDN U12388 ( .B(n11340), .A(n6419), .Z(n11338) );
  XNOR U12389 ( .A(n11341), .B(n11342), .Z(n6419) );
  IV U12390 ( .A(n11339), .Z(n11342) );
  XOR U12391 ( .A(n6418), .B(n11339), .Z(n11340) );
  XOR U12392 ( .A(n11343), .B(n11344), .Z(n11339) );
  ANDN U12393 ( .B(n11345), .A(n6434), .Z(n11343) );
  XNOR U12394 ( .A(n11346), .B(n11347), .Z(n6434) );
  IV U12395 ( .A(n11344), .Z(n11347) );
  XOR U12396 ( .A(n6433), .B(n11344), .Z(n11345) );
  XOR U12397 ( .A(n11348), .B(n11349), .Z(n11344) );
  ANDN U12398 ( .B(n11350), .A(n6439), .Z(n11348) );
  XNOR U12399 ( .A(n11351), .B(n11352), .Z(n6439) );
  IV U12400 ( .A(n11349), .Z(n11352) );
  XOR U12401 ( .A(n6438), .B(n11349), .Z(n11350) );
  XOR U12402 ( .A(n11353), .B(n11354), .Z(n11349) );
  ANDN U12403 ( .B(n11355), .A(n6444), .Z(n11353) );
  XNOR U12404 ( .A(n11356), .B(n11357), .Z(n6444) );
  IV U12405 ( .A(n11354), .Z(n11357) );
  XOR U12406 ( .A(n6443), .B(n11354), .Z(n11355) );
  XOR U12407 ( .A(n11358), .B(n11359), .Z(n11354) );
  ANDN U12408 ( .B(n11360), .A(n6449), .Z(n11358) );
  XNOR U12409 ( .A(n11361), .B(n11362), .Z(n6449) );
  IV U12410 ( .A(n11359), .Z(n11362) );
  XOR U12411 ( .A(n6448), .B(n11359), .Z(n11360) );
  XOR U12412 ( .A(n11363), .B(n11364), .Z(n11359) );
  ANDN U12413 ( .B(n11365), .A(n6454), .Z(n11363) );
  XNOR U12414 ( .A(n11366), .B(n11367), .Z(n6454) );
  IV U12415 ( .A(n11364), .Z(n11367) );
  XOR U12416 ( .A(n6453), .B(n11364), .Z(n11365) );
  XOR U12417 ( .A(n11368), .B(n11369), .Z(n11364) );
  ANDN U12418 ( .B(n11370), .A(n6459), .Z(n11368) );
  XNOR U12419 ( .A(n11371), .B(n11372), .Z(n6459) );
  IV U12420 ( .A(n11369), .Z(n11372) );
  XOR U12421 ( .A(n6458), .B(n11369), .Z(n11370) );
  XOR U12422 ( .A(n11373), .B(n11374), .Z(n11369) );
  ANDN U12423 ( .B(n11375), .A(n6464), .Z(n11373) );
  XNOR U12424 ( .A(n11376), .B(n11377), .Z(n6464) );
  IV U12425 ( .A(n11374), .Z(n11377) );
  XOR U12426 ( .A(n6463), .B(n11374), .Z(n11375) );
  XOR U12427 ( .A(n11378), .B(n11379), .Z(n11374) );
  ANDN U12428 ( .B(n11380), .A(n6469), .Z(n11378) );
  XNOR U12429 ( .A(n11381), .B(n11382), .Z(n6469) );
  IV U12430 ( .A(n11379), .Z(n11382) );
  XOR U12431 ( .A(n6468), .B(n11379), .Z(n11380) );
  XOR U12432 ( .A(n11383), .B(n11384), .Z(n11379) );
  ANDN U12433 ( .B(n11385), .A(n6474), .Z(n11383) );
  XNOR U12434 ( .A(n11386), .B(n11387), .Z(n6474) );
  IV U12435 ( .A(n11384), .Z(n11387) );
  XOR U12436 ( .A(n6473), .B(n11384), .Z(n11385) );
  XOR U12437 ( .A(n11388), .B(n11389), .Z(n11384) );
  ANDN U12438 ( .B(n11390), .A(n6479), .Z(n11388) );
  XNOR U12439 ( .A(n11391), .B(n11392), .Z(n6479) );
  IV U12440 ( .A(n11389), .Z(n11392) );
  XOR U12441 ( .A(n6478), .B(n11389), .Z(n11390) );
  XOR U12442 ( .A(n11393), .B(n11394), .Z(n11389) );
  ANDN U12443 ( .B(n11395), .A(n6489), .Z(n11393) );
  XNOR U12444 ( .A(n11396), .B(n11397), .Z(n6489) );
  IV U12445 ( .A(n11394), .Z(n11397) );
  XOR U12446 ( .A(n6488), .B(n11394), .Z(n11395) );
  XOR U12447 ( .A(n11398), .B(n11399), .Z(n11394) );
  ANDN U12448 ( .B(n11400), .A(n6494), .Z(n11398) );
  XNOR U12449 ( .A(n11401), .B(n11402), .Z(n6494) );
  IV U12450 ( .A(n11399), .Z(n11402) );
  XOR U12451 ( .A(n6493), .B(n11399), .Z(n11400) );
  XOR U12452 ( .A(n11403), .B(n11404), .Z(n11399) );
  ANDN U12453 ( .B(n11405), .A(n6499), .Z(n11403) );
  XNOR U12454 ( .A(n11406), .B(n11407), .Z(n6499) );
  IV U12455 ( .A(n11404), .Z(n11407) );
  XOR U12456 ( .A(n6498), .B(n11404), .Z(n11405) );
  XOR U12457 ( .A(n11408), .B(n11409), .Z(n11404) );
  ANDN U12458 ( .B(n11410), .A(n6504), .Z(n11408) );
  XNOR U12459 ( .A(n11411), .B(n11412), .Z(n6504) );
  IV U12460 ( .A(n11409), .Z(n11412) );
  XOR U12461 ( .A(n6503), .B(n11409), .Z(n11410) );
  XOR U12462 ( .A(n11413), .B(n11414), .Z(n11409) );
  ANDN U12463 ( .B(n11415), .A(n6509), .Z(n11413) );
  XNOR U12464 ( .A(n11416), .B(n11417), .Z(n6509) );
  IV U12465 ( .A(n11414), .Z(n11417) );
  XOR U12466 ( .A(n6508), .B(n11414), .Z(n11415) );
  XOR U12467 ( .A(n11418), .B(n11419), .Z(n11414) );
  ANDN U12468 ( .B(n11420), .A(n6514), .Z(n11418) );
  XNOR U12469 ( .A(n11421), .B(n11422), .Z(n6514) );
  IV U12470 ( .A(n11419), .Z(n11422) );
  XOR U12471 ( .A(n6513), .B(n11419), .Z(n11420) );
  XOR U12472 ( .A(n11423), .B(n11424), .Z(n11419) );
  ANDN U12473 ( .B(n11425), .A(n6519), .Z(n11423) );
  XNOR U12474 ( .A(n11426), .B(n11427), .Z(n6519) );
  IV U12475 ( .A(n11424), .Z(n11427) );
  XOR U12476 ( .A(n6518), .B(n11424), .Z(n11425) );
  XOR U12477 ( .A(n11428), .B(n11429), .Z(n11424) );
  ANDN U12478 ( .B(n11430), .A(n6524), .Z(n11428) );
  XNOR U12479 ( .A(n11431), .B(n11432), .Z(n6524) );
  IV U12480 ( .A(n11429), .Z(n11432) );
  XOR U12481 ( .A(n6523), .B(n11429), .Z(n11430) );
  XOR U12482 ( .A(n11433), .B(n11434), .Z(n11429) );
  ANDN U12483 ( .B(n11435), .A(n6529), .Z(n11433) );
  XNOR U12484 ( .A(n11436), .B(n11437), .Z(n6529) );
  IV U12485 ( .A(n11434), .Z(n11437) );
  XOR U12486 ( .A(n6528), .B(n11434), .Z(n11435) );
  XOR U12487 ( .A(n11438), .B(n11439), .Z(n11434) );
  ANDN U12488 ( .B(n11440), .A(n6534), .Z(n11438) );
  XNOR U12489 ( .A(n11441), .B(n11442), .Z(n6534) );
  IV U12490 ( .A(n11439), .Z(n11442) );
  XOR U12491 ( .A(n6533), .B(n11439), .Z(n11440) );
  XOR U12492 ( .A(n11443), .B(n11444), .Z(n11439) );
  ANDN U12493 ( .B(n11445), .A(n6544), .Z(n11443) );
  XNOR U12494 ( .A(n11446), .B(n11447), .Z(n6544) );
  IV U12495 ( .A(n11444), .Z(n11447) );
  XOR U12496 ( .A(n6543), .B(n11444), .Z(n11445) );
  XOR U12497 ( .A(n11448), .B(n11449), .Z(n11444) );
  ANDN U12498 ( .B(n11450), .A(n6549), .Z(n11448) );
  XNOR U12499 ( .A(n11451), .B(n11452), .Z(n6549) );
  IV U12500 ( .A(n11449), .Z(n11452) );
  XOR U12501 ( .A(n6548), .B(n11449), .Z(n11450) );
  XOR U12502 ( .A(n11453), .B(n11454), .Z(n11449) );
  ANDN U12503 ( .B(n11455), .A(n6554), .Z(n11453) );
  XNOR U12504 ( .A(n11456), .B(n11457), .Z(n6554) );
  IV U12505 ( .A(n11454), .Z(n11457) );
  XOR U12506 ( .A(n6553), .B(n11454), .Z(n11455) );
  XOR U12507 ( .A(n11458), .B(n11459), .Z(n11454) );
  ANDN U12508 ( .B(n11460), .A(n6559), .Z(n11458) );
  XNOR U12509 ( .A(n11461), .B(n11462), .Z(n6559) );
  IV U12510 ( .A(n11459), .Z(n11462) );
  XOR U12511 ( .A(n6558), .B(n11459), .Z(n11460) );
  XOR U12512 ( .A(n11463), .B(n11464), .Z(n11459) );
  ANDN U12513 ( .B(n11465), .A(n6564), .Z(n11463) );
  XNOR U12514 ( .A(n11466), .B(n11467), .Z(n6564) );
  IV U12515 ( .A(n11464), .Z(n11467) );
  XOR U12516 ( .A(n6563), .B(n11464), .Z(n11465) );
  XOR U12517 ( .A(n11468), .B(n11469), .Z(n11464) );
  ANDN U12518 ( .B(n11470), .A(n6569), .Z(n11468) );
  XNOR U12519 ( .A(n11471), .B(n11472), .Z(n6569) );
  IV U12520 ( .A(n11469), .Z(n11472) );
  XOR U12521 ( .A(n6568), .B(n11469), .Z(n11470) );
  XOR U12522 ( .A(n11473), .B(n11474), .Z(n11469) );
  ANDN U12523 ( .B(n11475), .A(n6574), .Z(n11473) );
  XNOR U12524 ( .A(n11476), .B(n11477), .Z(n6574) );
  IV U12525 ( .A(n11474), .Z(n11477) );
  XOR U12526 ( .A(n6573), .B(n11474), .Z(n11475) );
  XOR U12527 ( .A(n11478), .B(n11479), .Z(n11474) );
  ANDN U12528 ( .B(n11480), .A(n6579), .Z(n11478) );
  XNOR U12529 ( .A(n11481), .B(n11482), .Z(n6579) );
  IV U12530 ( .A(n11479), .Z(n11482) );
  XOR U12531 ( .A(n6578), .B(n11479), .Z(n11480) );
  XOR U12532 ( .A(n11483), .B(n11484), .Z(n11479) );
  ANDN U12533 ( .B(n11485), .A(n6584), .Z(n11483) );
  XNOR U12534 ( .A(n11486), .B(n11487), .Z(n6584) );
  IV U12535 ( .A(n11484), .Z(n11487) );
  XOR U12536 ( .A(n6583), .B(n11484), .Z(n11485) );
  XOR U12537 ( .A(n11488), .B(n11489), .Z(n11484) );
  ANDN U12538 ( .B(n11490), .A(n6589), .Z(n11488) );
  XNOR U12539 ( .A(n11491), .B(n11492), .Z(n6589) );
  IV U12540 ( .A(n11489), .Z(n11492) );
  XOR U12541 ( .A(n6588), .B(n11489), .Z(n11490) );
  XOR U12542 ( .A(n11493), .B(n11494), .Z(n11489) );
  ANDN U12543 ( .B(n11495), .A(n6599), .Z(n11493) );
  XNOR U12544 ( .A(n11496), .B(n11497), .Z(n6599) );
  IV U12545 ( .A(n11494), .Z(n11497) );
  XOR U12546 ( .A(n6598), .B(n11494), .Z(n11495) );
  XOR U12547 ( .A(n11498), .B(n11499), .Z(n11494) );
  ANDN U12548 ( .B(n11500), .A(n6604), .Z(n11498) );
  XNOR U12549 ( .A(n11501), .B(n11502), .Z(n6604) );
  IV U12550 ( .A(n11499), .Z(n11502) );
  XOR U12551 ( .A(n6603), .B(n11499), .Z(n11500) );
  XOR U12552 ( .A(n11503), .B(n11504), .Z(n11499) );
  ANDN U12553 ( .B(n11505), .A(n6609), .Z(n11503) );
  XNOR U12554 ( .A(n11506), .B(n11507), .Z(n6609) );
  IV U12555 ( .A(n11504), .Z(n11507) );
  XOR U12556 ( .A(n6608), .B(n11504), .Z(n11505) );
  XOR U12557 ( .A(n11508), .B(n11509), .Z(n11504) );
  ANDN U12558 ( .B(n11510), .A(n6614), .Z(n11508) );
  XNOR U12559 ( .A(n11511), .B(n11512), .Z(n6614) );
  IV U12560 ( .A(n11509), .Z(n11512) );
  XOR U12561 ( .A(n6613), .B(n11509), .Z(n11510) );
  XOR U12562 ( .A(n11513), .B(n11514), .Z(n11509) );
  ANDN U12563 ( .B(n11515), .A(n6619), .Z(n11513) );
  XNOR U12564 ( .A(n11516), .B(n11517), .Z(n6619) );
  IV U12565 ( .A(n11514), .Z(n11517) );
  XOR U12566 ( .A(n6618), .B(n11514), .Z(n11515) );
  XOR U12567 ( .A(n11518), .B(n11519), .Z(n11514) );
  ANDN U12568 ( .B(n11520), .A(n6624), .Z(n11518) );
  XNOR U12569 ( .A(n11521), .B(n11522), .Z(n6624) );
  IV U12570 ( .A(n11519), .Z(n11522) );
  XOR U12571 ( .A(n6623), .B(n11519), .Z(n11520) );
  XOR U12572 ( .A(n11523), .B(n11524), .Z(n11519) );
  ANDN U12573 ( .B(n11525), .A(n6629), .Z(n11523) );
  XNOR U12574 ( .A(n11526), .B(n11527), .Z(n6629) );
  IV U12575 ( .A(n11524), .Z(n11527) );
  XOR U12576 ( .A(n6628), .B(n11524), .Z(n11525) );
  XOR U12577 ( .A(n11528), .B(n11529), .Z(n11524) );
  ANDN U12578 ( .B(n11530), .A(n6634), .Z(n11528) );
  XNOR U12579 ( .A(n11531), .B(n11532), .Z(n6634) );
  IV U12580 ( .A(n11529), .Z(n11532) );
  XOR U12581 ( .A(n6633), .B(n11529), .Z(n11530) );
  XOR U12582 ( .A(n11533), .B(n11534), .Z(n11529) );
  ANDN U12583 ( .B(n11535), .A(n6639), .Z(n11533) );
  XNOR U12584 ( .A(n11536), .B(n11537), .Z(n6639) );
  IV U12585 ( .A(n11534), .Z(n11537) );
  XOR U12586 ( .A(n6638), .B(n11534), .Z(n11535) );
  XOR U12587 ( .A(n11538), .B(n11539), .Z(n11534) );
  ANDN U12588 ( .B(n11540), .A(n6644), .Z(n11538) );
  XNOR U12589 ( .A(n11541), .B(n11542), .Z(n6644) );
  IV U12590 ( .A(n11539), .Z(n11542) );
  XOR U12591 ( .A(n6643), .B(n11539), .Z(n11540) );
  XOR U12592 ( .A(n11543), .B(n11544), .Z(n11539) );
  ANDN U12593 ( .B(n11545), .A(n6654), .Z(n11543) );
  XNOR U12594 ( .A(n11546), .B(n11547), .Z(n6654) );
  IV U12595 ( .A(n11544), .Z(n11547) );
  XOR U12596 ( .A(n6653), .B(n11544), .Z(n11545) );
  XOR U12597 ( .A(n11548), .B(n11549), .Z(n11544) );
  ANDN U12598 ( .B(n11550), .A(n6659), .Z(n11548) );
  XNOR U12599 ( .A(n11551), .B(n11552), .Z(n6659) );
  IV U12600 ( .A(n11549), .Z(n11552) );
  XOR U12601 ( .A(n6658), .B(n11549), .Z(n11550) );
  XOR U12602 ( .A(n11553), .B(n11554), .Z(n11549) );
  ANDN U12603 ( .B(n11555), .A(n6664), .Z(n11553) );
  XNOR U12604 ( .A(n11556), .B(n11557), .Z(n6664) );
  IV U12605 ( .A(n11554), .Z(n11557) );
  XOR U12606 ( .A(n6663), .B(n11554), .Z(n11555) );
  XOR U12607 ( .A(n11558), .B(n11559), .Z(n11554) );
  ANDN U12608 ( .B(n11560), .A(n6669), .Z(n11558) );
  XNOR U12609 ( .A(n11561), .B(n11562), .Z(n6669) );
  IV U12610 ( .A(n11559), .Z(n11562) );
  XOR U12611 ( .A(n6668), .B(n11559), .Z(n11560) );
  XOR U12612 ( .A(n11563), .B(n11564), .Z(n11559) );
  ANDN U12613 ( .B(n11565), .A(n6674), .Z(n11563) );
  XNOR U12614 ( .A(n11566), .B(n11567), .Z(n6674) );
  IV U12615 ( .A(n11564), .Z(n11567) );
  XOR U12616 ( .A(n6673), .B(n11564), .Z(n11565) );
  XOR U12617 ( .A(n11568), .B(n11569), .Z(n11564) );
  ANDN U12618 ( .B(n11570), .A(n6679), .Z(n11568) );
  XNOR U12619 ( .A(n11571), .B(n11572), .Z(n6679) );
  IV U12620 ( .A(n11569), .Z(n11572) );
  XOR U12621 ( .A(n6678), .B(n11569), .Z(n11570) );
  XOR U12622 ( .A(n11573), .B(n11574), .Z(n11569) );
  ANDN U12623 ( .B(n11575), .A(n6684), .Z(n11573) );
  XNOR U12624 ( .A(n11576), .B(n11577), .Z(n6684) );
  IV U12625 ( .A(n11574), .Z(n11577) );
  XOR U12626 ( .A(n6683), .B(n11574), .Z(n11575) );
  XOR U12627 ( .A(n11578), .B(n11579), .Z(n11574) );
  ANDN U12628 ( .B(n11580), .A(n6689), .Z(n11578) );
  XNOR U12629 ( .A(n11581), .B(n11582), .Z(n6689) );
  IV U12630 ( .A(n11579), .Z(n11582) );
  XOR U12631 ( .A(n6688), .B(n11579), .Z(n11580) );
  XOR U12632 ( .A(n11583), .B(n11584), .Z(n11579) );
  ANDN U12633 ( .B(n11585), .A(n6694), .Z(n11583) );
  XNOR U12634 ( .A(n11586), .B(n11587), .Z(n6694) );
  IV U12635 ( .A(n11584), .Z(n11587) );
  XOR U12636 ( .A(n6693), .B(n11584), .Z(n11585) );
  XOR U12637 ( .A(n11588), .B(n11589), .Z(n11584) );
  ANDN U12638 ( .B(n11590), .A(n6699), .Z(n11588) );
  XNOR U12639 ( .A(n11591), .B(n11592), .Z(n6699) );
  IV U12640 ( .A(n11589), .Z(n11592) );
  XOR U12641 ( .A(n6698), .B(n11589), .Z(n11590) );
  XOR U12642 ( .A(n11593), .B(n11594), .Z(n11589) );
  ANDN U12643 ( .B(n11595), .A(n6709), .Z(n11593) );
  XNOR U12644 ( .A(n11596), .B(n11597), .Z(n6709) );
  IV U12645 ( .A(n11594), .Z(n11597) );
  XOR U12646 ( .A(n6708), .B(n11594), .Z(n11595) );
  XOR U12647 ( .A(n11598), .B(n11599), .Z(n11594) );
  ANDN U12648 ( .B(n11600), .A(n6714), .Z(n11598) );
  XNOR U12649 ( .A(n11601), .B(n11602), .Z(n6714) );
  IV U12650 ( .A(n11599), .Z(n11602) );
  XOR U12651 ( .A(n6713), .B(n11599), .Z(n11600) );
  XOR U12652 ( .A(n11603), .B(n11604), .Z(n11599) );
  ANDN U12653 ( .B(n11605), .A(n6719), .Z(n11603) );
  XNOR U12654 ( .A(n11606), .B(n11607), .Z(n6719) );
  IV U12655 ( .A(n11604), .Z(n11607) );
  XOR U12656 ( .A(n6718), .B(n11604), .Z(n11605) );
  XOR U12657 ( .A(n11608), .B(n11609), .Z(n11604) );
  ANDN U12658 ( .B(n11610), .A(n6724), .Z(n11608) );
  XNOR U12659 ( .A(n11611), .B(n11612), .Z(n6724) );
  IV U12660 ( .A(n11609), .Z(n11612) );
  XOR U12661 ( .A(n6723), .B(n11609), .Z(n11610) );
  XOR U12662 ( .A(n11613), .B(n11614), .Z(n11609) );
  ANDN U12663 ( .B(n11615), .A(n6729), .Z(n11613) );
  XNOR U12664 ( .A(n11616), .B(n11617), .Z(n6729) );
  IV U12665 ( .A(n11614), .Z(n11617) );
  XOR U12666 ( .A(n6728), .B(n11614), .Z(n11615) );
  XOR U12667 ( .A(n11618), .B(n11619), .Z(n11614) );
  ANDN U12668 ( .B(n11620), .A(n6734), .Z(n11618) );
  XNOR U12669 ( .A(n11621), .B(n11622), .Z(n6734) );
  IV U12670 ( .A(n11619), .Z(n11622) );
  XOR U12671 ( .A(n6733), .B(n11619), .Z(n11620) );
  XOR U12672 ( .A(n11623), .B(n11624), .Z(n11619) );
  ANDN U12673 ( .B(n11625), .A(n6739), .Z(n11623) );
  XNOR U12674 ( .A(n11626), .B(n11627), .Z(n6739) );
  IV U12675 ( .A(n11624), .Z(n11627) );
  XOR U12676 ( .A(n6738), .B(n11624), .Z(n11625) );
  XOR U12677 ( .A(n11628), .B(n11629), .Z(n11624) );
  ANDN U12678 ( .B(n11630), .A(n6744), .Z(n11628) );
  XNOR U12679 ( .A(n11631), .B(n11632), .Z(n6744) );
  IV U12680 ( .A(n11629), .Z(n11632) );
  XOR U12681 ( .A(n6743), .B(n11629), .Z(n11630) );
  XOR U12682 ( .A(n11633), .B(n11634), .Z(n11629) );
  ANDN U12683 ( .B(n11635), .A(n6749), .Z(n11633) );
  XNOR U12684 ( .A(n11636), .B(n11637), .Z(n6749) );
  IV U12685 ( .A(n11634), .Z(n11637) );
  XOR U12686 ( .A(n6748), .B(n11634), .Z(n11635) );
  XOR U12687 ( .A(n11638), .B(n11639), .Z(n11634) );
  ANDN U12688 ( .B(n11640), .A(n6754), .Z(n11638) );
  XNOR U12689 ( .A(n11641), .B(n11642), .Z(n6754) );
  IV U12690 ( .A(n11639), .Z(n11642) );
  XOR U12691 ( .A(n6753), .B(n11639), .Z(n11640) );
  XOR U12692 ( .A(n11643), .B(n11644), .Z(n11639) );
  ANDN U12693 ( .B(n11645), .A(n6764), .Z(n11643) );
  XNOR U12694 ( .A(n11646), .B(n11647), .Z(n6764) );
  IV U12695 ( .A(n11644), .Z(n11647) );
  XOR U12696 ( .A(n6763), .B(n11644), .Z(n11645) );
  XOR U12697 ( .A(n11648), .B(n11649), .Z(n11644) );
  ANDN U12698 ( .B(n11650), .A(n6769), .Z(n11648) );
  XNOR U12699 ( .A(n11651), .B(n11652), .Z(n6769) );
  IV U12700 ( .A(n11649), .Z(n11652) );
  XOR U12701 ( .A(n6768), .B(n11649), .Z(n11650) );
  XOR U12702 ( .A(n11653), .B(n11654), .Z(n11649) );
  ANDN U12703 ( .B(n11655), .A(n6774), .Z(n11653) );
  XNOR U12704 ( .A(n11656), .B(n11657), .Z(n6774) );
  IV U12705 ( .A(n11654), .Z(n11657) );
  XOR U12706 ( .A(n6773), .B(n11654), .Z(n11655) );
  XOR U12707 ( .A(n11658), .B(n11659), .Z(n11654) );
  ANDN U12708 ( .B(n11660), .A(n6779), .Z(n11658) );
  XNOR U12709 ( .A(n11661), .B(n11662), .Z(n6779) );
  IV U12710 ( .A(n11659), .Z(n11662) );
  XOR U12711 ( .A(n6778), .B(n11659), .Z(n11660) );
  XOR U12712 ( .A(n11663), .B(n11664), .Z(n11659) );
  ANDN U12713 ( .B(n11665), .A(n6784), .Z(n11663) );
  XNOR U12714 ( .A(n11666), .B(n11667), .Z(n6784) );
  IV U12715 ( .A(n11664), .Z(n11667) );
  XOR U12716 ( .A(n6783), .B(n11664), .Z(n11665) );
  XOR U12717 ( .A(n11668), .B(n11669), .Z(n11664) );
  ANDN U12718 ( .B(n11670), .A(n6789), .Z(n11668) );
  XNOR U12719 ( .A(n11671), .B(n11672), .Z(n6789) );
  IV U12720 ( .A(n11669), .Z(n11672) );
  XOR U12721 ( .A(n6788), .B(n11669), .Z(n11670) );
  XOR U12722 ( .A(n11673), .B(n11674), .Z(n11669) );
  ANDN U12723 ( .B(n11675), .A(n6794), .Z(n11673) );
  XNOR U12724 ( .A(n11676), .B(n11677), .Z(n6794) );
  IV U12725 ( .A(n11674), .Z(n11677) );
  XOR U12726 ( .A(n6793), .B(n11674), .Z(n11675) );
  XOR U12727 ( .A(n11678), .B(n11679), .Z(n11674) );
  ANDN U12728 ( .B(n11680), .A(n6799), .Z(n11678) );
  XNOR U12729 ( .A(n11681), .B(n11682), .Z(n6799) );
  IV U12730 ( .A(n11679), .Z(n11682) );
  XOR U12731 ( .A(n6798), .B(n11679), .Z(n11680) );
  XOR U12732 ( .A(n11683), .B(n11684), .Z(n11679) );
  ANDN U12733 ( .B(n11685), .A(n6804), .Z(n11683) );
  XNOR U12734 ( .A(n11686), .B(n11687), .Z(n6804) );
  IV U12735 ( .A(n11684), .Z(n11687) );
  XOR U12736 ( .A(n6803), .B(n11684), .Z(n11685) );
  XOR U12737 ( .A(n11688), .B(n11689), .Z(n11684) );
  ANDN U12738 ( .B(n11690), .A(n6809), .Z(n11688) );
  XNOR U12739 ( .A(n11691), .B(n11692), .Z(n6809) );
  IV U12740 ( .A(n11689), .Z(n11692) );
  XOR U12741 ( .A(n6808), .B(n11689), .Z(n11690) );
  XOR U12742 ( .A(n11693), .B(n11694), .Z(n11689) );
  ANDN U12743 ( .B(n11695), .A(n6819), .Z(n11693) );
  XNOR U12744 ( .A(n11696), .B(n11697), .Z(n6819) );
  IV U12745 ( .A(n11694), .Z(n11697) );
  XOR U12746 ( .A(n6818), .B(n11694), .Z(n11695) );
  XOR U12747 ( .A(n11698), .B(n11699), .Z(n11694) );
  ANDN U12748 ( .B(n11700), .A(n6824), .Z(n11698) );
  XNOR U12749 ( .A(n11701), .B(n11702), .Z(n6824) );
  IV U12750 ( .A(n11699), .Z(n11702) );
  XOR U12751 ( .A(n6823), .B(n11699), .Z(n11700) );
  XOR U12752 ( .A(n11703), .B(n11704), .Z(n11699) );
  ANDN U12753 ( .B(n11705), .A(n6829), .Z(n11703) );
  XNOR U12754 ( .A(n11706), .B(n11707), .Z(n6829) );
  IV U12755 ( .A(n11704), .Z(n11707) );
  XOR U12756 ( .A(n6828), .B(n11704), .Z(n11705) );
  XOR U12757 ( .A(n11708), .B(n11709), .Z(n11704) );
  ANDN U12758 ( .B(n11710), .A(n6834), .Z(n11708) );
  XNOR U12759 ( .A(n11711), .B(n11712), .Z(n6834) );
  IV U12760 ( .A(n11709), .Z(n11712) );
  XOR U12761 ( .A(n6833), .B(n11709), .Z(n11710) );
  XOR U12762 ( .A(n11713), .B(n11714), .Z(n11709) );
  ANDN U12763 ( .B(n11715), .A(n6839), .Z(n11713) );
  XNOR U12764 ( .A(n11716), .B(n11717), .Z(n6839) );
  IV U12765 ( .A(n11714), .Z(n11717) );
  XOR U12766 ( .A(n6838), .B(n11714), .Z(n11715) );
  XOR U12767 ( .A(n11718), .B(n11719), .Z(n11714) );
  ANDN U12768 ( .B(n11720), .A(n6844), .Z(n11718) );
  XNOR U12769 ( .A(n11721), .B(n11722), .Z(n6844) );
  IV U12770 ( .A(n11719), .Z(n11722) );
  XOR U12771 ( .A(n6843), .B(n11719), .Z(n11720) );
  XOR U12772 ( .A(n11723), .B(n11724), .Z(n11719) );
  ANDN U12773 ( .B(n11725), .A(n6849), .Z(n11723) );
  XNOR U12774 ( .A(n11726), .B(n11727), .Z(n6849) );
  IV U12775 ( .A(n11724), .Z(n11727) );
  XOR U12776 ( .A(n6848), .B(n11724), .Z(n11725) );
  XOR U12777 ( .A(n11728), .B(n11729), .Z(n11724) );
  ANDN U12778 ( .B(n11730), .A(n6854), .Z(n11728) );
  XNOR U12779 ( .A(n11731), .B(n11732), .Z(n6854) );
  IV U12780 ( .A(n11729), .Z(n11732) );
  XOR U12781 ( .A(n6853), .B(n11729), .Z(n11730) );
  XOR U12782 ( .A(n11733), .B(n11734), .Z(n11729) );
  ANDN U12783 ( .B(n11735), .A(n6859), .Z(n11733) );
  XNOR U12784 ( .A(n11736), .B(n11737), .Z(n6859) );
  IV U12785 ( .A(n11734), .Z(n11737) );
  XOR U12786 ( .A(n6858), .B(n11734), .Z(n11735) );
  XOR U12787 ( .A(n11738), .B(n11739), .Z(n11734) );
  ANDN U12788 ( .B(n11740), .A(n6864), .Z(n11738) );
  XNOR U12789 ( .A(n11741), .B(n11742), .Z(n6864) );
  IV U12790 ( .A(n11739), .Z(n11742) );
  XOR U12791 ( .A(n6863), .B(n11739), .Z(n11740) );
  XOR U12792 ( .A(n11743), .B(n11744), .Z(n11739) );
  ANDN U12793 ( .B(n11745), .A(n6874), .Z(n11743) );
  XNOR U12794 ( .A(n11746), .B(n11747), .Z(n6874) );
  IV U12795 ( .A(n11744), .Z(n11747) );
  XOR U12796 ( .A(n6873), .B(n11744), .Z(n11745) );
  XOR U12797 ( .A(n11748), .B(n11749), .Z(n11744) );
  ANDN U12798 ( .B(n11750), .A(n6879), .Z(n11748) );
  XNOR U12799 ( .A(n11751), .B(n11752), .Z(n6879) );
  IV U12800 ( .A(n11749), .Z(n11752) );
  XOR U12801 ( .A(n6878), .B(n11749), .Z(n11750) );
  XOR U12802 ( .A(n11753), .B(n11754), .Z(n11749) );
  ANDN U12803 ( .B(n11755), .A(n6884), .Z(n11753) );
  XNOR U12804 ( .A(n11756), .B(n11757), .Z(n6884) );
  IV U12805 ( .A(n11754), .Z(n11757) );
  XOR U12806 ( .A(n6883), .B(n11754), .Z(n11755) );
  XOR U12807 ( .A(n11758), .B(n11759), .Z(n11754) );
  ANDN U12808 ( .B(n11760), .A(n6889), .Z(n11758) );
  XNOR U12809 ( .A(n11761), .B(n11762), .Z(n6889) );
  IV U12810 ( .A(n11759), .Z(n11762) );
  XOR U12811 ( .A(n6888), .B(n11759), .Z(n11760) );
  XOR U12812 ( .A(n11763), .B(n11764), .Z(n11759) );
  ANDN U12813 ( .B(n11765), .A(n6894), .Z(n11763) );
  XNOR U12814 ( .A(n11766), .B(n11767), .Z(n6894) );
  IV U12815 ( .A(n11764), .Z(n11767) );
  XOR U12816 ( .A(n6893), .B(n11764), .Z(n11765) );
  XOR U12817 ( .A(n11768), .B(n11769), .Z(n11764) );
  ANDN U12818 ( .B(n11770), .A(n6899), .Z(n11768) );
  XNOR U12819 ( .A(n11771), .B(n11772), .Z(n6899) );
  IV U12820 ( .A(n11769), .Z(n11772) );
  XOR U12821 ( .A(n6898), .B(n11769), .Z(n11770) );
  XOR U12822 ( .A(n11773), .B(n11774), .Z(n11769) );
  ANDN U12823 ( .B(n11775), .A(n6904), .Z(n11773) );
  XNOR U12824 ( .A(n11776), .B(n11777), .Z(n6904) );
  IV U12825 ( .A(n11774), .Z(n11777) );
  XOR U12826 ( .A(n6903), .B(n11774), .Z(n11775) );
  XOR U12827 ( .A(n11778), .B(n11779), .Z(n11774) );
  ANDN U12828 ( .B(n11780), .A(n6909), .Z(n11778) );
  XNOR U12829 ( .A(n11781), .B(n11782), .Z(n6909) );
  IV U12830 ( .A(n11779), .Z(n11782) );
  XOR U12831 ( .A(n6908), .B(n11779), .Z(n11780) );
  XOR U12832 ( .A(n11783), .B(n11784), .Z(n11779) );
  ANDN U12833 ( .B(n11785), .A(n6914), .Z(n11783) );
  XNOR U12834 ( .A(n11786), .B(n11787), .Z(n6914) );
  IV U12835 ( .A(n11784), .Z(n11787) );
  XOR U12836 ( .A(n6913), .B(n11784), .Z(n11785) );
  XOR U12837 ( .A(n11788), .B(n11789), .Z(n11784) );
  ANDN U12838 ( .B(n11790), .A(n6919), .Z(n11788) );
  XNOR U12839 ( .A(n11791), .B(n11792), .Z(n6919) );
  IV U12840 ( .A(n11789), .Z(n11792) );
  XOR U12841 ( .A(n6918), .B(n11789), .Z(n11790) );
  XOR U12842 ( .A(n11793), .B(n11794), .Z(n11789) );
  ANDN U12843 ( .B(n11795), .A(n6929), .Z(n11793) );
  XNOR U12844 ( .A(n11796), .B(n11797), .Z(n6929) );
  IV U12845 ( .A(n11794), .Z(n11797) );
  XOR U12846 ( .A(n6928), .B(n11794), .Z(n11795) );
  XOR U12847 ( .A(n11798), .B(n11799), .Z(n11794) );
  ANDN U12848 ( .B(n11800), .A(n6934), .Z(n11798) );
  XNOR U12849 ( .A(n11801), .B(n11802), .Z(n6934) );
  IV U12850 ( .A(n11799), .Z(n11802) );
  XOR U12851 ( .A(n6933), .B(n11799), .Z(n11800) );
  XOR U12852 ( .A(n11803), .B(n11804), .Z(n11799) );
  ANDN U12853 ( .B(n11805), .A(n6939), .Z(n11803) );
  XNOR U12854 ( .A(n11806), .B(n11807), .Z(n6939) );
  IV U12855 ( .A(n11804), .Z(n11807) );
  XOR U12856 ( .A(n6938), .B(n11804), .Z(n11805) );
  XOR U12857 ( .A(n11808), .B(n11809), .Z(n11804) );
  ANDN U12858 ( .B(n11810), .A(n6944), .Z(n11808) );
  XNOR U12859 ( .A(n11811), .B(n11812), .Z(n6944) );
  IV U12860 ( .A(n11809), .Z(n11812) );
  XOR U12861 ( .A(n6943), .B(n11809), .Z(n11810) );
  XOR U12862 ( .A(n11813), .B(n11814), .Z(n11809) );
  ANDN U12863 ( .B(n11815), .A(n6949), .Z(n11813) );
  XNOR U12864 ( .A(n11816), .B(n11817), .Z(n6949) );
  IV U12865 ( .A(n11814), .Z(n11817) );
  XOR U12866 ( .A(n6948), .B(n11814), .Z(n11815) );
  XOR U12867 ( .A(n11818), .B(n11819), .Z(n11814) );
  ANDN U12868 ( .B(n11820), .A(n6954), .Z(n11818) );
  XNOR U12869 ( .A(n11821), .B(n11822), .Z(n6954) );
  IV U12870 ( .A(n11819), .Z(n11822) );
  XOR U12871 ( .A(n6953), .B(n11819), .Z(n11820) );
  XOR U12872 ( .A(n11823), .B(n11824), .Z(n11819) );
  ANDN U12873 ( .B(n11825), .A(n6959), .Z(n11823) );
  XNOR U12874 ( .A(n11826), .B(n11827), .Z(n6959) );
  IV U12875 ( .A(n11824), .Z(n11827) );
  XOR U12876 ( .A(n6958), .B(n11824), .Z(n11825) );
  XOR U12877 ( .A(n11828), .B(n11829), .Z(n11824) );
  ANDN U12878 ( .B(n11830), .A(n6964), .Z(n11828) );
  XNOR U12879 ( .A(n11831), .B(n11832), .Z(n6964) );
  IV U12880 ( .A(n11829), .Z(n11832) );
  XOR U12881 ( .A(n6963), .B(n11829), .Z(n11830) );
  XOR U12882 ( .A(n11833), .B(n11834), .Z(n11829) );
  ANDN U12883 ( .B(n11835), .A(n6969), .Z(n11833) );
  XNOR U12884 ( .A(n11836), .B(n11837), .Z(n6969) );
  IV U12885 ( .A(n11834), .Z(n11837) );
  XOR U12886 ( .A(n6968), .B(n11834), .Z(n11835) );
  XOR U12887 ( .A(n11838), .B(n11839), .Z(n11834) );
  ANDN U12888 ( .B(n11840), .A(n6974), .Z(n11838) );
  XNOR U12889 ( .A(n11841), .B(n11842), .Z(n6974) );
  IV U12890 ( .A(n11839), .Z(n11842) );
  XOR U12891 ( .A(n6973), .B(n11839), .Z(n11840) );
  XOR U12892 ( .A(n11843), .B(n11844), .Z(n11839) );
  ANDN U12893 ( .B(n11845), .A(n6989), .Z(n11843) );
  XNOR U12894 ( .A(n11846), .B(n11847), .Z(n6989) );
  IV U12895 ( .A(n11844), .Z(n11847) );
  XOR U12896 ( .A(n6988), .B(n11844), .Z(n11845) );
  XOR U12897 ( .A(n11848), .B(n11849), .Z(n11844) );
  ANDN U12898 ( .B(n11850), .A(n6994), .Z(n11848) );
  XNOR U12899 ( .A(n11851), .B(n11852), .Z(n6994) );
  IV U12900 ( .A(n11849), .Z(n11852) );
  XOR U12901 ( .A(n6993), .B(n11849), .Z(n11850) );
  XOR U12902 ( .A(n11853), .B(n11854), .Z(n11849) );
  ANDN U12903 ( .B(n11855), .A(n6999), .Z(n11853) );
  XNOR U12904 ( .A(n11856), .B(n11857), .Z(n6999) );
  IV U12905 ( .A(n11854), .Z(n11857) );
  XOR U12906 ( .A(n6998), .B(n11854), .Z(n11855) );
  XOR U12907 ( .A(n11858), .B(n11859), .Z(n11854) );
  ANDN U12908 ( .B(n11860), .A(n7004), .Z(n11858) );
  XNOR U12909 ( .A(n11861), .B(n11862), .Z(n7004) );
  IV U12910 ( .A(n11859), .Z(n11862) );
  XOR U12911 ( .A(n7003), .B(n11859), .Z(n11860) );
  XOR U12912 ( .A(n11863), .B(n11864), .Z(n11859) );
  ANDN U12913 ( .B(n11865), .A(n7009), .Z(n11863) );
  XNOR U12914 ( .A(n11866), .B(n11867), .Z(n7009) );
  IV U12915 ( .A(n11864), .Z(n11867) );
  XOR U12916 ( .A(n7008), .B(n11864), .Z(n11865) );
  XOR U12917 ( .A(n11868), .B(n11869), .Z(n11864) );
  ANDN U12918 ( .B(n11870), .A(n7014), .Z(n11868) );
  XNOR U12919 ( .A(n11871), .B(n11872), .Z(n7014) );
  IV U12920 ( .A(n11869), .Z(n11872) );
  XOR U12921 ( .A(n7013), .B(n11869), .Z(n11870) );
  XOR U12922 ( .A(n11873), .B(n11874), .Z(n11869) );
  ANDN U12923 ( .B(n11875), .A(n7019), .Z(n11873) );
  XNOR U12924 ( .A(n11876), .B(n11877), .Z(n7019) );
  IV U12925 ( .A(n11874), .Z(n11877) );
  XOR U12926 ( .A(n7018), .B(n11874), .Z(n11875) );
  XOR U12927 ( .A(n11878), .B(n11879), .Z(n11874) );
  ANDN U12928 ( .B(n11880), .A(n7024), .Z(n11878) );
  XNOR U12929 ( .A(n11881), .B(n11882), .Z(n7024) );
  IV U12930 ( .A(n11879), .Z(n11882) );
  XOR U12931 ( .A(n7023), .B(n11879), .Z(n11880) );
  XOR U12932 ( .A(n11883), .B(n11884), .Z(n11879) );
  ANDN U12933 ( .B(n11885), .A(n7029), .Z(n11883) );
  XNOR U12934 ( .A(n11886), .B(n11887), .Z(n7029) );
  IV U12935 ( .A(n11884), .Z(n11887) );
  XOR U12936 ( .A(n7028), .B(n11884), .Z(n11885) );
  XOR U12937 ( .A(n11888), .B(n11889), .Z(n11884) );
  ANDN U12938 ( .B(n11890), .A(n7034), .Z(n11888) );
  XNOR U12939 ( .A(n11891), .B(n11892), .Z(n7034) );
  IV U12940 ( .A(n11889), .Z(n11892) );
  XOR U12941 ( .A(n7033), .B(n11889), .Z(n11890) );
  XOR U12942 ( .A(n11893), .B(n11894), .Z(n11889) );
  ANDN U12943 ( .B(n11895), .A(n7044), .Z(n11893) );
  XNOR U12944 ( .A(n11896), .B(n11897), .Z(n7044) );
  IV U12945 ( .A(n11894), .Z(n11897) );
  XOR U12946 ( .A(n7043), .B(n11894), .Z(n11895) );
  XOR U12947 ( .A(n11898), .B(n11899), .Z(n11894) );
  ANDN U12948 ( .B(n11900), .A(n7049), .Z(n11898) );
  XNOR U12949 ( .A(n11901), .B(n11902), .Z(n7049) );
  IV U12950 ( .A(n11899), .Z(n11902) );
  XOR U12951 ( .A(n7048), .B(n11899), .Z(n11900) );
  XOR U12952 ( .A(n11903), .B(n11904), .Z(n11899) );
  ANDN U12953 ( .B(n11905), .A(n7054), .Z(n11903) );
  XNOR U12954 ( .A(n11906), .B(n11907), .Z(n7054) );
  IV U12955 ( .A(n11904), .Z(n11907) );
  XOR U12956 ( .A(n7053), .B(n11904), .Z(n11905) );
  XOR U12957 ( .A(n11908), .B(n11909), .Z(n11904) );
  ANDN U12958 ( .B(n11910), .A(n7059), .Z(n11908) );
  XNOR U12959 ( .A(n11911), .B(n11912), .Z(n7059) );
  IV U12960 ( .A(n11909), .Z(n11912) );
  XOR U12961 ( .A(n7058), .B(n11909), .Z(n11910) );
  XOR U12962 ( .A(n11913), .B(n11914), .Z(n11909) );
  ANDN U12963 ( .B(n11915), .A(n7064), .Z(n11913) );
  XNOR U12964 ( .A(n11916), .B(n11917), .Z(n7064) );
  IV U12965 ( .A(n11914), .Z(n11917) );
  XOR U12966 ( .A(n7063), .B(n11914), .Z(n11915) );
  XOR U12967 ( .A(n11918), .B(n11919), .Z(n11914) );
  ANDN U12968 ( .B(n11920), .A(n7069), .Z(n11918) );
  XNOR U12969 ( .A(n11921), .B(n11922), .Z(n7069) );
  IV U12970 ( .A(n11919), .Z(n11922) );
  XOR U12971 ( .A(n7068), .B(n11919), .Z(n11920) );
  XOR U12972 ( .A(n11923), .B(n11924), .Z(n11919) );
  ANDN U12973 ( .B(n11925), .A(n7074), .Z(n11923) );
  XNOR U12974 ( .A(n11926), .B(n11927), .Z(n7074) );
  IV U12975 ( .A(n11924), .Z(n11927) );
  XOR U12976 ( .A(n7073), .B(n11924), .Z(n11925) );
  XOR U12977 ( .A(n11928), .B(n11929), .Z(n11924) );
  ANDN U12978 ( .B(n11930), .A(n7079), .Z(n11928) );
  XNOR U12979 ( .A(n11931), .B(n11932), .Z(n7079) );
  IV U12980 ( .A(n11929), .Z(n11932) );
  XOR U12981 ( .A(n7078), .B(n11929), .Z(n11930) );
  XOR U12982 ( .A(n11933), .B(n11934), .Z(n11929) );
  ANDN U12983 ( .B(n11935), .A(n7084), .Z(n11933) );
  XNOR U12984 ( .A(n11936), .B(n11937), .Z(n7084) );
  IV U12985 ( .A(n11934), .Z(n11937) );
  XOR U12986 ( .A(n7083), .B(n11934), .Z(n11935) );
  XOR U12987 ( .A(n11938), .B(n11939), .Z(n11934) );
  ANDN U12988 ( .B(n11940), .A(n7089), .Z(n11938) );
  XNOR U12989 ( .A(n11941), .B(n11942), .Z(n7089) );
  IV U12990 ( .A(n11939), .Z(n11942) );
  XOR U12991 ( .A(n7088), .B(n11939), .Z(n11940) );
  XOR U12992 ( .A(n11943), .B(n11944), .Z(n11939) );
  ANDN U12993 ( .B(n11945), .A(n7099), .Z(n11943) );
  XNOR U12994 ( .A(n11946), .B(n11947), .Z(n7099) );
  IV U12995 ( .A(n11944), .Z(n11947) );
  XOR U12996 ( .A(n7098), .B(n11944), .Z(n11945) );
  XOR U12997 ( .A(n11948), .B(n11949), .Z(n11944) );
  ANDN U12998 ( .B(n11950), .A(n7104), .Z(n11948) );
  XNOR U12999 ( .A(n11951), .B(n11952), .Z(n7104) );
  IV U13000 ( .A(n11949), .Z(n11952) );
  XOR U13001 ( .A(n7103), .B(n11949), .Z(n11950) );
  XOR U13002 ( .A(n11953), .B(n11954), .Z(n11949) );
  ANDN U13003 ( .B(n11955), .A(n7109), .Z(n11953) );
  XNOR U13004 ( .A(n11956), .B(n11957), .Z(n7109) );
  IV U13005 ( .A(n11954), .Z(n11957) );
  XOR U13006 ( .A(n7108), .B(n11954), .Z(n11955) );
  XOR U13007 ( .A(n11958), .B(n11959), .Z(n11954) );
  ANDN U13008 ( .B(n11960), .A(n7114), .Z(n11958) );
  XNOR U13009 ( .A(n11961), .B(n11962), .Z(n7114) );
  IV U13010 ( .A(n11959), .Z(n11962) );
  XOR U13011 ( .A(n7113), .B(n11959), .Z(n11960) );
  XOR U13012 ( .A(n11963), .B(n11964), .Z(n11959) );
  ANDN U13013 ( .B(n11965), .A(n7119), .Z(n11963) );
  XNOR U13014 ( .A(n11966), .B(n11967), .Z(n7119) );
  IV U13015 ( .A(n11964), .Z(n11967) );
  XOR U13016 ( .A(n7118), .B(n11964), .Z(n11965) );
  XOR U13017 ( .A(n11968), .B(n11969), .Z(n11964) );
  ANDN U13018 ( .B(n11970), .A(n7124), .Z(n11968) );
  XNOR U13019 ( .A(n11971), .B(n11972), .Z(n7124) );
  IV U13020 ( .A(n11969), .Z(n11972) );
  XOR U13021 ( .A(n7123), .B(n11969), .Z(n11970) );
  XOR U13022 ( .A(n11973), .B(n11974), .Z(n11969) );
  ANDN U13023 ( .B(n11975), .A(n7129), .Z(n11973) );
  XNOR U13024 ( .A(n11976), .B(n11977), .Z(n7129) );
  IV U13025 ( .A(n11974), .Z(n11977) );
  XOR U13026 ( .A(n7128), .B(n11974), .Z(n11975) );
  XOR U13027 ( .A(n11978), .B(n11979), .Z(n11974) );
  ANDN U13028 ( .B(n11980), .A(n7134), .Z(n11978) );
  XNOR U13029 ( .A(n11981), .B(n11982), .Z(n7134) );
  IV U13030 ( .A(n11979), .Z(n11982) );
  XOR U13031 ( .A(n7133), .B(n11979), .Z(n11980) );
  XOR U13032 ( .A(n11983), .B(n11984), .Z(n11979) );
  ANDN U13033 ( .B(n11985), .A(n7139), .Z(n11983) );
  XNOR U13034 ( .A(n11986), .B(n11987), .Z(n7139) );
  IV U13035 ( .A(n11984), .Z(n11987) );
  XOR U13036 ( .A(n7138), .B(n11984), .Z(n11985) );
  XOR U13037 ( .A(n11988), .B(n11989), .Z(n11984) );
  ANDN U13038 ( .B(n11990), .A(n7144), .Z(n11988) );
  XNOR U13039 ( .A(n11991), .B(n11992), .Z(n7144) );
  IV U13040 ( .A(n11989), .Z(n11992) );
  XOR U13041 ( .A(n7143), .B(n11989), .Z(n11990) );
  XOR U13042 ( .A(n11993), .B(n11994), .Z(n11989) );
  ANDN U13043 ( .B(n11995), .A(n7154), .Z(n11993) );
  XNOR U13044 ( .A(n11996), .B(n11997), .Z(n7154) );
  IV U13045 ( .A(n11994), .Z(n11997) );
  XOR U13046 ( .A(n7153), .B(n11994), .Z(n11995) );
  XOR U13047 ( .A(n11998), .B(n11999), .Z(n11994) );
  ANDN U13048 ( .B(n12000), .A(n7159), .Z(n11998) );
  XNOR U13049 ( .A(n12001), .B(n12002), .Z(n7159) );
  IV U13050 ( .A(n11999), .Z(n12002) );
  XOR U13051 ( .A(n7158), .B(n11999), .Z(n12000) );
  XOR U13052 ( .A(n12003), .B(n12004), .Z(n11999) );
  ANDN U13053 ( .B(n12005), .A(n7164), .Z(n12003) );
  XNOR U13054 ( .A(n12006), .B(n12007), .Z(n7164) );
  IV U13055 ( .A(n12004), .Z(n12007) );
  XOR U13056 ( .A(n7163), .B(n12004), .Z(n12005) );
  XOR U13057 ( .A(n12008), .B(n12009), .Z(n12004) );
  ANDN U13058 ( .B(n12010), .A(n7169), .Z(n12008) );
  XNOR U13059 ( .A(n12011), .B(n12012), .Z(n7169) );
  IV U13060 ( .A(n12009), .Z(n12012) );
  XOR U13061 ( .A(n7168), .B(n12009), .Z(n12010) );
  XOR U13062 ( .A(n12013), .B(n12014), .Z(n12009) );
  ANDN U13063 ( .B(n12015), .A(n7174), .Z(n12013) );
  XNOR U13064 ( .A(n12016), .B(n12017), .Z(n7174) );
  IV U13065 ( .A(n12014), .Z(n12017) );
  XOR U13066 ( .A(n7173), .B(n12014), .Z(n12015) );
  XOR U13067 ( .A(n12018), .B(n12019), .Z(n12014) );
  ANDN U13068 ( .B(n12020), .A(n7179), .Z(n12018) );
  XNOR U13069 ( .A(n12021), .B(n12022), .Z(n7179) );
  IV U13070 ( .A(n12019), .Z(n12022) );
  XOR U13071 ( .A(n7178), .B(n12019), .Z(n12020) );
  XOR U13072 ( .A(n12023), .B(n12024), .Z(n12019) );
  ANDN U13073 ( .B(n12025), .A(n7184), .Z(n12023) );
  XNOR U13074 ( .A(n12026), .B(n12027), .Z(n7184) );
  IV U13075 ( .A(n12024), .Z(n12027) );
  XOR U13076 ( .A(n7183), .B(n12024), .Z(n12025) );
  XOR U13077 ( .A(n12028), .B(n12029), .Z(n12024) );
  ANDN U13078 ( .B(n12030), .A(n7189), .Z(n12028) );
  XNOR U13079 ( .A(n12031), .B(n12032), .Z(n7189) );
  IV U13080 ( .A(n12029), .Z(n12032) );
  XOR U13081 ( .A(n7188), .B(n12029), .Z(n12030) );
  XOR U13082 ( .A(n12033), .B(n12034), .Z(n12029) );
  ANDN U13083 ( .B(n12035), .A(n7194), .Z(n12033) );
  XNOR U13084 ( .A(n12036), .B(n12037), .Z(n7194) );
  IV U13085 ( .A(n12034), .Z(n12037) );
  XOR U13086 ( .A(n7193), .B(n12034), .Z(n12035) );
  XOR U13087 ( .A(n12038), .B(n12039), .Z(n12034) );
  ANDN U13088 ( .B(n12040), .A(n7199), .Z(n12038) );
  XNOR U13089 ( .A(n12041), .B(n12042), .Z(n7199) );
  IV U13090 ( .A(n12039), .Z(n12042) );
  XOR U13091 ( .A(n7198), .B(n12039), .Z(n12040) );
  XOR U13092 ( .A(n12043), .B(n12044), .Z(n12039) );
  ANDN U13093 ( .B(n12045), .A(n7209), .Z(n12043) );
  XNOR U13094 ( .A(n12046), .B(n12047), .Z(n7209) );
  IV U13095 ( .A(n12044), .Z(n12047) );
  XOR U13096 ( .A(n7208), .B(n12044), .Z(n12045) );
  XOR U13097 ( .A(n12048), .B(n12049), .Z(n12044) );
  ANDN U13098 ( .B(n12050), .A(n7214), .Z(n12048) );
  XNOR U13099 ( .A(n12051), .B(n12052), .Z(n7214) );
  IV U13100 ( .A(n12049), .Z(n12052) );
  XOR U13101 ( .A(n7213), .B(n12049), .Z(n12050) );
  XOR U13102 ( .A(n12053), .B(n12054), .Z(n12049) );
  ANDN U13103 ( .B(n12055), .A(n7219), .Z(n12053) );
  XNOR U13104 ( .A(n12056), .B(n12057), .Z(n7219) );
  IV U13105 ( .A(n12054), .Z(n12057) );
  XOR U13106 ( .A(n7218), .B(n12054), .Z(n12055) );
  XOR U13107 ( .A(n12058), .B(n12059), .Z(n12054) );
  ANDN U13108 ( .B(n12060), .A(n7224), .Z(n12058) );
  XNOR U13109 ( .A(n12061), .B(n12062), .Z(n7224) );
  IV U13110 ( .A(n12059), .Z(n12062) );
  XOR U13111 ( .A(n7223), .B(n12059), .Z(n12060) );
  XOR U13112 ( .A(n12063), .B(n12064), .Z(n12059) );
  ANDN U13113 ( .B(n12065), .A(n7229), .Z(n12063) );
  XNOR U13114 ( .A(n12066), .B(n12067), .Z(n7229) );
  IV U13115 ( .A(n12064), .Z(n12067) );
  XOR U13116 ( .A(n7228), .B(n12064), .Z(n12065) );
  XOR U13117 ( .A(n12068), .B(n12069), .Z(n12064) );
  ANDN U13118 ( .B(n12070), .A(n7234), .Z(n12068) );
  XNOR U13119 ( .A(n12071), .B(n12072), .Z(n7234) );
  IV U13120 ( .A(n12069), .Z(n12072) );
  XOR U13121 ( .A(n7233), .B(n12069), .Z(n12070) );
  XOR U13122 ( .A(n12073), .B(n12074), .Z(n12069) );
  ANDN U13123 ( .B(n12075), .A(n7239), .Z(n12073) );
  XNOR U13124 ( .A(n12076), .B(n12077), .Z(n7239) );
  IV U13125 ( .A(n12074), .Z(n12077) );
  XOR U13126 ( .A(n7238), .B(n12074), .Z(n12075) );
  XOR U13127 ( .A(n12078), .B(n12079), .Z(n12074) );
  ANDN U13128 ( .B(n12080), .A(n7244), .Z(n12078) );
  XNOR U13129 ( .A(n12081), .B(n12082), .Z(n7244) );
  IV U13130 ( .A(n12079), .Z(n12082) );
  XOR U13131 ( .A(n7243), .B(n12079), .Z(n12080) );
  XOR U13132 ( .A(n12083), .B(n12084), .Z(n12079) );
  ANDN U13133 ( .B(n12085), .A(n7249), .Z(n12083) );
  XNOR U13134 ( .A(n12086), .B(n12087), .Z(n7249) );
  IV U13135 ( .A(n12084), .Z(n12087) );
  XOR U13136 ( .A(n7248), .B(n12084), .Z(n12085) );
  XOR U13137 ( .A(n12088), .B(n12089), .Z(n12084) );
  ANDN U13138 ( .B(n12090), .A(n7254), .Z(n12088) );
  XNOR U13139 ( .A(n12091), .B(n12092), .Z(n7254) );
  IV U13140 ( .A(n12089), .Z(n12092) );
  XOR U13141 ( .A(n7253), .B(n12089), .Z(n12090) );
  XOR U13142 ( .A(n12093), .B(n12094), .Z(n12089) );
  ANDN U13143 ( .B(n12095), .A(n7264), .Z(n12093) );
  XNOR U13144 ( .A(n12096), .B(n12097), .Z(n7264) );
  IV U13145 ( .A(n12094), .Z(n12097) );
  XOR U13146 ( .A(n7263), .B(n12094), .Z(n12095) );
  XOR U13147 ( .A(n12098), .B(n12099), .Z(n12094) );
  ANDN U13148 ( .B(n12100), .A(n7269), .Z(n12098) );
  XNOR U13149 ( .A(n12101), .B(n12102), .Z(n7269) );
  IV U13150 ( .A(n12099), .Z(n12102) );
  XOR U13151 ( .A(n7268), .B(n12099), .Z(n12100) );
  XOR U13152 ( .A(n12103), .B(n12104), .Z(n12099) );
  ANDN U13153 ( .B(n12105), .A(n7274), .Z(n12103) );
  XNOR U13154 ( .A(n12106), .B(n12107), .Z(n7274) );
  IV U13155 ( .A(n12104), .Z(n12107) );
  XOR U13156 ( .A(n7273), .B(n12104), .Z(n12105) );
  XOR U13157 ( .A(n12108), .B(n12109), .Z(n12104) );
  ANDN U13158 ( .B(n12110), .A(n7279), .Z(n12108) );
  XNOR U13159 ( .A(n12111), .B(n12112), .Z(n7279) );
  IV U13160 ( .A(n12109), .Z(n12112) );
  XOR U13161 ( .A(n7278), .B(n12109), .Z(n12110) );
  XOR U13162 ( .A(n12113), .B(n12114), .Z(n12109) );
  ANDN U13163 ( .B(n12115), .A(n7284), .Z(n12113) );
  XNOR U13164 ( .A(n12116), .B(n12117), .Z(n7284) );
  IV U13165 ( .A(n12114), .Z(n12117) );
  XOR U13166 ( .A(n7283), .B(n12114), .Z(n12115) );
  XOR U13167 ( .A(n12118), .B(n12119), .Z(n12114) );
  ANDN U13168 ( .B(n12120), .A(n7289), .Z(n12118) );
  XNOR U13169 ( .A(n12121), .B(n12122), .Z(n7289) );
  IV U13170 ( .A(n12119), .Z(n12122) );
  XOR U13171 ( .A(n7288), .B(n12119), .Z(n12120) );
  XOR U13172 ( .A(n12123), .B(n12124), .Z(n12119) );
  ANDN U13173 ( .B(n12125), .A(n7294), .Z(n12123) );
  XNOR U13174 ( .A(n12126), .B(n12127), .Z(n7294) );
  IV U13175 ( .A(n12124), .Z(n12127) );
  XOR U13176 ( .A(n7293), .B(n12124), .Z(n12125) );
  XOR U13177 ( .A(n12128), .B(n12129), .Z(n12124) );
  ANDN U13178 ( .B(n12130), .A(n7299), .Z(n12128) );
  XNOR U13179 ( .A(n12131), .B(n12132), .Z(n7299) );
  IV U13180 ( .A(n12129), .Z(n12132) );
  XOR U13181 ( .A(n7298), .B(n12129), .Z(n12130) );
  XOR U13182 ( .A(n12133), .B(n12134), .Z(n12129) );
  ANDN U13183 ( .B(n12135), .A(n7304), .Z(n12133) );
  XNOR U13184 ( .A(n12136), .B(n12137), .Z(n7304) );
  IV U13185 ( .A(n12134), .Z(n12137) );
  XOR U13186 ( .A(n7303), .B(n12134), .Z(n12135) );
  XOR U13187 ( .A(n12138), .B(n12139), .Z(n12134) );
  ANDN U13188 ( .B(n12140), .A(n7309), .Z(n12138) );
  XNOR U13189 ( .A(n12141), .B(n12142), .Z(n7309) );
  IV U13190 ( .A(n12139), .Z(n12142) );
  XOR U13191 ( .A(n7308), .B(n12139), .Z(n12140) );
  XOR U13192 ( .A(n12143), .B(n12144), .Z(n12139) );
  ANDN U13193 ( .B(n12145), .A(n7319), .Z(n12143) );
  XNOR U13194 ( .A(n12146), .B(n12147), .Z(n7319) );
  IV U13195 ( .A(n12144), .Z(n12147) );
  XOR U13196 ( .A(n7318), .B(n12144), .Z(n12145) );
  XOR U13197 ( .A(n12148), .B(n12149), .Z(n12144) );
  ANDN U13198 ( .B(n12150), .A(n7324), .Z(n12148) );
  XNOR U13199 ( .A(n12151), .B(n12152), .Z(n7324) );
  IV U13200 ( .A(n12149), .Z(n12152) );
  XOR U13201 ( .A(n7323), .B(n12149), .Z(n12150) );
  XOR U13202 ( .A(n12153), .B(n12154), .Z(n12149) );
  ANDN U13203 ( .B(n12155), .A(n7329), .Z(n12153) );
  XNOR U13204 ( .A(n12156), .B(n12157), .Z(n7329) );
  IV U13205 ( .A(n12154), .Z(n12157) );
  XOR U13206 ( .A(n7328), .B(n12154), .Z(n12155) );
  XOR U13207 ( .A(n12158), .B(n12159), .Z(n12154) );
  ANDN U13208 ( .B(n12160), .A(n7334), .Z(n12158) );
  XNOR U13209 ( .A(n12161), .B(n12162), .Z(n7334) );
  IV U13210 ( .A(n12159), .Z(n12162) );
  XOR U13211 ( .A(n7333), .B(n12159), .Z(n12160) );
  XOR U13212 ( .A(n12163), .B(n12164), .Z(n12159) );
  ANDN U13213 ( .B(n12165), .A(n7339), .Z(n12163) );
  XNOR U13214 ( .A(n12166), .B(n12167), .Z(n7339) );
  IV U13215 ( .A(n12164), .Z(n12167) );
  XOR U13216 ( .A(n7338), .B(n12164), .Z(n12165) );
  XOR U13217 ( .A(n12168), .B(n12169), .Z(n12164) );
  ANDN U13218 ( .B(n12170), .A(n7344), .Z(n12168) );
  XNOR U13219 ( .A(n12171), .B(n12172), .Z(n7344) );
  IV U13220 ( .A(n12169), .Z(n12172) );
  XOR U13221 ( .A(n7343), .B(n12169), .Z(n12170) );
  XOR U13222 ( .A(n12173), .B(n12174), .Z(n12169) );
  ANDN U13223 ( .B(n12175), .A(n7349), .Z(n12173) );
  XNOR U13224 ( .A(n12176), .B(n12177), .Z(n7349) );
  IV U13225 ( .A(n12174), .Z(n12177) );
  XOR U13226 ( .A(n7348), .B(n12174), .Z(n12175) );
  XOR U13227 ( .A(n12178), .B(n12179), .Z(n12174) );
  ANDN U13228 ( .B(n12180), .A(n7354), .Z(n12178) );
  XNOR U13229 ( .A(n12181), .B(n12182), .Z(n7354) );
  IV U13230 ( .A(n12179), .Z(n12182) );
  XOR U13231 ( .A(n7353), .B(n12179), .Z(n12180) );
  XOR U13232 ( .A(n12183), .B(n12184), .Z(n12179) );
  ANDN U13233 ( .B(n12185), .A(n7359), .Z(n12183) );
  XNOR U13234 ( .A(n12186), .B(n12187), .Z(n7359) );
  IV U13235 ( .A(n12184), .Z(n12187) );
  XOR U13236 ( .A(n7358), .B(n12184), .Z(n12185) );
  XOR U13237 ( .A(n12188), .B(n12189), .Z(n12184) );
  ANDN U13238 ( .B(n12190), .A(n7364), .Z(n12188) );
  XNOR U13239 ( .A(n12191), .B(n12192), .Z(n7364) );
  IV U13240 ( .A(n12189), .Z(n12192) );
  XOR U13241 ( .A(n7363), .B(n12189), .Z(n12190) );
  XOR U13242 ( .A(n12193), .B(n12194), .Z(n12189) );
  ANDN U13243 ( .B(n12195), .A(n7374), .Z(n12193) );
  XNOR U13244 ( .A(n12196), .B(n12197), .Z(n7374) );
  IV U13245 ( .A(n12194), .Z(n12197) );
  XOR U13246 ( .A(n7373), .B(n12194), .Z(n12195) );
  XOR U13247 ( .A(n12198), .B(n12199), .Z(n12194) );
  ANDN U13248 ( .B(n12200), .A(n7379), .Z(n12198) );
  XNOR U13249 ( .A(n12201), .B(n12202), .Z(n7379) );
  IV U13250 ( .A(n12199), .Z(n12202) );
  XOR U13251 ( .A(n7378), .B(n12199), .Z(n12200) );
  XOR U13252 ( .A(n12203), .B(n12204), .Z(n12199) );
  ANDN U13253 ( .B(n12205), .A(n7384), .Z(n12203) );
  XNOR U13254 ( .A(n12206), .B(n12207), .Z(n7384) );
  IV U13255 ( .A(n12204), .Z(n12207) );
  XOR U13256 ( .A(n7383), .B(n12204), .Z(n12205) );
  XOR U13257 ( .A(n12208), .B(n12209), .Z(n12204) );
  ANDN U13258 ( .B(n12210), .A(n7389), .Z(n12208) );
  XNOR U13259 ( .A(n12211), .B(n12212), .Z(n7389) );
  IV U13260 ( .A(n12209), .Z(n12212) );
  XOR U13261 ( .A(n7388), .B(n12209), .Z(n12210) );
  XOR U13262 ( .A(n12213), .B(n12214), .Z(n12209) );
  ANDN U13263 ( .B(n12215), .A(n7394), .Z(n12213) );
  XNOR U13264 ( .A(n12216), .B(n12217), .Z(n7394) );
  IV U13265 ( .A(n12214), .Z(n12217) );
  XOR U13266 ( .A(n7393), .B(n12214), .Z(n12215) );
  XOR U13267 ( .A(n12218), .B(n12219), .Z(n12214) );
  ANDN U13268 ( .B(n12220), .A(n7399), .Z(n12218) );
  XNOR U13269 ( .A(n12221), .B(n12222), .Z(n7399) );
  IV U13270 ( .A(n12219), .Z(n12222) );
  XOR U13271 ( .A(n7398), .B(n12219), .Z(n12220) );
  XOR U13272 ( .A(n12223), .B(n12224), .Z(n12219) );
  ANDN U13273 ( .B(n12225), .A(n7404), .Z(n12223) );
  XNOR U13274 ( .A(n12226), .B(n12227), .Z(n7404) );
  IV U13275 ( .A(n12224), .Z(n12227) );
  XOR U13276 ( .A(n7403), .B(n12224), .Z(n12225) );
  XOR U13277 ( .A(n12228), .B(n12229), .Z(n12224) );
  ANDN U13278 ( .B(n12230), .A(n7409), .Z(n12228) );
  XNOR U13279 ( .A(n12231), .B(n12232), .Z(n7409) );
  IV U13280 ( .A(n12229), .Z(n12232) );
  XOR U13281 ( .A(n7408), .B(n12229), .Z(n12230) );
  XOR U13282 ( .A(n12233), .B(n12234), .Z(n12229) );
  ANDN U13283 ( .B(n12235), .A(n7414), .Z(n12233) );
  XNOR U13284 ( .A(n12236), .B(n12237), .Z(n7414) );
  IV U13285 ( .A(n12234), .Z(n12237) );
  XOR U13286 ( .A(n7413), .B(n12234), .Z(n12235) );
  XOR U13287 ( .A(n12238), .B(n12239), .Z(n12234) );
  ANDN U13288 ( .B(n12240), .A(n7419), .Z(n12238) );
  XNOR U13289 ( .A(n12241), .B(n12242), .Z(n7419) );
  IV U13290 ( .A(n12239), .Z(n12242) );
  XOR U13291 ( .A(n7418), .B(n12239), .Z(n12240) );
  XOR U13292 ( .A(n12243), .B(n12244), .Z(n12239) );
  ANDN U13293 ( .B(n12245), .A(n7429), .Z(n12243) );
  XNOR U13294 ( .A(n12246), .B(n12247), .Z(n7429) );
  IV U13295 ( .A(n12244), .Z(n12247) );
  XOR U13296 ( .A(n7428), .B(n12244), .Z(n12245) );
  XOR U13297 ( .A(n12248), .B(n12249), .Z(n12244) );
  ANDN U13298 ( .B(n12250), .A(n7434), .Z(n12248) );
  XNOR U13299 ( .A(n12251), .B(n12252), .Z(n7434) );
  IV U13300 ( .A(n12249), .Z(n12252) );
  XOR U13301 ( .A(n7433), .B(n12249), .Z(n12250) );
  XOR U13302 ( .A(n12253), .B(n12254), .Z(n12249) );
  ANDN U13303 ( .B(n12255), .A(n7439), .Z(n12253) );
  XNOR U13304 ( .A(n12256), .B(n12257), .Z(n7439) );
  IV U13305 ( .A(n12254), .Z(n12257) );
  XOR U13306 ( .A(n7438), .B(n12254), .Z(n12255) );
  XOR U13307 ( .A(n12258), .B(n12259), .Z(n12254) );
  ANDN U13308 ( .B(n12260), .A(n7444), .Z(n12258) );
  XNOR U13309 ( .A(n12261), .B(n12262), .Z(n7444) );
  IV U13310 ( .A(n12259), .Z(n12262) );
  XOR U13311 ( .A(n7443), .B(n12259), .Z(n12260) );
  XOR U13312 ( .A(n12263), .B(n12264), .Z(n12259) );
  ANDN U13313 ( .B(n12265), .A(n7449), .Z(n12263) );
  XNOR U13314 ( .A(n12266), .B(n12267), .Z(n7449) );
  IV U13315 ( .A(n12264), .Z(n12267) );
  XOR U13316 ( .A(n7448), .B(n12264), .Z(n12265) );
  XOR U13317 ( .A(n12268), .B(n12269), .Z(n12264) );
  ANDN U13318 ( .B(n12270), .A(n7454), .Z(n12268) );
  XNOR U13319 ( .A(n12271), .B(n12272), .Z(n7454) );
  IV U13320 ( .A(n12269), .Z(n12272) );
  XOR U13321 ( .A(n7453), .B(n12269), .Z(n12270) );
  XOR U13322 ( .A(n12273), .B(n12274), .Z(n12269) );
  ANDN U13323 ( .B(n12275), .A(n7459), .Z(n12273) );
  XNOR U13324 ( .A(n12276), .B(n12277), .Z(n7459) );
  IV U13325 ( .A(n12274), .Z(n12277) );
  XOR U13326 ( .A(n7458), .B(n12274), .Z(n12275) );
  XOR U13327 ( .A(n12278), .B(n12279), .Z(n12274) );
  ANDN U13328 ( .B(n12280), .A(n7464), .Z(n12278) );
  XNOR U13329 ( .A(n12281), .B(n12282), .Z(n7464) );
  IV U13330 ( .A(n12279), .Z(n12282) );
  XOR U13331 ( .A(n7463), .B(n12279), .Z(n12280) );
  XOR U13332 ( .A(n12283), .B(n12284), .Z(n12279) );
  ANDN U13333 ( .B(n12285), .A(n7469), .Z(n12283) );
  XNOR U13334 ( .A(n12286), .B(n12287), .Z(n7469) );
  IV U13335 ( .A(n12284), .Z(n12287) );
  XOR U13336 ( .A(n7468), .B(n12284), .Z(n12285) );
  XOR U13337 ( .A(n12288), .B(n12289), .Z(n12284) );
  ANDN U13338 ( .B(n12290), .A(n7474), .Z(n12288) );
  XNOR U13339 ( .A(n12291), .B(n12292), .Z(n7474) );
  IV U13340 ( .A(n12289), .Z(n12292) );
  XOR U13341 ( .A(n7473), .B(n12289), .Z(n12290) );
  XOR U13342 ( .A(n12293), .B(n12294), .Z(n12289) );
  ANDN U13343 ( .B(n12295), .A(n7484), .Z(n12293) );
  XNOR U13344 ( .A(n12296), .B(n12297), .Z(n7484) );
  IV U13345 ( .A(n12294), .Z(n12297) );
  XOR U13346 ( .A(n7483), .B(n12294), .Z(n12295) );
  XOR U13347 ( .A(n12298), .B(n12299), .Z(n12294) );
  ANDN U13348 ( .B(n12300), .A(n7489), .Z(n12298) );
  XNOR U13349 ( .A(n12301), .B(n12302), .Z(n7489) );
  IV U13350 ( .A(n12299), .Z(n12302) );
  XOR U13351 ( .A(n7488), .B(n12299), .Z(n12300) );
  XOR U13352 ( .A(n12303), .B(n12304), .Z(n12299) );
  ANDN U13353 ( .B(n12305), .A(n7494), .Z(n12303) );
  XNOR U13354 ( .A(n12306), .B(n12307), .Z(n7494) );
  IV U13355 ( .A(n12304), .Z(n12307) );
  XOR U13356 ( .A(n7493), .B(n12304), .Z(n12305) );
  XOR U13357 ( .A(n12308), .B(n12309), .Z(n12304) );
  ANDN U13358 ( .B(n12310), .A(n7499), .Z(n12308) );
  XNOR U13359 ( .A(n12311), .B(n12312), .Z(n7499) );
  IV U13360 ( .A(n12309), .Z(n12312) );
  XOR U13361 ( .A(n7498), .B(n12309), .Z(n12310) );
  XOR U13362 ( .A(n12313), .B(n12314), .Z(n12309) );
  ANDN U13363 ( .B(n12315), .A(n7504), .Z(n12313) );
  XNOR U13364 ( .A(n12316), .B(n12317), .Z(n7504) );
  IV U13365 ( .A(n12314), .Z(n12317) );
  XOR U13366 ( .A(n7503), .B(n12314), .Z(n12315) );
  XOR U13367 ( .A(n12318), .B(n12319), .Z(n12314) );
  ANDN U13368 ( .B(n12320), .A(n7509), .Z(n12318) );
  XNOR U13369 ( .A(n12321), .B(n12322), .Z(n7509) );
  IV U13370 ( .A(n12319), .Z(n12322) );
  XOR U13371 ( .A(n7508), .B(n12319), .Z(n12320) );
  XOR U13372 ( .A(n12323), .B(n12324), .Z(n12319) );
  ANDN U13373 ( .B(n12325), .A(n7514), .Z(n12323) );
  XNOR U13374 ( .A(n12326), .B(n12327), .Z(n7514) );
  IV U13375 ( .A(n12324), .Z(n12327) );
  XOR U13376 ( .A(n7513), .B(n12324), .Z(n12325) );
  XOR U13377 ( .A(n12328), .B(n12329), .Z(n12324) );
  ANDN U13378 ( .B(n12330), .A(n7519), .Z(n12328) );
  XNOR U13379 ( .A(n12331), .B(n12332), .Z(n7519) );
  IV U13380 ( .A(n12329), .Z(n12332) );
  XOR U13381 ( .A(n7518), .B(n12329), .Z(n12330) );
  XOR U13382 ( .A(n12333), .B(n12334), .Z(n12329) );
  ANDN U13383 ( .B(n12335), .A(n7524), .Z(n12333) );
  XNOR U13384 ( .A(n12336), .B(n12337), .Z(n7524) );
  IV U13385 ( .A(n12334), .Z(n12337) );
  XOR U13386 ( .A(n7523), .B(n12334), .Z(n12335) );
  XOR U13387 ( .A(n12338), .B(n12339), .Z(n12334) );
  ANDN U13388 ( .B(n12340), .A(n7529), .Z(n12338) );
  XNOR U13389 ( .A(n12341), .B(n12342), .Z(n7529) );
  IV U13390 ( .A(n12339), .Z(n12342) );
  XOR U13391 ( .A(n7528), .B(n12339), .Z(n12340) );
  XOR U13392 ( .A(n12343), .B(n12344), .Z(n12339) );
  ANDN U13393 ( .B(n12345), .A(n7544), .Z(n12343) );
  XNOR U13394 ( .A(n12346), .B(n12347), .Z(n7544) );
  IV U13395 ( .A(n12344), .Z(n12347) );
  XOR U13396 ( .A(n7543), .B(n12344), .Z(n12345) );
  XOR U13397 ( .A(n12348), .B(n12349), .Z(n12344) );
  ANDN U13398 ( .B(n12350), .A(n7549), .Z(n12348) );
  XNOR U13399 ( .A(n12351), .B(n12352), .Z(n7549) );
  IV U13400 ( .A(n12349), .Z(n12352) );
  XOR U13401 ( .A(n7548), .B(n12349), .Z(n12350) );
  XOR U13402 ( .A(n12353), .B(n12354), .Z(n12349) );
  ANDN U13403 ( .B(n12355), .A(n7554), .Z(n12353) );
  XNOR U13404 ( .A(n12356), .B(n12357), .Z(n7554) );
  IV U13405 ( .A(n12354), .Z(n12357) );
  XOR U13406 ( .A(n7553), .B(n12354), .Z(n12355) );
  XOR U13407 ( .A(n12358), .B(n12359), .Z(n12354) );
  ANDN U13408 ( .B(n12360), .A(n7559), .Z(n12358) );
  XNOR U13409 ( .A(n12361), .B(n12362), .Z(n7559) );
  IV U13410 ( .A(n12359), .Z(n12362) );
  XOR U13411 ( .A(n7558), .B(n12359), .Z(n12360) );
  XOR U13412 ( .A(n12363), .B(n12364), .Z(n12359) );
  ANDN U13413 ( .B(n12365), .A(n7564), .Z(n12363) );
  XNOR U13414 ( .A(n12366), .B(n12367), .Z(n7564) );
  IV U13415 ( .A(n12364), .Z(n12367) );
  XOR U13416 ( .A(n7563), .B(n12364), .Z(n12365) );
  XOR U13417 ( .A(n12368), .B(n12369), .Z(n12364) );
  ANDN U13418 ( .B(n12370), .A(n7569), .Z(n12368) );
  XNOR U13419 ( .A(n12371), .B(n12372), .Z(n7569) );
  IV U13420 ( .A(n12369), .Z(n12372) );
  XOR U13421 ( .A(n7568), .B(n12369), .Z(n12370) );
  XOR U13422 ( .A(n12373), .B(n12374), .Z(n12369) );
  ANDN U13423 ( .B(n12375), .A(n7574), .Z(n12373) );
  XNOR U13424 ( .A(n12376), .B(n12377), .Z(n7574) );
  IV U13425 ( .A(n12374), .Z(n12377) );
  XOR U13426 ( .A(n7573), .B(n12374), .Z(n12375) );
  XOR U13427 ( .A(n12378), .B(n12379), .Z(n12374) );
  ANDN U13428 ( .B(n12380), .A(n7579), .Z(n12378) );
  XNOR U13429 ( .A(n12381), .B(n12382), .Z(n7579) );
  IV U13430 ( .A(n12379), .Z(n12382) );
  XOR U13431 ( .A(n7578), .B(n12379), .Z(n12380) );
  XOR U13432 ( .A(n12383), .B(n12384), .Z(n12379) );
  ANDN U13433 ( .B(n12385), .A(n7584), .Z(n12383) );
  XNOR U13434 ( .A(n12386), .B(n12387), .Z(n7584) );
  IV U13435 ( .A(n12384), .Z(n12387) );
  XOR U13436 ( .A(n7583), .B(n12384), .Z(n12385) );
  XOR U13437 ( .A(n12388), .B(n12389), .Z(n12384) );
  ANDN U13438 ( .B(n12390), .A(n7589), .Z(n12388) );
  XNOR U13439 ( .A(n12391), .B(n12392), .Z(n7589) );
  IV U13440 ( .A(n12389), .Z(n12392) );
  XOR U13441 ( .A(n7588), .B(n12389), .Z(n12390) );
  XOR U13442 ( .A(n12393), .B(n12394), .Z(n12389) );
  ANDN U13443 ( .B(n12395), .A(n7599), .Z(n12393) );
  XNOR U13444 ( .A(n12396), .B(n12397), .Z(n7599) );
  IV U13445 ( .A(n12394), .Z(n12397) );
  XOR U13446 ( .A(n7598), .B(n12394), .Z(n12395) );
  XOR U13447 ( .A(n12398), .B(n12399), .Z(n12394) );
  ANDN U13448 ( .B(n12400), .A(n7604), .Z(n12398) );
  XNOR U13449 ( .A(n12401), .B(n12402), .Z(n7604) );
  IV U13450 ( .A(n12399), .Z(n12402) );
  XOR U13451 ( .A(n7603), .B(n12399), .Z(n12400) );
  XOR U13452 ( .A(n12403), .B(n12404), .Z(n12399) );
  ANDN U13453 ( .B(n12405), .A(n7609), .Z(n12403) );
  XNOR U13454 ( .A(n12406), .B(n12407), .Z(n7609) );
  IV U13455 ( .A(n12404), .Z(n12407) );
  XOR U13456 ( .A(n7608), .B(n12404), .Z(n12405) );
  XOR U13457 ( .A(n12408), .B(n12409), .Z(n12404) );
  ANDN U13458 ( .B(n12410), .A(n7614), .Z(n12408) );
  XNOR U13459 ( .A(n12411), .B(n12412), .Z(n7614) );
  IV U13460 ( .A(n12409), .Z(n12412) );
  XOR U13461 ( .A(n7613), .B(n12409), .Z(n12410) );
  XOR U13462 ( .A(n12413), .B(n12414), .Z(n12409) );
  ANDN U13463 ( .B(n12415), .A(n7619), .Z(n12413) );
  XNOR U13464 ( .A(n12416), .B(n12417), .Z(n7619) );
  IV U13465 ( .A(n12414), .Z(n12417) );
  XOR U13466 ( .A(n7618), .B(n12414), .Z(n12415) );
  XOR U13467 ( .A(n12418), .B(n12419), .Z(n12414) );
  ANDN U13468 ( .B(n12420), .A(n7624), .Z(n12418) );
  XNOR U13469 ( .A(n12421), .B(n12422), .Z(n7624) );
  IV U13470 ( .A(n12419), .Z(n12422) );
  XOR U13471 ( .A(n7623), .B(n12419), .Z(n12420) );
  XOR U13472 ( .A(n12423), .B(n12424), .Z(n12419) );
  ANDN U13473 ( .B(n12425), .A(n7629), .Z(n12423) );
  XNOR U13474 ( .A(n12426), .B(n12427), .Z(n7629) );
  IV U13475 ( .A(n12424), .Z(n12427) );
  XOR U13476 ( .A(n7628), .B(n12424), .Z(n12425) );
  XOR U13477 ( .A(n12428), .B(n12429), .Z(n12424) );
  ANDN U13478 ( .B(n12430), .A(n7634), .Z(n12428) );
  XNOR U13479 ( .A(n12431), .B(n12432), .Z(n7634) );
  IV U13480 ( .A(n12429), .Z(n12432) );
  XOR U13481 ( .A(n7633), .B(n12429), .Z(n12430) );
  XOR U13482 ( .A(n12433), .B(n12434), .Z(n12429) );
  ANDN U13483 ( .B(n12435), .A(n7639), .Z(n12433) );
  XNOR U13484 ( .A(n12436), .B(n12437), .Z(n7639) );
  IV U13485 ( .A(n12434), .Z(n12437) );
  XOR U13486 ( .A(n7638), .B(n12434), .Z(n12435) );
  XOR U13487 ( .A(n12438), .B(n12439), .Z(n12434) );
  ANDN U13488 ( .B(n12440), .A(n7644), .Z(n12438) );
  XNOR U13489 ( .A(n12441), .B(n12442), .Z(n7644) );
  IV U13490 ( .A(n12439), .Z(n12442) );
  XOR U13491 ( .A(n7643), .B(n12439), .Z(n12440) );
  XOR U13492 ( .A(n12443), .B(n12444), .Z(n12439) );
  ANDN U13493 ( .B(n12445), .A(n7654), .Z(n12443) );
  XNOR U13494 ( .A(n12446), .B(n12447), .Z(n7654) );
  IV U13495 ( .A(n12444), .Z(n12447) );
  XOR U13496 ( .A(n7653), .B(n12444), .Z(n12445) );
  XOR U13497 ( .A(n12448), .B(n12449), .Z(n12444) );
  ANDN U13498 ( .B(n12450), .A(n7659), .Z(n12448) );
  XNOR U13499 ( .A(n12451), .B(n12452), .Z(n7659) );
  IV U13500 ( .A(n12449), .Z(n12452) );
  XOR U13501 ( .A(n7658), .B(n12449), .Z(n12450) );
  XOR U13502 ( .A(n12453), .B(n12454), .Z(n12449) );
  ANDN U13503 ( .B(n12455), .A(n7664), .Z(n12453) );
  XNOR U13504 ( .A(n12456), .B(n12457), .Z(n7664) );
  IV U13505 ( .A(n12454), .Z(n12457) );
  XOR U13506 ( .A(n7663), .B(n12454), .Z(n12455) );
  XOR U13507 ( .A(n12458), .B(n12459), .Z(n12454) );
  ANDN U13508 ( .B(n12460), .A(n7669), .Z(n12458) );
  XNOR U13509 ( .A(n12461), .B(n12462), .Z(n7669) );
  IV U13510 ( .A(n12459), .Z(n12462) );
  XOR U13511 ( .A(n7668), .B(n12459), .Z(n12460) );
  XOR U13512 ( .A(n12463), .B(n12464), .Z(n12459) );
  ANDN U13513 ( .B(n12465), .A(n7674), .Z(n12463) );
  XNOR U13514 ( .A(n12466), .B(n12467), .Z(n7674) );
  IV U13515 ( .A(n12464), .Z(n12467) );
  XOR U13516 ( .A(n7673), .B(n12464), .Z(n12465) );
  XOR U13517 ( .A(n12468), .B(n12469), .Z(n12464) );
  ANDN U13518 ( .B(n12470), .A(n7679), .Z(n12468) );
  XNOR U13519 ( .A(n12471), .B(n12472), .Z(n7679) );
  IV U13520 ( .A(n12469), .Z(n12472) );
  XOR U13521 ( .A(n7678), .B(n12469), .Z(n12470) );
  XOR U13522 ( .A(n12473), .B(n12474), .Z(n12469) );
  ANDN U13523 ( .B(n12475), .A(n7684), .Z(n12473) );
  XNOR U13524 ( .A(n12476), .B(n12477), .Z(n7684) );
  IV U13525 ( .A(n12474), .Z(n12477) );
  XOR U13526 ( .A(n7683), .B(n12474), .Z(n12475) );
  XOR U13527 ( .A(n12478), .B(n12479), .Z(n12474) );
  ANDN U13528 ( .B(n12480), .A(n7689), .Z(n12478) );
  XNOR U13529 ( .A(n12481), .B(n12482), .Z(n7689) );
  IV U13530 ( .A(n12479), .Z(n12482) );
  XOR U13531 ( .A(n7688), .B(n12479), .Z(n12480) );
  XOR U13532 ( .A(n12483), .B(n12484), .Z(n12479) );
  ANDN U13533 ( .B(n12485), .A(n7694), .Z(n12483) );
  XNOR U13534 ( .A(n12486), .B(n12487), .Z(n7694) );
  IV U13535 ( .A(n12484), .Z(n12487) );
  XOR U13536 ( .A(n7693), .B(n12484), .Z(n12485) );
  XOR U13537 ( .A(n12488), .B(n12489), .Z(n12484) );
  ANDN U13538 ( .B(n12490), .A(n7699), .Z(n12488) );
  XNOR U13539 ( .A(n12491), .B(n12492), .Z(n7699) );
  IV U13540 ( .A(n12489), .Z(n12492) );
  XOR U13541 ( .A(n7698), .B(n12489), .Z(n12490) );
  XOR U13542 ( .A(n12493), .B(n12494), .Z(n12489) );
  ANDN U13543 ( .B(n12495), .A(n7709), .Z(n12493) );
  XNOR U13544 ( .A(n12496), .B(n12497), .Z(n7709) );
  IV U13545 ( .A(n12494), .Z(n12497) );
  XOR U13546 ( .A(n7708), .B(n12494), .Z(n12495) );
  XOR U13547 ( .A(n12498), .B(n12499), .Z(n12494) );
  ANDN U13548 ( .B(n12500), .A(n7714), .Z(n12498) );
  XNOR U13549 ( .A(n12501), .B(n12502), .Z(n7714) );
  IV U13550 ( .A(n12499), .Z(n12502) );
  XOR U13551 ( .A(n7713), .B(n12499), .Z(n12500) );
  XOR U13552 ( .A(n12503), .B(n12504), .Z(n12499) );
  ANDN U13553 ( .B(n12505), .A(n7719), .Z(n12503) );
  XNOR U13554 ( .A(n12506), .B(n12507), .Z(n7719) );
  IV U13555 ( .A(n12504), .Z(n12507) );
  XOR U13556 ( .A(n7718), .B(n12504), .Z(n12505) );
  XOR U13557 ( .A(n12508), .B(n12509), .Z(n12504) );
  ANDN U13558 ( .B(n12510), .A(n7724), .Z(n12508) );
  XNOR U13559 ( .A(n12511), .B(n12512), .Z(n7724) );
  IV U13560 ( .A(n12509), .Z(n12512) );
  XOR U13561 ( .A(n7723), .B(n12509), .Z(n12510) );
  XOR U13562 ( .A(n12513), .B(n12514), .Z(n12509) );
  ANDN U13563 ( .B(n12515), .A(n7729), .Z(n12513) );
  XNOR U13564 ( .A(n12516), .B(n12517), .Z(n7729) );
  IV U13565 ( .A(n12514), .Z(n12517) );
  XOR U13566 ( .A(n7728), .B(n12514), .Z(n12515) );
  XOR U13567 ( .A(n12518), .B(n12519), .Z(n12514) );
  ANDN U13568 ( .B(n12520), .A(n7734), .Z(n12518) );
  XNOR U13569 ( .A(n12521), .B(n12522), .Z(n7734) );
  IV U13570 ( .A(n12519), .Z(n12522) );
  XOR U13571 ( .A(n7733), .B(n12519), .Z(n12520) );
  XOR U13572 ( .A(n12523), .B(n12524), .Z(n12519) );
  ANDN U13573 ( .B(n12525), .A(n7739), .Z(n12523) );
  XNOR U13574 ( .A(n12526), .B(n12527), .Z(n7739) );
  IV U13575 ( .A(n12524), .Z(n12527) );
  XOR U13576 ( .A(n7738), .B(n12524), .Z(n12525) );
  XOR U13577 ( .A(n12528), .B(n12529), .Z(n12524) );
  ANDN U13578 ( .B(n12530), .A(n7744), .Z(n12528) );
  XNOR U13579 ( .A(n12531), .B(n12532), .Z(n7744) );
  IV U13580 ( .A(n12529), .Z(n12532) );
  XOR U13581 ( .A(n7743), .B(n12529), .Z(n12530) );
  XOR U13582 ( .A(n12533), .B(n12534), .Z(n12529) );
  ANDN U13583 ( .B(n12535), .A(n7749), .Z(n12533) );
  XNOR U13584 ( .A(n12536), .B(n12537), .Z(n7749) );
  IV U13585 ( .A(n12534), .Z(n12537) );
  XOR U13586 ( .A(n7748), .B(n12534), .Z(n12535) );
  XOR U13587 ( .A(n12538), .B(n12539), .Z(n12534) );
  ANDN U13588 ( .B(n12540), .A(n7754), .Z(n12538) );
  XNOR U13589 ( .A(n12541), .B(n12542), .Z(n7754) );
  IV U13590 ( .A(n12539), .Z(n12542) );
  XOR U13591 ( .A(n7753), .B(n12539), .Z(n12540) );
  XOR U13592 ( .A(n12543), .B(n12544), .Z(n12539) );
  ANDN U13593 ( .B(n12545), .A(n7764), .Z(n12543) );
  XNOR U13594 ( .A(n12546), .B(n12547), .Z(n7764) );
  IV U13595 ( .A(n12544), .Z(n12547) );
  XOR U13596 ( .A(n7763), .B(n12544), .Z(n12545) );
  XOR U13597 ( .A(n12548), .B(n12549), .Z(n12544) );
  ANDN U13598 ( .B(n12550), .A(n7769), .Z(n12548) );
  XNOR U13599 ( .A(n12551), .B(n12552), .Z(n7769) );
  IV U13600 ( .A(n12549), .Z(n12552) );
  XOR U13601 ( .A(n7768), .B(n12549), .Z(n12550) );
  XOR U13602 ( .A(n12553), .B(n12554), .Z(n12549) );
  ANDN U13603 ( .B(n12555), .A(n7774), .Z(n12553) );
  XNOR U13604 ( .A(n12556), .B(n12557), .Z(n7774) );
  IV U13605 ( .A(n12554), .Z(n12557) );
  XOR U13606 ( .A(n7773), .B(n12554), .Z(n12555) );
  XOR U13607 ( .A(n12558), .B(n12559), .Z(n12554) );
  ANDN U13608 ( .B(n12560), .A(n7779), .Z(n12558) );
  XNOR U13609 ( .A(n12561), .B(n12562), .Z(n7779) );
  IV U13610 ( .A(n12559), .Z(n12562) );
  XOR U13611 ( .A(n7778), .B(n12559), .Z(n12560) );
  XOR U13612 ( .A(n12563), .B(n12564), .Z(n12559) );
  ANDN U13613 ( .B(n12565), .A(n7784), .Z(n12563) );
  XNOR U13614 ( .A(n12566), .B(n12567), .Z(n7784) );
  IV U13615 ( .A(n12564), .Z(n12567) );
  XOR U13616 ( .A(n7783), .B(n12564), .Z(n12565) );
  XOR U13617 ( .A(n12568), .B(n12569), .Z(n12564) );
  ANDN U13618 ( .B(n12570), .A(n7789), .Z(n12568) );
  XNOR U13619 ( .A(n12571), .B(n12572), .Z(n7789) );
  IV U13620 ( .A(n12569), .Z(n12572) );
  XOR U13621 ( .A(n7788), .B(n12569), .Z(n12570) );
  XOR U13622 ( .A(n12573), .B(n12574), .Z(n12569) );
  ANDN U13623 ( .B(n12575), .A(n7794), .Z(n12573) );
  XNOR U13624 ( .A(n12576), .B(n12577), .Z(n7794) );
  IV U13625 ( .A(n12574), .Z(n12577) );
  XOR U13626 ( .A(n7793), .B(n12574), .Z(n12575) );
  XOR U13627 ( .A(n12578), .B(n12579), .Z(n12574) );
  ANDN U13628 ( .B(n12580), .A(n7799), .Z(n12578) );
  XNOR U13629 ( .A(n12581), .B(n12582), .Z(n7799) );
  IV U13630 ( .A(n12579), .Z(n12582) );
  XOR U13631 ( .A(n7798), .B(n12579), .Z(n12580) );
  XOR U13632 ( .A(n12583), .B(n12584), .Z(n12579) );
  ANDN U13633 ( .B(n12585), .A(n7804), .Z(n12583) );
  XNOR U13634 ( .A(n12586), .B(n12587), .Z(n7804) );
  IV U13635 ( .A(n12584), .Z(n12587) );
  XOR U13636 ( .A(n7803), .B(n12584), .Z(n12585) );
  XOR U13637 ( .A(n12588), .B(n12589), .Z(n12584) );
  ANDN U13638 ( .B(n12590), .A(n7809), .Z(n12588) );
  XNOR U13639 ( .A(n12591), .B(n12592), .Z(n7809) );
  IV U13640 ( .A(n12589), .Z(n12592) );
  XOR U13641 ( .A(n7808), .B(n12589), .Z(n12590) );
  XOR U13642 ( .A(n12593), .B(n12594), .Z(n12589) );
  ANDN U13643 ( .B(n12595), .A(n7819), .Z(n12593) );
  XNOR U13644 ( .A(n12596), .B(n12597), .Z(n7819) );
  IV U13645 ( .A(n12594), .Z(n12597) );
  XOR U13646 ( .A(n7818), .B(n12594), .Z(n12595) );
  XOR U13647 ( .A(n12598), .B(n12599), .Z(n12594) );
  ANDN U13648 ( .B(n12600), .A(n7824), .Z(n12598) );
  XNOR U13649 ( .A(n12601), .B(n12602), .Z(n7824) );
  IV U13650 ( .A(n12599), .Z(n12602) );
  XOR U13651 ( .A(n7823), .B(n12599), .Z(n12600) );
  XOR U13652 ( .A(n12603), .B(n12604), .Z(n12599) );
  ANDN U13653 ( .B(n12605), .A(n7829), .Z(n12603) );
  XNOR U13654 ( .A(n12606), .B(n12607), .Z(n7829) );
  IV U13655 ( .A(n12604), .Z(n12607) );
  XOR U13656 ( .A(n7828), .B(n12604), .Z(n12605) );
  XOR U13657 ( .A(n12608), .B(n12609), .Z(n12604) );
  ANDN U13658 ( .B(n12610), .A(n7834), .Z(n12608) );
  XNOR U13659 ( .A(n12611), .B(n12612), .Z(n7834) );
  IV U13660 ( .A(n12609), .Z(n12612) );
  XOR U13661 ( .A(n7833), .B(n12609), .Z(n12610) );
  XOR U13662 ( .A(n12613), .B(n12614), .Z(n12609) );
  ANDN U13663 ( .B(n12615), .A(n7839), .Z(n12613) );
  XNOR U13664 ( .A(n12616), .B(n12617), .Z(n7839) );
  IV U13665 ( .A(n12614), .Z(n12617) );
  XOR U13666 ( .A(n7838), .B(n12614), .Z(n12615) );
  XOR U13667 ( .A(n12618), .B(n12619), .Z(n12614) );
  ANDN U13668 ( .B(n12620), .A(n7844), .Z(n12618) );
  XNOR U13669 ( .A(n12621), .B(n12622), .Z(n7844) );
  IV U13670 ( .A(n12619), .Z(n12622) );
  XOR U13671 ( .A(n7843), .B(n12619), .Z(n12620) );
  XOR U13672 ( .A(n12623), .B(n12624), .Z(n12619) );
  ANDN U13673 ( .B(n12625), .A(n7849), .Z(n12623) );
  XNOR U13674 ( .A(n12626), .B(n12627), .Z(n7849) );
  IV U13675 ( .A(n12624), .Z(n12627) );
  XOR U13676 ( .A(n7848), .B(n12624), .Z(n12625) );
  XOR U13677 ( .A(n12628), .B(n12629), .Z(n12624) );
  ANDN U13678 ( .B(n12630), .A(n7854), .Z(n12628) );
  XNOR U13679 ( .A(n12631), .B(n12632), .Z(n7854) );
  IV U13680 ( .A(n12629), .Z(n12632) );
  XOR U13681 ( .A(n7853), .B(n12629), .Z(n12630) );
  XOR U13682 ( .A(n12633), .B(n12634), .Z(n12629) );
  ANDN U13683 ( .B(n12635), .A(n7859), .Z(n12633) );
  XNOR U13684 ( .A(n12636), .B(n12637), .Z(n7859) );
  IV U13685 ( .A(n12634), .Z(n12637) );
  XOR U13686 ( .A(n7858), .B(n12634), .Z(n12635) );
  XOR U13687 ( .A(n12638), .B(n12639), .Z(n12634) );
  ANDN U13688 ( .B(n12640), .A(n7864), .Z(n12638) );
  XNOR U13689 ( .A(n12641), .B(n12642), .Z(n7864) );
  IV U13690 ( .A(n12639), .Z(n12642) );
  XOR U13691 ( .A(n7863), .B(n12639), .Z(n12640) );
  XOR U13692 ( .A(n12643), .B(n12644), .Z(n12639) );
  ANDN U13693 ( .B(n12645), .A(n7874), .Z(n12643) );
  XNOR U13694 ( .A(n12646), .B(n12647), .Z(n7874) );
  IV U13695 ( .A(n12644), .Z(n12647) );
  XOR U13696 ( .A(n7873), .B(n12644), .Z(n12645) );
  XOR U13697 ( .A(n12648), .B(n12649), .Z(n12644) );
  ANDN U13698 ( .B(n12650), .A(n7879), .Z(n12648) );
  XNOR U13699 ( .A(n12651), .B(n12652), .Z(n7879) );
  IV U13700 ( .A(n12649), .Z(n12652) );
  XOR U13701 ( .A(n7878), .B(n12649), .Z(n12650) );
  XOR U13702 ( .A(n12653), .B(n12654), .Z(n12649) );
  ANDN U13703 ( .B(n12655), .A(n7884), .Z(n12653) );
  XNOR U13704 ( .A(n12656), .B(n12657), .Z(n7884) );
  IV U13705 ( .A(n12654), .Z(n12657) );
  XOR U13706 ( .A(n7883), .B(n12654), .Z(n12655) );
  XOR U13707 ( .A(n12658), .B(n12659), .Z(n12654) );
  ANDN U13708 ( .B(n12660), .A(n7889), .Z(n12658) );
  XNOR U13709 ( .A(n12661), .B(n12662), .Z(n7889) );
  IV U13710 ( .A(n12659), .Z(n12662) );
  XOR U13711 ( .A(n7888), .B(n12659), .Z(n12660) );
  XOR U13712 ( .A(n12663), .B(n12664), .Z(n12659) );
  ANDN U13713 ( .B(n12665), .A(n7894), .Z(n12663) );
  XNOR U13714 ( .A(n12666), .B(n12667), .Z(n7894) );
  IV U13715 ( .A(n12664), .Z(n12667) );
  XOR U13716 ( .A(n7893), .B(n12664), .Z(n12665) );
  XOR U13717 ( .A(n12668), .B(n12669), .Z(n12664) );
  ANDN U13718 ( .B(n12670), .A(n7899), .Z(n12668) );
  XNOR U13719 ( .A(n12671), .B(n12672), .Z(n7899) );
  IV U13720 ( .A(n12669), .Z(n12672) );
  XOR U13721 ( .A(n7898), .B(n12669), .Z(n12670) );
  XOR U13722 ( .A(n12673), .B(n12674), .Z(n12669) );
  ANDN U13723 ( .B(n12675), .A(n7904), .Z(n12673) );
  XNOR U13724 ( .A(n12676), .B(n12677), .Z(n7904) );
  IV U13725 ( .A(n12674), .Z(n12677) );
  XOR U13726 ( .A(n7903), .B(n12674), .Z(n12675) );
  XOR U13727 ( .A(n12678), .B(n12679), .Z(n12674) );
  ANDN U13728 ( .B(n12680), .A(n7909), .Z(n12678) );
  XNOR U13729 ( .A(n12681), .B(n12682), .Z(n7909) );
  IV U13730 ( .A(n12679), .Z(n12682) );
  XOR U13731 ( .A(n7908), .B(n12679), .Z(n12680) );
  XOR U13732 ( .A(n12683), .B(n12684), .Z(n12679) );
  ANDN U13733 ( .B(n12685), .A(n7914), .Z(n12683) );
  XNOR U13734 ( .A(n12686), .B(n12687), .Z(n7914) );
  IV U13735 ( .A(n12684), .Z(n12687) );
  XOR U13736 ( .A(n7913), .B(n12684), .Z(n12685) );
  XOR U13737 ( .A(n12688), .B(n12689), .Z(n12684) );
  ANDN U13738 ( .B(n12690), .A(n7919), .Z(n12688) );
  XNOR U13739 ( .A(n12691), .B(n12692), .Z(n7919) );
  IV U13740 ( .A(n12689), .Z(n12692) );
  XOR U13741 ( .A(n7918), .B(n12689), .Z(n12690) );
  XOR U13742 ( .A(n12693), .B(n12694), .Z(n12689) );
  ANDN U13743 ( .B(n12695), .A(n7929), .Z(n12693) );
  XNOR U13744 ( .A(n12696), .B(n12697), .Z(n7929) );
  IV U13745 ( .A(n12694), .Z(n12697) );
  XOR U13746 ( .A(n7928), .B(n12694), .Z(n12695) );
  XOR U13747 ( .A(n12698), .B(n12699), .Z(n12694) );
  ANDN U13748 ( .B(n12700), .A(n7934), .Z(n12698) );
  XNOR U13749 ( .A(n12701), .B(n12702), .Z(n7934) );
  IV U13750 ( .A(n12699), .Z(n12702) );
  XOR U13751 ( .A(n7933), .B(n12699), .Z(n12700) );
  XOR U13752 ( .A(n12703), .B(n12704), .Z(n12699) );
  ANDN U13753 ( .B(n12705), .A(n7939), .Z(n12703) );
  XNOR U13754 ( .A(n12706), .B(n12707), .Z(n7939) );
  IV U13755 ( .A(n12704), .Z(n12707) );
  XOR U13756 ( .A(n7938), .B(n12704), .Z(n12705) );
  XOR U13757 ( .A(n12708), .B(n12709), .Z(n12704) );
  ANDN U13758 ( .B(n12710), .A(n7944), .Z(n12708) );
  XNOR U13759 ( .A(n12711), .B(n12712), .Z(n7944) );
  IV U13760 ( .A(n12709), .Z(n12712) );
  XOR U13761 ( .A(n7943), .B(n12709), .Z(n12710) );
  XOR U13762 ( .A(n12713), .B(n12714), .Z(n12709) );
  ANDN U13763 ( .B(n12715), .A(n7949), .Z(n12713) );
  XNOR U13764 ( .A(n12716), .B(n12717), .Z(n7949) );
  IV U13765 ( .A(n12714), .Z(n12717) );
  XOR U13766 ( .A(n7948), .B(n12714), .Z(n12715) );
  XOR U13767 ( .A(n12718), .B(n12719), .Z(n12714) );
  ANDN U13768 ( .B(n12720), .A(n7954), .Z(n12718) );
  XNOR U13769 ( .A(n12721), .B(n12722), .Z(n7954) );
  IV U13770 ( .A(n12719), .Z(n12722) );
  XOR U13771 ( .A(n7953), .B(n12719), .Z(n12720) );
  XOR U13772 ( .A(n12723), .B(n12724), .Z(n12719) );
  ANDN U13773 ( .B(n12725), .A(n7959), .Z(n12723) );
  XNOR U13774 ( .A(n12726), .B(n12727), .Z(n7959) );
  IV U13775 ( .A(n12724), .Z(n12727) );
  XOR U13776 ( .A(n7958), .B(n12724), .Z(n12725) );
  XOR U13777 ( .A(n12728), .B(n12729), .Z(n12724) );
  ANDN U13778 ( .B(n12730), .A(n7964), .Z(n12728) );
  XNOR U13779 ( .A(n12731), .B(n12732), .Z(n7964) );
  IV U13780 ( .A(n12729), .Z(n12732) );
  XOR U13781 ( .A(n7963), .B(n12729), .Z(n12730) );
  XOR U13782 ( .A(n12733), .B(n12734), .Z(n12729) );
  ANDN U13783 ( .B(n12735), .A(n7969), .Z(n12733) );
  XNOR U13784 ( .A(n12736), .B(n12737), .Z(n7969) );
  IV U13785 ( .A(n12734), .Z(n12737) );
  XOR U13786 ( .A(n7968), .B(n12734), .Z(n12735) );
  XOR U13787 ( .A(n12738), .B(n12739), .Z(n12734) );
  ANDN U13788 ( .B(n12740), .A(n7974), .Z(n12738) );
  XNOR U13789 ( .A(n12741), .B(n12742), .Z(n7974) );
  IV U13790 ( .A(n12739), .Z(n12742) );
  XOR U13791 ( .A(n7973), .B(n12739), .Z(n12740) );
  XOR U13792 ( .A(n12743), .B(n12744), .Z(n12739) );
  ANDN U13793 ( .B(n12745), .A(n7984), .Z(n12743) );
  XNOR U13794 ( .A(n12746), .B(n12747), .Z(n7984) );
  IV U13795 ( .A(n12744), .Z(n12747) );
  XOR U13796 ( .A(n7983), .B(n12744), .Z(n12745) );
  XOR U13797 ( .A(n12748), .B(n12749), .Z(n12744) );
  ANDN U13798 ( .B(n12750), .A(n7989), .Z(n12748) );
  XNOR U13799 ( .A(n12751), .B(n12752), .Z(n7989) );
  IV U13800 ( .A(n12749), .Z(n12752) );
  XOR U13801 ( .A(n7988), .B(n12749), .Z(n12750) );
  XOR U13802 ( .A(n12753), .B(n12754), .Z(n12749) );
  ANDN U13803 ( .B(n12755), .A(n7994), .Z(n12753) );
  XNOR U13804 ( .A(n12756), .B(n12757), .Z(n7994) );
  IV U13805 ( .A(n12754), .Z(n12757) );
  XOR U13806 ( .A(n7993), .B(n12754), .Z(n12755) );
  XOR U13807 ( .A(n12758), .B(n12759), .Z(n12754) );
  ANDN U13808 ( .B(n12760), .A(n7999), .Z(n12758) );
  XNOR U13809 ( .A(n12761), .B(n12762), .Z(n7999) );
  IV U13810 ( .A(n12759), .Z(n12762) );
  XOR U13811 ( .A(n7998), .B(n12759), .Z(n12760) );
  XOR U13812 ( .A(n12763), .B(n12764), .Z(n12759) );
  ANDN U13813 ( .B(n12765), .A(n8004), .Z(n12763) );
  XNOR U13814 ( .A(n12766), .B(n12767), .Z(n8004) );
  IV U13815 ( .A(n12764), .Z(n12767) );
  XOR U13816 ( .A(n8003), .B(n12764), .Z(n12765) );
  XOR U13817 ( .A(n12768), .B(n12769), .Z(n12764) );
  ANDN U13818 ( .B(n12770), .A(n8009), .Z(n12768) );
  XNOR U13819 ( .A(n12771), .B(n12772), .Z(n8009) );
  IV U13820 ( .A(n12769), .Z(n12772) );
  XOR U13821 ( .A(n8008), .B(n12769), .Z(n12770) );
  XOR U13822 ( .A(n12773), .B(n12774), .Z(n12769) );
  ANDN U13823 ( .B(n12775), .A(n8014), .Z(n12773) );
  XNOR U13824 ( .A(n12776), .B(n12777), .Z(n8014) );
  IV U13825 ( .A(n12774), .Z(n12777) );
  XOR U13826 ( .A(n8013), .B(n12774), .Z(n12775) );
  XOR U13827 ( .A(n12778), .B(n12779), .Z(n12774) );
  ANDN U13828 ( .B(n12780), .A(n8019), .Z(n12778) );
  XNOR U13829 ( .A(n12781), .B(n12782), .Z(n8019) );
  IV U13830 ( .A(n12779), .Z(n12782) );
  XOR U13831 ( .A(n8018), .B(n12779), .Z(n12780) );
  XOR U13832 ( .A(n12783), .B(n12784), .Z(n12779) );
  ANDN U13833 ( .B(n12785), .A(n8024), .Z(n12783) );
  XNOR U13834 ( .A(n12786), .B(n12787), .Z(n8024) );
  IV U13835 ( .A(n12784), .Z(n12787) );
  XOR U13836 ( .A(n8023), .B(n12784), .Z(n12785) );
  XOR U13837 ( .A(n12788), .B(n12789), .Z(n12784) );
  ANDN U13838 ( .B(n12790), .A(n8029), .Z(n12788) );
  XNOR U13839 ( .A(n12791), .B(n12792), .Z(n8029) );
  IV U13840 ( .A(n12789), .Z(n12792) );
  XOR U13841 ( .A(n8028), .B(n12789), .Z(n12790) );
  XOR U13842 ( .A(n12793), .B(n12794), .Z(n12789) );
  ANDN U13843 ( .B(n12795), .A(n8039), .Z(n12793) );
  XNOR U13844 ( .A(n12796), .B(n12797), .Z(n8039) );
  IV U13845 ( .A(n12794), .Z(n12797) );
  XOR U13846 ( .A(n8038), .B(n12794), .Z(n12795) );
  XOR U13847 ( .A(n12798), .B(n12799), .Z(n12794) );
  ANDN U13848 ( .B(n12800), .A(n8044), .Z(n12798) );
  XNOR U13849 ( .A(n12801), .B(n12802), .Z(n8044) );
  IV U13850 ( .A(n12799), .Z(n12802) );
  XOR U13851 ( .A(n8043), .B(n12799), .Z(n12800) );
  XOR U13852 ( .A(n12803), .B(n12804), .Z(n12799) );
  ANDN U13853 ( .B(n12805), .A(n8049), .Z(n12803) );
  XNOR U13854 ( .A(n12806), .B(n12807), .Z(n8049) );
  IV U13855 ( .A(n12804), .Z(n12807) );
  XOR U13856 ( .A(n8048), .B(n12804), .Z(n12805) );
  XOR U13857 ( .A(n12808), .B(n12809), .Z(n12804) );
  ANDN U13858 ( .B(n12810), .A(n8054), .Z(n12808) );
  XNOR U13859 ( .A(n12811), .B(n12812), .Z(n8054) );
  IV U13860 ( .A(n12809), .Z(n12812) );
  XOR U13861 ( .A(n8053), .B(n12809), .Z(n12810) );
  XOR U13862 ( .A(n12813), .B(n12814), .Z(n12809) );
  ANDN U13863 ( .B(n12815), .A(n8059), .Z(n12813) );
  XNOR U13864 ( .A(n12816), .B(n12817), .Z(n8059) );
  IV U13865 ( .A(n12814), .Z(n12817) );
  XOR U13866 ( .A(n8058), .B(n12814), .Z(n12815) );
  XOR U13867 ( .A(n12818), .B(n12819), .Z(n12814) );
  ANDN U13868 ( .B(n12820), .A(n8064), .Z(n12818) );
  XNOR U13869 ( .A(n12821), .B(n12822), .Z(n8064) );
  IV U13870 ( .A(n12819), .Z(n12822) );
  XOR U13871 ( .A(n8063), .B(n12819), .Z(n12820) );
  XOR U13872 ( .A(n12823), .B(n12824), .Z(n12819) );
  ANDN U13873 ( .B(n12825), .A(n8069), .Z(n12823) );
  XNOR U13874 ( .A(n12826), .B(n12827), .Z(n8069) );
  IV U13875 ( .A(n12824), .Z(n12827) );
  XOR U13876 ( .A(n8068), .B(n12824), .Z(n12825) );
  XOR U13877 ( .A(n12828), .B(n12829), .Z(n12824) );
  ANDN U13878 ( .B(n12830), .A(n8074), .Z(n12828) );
  XNOR U13879 ( .A(n12831), .B(n12832), .Z(n8074) );
  IV U13880 ( .A(n12829), .Z(n12832) );
  XOR U13881 ( .A(n8073), .B(n12829), .Z(n12830) );
  XOR U13882 ( .A(n12833), .B(n12834), .Z(n12829) );
  ANDN U13883 ( .B(n12835), .A(n8123), .Z(n12833) );
  XNOR U13884 ( .A(n12836), .B(n12837), .Z(n8123) );
  IV U13885 ( .A(n12834), .Z(n12837) );
  XOR U13886 ( .A(n8122), .B(n12834), .Z(n12835) );
  XOR U13887 ( .A(n12838), .B(n12839), .Z(n12834) );
  ANDN U13888 ( .B(n12840), .A(n8238), .Z(n12838) );
  XNOR U13889 ( .A(n12841), .B(n12842), .Z(n8238) );
  IV U13890 ( .A(n12839), .Z(n12842) );
  XOR U13891 ( .A(n8237), .B(n12839), .Z(n12840) );
  XOR U13892 ( .A(n12843), .B(n12844), .Z(n12839) );
  ANDN U13893 ( .B(n12845), .A(n3099), .Z(n12843) );
  XNOR U13894 ( .A(n12846), .B(n12847), .Z(n3099) );
  IV U13895 ( .A(n12844), .Z(n12847) );
  XOR U13896 ( .A(n3098), .B(n12844), .Z(n12845) );
  XOR U13897 ( .A(n12848), .B(n12849), .Z(n12844) );
  ANDN U13898 ( .B(n12850), .A(n3154), .Z(n12848) );
  XNOR U13899 ( .A(n12851), .B(n12852), .Z(n3154) );
  IV U13900 ( .A(n12849), .Z(n12852) );
  XOR U13901 ( .A(n3153), .B(n12849), .Z(n12850) );
  XOR U13902 ( .A(n12853), .B(n12854), .Z(n12849) );
  ANDN U13903 ( .B(n12855), .A(n3209), .Z(n12853) );
  XNOR U13904 ( .A(n12856), .B(n12857), .Z(n3209) );
  IV U13905 ( .A(n12854), .Z(n12857) );
  XOR U13906 ( .A(n3208), .B(n12854), .Z(n12855) );
  XOR U13907 ( .A(n12858), .B(n12859), .Z(n12854) );
  ANDN U13908 ( .B(n12860), .A(n3264), .Z(n12858) );
  XNOR U13909 ( .A(n12861), .B(n12862), .Z(n3264) );
  IV U13910 ( .A(n12859), .Z(n12862) );
  XOR U13911 ( .A(n3263), .B(n12859), .Z(n12860) );
  XOR U13912 ( .A(n12863), .B(n12864), .Z(n12859) );
  ANDN U13913 ( .B(n12865), .A(n3319), .Z(n12863) );
  XNOR U13914 ( .A(n12866), .B(n12867), .Z(n3319) );
  IV U13915 ( .A(n12864), .Z(n12867) );
  XOR U13916 ( .A(n3318), .B(n12864), .Z(n12865) );
  XOR U13917 ( .A(n12868), .B(n12869), .Z(n12864) );
  ANDN U13918 ( .B(n12870), .A(n3374), .Z(n12868) );
  XNOR U13919 ( .A(n12871), .B(n12872), .Z(n3374) );
  IV U13920 ( .A(n12869), .Z(n12872) );
  XOR U13921 ( .A(n3373), .B(n12869), .Z(n12870) );
  XOR U13922 ( .A(n12873), .B(n12874), .Z(n12869) );
  ANDN U13923 ( .B(n12875), .A(n3429), .Z(n12873) );
  XNOR U13924 ( .A(n12876), .B(n12877), .Z(n3429) );
  IV U13925 ( .A(n12874), .Z(n12877) );
  XOR U13926 ( .A(n3428), .B(n12874), .Z(n12875) );
  XOR U13927 ( .A(n12878), .B(n12879), .Z(n12874) );
  ANDN U13928 ( .B(n12880), .A(n3484), .Z(n12878) );
  XNOR U13929 ( .A(n12881), .B(n12882), .Z(n3484) );
  IV U13930 ( .A(n12879), .Z(n12882) );
  XOR U13931 ( .A(n3483), .B(n12879), .Z(n12880) );
  XOR U13932 ( .A(n12883), .B(n12884), .Z(n12879) );
  ANDN U13933 ( .B(n12885), .A(n3539), .Z(n12883) );
  XNOR U13934 ( .A(n12886), .B(n12887), .Z(n3539) );
  IV U13935 ( .A(n12884), .Z(n12887) );
  XOR U13936 ( .A(n3538), .B(n12884), .Z(n12885) );
  XOR U13937 ( .A(n12888), .B(n12889), .Z(n12884) );
  ANDN U13938 ( .B(n12890), .A(n3594), .Z(n12888) );
  XNOR U13939 ( .A(n12891), .B(n12892), .Z(n3594) );
  IV U13940 ( .A(n12889), .Z(n12892) );
  XOR U13941 ( .A(n3593), .B(n12889), .Z(n12890) );
  XOR U13942 ( .A(n12893), .B(n12894), .Z(n12889) );
  ANDN U13943 ( .B(n12895), .A(n3654), .Z(n12893) );
  XNOR U13944 ( .A(n12896), .B(n12897), .Z(n3654) );
  IV U13945 ( .A(n12894), .Z(n12897) );
  XOR U13946 ( .A(n3653), .B(n12894), .Z(n12895) );
  XOR U13947 ( .A(n12898), .B(n12899), .Z(n12894) );
  ANDN U13948 ( .B(n12900), .A(n3709), .Z(n12898) );
  XNOR U13949 ( .A(n12901), .B(n12902), .Z(n3709) );
  IV U13950 ( .A(n12899), .Z(n12902) );
  XOR U13951 ( .A(n3708), .B(n12899), .Z(n12900) );
  XOR U13952 ( .A(n12903), .B(n12904), .Z(n12899) );
  ANDN U13953 ( .B(n12905), .A(n3764), .Z(n12903) );
  XNOR U13954 ( .A(n12906), .B(n12907), .Z(n3764) );
  IV U13955 ( .A(n12904), .Z(n12907) );
  XOR U13956 ( .A(n3763), .B(n12904), .Z(n12905) );
  XOR U13957 ( .A(n12908), .B(n12909), .Z(n12904) );
  ANDN U13958 ( .B(n12910), .A(n3819), .Z(n12908) );
  XNOR U13959 ( .A(n12911), .B(n12912), .Z(n3819) );
  IV U13960 ( .A(n12909), .Z(n12912) );
  XOR U13961 ( .A(n3818), .B(n12909), .Z(n12910) );
  XOR U13962 ( .A(n12913), .B(n12914), .Z(n12909) );
  ANDN U13963 ( .B(n12915), .A(n3874), .Z(n12913) );
  XNOR U13964 ( .A(n12916), .B(n12917), .Z(n3874) );
  IV U13965 ( .A(n12914), .Z(n12917) );
  XOR U13966 ( .A(n3873), .B(n12914), .Z(n12915) );
  XOR U13967 ( .A(n12918), .B(n12919), .Z(n12914) );
  ANDN U13968 ( .B(n12920), .A(n3929), .Z(n12918) );
  XNOR U13969 ( .A(n12921), .B(n12922), .Z(n3929) );
  IV U13970 ( .A(n12919), .Z(n12922) );
  XOR U13971 ( .A(n3928), .B(n12919), .Z(n12920) );
  XOR U13972 ( .A(n12923), .B(n12924), .Z(n12919) );
  ANDN U13973 ( .B(n12925), .A(n3984), .Z(n12923) );
  XNOR U13974 ( .A(n12926), .B(n12927), .Z(n3984) );
  IV U13975 ( .A(n12924), .Z(n12927) );
  XOR U13976 ( .A(n3983), .B(n12924), .Z(n12925) );
  XOR U13977 ( .A(n12928), .B(n12929), .Z(n12924) );
  ANDN U13978 ( .B(n12930), .A(n4039), .Z(n12928) );
  XNOR U13979 ( .A(n12931), .B(n12932), .Z(n4039) );
  IV U13980 ( .A(n12929), .Z(n12932) );
  XOR U13981 ( .A(n4038), .B(n12929), .Z(n12930) );
  XOR U13982 ( .A(n12933), .B(n12934), .Z(n12929) );
  ANDN U13983 ( .B(n12935), .A(n4094), .Z(n12933) );
  XNOR U13984 ( .A(n12936), .B(n12937), .Z(n4094) );
  IV U13985 ( .A(n12934), .Z(n12937) );
  XOR U13986 ( .A(n4093), .B(n12934), .Z(n12935) );
  XOR U13987 ( .A(n12938), .B(n12939), .Z(n12934) );
  ANDN U13988 ( .B(n12940), .A(n4149), .Z(n12938) );
  XNOR U13989 ( .A(n12941), .B(n12942), .Z(n4149) );
  IV U13990 ( .A(n12939), .Z(n12942) );
  XOR U13991 ( .A(n4148), .B(n12939), .Z(n12940) );
  XOR U13992 ( .A(n12943), .B(n12944), .Z(n12939) );
  ANDN U13993 ( .B(n12945), .A(n4209), .Z(n12943) );
  XNOR U13994 ( .A(n12946), .B(n12947), .Z(n4209) );
  IV U13995 ( .A(n12944), .Z(n12947) );
  XOR U13996 ( .A(n4208), .B(n12944), .Z(n12945) );
  XOR U13997 ( .A(n12948), .B(n12949), .Z(n12944) );
  ANDN U13998 ( .B(n12950), .A(n4264), .Z(n12948) );
  XNOR U13999 ( .A(n12951), .B(n12952), .Z(n4264) );
  IV U14000 ( .A(n12949), .Z(n12952) );
  XOR U14001 ( .A(n4263), .B(n12949), .Z(n12950) );
  XOR U14002 ( .A(n12953), .B(n12954), .Z(n12949) );
  ANDN U14003 ( .B(n12955), .A(n4319), .Z(n12953) );
  XNOR U14004 ( .A(n12956), .B(n12957), .Z(n4319) );
  IV U14005 ( .A(n12954), .Z(n12957) );
  XOR U14006 ( .A(n4318), .B(n12954), .Z(n12955) );
  XOR U14007 ( .A(n12958), .B(n12959), .Z(n12954) );
  ANDN U14008 ( .B(n12960), .A(n4374), .Z(n12958) );
  XNOR U14009 ( .A(n12961), .B(n12962), .Z(n4374) );
  IV U14010 ( .A(n12959), .Z(n12962) );
  XOR U14011 ( .A(n4373), .B(n12959), .Z(n12960) );
  XOR U14012 ( .A(n12963), .B(n12964), .Z(n12959) );
  ANDN U14013 ( .B(n12965), .A(n4429), .Z(n12963) );
  XNOR U14014 ( .A(n12966), .B(n12967), .Z(n4429) );
  IV U14015 ( .A(n12964), .Z(n12967) );
  XOR U14016 ( .A(n4428), .B(n12964), .Z(n12965) );
  XOR U14017 ( .A(n12968), .B(n12969), .Z(n12964) );
  ANDN U14018 ( .B(n12970), .A(n4484), .Z(n12968) );
  XNOR U14019 ( .A(n12971), .B(n12972), .Z(n4484) );
  IV U14020 ( .A(n12969), .Z(n12972) );
  XOR U14021 ( .A(n4483), .B(n12969), .Z(n12970) );
  XOR U14022 ( .A(n12973), .B(n12974), .Z(n12969) );
  ANDN U14023 ( .B(n12975), .A(n4539), .Z(n12973) );
  XNOR U14024 ( .A(n12976), .B(n12977), .Z(n4539) );
  IV U14025 ( .A(n12974), .Z(n12977) );
  XOR U14026 ( .A(n4538), .B(n12974), .Z(n12975) );
  XOR U14027 ( .A(n12978), .B(n12979), .Z(n12974) );
  ANDN U14028 ( .B(n12980), .A(n4594), .Z(n12978) );
  XNOR U14029 ( .A(n12981), .B(n12982), .Z(n4594) );
  IV U14030 ( .A(n12979), .Z(n12982) );
  XOR U14031 ( .A(n4593), .B(n12979), .Z(n12980) );
  XOR U14032 ( .A(n12983), .B(n12984), .Z(n12979) );
  ANDN U14033 ( .B(n12985), .A(n4649), .Z(n12983) );
  XNOR U14034 ( .A(n12986), .B(n12987), .Z(n4649) );
  IV U14035 ( .A(n12984), .Z(n12987) );
  XOR U14036 ( .A(n4648), .B(n12984), .Z(n12985) );
  XOR U14037 ( .A(n12988), .B(n12989), .Z(n12984) );
  ANDN U14038 ( .B(n12990), .A(n4704), .Z(n12988) );
  XNOR U14039 ( .A(n12991), .B(n12992), .Z(n4704) );
  IV U14040 ( .A(n12989), .Z(n12992) );
  XOR U14041 ( .A(n4703), .B(n12989), .Z(n12990) );
  XOR U14042 ( .A(n12993), .B(n12994), .Z(n12989) );
  ANDN U14043 ( .B(n12995), .A(n4764), .Z(n12993) );
  XNOR U14044 ( .A(n12996), .B(n12997), .Z(n4764) );
  IV U14045 ( .A(n12994), .Z(n12997) );
  XOR U14046 ( .A(n4763), .B(n12994), .Z(n12995) );
  XOR U14047 ( .A(n12998), .B(n12999), .Z(n12994) );
  ANDN U14048 ( .B(n13000), .A(n4819), .Z(n12998) );
  XNOR U14049 ( .A(n13001), .B(n13002), .Z(n4819) );
  IV U14050 ( .A(n12999), .Z(n13002) );
  XOR U14051 ( .A(n4818), .B(n12999), .Z(n13000) );
  XOR U14052 ( .A(n13003), .B(n13004), .Z(n12999) );
  ANDN U14053 ( .B(n13005), .A(n4874), .Z(n13003) );
  XNOR U14054 ( .A(n13006), .B(n13007), .Z(n4874) );
  IV U14055 ( .A(n13004), .Z(n13007) );
  XOR U14056 ( .A(n4873), .B(n13004), .Z(n13005) );
  XOR U14057 ( .A(n13008), .B(n13009), .Z(n13004) );
  ANDN U14058 ( .B(n13010), .A(n4929), .Z(n13008) );
  XNOR U14059 ( .A(n13011), .B(n13012), .Z(n4929) );
  IV U14060 ( .A(n13009), .Z(n13012) );
  XOR U14061 ( .A(n4928), .B(n13009), .Z(n13010) );
  XOR U14062 ( .A(n13013), .B(n13014), .Z(n13009) );
  ANDN U14063 ( .B(n13015), .A(n4984), .Z(n13013) );
  XNOR U14064 ( .A(n13016), .B(n13017), .Z(n4984) );
  IV U14065 ( .A(n13014), .Z(n13017) );
  XOR U14066 ( .A(n4983), .B(n13014), .Z(n13015) );
  XOR U14067 ( .A(n13018), .B(n13019), .Z(n13014) );
  ANDN U14068 ( .B(n13020), .A(n5039), .Z(n13018) );
  XNOR U14069 ( .A(n13021), .B(n13022), .Z(n5039) );
  IV U14070 ( .A(n13019), .Z(n13022) );
  XOR U14071 ( .A(n5038), .B(n13019), .Z(n13020) );
  XOR U14072 ( .A(n13023), .B(n13024), .Z(n13019) );
  ANDN U14073 ( .B(n13025), .A(n5094), .Z(n13023) );
  XNOR U14074 ( .A(n13026), .B(n13027), .Z(n5094) );
  IV U14075 ( .A(n13024), .Z(n13027) );
  XOR U14076 ( .A(n5093), .B(n13024), .Z(n13025) );
  XOR U14077 ( .A(n13028), .B(n13029), .Z(n13024) );
  ANDN U14078 ( .B(n13030), .A(n5149), .Z(n13028) );
  XNOR U14079 ( .A(n13031), .B(n13032), .Z(n5149) );
  IV U14080 ( .A(n13029), .Z(n13032) );
  XOR U14081 ( .A(n5148), .B(n13029), .Z(n13030) );
  XOR U14082 ( .A(n13033), .B(n13034), .Z(n13029) );
  ANDN U14083 ( .B(n13035), .A(n5204), .Z(n13033) );
  XNOR U14084 ( .A(n13036), .B(n13037), .Z(n5204) );
  IV U14085 ( .A(n13034), .Z(n13037) );
  XOR U14086 ( .A(n5203), .B(n13034), .Z(n13035) );
  XOR U14087 ( .A(n13038), .B(n13039), .Z(n13034) );
  ANDN U14088 ( .B(n13040), .A(n5259), .Z(n13038) );
  XNOR U14089 ( .A(n13041), .B(n13042), .Z(n5259) );
  IV U14090 ( .A(n13039), .Z(n13042) );
  XOR U14091 ( .A(n5258), .B(n13039), .Z(n13040) );
  XOR U14092 ( .A(n13043), .B(n13044), .Z(n13039) );
  ANDN U14093 ( .B(n13045), .A(n5319), .Z(n13043) );
  XNOR U14094 ( .A(n13046), .B(n13047), .Z(n5319) );
  IV U14095 ( .A(n13044), .Z(n13047) );
  XOR U14096 ( .A(n5318), .B(n13044), .Z(n13045) );
  XOR U14097 ( .A(n13048), .B(n13049), .Z(n13044) );
  ANDN U14098 ( .B(n13050), .A(n5374), .Z(n13048) );
  XNOR U14099 ( .A(n13051), .B(n13052), .Z(n5374) );
  IV U14100 ( .A(n13049), .Z(n13052) );
  XOR U14101 ( .A(n5373), .B(n13049), .Z(n13050) );
  XOR U14102 ( .A(n13053), .B(n13054), .Z(n13049) );
  ANDN U14103 ( .B(n13055), .A(n5429), .Z(n13053) );
  XNOR U14104 ( .A(n13056), .B(n13057), .Z(n5429) );
  IV U14105 ( .A(n13054), .Z(n13057) );
  XOR U14106 ( .A(n5428), .B(n13054), .Z(n13055) );
  XOR U14107 ( .A(n13058), .B(n13059), .Z(n13054) );
  ANDN U14108 ( .B(n13060), .A(n5484), .Z(n13058) );
  XNOR U14109 ( .A(n13061), .B(n13062), .Z(n5484) );
  IV U14110 ( .A(n13059), .Z(n13062) );
  XOR U14111 ( .A(n5483), .B(n13059), .Z(n13060) );
  XOR U14112 ( .A(n13063), .B(n13064), .Z(n13059) );
  ANDN U14113 ( .B(n13065), .A(n5539), .Z(n13063) );
  XNOR U14114 ( .A(n13066), .B(n13067), .Z(n5539) );
  IV U14115 ( .A(n13064), .Z(n13067) );
  XOR U14116 ( .A(n5538), .B(n13064), .Z(n13065) );
  XOR U14117 ( .A(n13068), .B(n13069), .Z(n13064) );
  ANDN U14118 ( .B(n13070), .A(n5594), .Z(n13068) );
  XNOR U14119 ( .A(n13071), .B(n13072), .Z(n5594) );
  IV U14120 ( .A(n13069), .Z(n13072) );
  XOR U14121 ( .A(n5593), .B(n13069), .Z(n13070) );
  XOR U14122 ( .A(n13073), .B(n13074), .Z(n13069) );
  ANDN U14123 ( .B(n13075), .A(n5649), .Z(n13073) );
  XNOR U14124 ( .A(n13076), .B(n13077), .Z(n5649) );
  IV U14125 ( .A(n13074), .Z(n13077) );
  XOR U14126 ( .A(n5648), .B(n13074), .Z(n13075) );
  XOR U14127 ( .A(n13078), .B(n13079), .Z(n13074) );
  ANDN U14128 ( .B(n13080), .A(n5704), .Z(n13078) );
  XNOR U14129 ( .A(n13081), .B(n13082), .Z(n5704) );
  IV U14130 ( .A(n13079), .Z(n13082) );
  XOR U14131 ( .A(n5703), .B(n13079), .Z(n13080) );
  XOR U14132 ( .A(n13083), .B(n13084), .Z(n13079) );
  ANDN U14133 ( .B(n13085), .A(n5759), .Z(n13083) );
  XNOR U14134 ( .A(n13086), .B(n13087), .Z(n5759) );
  IV U14135 ( .A(n13084), .Z(n13087) );
  XOR U14136 ( .A(n5758), .B(n13084), .Z(n13085) );
  XOR U14137 ( .A(n13088), .B(n13089), .Z(n13084) );
  ANDN U14138 ( .B(n13090), .A(n5814), .Z(n13088) );
  XNOR U14139 ( .A(n13091), .B(n13092), .Z(n5814) );
  IV U14140 ( .A(n13089), .Z(n13092) );
  XOR U14141 ( .A(n5813), .B(n13089), .Z(n13090) );
  XOR U14142 ( .A(n13093), .B(n13094), .Z(n13089) );
  ANDN U14143 ( .B(n13095), .A(n5874), .Z(n13093) );
  XNOR U14144 ( .A(n13096), .B(n13097), .Z(n5874) );
  IV U14145 ( .A(n13094), .Z(n13097) );
  XOR U14146 ( .A(n5873), .B(n13094), .Z(n13095) );
  XOR U14147 ( .A(n13098), .B(n13099), .Z(n13094) );
  ANDN U14148 ( .B(n13100), .A(n5929), .Z(n13098) );
  XNOR U14149 ( .A(n13101), .B(n13102), .Z(n5929) );
  IV U14150 ( .A(n13099), .Z(n13102) );
  XOR U14151 ( .A(n5928), .B(n13099), .Z(n13100) );
  XOR U14152 ( .A(n13103), .B(n13104), .Z(n13099) );
  ANDN U14153 ( .B(n13105), .A(n5984), .Z(n13103) );
  XNOR U14154 ( .A(n13106), .B(n13107), .Z(n5984) );
  IV U14155 ( .A(n13104), .Z(n13107) );
  XOR U14156 ( .A(n5983), .B(n13104), .Z(n13105) );
  XOR U14157 ( .A(n13108), .B(n13109), .Z(n13104) );
  ANDN U14158 ( .B(n13110), .A(n6039), .Z(n13108) );
  XNOR U14159 ( .A(n13111), .B(n13112), .Z(n6039) );
  IV U14160 ( .A(n13109), .Z(n13112) );
  XOR U14161 ( .A(n6038), .B(n13109), .Z(n13110) );
  XOR U14162 ( .A(n13113), .B(n13114), .Z(n13109) );
  ANDN U14163 ( .B(n13115), .A(n6094), .Z(n13113) );
  XNOR U14164 ( .A(n13116), .B(n13117), .Z(n6094) );
  IV U14165 ( .A(n13114), .Z(n13117) );
  XOR U14166 ( .A(n6093), .B(n13114), .Z(n13115) );
  XOR U14167 ( .A(n13118), .B(n13119), .Z(n13114) );
  ANDN U14168 ( .B(n13120), .A(n6149), .Z(n13118) );
  XNOR U14169 ( .A(n13121), .B(n13122), .Z(n6149) );
  IV U14170 ( .A(n13119), .Z(n13122) );
  XOR U14171 ( .A(n6148), .B(n13119), .Z(n13120) );
  XOR U14172 ( .A(n13123), .B(n13124), .Z(n13119) );
  ANDN U14173 ( .B(n13125), .A(n6204), .Z(n13123) );
  XNOR U14174 ( .A(n13126), .B(n13127), .Z(n6204) );
  IV U14175 ( .A(n13124), .Z(n13127) );
  XOR U14176 ( .A(n6203), .B(n13124), .Z(n13125) );
  XOR U14177 ( .A(n13128), .B(n13129), .Z(n13124) );
  ANDN U14178 ( .B(n13130), .A(n6259), .Z(n13128) );
  XNOR U14179 ( .A(n13131), .B(n13132), .Z(n6259) );
  IV U14180 ( .A(n13129), .Z(n13132) );
  XOR U14181 ( .A(n6258), .B(n13129), .Z(n13130) );
  XOR U14182 ( .A(n13133), .B(n13134), .Z(n13129) );
  ANDN U14183 ( .B(n13135), .A(n6314), .Z(n13133) );
  XNOR U14184 ( .A(n13136), .B(n13137), .Z(n6314) );
  IV U14185 ( .A(n13134), .Z(n13137) );
  XOR U14186 ( .A(n6313), .B(n13134), .Z(n13135) );
  XOR U14187 ( .A(n13138), .B(n13139), .Z(n13134) );
  ANDN U14188 ( .B(n13140), .A(n6369), .Z(n13138) );
  XNOR U14189 ( .A(n13141), .B(n13142), .Z(n6369) );
  IV U14190 ( .A(n13139), .Z(n13142) );
  XOR U14191 ( .A(n6368), .B(n13139), .Z(n13140) );
  XOR U14192 ( .A(n13143), .B(n13144), .Z(n13139) );
  ANDN U14193 ( .B(n13145), .A(n6429), .Z(n13143) );
  XNOR U14194 ( .A(n13146), .B(n13147), .Z(n6429) );
  IV U14195 ( .A(n13144), .Z(n13147) );
  XOR U14196 ( .A(n6428), .B(n13144), .Z(n13145) );
  XOR U14197 ( .A(n13148), .B(n13149), .Z(n13144) );
  ANDN U14198 ( .B(n13150), .A(n6484), .Z(n13148) );
  XNOR U14199 ( .A(n13151), .B(n13152), .Z(n6484) );
  IV U14200 ( .A(n13149), .Z(n13152) );
  XOR U14201 ( .A(n6483), .B(n13149), .Z(n13150) );
  XOR U14202 ( .A(n13153), .B(n13154), .Z(n13149) );
  ANDN U14203 ( .B(n13155), .A(n6539), .Z(n13153) );
  XNOR U14204 ( .A(n13156), .B(n13157), .Z(n6539) );
  IV U14205 ( .A(n13154), .Z(n13157) );
  XOR U14206 ( .A(n6538), .B(n13154), .Z(n13155) );
  XOR U14207 ( .A(n13158), .B(n13159), .Z(n13154) );
  ANDN U14208 ( .B(n13160), .A(n6594), .Z(n13158) );
  XNOR U14209 ( .A(n13161), .B(n13162), .Z(n6594) );
  IV U14210 ( .A(n13159), .Z(n13162) );
  XOR U14211 ( .A(n6593), .B(n13159), .Z(n13160) );
  XOR U14212 ( .A(n13163), .B(n13164), .Z(n13159) );
  ANDN U14213 ( .B(n13165), .A(n6649), .Z(n13163) );
  XNOR U14214 ( .A(n13166), .B(n13167), .Z(n6649) );
  IV U14215 ( .A(n13164), .Z(n13167) );
  XOR U14216 ( .A(n6648), .B(n13164), .Z(n13165) );
  XOR U14217 ( .A(n13168), .B(n13169), .Z(n13164) );
  ANDN U14218 ( .B(n13170), .A(n6704), .Z(n13168) );
  XNOR U14219 ( .A(n13171), .B(n13172), .Z(n6704) );
  IV U14220 ( .A(n13169), .Z(n13172) );
  XOR U14221 ( .A(n6703), .B(n13169), .Z(n13170) );
  XOR U14222 ( .A(n13173), .B(n13174), .Z(n13169) );
  ANDN U14223 ( .B(n13175), .A(n6759), .Z(n13173) );
  XNOR U14224 ( .A(n13176), .B(n13177), .Z(n6759) );
  IV U14225 ( .A(n13174), .Z(n13177) );
  XOR U14226 ( .A(n6758), .B(n13174), .Z(n13175) );
  XOR U14227 ( .A(n13178), .B(n13179), .Z(n13174) );
  ANDN U14228 ( .B(n13180), .A(n6814), .Z(n13178) );
  XNOR U14229 ( .A(n13181), .B(n13182), .Z(n6814) );
  IV U14230 ( .A(n13179), .Z(n13182) );
  XOR U14231 ( .A(n6813), .B(n13179), .Z(n13180) );
  XOR U14232 ( .A(n13183), .B(n13184), .Z(n13179) );
  ANDN U14233 ( .B(n13185), .A(n6869), .Z(n13183) );
  XNOR U14234 ( .A(n13186), .B(n13187), .Z(n6869) );
  IV U14235 ( .A(n13184), .Z(n13187) );
  XOR U14236 ( .A(n6868), .B(n13184), .Z(n13185) );
  XOR U14237 ( .A(n13188), .B(n13189), .Z(n13184) );
  ANDN U14238 ( .B(n13190), .A(n6924), .Z(n13188) );
  XNOR U14239 ( .A(n13191), .B(n13192), .Z(n6924) );
  IV U14240 ( .A(n13189), .Z(n13192) );
  XOR U14241 ( .A(n6923), .B(n13189), .Z(n13190) );
  XOR U14242 ( .A(n13193), .B(n13194), .Z(n13189) );
  ANDN U14243 ( .B(n13195), .A(n6984), .Z(n13193) );
  XNOR U14244 ( .A(n13196), .B(n13197), .Z(n6984) );
  IV U14245 ( .A(n13194), .Z(n13197) );
  XOR U14246 ( .A(n6983), .B(n13194), .Z(n13195) );
  XOR U14247 ( .A(n13198), .B(n13199), .Z(n13194) );
  ANDN U14248 ( .B(n13200), .A(n7039), .Z(n13198) );
  XNOR U14249 ( .A(n13201), .B(n13202), .Z(n7039) );
  IV U14250 ( .A(n13199), .Z(n13202) );
  XOR U14251 ( .A(n7038), .B(n13199), .Z(n13200) );
  XOR U14252 ( .A(n13203), .B(n13204), .Z(n13199) );
  ANDN U14253 ( .B(n13205), .A(n7094), .Z(n13203) );
  XNOR U14254 ( .A(n13206), .B(n13207), .Z(n7094) );
  IV U14255 ( .A(n13204), .Z(n13207) );
  XOR U14256 ( .A(n7093), .B(n13204), .Z(n13205) );
  XOR U14257 ( .A(n13208), .B(n13209), .Z(n13204) );
  ANDN U14258 ( .B(n13210), .A(n7149), .Z(n13208) );
  XNOR U14259 ( .A(n13211), .B(n13212), .Z(n7149) );
  IV U14260 ( .A(n13209), .Z(n13212) );
  XOR U14261 ( .A(n7148), .B(n13209), .Z(n13210) );
  XOR U14262 ( .A(n13213), .B(n13214), .Z(n13209) );
  ANDN U14263 ( .B(n13215), .A(n7204), .Z(n13213) );
  XNOR U14264 ( .A(n13216), .B(n13217), .Z(n7204) );
  IV U14265 ( .A(n13214), .Z(n13217) );
  XOR U14266 ( .A(n7203), .B(n13214), .Z(n13215) );
  XOR U14267 ( .A(n13218), .B(n13219), .Z(n13214) );
  ANDN U14268 ( .B(n13220), .A(n7259), .Z(n13218) );
  XNOR U14269 ( .A(n13221), .B(n13222), .Z(n7259) );
  IV U14270 ( .A(n13219), .Z(n13222) );
  XOR U14271 ( .A(n7258), .B(n13219), .Z(n13220) );
  XOR U14272 ( .A(n13223), .B(n13224), .Z(n13219) );
  ANDN U14273 ( .B(n13225), .A(n7314), .Z(n13223) );
  XNOR U14274 ( .A(n13226), .B(n13227), .Z(n7314) );
  IV U14275 ( .A(n13224), .Z(n13227) );
  XOR U14276 ( .A(n7313), .B(n13224), .Z(n13225) );
  XOR U14277 ( .A(n13228), .B(n13229), .Z(n13224) );
  ANDN U14278 ( .B(n13230), .A(n7369), .Z(n13228) );
  XNOR U14279 ( .A(n13231), .B(n13232), .Z(n7369) );
  IV U14280 ( .A(n13229), .Z(n13232) );
  XOR U14281 ( .A(n7368), .B(n13229), .Z(n13230) );
  XOR U14282 ( .A(n13233), .B(n13234), .Z(n13229) );
  ANDN U14283 ( .B(n13235), .A(n7424), .Z(n13233) );
  XNOR U14284 ( .A(n13236), .B(n13237), .Z(n7424) );
  IV U14285 ( .A(n13234), .Z(n13237) );
  XOR U14286 ( .A(n7423), .B(n13234), .Z(n13235) );
  XOR U14287 ( .A(n13238), .B(n13239), .Z(n13234) );
  ANDN U14288 ( .B(n13240), .A(n7479), .Z(n13238) );
  XNOR U14289 ( .A(n13241), .B(n13242), .Z(n7479) );
  IV U14290 ( .A(n13239), .Z(n13242) );
  XOR U14291 ( .A(n7478), .B(n13239), .Z(n13240) );
  XOR U14292 ( .A(n13243), .B(n13244), .Z(n13239) );
  ANDN U14293 ( .B(n13245), .A(n7539), .Z(n13243) );
  XNOR U14294 ( .A(n13246), .B(n13247), .Z(n7539) );
  IV U14295 ( .A(n13244), .Z(n13247) );
  XOR U14296 ( .A(n7538), .B(n13244), .Z(n13245) );
  XOR U14297 ( .A(n13248), .B(n13249), .Z(n13244) );
  ANDN U14298 ( .B(n13250), .A(n7594), .Z(n13248) );
  XNOR U14299 ( .A(n13251), .B(n13252), .Z(n7594) );
  IV U14300 ( .A(n13249), .Z(n13252) );
  XOR U14301 ( .A(n7593), .B(n13249), .Z(n13250) );
  XOR U14302 ( .A(n13253), .B(n13254), .Z(n13249) );
  ANDN U14303 ( .B(n13255), .A(n7649), .Z(n13253) );
  XNOR U14304 ( .A(n13256), .B(n13257), .Z(n7649) );
  IV U14305 ( .A(n13254), .Z(n13257) );
  XOR U14306 ( .A(n7648), .B(n13254), .Z(n13255) );
  XOR U14307 ( .A(n13258), .B(n13259), .Z(n13254) );
  ANDN U14308 ( .B(n13260), .A(n7704), .Z(n13258) );
  XNOR U14309 ( .A(n13261), .B(n13262), .Z(n7704) );
  IV U14310 ( .A(n13259), .Z(n13262) );
  XOR U14311 ( .A(n7703), .B(n13259), .Z(n13260) );
  XOR U14312 ( .A(n13263), .B(n13264), .Z(n13259) );
  ANDN U14313 ( .B(n13265), .A(n7759), .Z(n13263) );
  XNOR U14314 ( .A(n13266), .B(n13267), .Z(n7759) );
  IV U14315 ( .A(n13264), .Z(n13267) );
  XOR U14316 ( .A(n7758), .B(n13264), .Z(n13265) );
  XOR U14317 ( .A(n13268), .B(n13269), .Z(n13264) );
  ANDN U14318 ( .B(n13270), .A(n7814), .Z(n13268) );
  XNOR U14319 ( .A(n13271), .B(n13272), .Z(n7814) );
  IV U14320 ( .A(n13269), .Z(n13272) );
  XOR U14321 ( .A(n7813), .B(n13269), .Z(n13270) );
  XOR U14322 ( .A(n13273), .B(n13274), .Z(n13269) );
  ANDN U14323 ( .B(n13275), .A(n7869), .Z(n13273) );
  XNOR U14324 ( .A(n13276), .B(n13277), .Z(n7869) );
  IV U14325 ( .A(n13274), .Z(n13277) );
  XOR U14326 ( .A(n7868), .B(n13274), .Z(n13275) );
  XOR U14327 ( .A(n13278), .B(n13279), .Z(n13274) );
  ANDN U14328 ( .B(n13280), .A(n7924), .Z(n13278) );
  XNOR U14329 ( .A(n13281), .B(n13282), .Z(n7924) );
  IV U14330 ( .A(n13279), .Z(n13282) );
  XOR U14331 ( .A(n7923), .B(n13279), .Z(n13280) );
  XOR U14332 ( .A(n13283), .B(n13284), .Z(n13279) );
  ANDN U14333 ( .B(n13285), .A(n7979), .Z(n13283) );
  XNOR U14334 ( .A(n13286), .B(n13287), .Z(n7979) );
  IV U14335 ( .A(n13284), .Z(n13287) );
  XOR U14336 ( .A(n7978), .B(n13284), .Z(n13285) );
  XOR U14337 ( .A(n13288), .B(n13289), .Z(n13284) );
  ANDN U14338 ( .B(n13290), .A(n8034), .Z(n13288) );
  XNOR U14339 ( .A(n13291), .B(n13292), .Z(n8034) );
  IV U14340 ( .A(n13289), .Z(n13292) );
  XOR U14341 ( .A(n8033), .B(n13289), .Z(n13290) );
  XOR U14342 ( .A(n13293), .B(n13294), .Z(n13289) );
  ANDN U14343 ( .B(n13295), .A(n3094), .Z(n13293) );
  XNOR U14344 ( .A(n13296), .B(n13297), .Z(n3094) );
  IV U14345 ( .A(n13294), .Z(n13297) );
  XOR U14346 ( .A(n3093), .B(n13294), .Z(n13295) );
  XOR U14347 ( .A(n13298), .B(n13299), .Z(n13294) );
  ANDN U14348 ( .B(n13300), .A(n3649), .Z(n13298) );
  XNOR U14349 ( .A(n13301), .B(n13302), .Z(n3649) );
  IV U14350 ( .A(n13299), .Z(n13302) );
  XOR U14351 ( .A(n3648), .B(n13299), .Z(n13300) );
  XOR U14352 ( .A(n13303), .B(n13304), .Z(n13299) );
  ANDN U14353 ( .B(n13305), .A(n4204), .Z(n13303) );
  XNOR U14354 ( .A(n13306), .B(n13307), .Z(n4204) );
  IV U14355 ( .A(n13304), .Z(n13307) );
  XOR U14356 ( .A(n4203), .B(n13304), .Z(n13305) );
  XOR U14357 ( .A(n13308), .B(n13309), .Z(n13304) );
  ANDN U14358 ( .B(n13310), .A(n4759), .Z(n13308) );
  XNOR U14359 ( .A(n13311), .B(n13312), .Z(n4759) );
  IV U14360 ( .A(n13309), .Z(n13312) );
  XOR U14361 ( .A(n4758), .B(n13309), .Z(n13310) );
  XOR U14362 ( .A(n13313), .B(n13314), .Z(n13309) );
  ANDN U14363 ( .B(n13315), .A(n5314), .Z(n13313) );
  XNOR U14364 ( .A(n13316), .B(n13317), .Z(n5314) );
  IV U14365 ( .A(n13314), .Z(n13317) );
  XOR U14366 ( .A(n5313), .B(n13314), .Z(n13315) );
  XOR U14367 ( .A(n13318), .B(n13319), .Z(n13314) );
  ANDN U14368 ( .B(n13320), .A(n5869), .Z(n13318) );
  XNOR U14369 ( .A(n13321), .B(n13322), .Z(n5869) );
  IV U14370 ( .A(n13319), .Z(n13322) );
  XOR U14371 ( .A(n5868), .B(n13319), .Z(n13320) );
  XOR U14372 ( .A(n13323), .B(n13324), .Z(n13319) );
  ANDN U14373 ( .B(n13325), .A(n6424), .Z(n13323) );
  XNOR U14374 ( .A(n13326), .B(n13327), .Z(n6424) );
  IV U14375 ( .A(n13324), .Z(n13327) );
  XOR U14376 ( .A(n6423), .B(n13324), .Z(n13325) );
  XOR U14377 ( .A(n13328), .B(n13329), .Z(n13324) );
  ANDN U14378 ( .B(n13330), .A(n6979), .Z(n13328) );
  XOR U14379 ( .A(n13331), .B(n13329), .Z(n6979) );
  XOR U14380 ( .A(n6978), .B(n13329), .Z(n13330) );
  XNOR U14381 ( .A(n13332), .B(n13333), .Z(n13329) );
  NANDN U14382 ( .A(n7534), .B(n13334), .Z(n13333) );
  XNOR U14383 ( .A(n13335), .B(n7533), .Z(n13334) );
  NAND U14384 ( .A(n13336), .B(n[1]), .Z(n7533) );
  NAND U14385 ( .A(n8085), .B(n[1]), .Z(n13336) );
  XOR U14386 ( .A(n13335), .B(n13337), .Z(n7534) );
  IV U14387 ( .A(n13332), .Z(n13335) );
  NANDN U14388 ( .A(n13338), .B(n13339), .Z(n13332) );
  NAND U14389 ( .A(n13340), .B(n[2]), .Z(n6978) );
  NAND U14390 ( .A(n8085), .B(n[2]), .Z(n13340) );
  NAND U14391 ( .A(n13341), .B(n[3]), .Z(n6423) );
  NAND U14392 ( .A(n8085), .B(n[3]), .Z(n13341) );
  NAND U14393 ( .A(n13342), .B(n[4]), .Z(n5868) );
  NAND U14394 ( .A(n8085), .B(n[4]), .Z(n13342) );
  NAND U14395 ( .A(n13343), .B(n[5]), .Z(n5313) );
  NAND U14396 ( .A(n8085), .B(n[5]), .Z(n13343) );
  NAND U14397 ( .A(n13344), .B(n[6]), .Z(n4758) );
  NAND U14398 ( .A(n8085), .B(n[6]), .Z(n13344) );
  NAND U14399 ( .A(n13345), .B(n[7]), .Z(n4203) );
  NAND U14400 ( .A(n8085), .B(n[7]), .Z(n13345) );
  NAND U14401 ( .A(n13346), .B(n[8]), .Z(n3648) );
  NAND U14402 ( .A(n8085), .B(n[8]), .Z(n13346) );
  NAND U14403 ( .A(n13347), .B(n[9]), .Z(n3093) );
  NAND U14404 ( .A(n8085), .B(n[9]), .Z(n13347) );
  NAND U14405 ( .A(n13348), .B(n[10]), .Z(n8033) );
  NAND U14406 ( .A(n8085), .B(n[10]), .Z(n13348) );
  NAND U14407 ( .A(n13349), .B(n[11]), .Z(n7978) );
  NAND U14408 ( .A(n8085), .B(n[11]), .Z(n13349) );
  NAND U14409 ( .A(n13350), .B(n[12]), .Z(n7923) );
  NAND U14410 ( .A(n8085), .B(n[12]), .Z(n13350) );
  NAND U14411 ( .A(n13351), .B(n[13]), .Z(n7868) );
  NAND U14412 ( .A(n8085), .B(n[13]), .Z(n13351) );
  NAND U14413 ( .A(n13352), .B(n[14]), .Z(n7813) );
  NAND U14414 ( .A(n8085), .B(n[14]), .Z(n13352) );
  NAND U14415 ( .A(n13353), .B(n[15]), .Z(n7758) );
  NAND U14416 ( .A(n8085), .B(n[15]), .Z(n13353) );
  NAND U14417 ( .A(n13354), .B(n[16]), .Z(n7703) );
  NAND U14418 ( .A(n8085), .B(n[16]), .Z(n13354) );
  NAND U14419 ( .A(n13355), .B(n[17]), .Z(n7648) );
  NAND U14420 ( .A(n8085), .B(n[17]), .Z(n13355) );
  NAND U14421 ( .A(n13356), .B(n[18]), .Z(n7593) );
  NAND U14422 ( .A(n8085), .B(n[18]), .Z(n13356) );
  NAND U14423 ( .A(n13357), .B(n[19]), .Z(n7538) );
  NAND U14424 ( .A(n8085), .B(n[19]), .Z(n13357) );
  NAND U14425 ( .A(n13358), .B(n[20]), .Z(n7478) );
  NAND U14426 ( .A(n8085), .B(n[20]), .Z(n13358) );
  NAND U14427 ( .A(n13359), .B(n[21]), .Z(n7423) );
  NAND U14428 ( .A(n8085), .B(n[21]), .Z(n13359) );
  NAND U14429 ( .A(n13360), .B(n[22]), .Z(n7368) );
  NAND U14430 ( .A(n8085), .B(n[22]), .Z(n13360) );
  NAND U14431 ( .A(n13361), .B(n[23]), .Z(n7313) );
  NAND U14432 ( .A(n8085), .B(n[23]), .Z(n13361) );
  NAND U14433 ( .A(n13362), .B(n[24]), .Z(n7258) );
  NAND U14434 ( .A(n8085), .B(n[24]), .Z(n13362) );
  NAND U14435 ( .A(n13363), .B(n[25]), .Z(n7203) );
  NAND U14436 ( .A(n8085), .B(n[25]), .Z(n13363) );
  NAND U14437 ( .A(n13364), .B(n[26]), .Z(n7148) );
  NAND U14438 ( .A(n8085), .B(n[26]), .Z(n13364) );
  NAND U14439 ( .A(n13365), .B(n[27]), .Z(n7093) );
  NAND U14440 ( .A(n8085), .B(n[27]), .Z(n13365) );
  NAND U14441 ( .A(n13366), .B(n[28]), .Z(n7038) );
  NAND U14442 ( .A(n8085), .B(n[28]), .Z(n13366) );
  NAND U14443 ( .A(n13367), .B(n[29]), .Z(n6983) );
  NAND U14444 ( .A(n8085), .B(n[29]), .Z(n13367) );
  NAND U14445 ( .A(n13368), .B(n[30]), .Z(n6923) );
  NAND U14446 ( .A(n8085), .B(n[30]), .Z(n13368) );
  NAND U14447 ( .A(n13369), .B(n[31]), .Z(n6868) );
  NAND U14448 ( .A(n8085), .B(n[31]), .Z(n13369) );
  NAND U14449 ( .A(n13370), .B(n[32]), .Z(n6813) );
  NAND U14450 ( .A(n8085), .B(n[32]), .Z(n13370) );
  NAND U14451 ( .A(n13371), .B(n[33]), .Z(n6758) );
  NAND U14452 ( .A(n8085), .B(n[33]), .Z(n13371) );
  NAND U14453 ( .A(n13372), .B(n[34]), .Z(n6703) );
  NAND U14454 ( .A(n8085), .B(n[34]), .Z(n13372) );
  NAND U14455 ( .A(n13373), .B(n[35]), .Z(n6648) );
  NAND U14456 ( .A(n8085), .B(n[35]), .Z(n13373) );
  NAND U14457 ( .A(n13374), .B(n[36]), .Z(n6593) );
  NAND U14458 ( .A(n8085), .B(n[36]), .Z(n13374) );
  NAND U14459 ( .A(n13375), .B(n[37]), .Z(n6538) );
  NAND U14460 ( .A(n8085), .B(n[37]), .Z(n13375) );
  NAND U14461 ( .A(n13376), .B(n[38]), .Z(n6483) );
  NAND U14462 ( .A(n8085), .B(n[38]), .Z(n13376) );
  NAND U14463 ( .A(n13377), .B(n[39]), .Z(n6428) );
  NAND U14464 ( .A(n8085), .B(n[39]), .Z(n13377) );
  NAND U14465 ( .A(n13378), .B(n[40]), .Z(n6368) );
  NAND U14466 ( .A(n8085), .B(n[40]), .Z(n13378) );
  NAND U14467 ( .A(n13379), .B(n[41]), .Z(n6313) );
  NAND U14468 ( .A(n8085), .B(n[41]), .Z(n13379) );
  NAND U14469 ( .A(n13380), .B(n[42]), .Z(n6258) );
  NAND U14470 ( .A(n8085), .B(n[42]), .Z(n13380) );
  NAND U14471 ( .A(n13381), .B(n[43]), .Z(n6203) );
  NAND U14472 ( .A(n8085), .B(n[43]), .Z(n13381) );
  NAND U14473 ( .A(n13382), .B(n[44]), .Z(n6148) );
  NAND U14474 ( .A(n8085), .B(n[44]), .Z(n13382) );
  NAND U14475 ( .A(n13383), .B(n[45]), .Z(n6093) );
  NAND U14476 ( .A(n8085), .B(n[45]), .Z(n13383) );
  NAND U14477 ( .A(n13384), .B(n[46]), .Z(n6038) );
  NAND U14478 ( .A(n8085), .B(n[46]), .Z(n13384) );
  NAND U14479 ( .A(n13385), .B(n[47]), .Z(n5983) );
  NAND U14480 ( .A(n8085), .B(n[47]), .Z(n13385) );
  NAND U14481 ( .A(n13386), .B(n[48]), .Z(n5928) );
  NAND U14482 ( .A(n8085), .B(n[48]), .Z(n13386) );
  NAND U14483 ( .A(n13387), .B(n[49]), .Z(n5873) );
  NAND U14484 ( .A(n8085), .B(n[49]), .Z(n13387) );
  NAND U14485 ( .A(n13388), .B(n[50]), .Z(n5813) );
  NAND U14486 ( .A(n8085), .B(n[50]), .Z(n13388) );
  NAND U14487 ( .A(n13389), .B(n[51]), .Z(n5758) );
  NAND U14488 ( .A(n8085), .B(n[51]), .Z(n13389) );
  NAND U14489 ( .A(n13390), .B(n[52]), .Z(n5703) );
  NAND U14490 ( .A(n8085), .B(n[52]), .Z(n13390) );
  NAND U14491 ( .A(n13391), .B(n[53]), .Z(n5648) );
  NAND U14492 ( .A(n8085), .B(n[53]), .Z(n13391) );
  NAND U14493 ( .A(n13392), .B(n[54]), .Z(n5593) );
  NAND U14494 ( .A(n8085), .B(n[54]), .Z(n13392) );
  NAND U14495 ( .A(n13393), .B(n[55]), .Z(n5538) );
  NAND U14496 ( .A(n8085), .B(n[55]), .Z(n13393) );
  NAND U14497 ( .A(n13394), .B(n[56]), .Z(n5483) );
  NAND U14498 ( .A(n8085), .B(n[56]), .Z(n13394) );
  NAND U14499 ( .A(n13395), .B(n[57]), .Z(n5428) );
  NAND U14500 ( .A(n8085), .B(n[57]), .Z(n13395) );
  NAND U14501 ( .A(n13396), .B(n[58]), .Z(n5373) );
  NAND U14502 ( .A(n8085), .B(n[58]), .Z(n13396) );
  NAND U14503 ( .A(n13397), .B(n[59]), .Z(n5318) );
  NAND U14504 ( .A(n8085), .B(n[59]), .Z(n13397) );
  NAND U14505 ( .A(n13398), .B(n[60]), .Z(n5258) );
  NAND U14506 ( .A(n8085), .B(n[60]), .Z(n13398) );
  NAND U14507 ( .A(n13399), .B(n[61]), .Z(n5203) );
  NAND U14508 ( .A(n8085), .B(n[61]), .Z(n13399) );
  NAND U14509 ( .A(n13400), .B(n[62]), .Z(n5148) );
  NAND U14510 ( .A(n8085), .B(n[62]), .Z(n13400) );
  NAND U14511 ( .A(n13401), .B(n[63]), .Z(n5093) );
  NAND U14512 ( .A(n8085), .B(n[63]), .Z(n13401) );
  NAND U14513 ( .A(n13402), .B(n[64]), .Z(n5038) );
  NAND U14514 ( .A(n8085), .B(n[64]), .Z(n13402) );
  NAND U14515 ( .A(n13403), .B(n[65]), .Z(n4983) );
  NAND U14516 ( .A(n8085), .B(n[65]), .Z(n13403) );
  NAND U14517 ( .A(n13404), .B(n[66]), .Z(n4928) );
  NAND U14518 ( .A(n8085), .B(n[66]), .Z(n13404) );
  NAND U14519 ( .A(n13405), .B(n[67]), .Z(n4873) );
  NAND U14520 ( .A(n8085), .B(n[67]), .Z(n13405) );
  NAND U14521 ( .A(n13406), .B(n[68]), .Z(n4818) );
  NAND U14522 ( .A(n8085), .B(n[68]), .Z(n13406) );
  NAND U14523 ( .A(n13407), .B(n[69]), .Z(n4763) );
  NAND U14524 ( .A(n8085), .B(n[69]), .Z(n13407) );
  NAND U14525 ( .A(n13408), .B(n[70]), .Z(n4703) );
  NAND U14526 ( .A(n8085), .B(n[70]), .Z(n13408) );
  NAND U14527 ( .A(n13409), .B(n[71]), .Z(n4648) );
  NAND U14528 ( .A(n8085), .B(n[71]), .Z(n13409) );
  NAND U14529 ( .A(n13410), .B(n[72]), .Z(n4593) );
  NAND U14530 ( .A(n8085), .B(n[72]), .Z(n13410) );
  NAND U14531 ( .A(n13411), .B(n[73]), .Z(n4538) );
  NAND U14532 ( .A(n8085), .B(n[73]), .Z(n13411) );
  NAND U14533 ( .A(n13412), .B(n[74]), .Z(n4483) );
  NAND U14534 ( .A(n8085), .B(n[74]), .Z(n13412) );
  NAND U14535 ( .A(n13413), .B(n[75]), .Z(n4428) );
  NAND U14536 ( .A(n8085), .B(n[75]), .Z(n13413) );
  NAND U14537 ( .A(n13414), .B(n[76]), .Z(n4373) );
  NAND U14538 ( .A(n8085), .B(n[76]), .Z(n13414) );
  NAND U14539 ( .A(n13415), .B(n[77]), .Z(n4318) );
  NAND U14540 ( .A(n8085), .B(n[77]), .Z(n13415) );
  NAND U14541 ( .A(n13416), .B(n[78]), .Z(n4263) );
  NAND U14542 ( .A(n8085), .B(n[78]), .Z(n13416) );
  NAND U14543 ( .A(n13417), .B(n[79]), .Z(n4208) );
  NAND U14544 ( .A(n8085), .B(n[79]), .Z(n13417) );
  NAND U14545 ( .A(n13418), .B(n[80]), .Z(n4148) );
  NAND U14546 ( .A(n8085), .B(n[80]), .Z(n13418) );
  NAND U14547 ( .A(n13419), .B(n[81]), .Z(n4093) );
  NAND U14548 ( .A(n8085), .B(n[81]), .Z(n13419) );
  NAND U14549 ( .A(n13420), .B(n[82]), .Z(n4038) );
  NAND U14550 ( .A(n8085), .B(n[82]), .Z(n13420) );
  NAND U14551 ( .A(n13421), .B(n[83]), .Z(n3983) );
  NAND U14552 ( .A(n8085), .B(n[83]), .Z(n13421) );
  NAND U14553 ( .A(n13422), .B(n[84]), .Z(n3928) );
  NAND U14554 ( .A(n8085), .B(n[84]), .Z(n13422) );
  NAND U14555 ( .A(n13423), .B(n[85]), .Z(n3873) );
  NAND U14556 ( .A(n8085), .B(n[85]), .Z(n13423) );
  NAND U14557 ( .A(n13424), .B(n[86]), .Z(n3818) );
  NAND U14558 ( .A(n8085), .B(n[86]), .Z(n13424) );
  NAND U14559 ( .A(n13425), .B(n[87]), .Z(n3763) );
  NAND U14560 ( .A(n8085), .B(n[87]), .Z(n13425) );
  NAND U14561 ( .A(n13426), .B(n[88]), .Z(n3708) );
  NAND U14562 ( .A(n8085), .B(n[88]), .Z(n13426) );
  NAND U14563 ( .A(n13427), .B(n[89]), .Z(n3653) );
  NAND U14564 ( .A(n8085), .B(n[89]), .Z(n13427) );
  NAND U14565 ( .A(n13428), .B(n[90]), .Z(n3593) );
  NAND U14566 ( .A(n8085), .B(n[90]), .Z(n13428) );
  NAND U14567 ( .A(n13429), .B(n[91]), .Z(n3538) );
  NAND U14568 ( .A(n8085), .B(n[91]), .Z(n13429) );
  NAND U14569 ( .A(n13430), .B(n[92]), .Z(n3483) );
  NAND U14570 ( .A(n8085), .B(n[92]), .Z(n13430) );
  NAND U14571 ( .A(n13431), .B(n[93]), .Z(n3428) );
  NAND U14572 ( .A(n8085), .B(n[93]), .Z(n13431) );
  NAND U14573 ( .A(n13432), .B(n[94]), .Z(n3373) );
  NAND U14574 ( .A(n8085), .B(n[94]), .Z(n13432) );
  NAND U14575 ( .A(n13433), .B(n[95]), .Z(n3318) );
  NAND U14576 ( .A(n8085), .B(n[95]), .Z(n13433) );
  NAND U14577 ( .A(n13434), .B(n[96]), .Z(n3263) );
  NAND U14578 ( .A(n8085), .B(n[96]), .Z(n13434) );
  NAND U14579 ( .A(n13435), .B(n[97]), .Z(n3208) );
  NAND U14580 ( .A(n8085), .B(n[97]), .Z(n13435) );
  NAND U14581 ( .A(n13436), .B(n[98]), .Z(n3153) );
  NAND U14582 ( .A(n8085), .B(n[98]), .Z(n13436) );
  NAND U14583 ( .A(n13437), .B(n[99]), .Z(n3098) );
  NAND U14584 ( .A(n8085), .B(n[99]), .Z(n13437) );
  NAND U14585 ( .A(n13438), .B(n[100]), .Z(n8237) );
  NAND U14586 ( .A(n8085), .B(n[100]), .Z(n13438) );
  NAND U14587 ( .A(n13439), .B(n[101]), .Z(n8122) );
  NAND U14588 ( .A(n8085), .B(n[101]), .Z(n13439) );
  NAND U14589 ( .A(n13440), .B(n[102]), .Z(n8073) );
  NAND U14590 ( .A(n8085), .B(n[102]), .Z(n13440) );
  NAND U14591 ( .A(n13441), .B(n[103]), .Z(n8068) );
  NAND U14592 ( .A(n8085), .B(n[103]), .Z(n13441) );
  NAND U14593 ( .A(n13442), .B(n[104]), .Z(n8063) );
  NAND U14594 ( .A(n8085), .B(n[104]), .Z(n13442) );
  NAND U14595 ( .A(n13443), .B(n[105]), .Z(n8058) );
  NAND U14596 ( .A(n8085), .B(n[105]), .Z(n13443) );
  NAND U14597 ( .A(n13444), .B(n[106]), .Z(n8053) );
  NAND U14598 ( .A(n8085), .B(n[106]), .Z(n13444) );
  NAND U14599 ( .A(n13445), .B(n[107]), .Z(n8048) );
  NAND U14600 ( .A(n8085), .B(n[107]), .Z(n13445) );
  NAND U14601 ( .A(n13446), .B(n[108]), .Z(n8043) );
  NAND U14602 ( .A(n8085), .B(n[108]), .Z(n13446) );
  NAND U14603 ( .A(n13447), .B(n[109]), .Z(n8038) );
  NAND U14604 ( .A(n8085), .B(n[109]), .Z(n13447) );
  NAND U14605 ( .A(n13448), .B(n[110]), .Z(n8028) );
  NAND U14606 ( .A(n8085), .B(n[110]), .Z(n13448) );
  NAND U14607 ( .A(n13449), .B(n[111]), .Z(n8023) );
  NAND U14608 ( .A(n8085), .B(n[111]), .Z(n13449) );
  NAND U14609 ( .A(n13450), .B(n[112]), .Z(n8018) );
  NAND U14610 ( .A(n8085), .B(n[112]), .Z(n13450) );
  NAND U14611 ( .A(n13451), .B(n[113]), .Z(n8013) );
  NAND U14612 ( .A(n8085), .B(n[113]), .Z(n13451) );
  NAND U14613 ( .A(n13452), .B(n[114]), .Z(n8008) );
  NAND U14614 ( .A(n8085), .B(n[114]), .Z(n13452) );
  NAND U14615 ( .A(n13453), .B(n[115]), .Z(n8003) );
  NAND U14616 ( .A(n8085), .B(n[115]), .Z(n13453) );
  NAND U14617 ( .A(n13454), .B(n[116]), .Z(n7998) );
  NAND U14618 ( .A(n8085), .B(n[116]), .Z(n13454) );
  NAND U14619 ( .A(n13455), .B(n[117]), .Z(n7993) );
  NAND U14620 ( .A(n8085), .B(n[117]), .Z(n13455) );
  NAND U14621 ( .A(n13456), .B(n[118]), .Z(n7988) );
  NAND U14622 ( .A(n8085), .B(n[118]), .Z(n13456) );
  NAND U14623 ( .A(n13457), .B(n[119]), .Z(n7983) );
  NAND U14624 ( .A(n8085), .B(n[119]), .Z(n13457) );
  NAND U14625 ( .A(n13458), .B(n[120]), .Z(n7973) );
  NAND U14626 ( .A(n8085), .B(n[120]), .Z(n13458) );
  NAND U14627 ( .A(n13459), .B(n[121]), .Z(n7968) );
  NAND U14628 ( .A(n8085), .B(n[121]), .Z(n13459) );
  NAND U14629 ( .A(n13460), .B(n[122]), .Z(n7963) );
  NAND U14630 ( .A(n8085), .B(n[122]), .Z(n13460) );
  NAND U14631 ( .A(n13461), .B(n[123]), .Z(n7958) );
  NAND U14632 ( .A(n8085), .B(n[123]), .Z(n13461) );
  NAND U14633 ( .A(n13462), .B(n[124]), .Z(n7953) );
  NAND U14634 ( .A(n8085), .B(n[124]), .Z(n13462) );
  NAND U14635 ( .A(n13463), .B(n[125]), .Z(n7948) );
  NAND U14636 ( .A(n8085), .B(n[125]), .Z(n13463) );
  NAND U14637 ( .A(n13464), .B(n[126]), .Z(n7943) );
  NAND U14638 ( .A(n8085), .B(n[126]), .Z(n13464) );
  NAND U14639 ( .A(n13465), .B(n[127]), .Z(n7938) );
  NAND U14640 ( .A(n8085), .B(n[127]), .Z(n13465) );
  NAND U14641 ( .A(n13466), .B(n[128]), .Z(n7933) );
  NAND U14642 ( .A(n8085), .B(n[128]), .Z(n13466) );
  NAND U14643 ( .A(n13467), .B(n[129]), .Z(n7928) );
  NAND U14644 ( .A(n8085), .B(n[129]), .Z(n13467) );
  NAND U14645 ( .A(n13468), .B(n[130]), .Z(n7918) );
  NAND U14646 ( .A(n8085), .B(n[130]), .Z(n13468) );
  NAND U14647 ( .A(n13469), .B(n[131]), .Z(n7913) );
  NAND U14648 ( .A(n8085), .B(n[131]), .Z(n13469) );
  NAND U14649 ( .A(n13470), .B(n[132]), .Z(n7908) );
  NAND U14650 ( .A(n8085), .B(n[132]), .Z(n13470) );
  NAND U14651 ( .A(n13471), .B(n[133]), .Z(n7903) );
  NAND U14652 ( .A(n8085), .B(n[133]), .Z(n13471) );
  NAND U14653 ( .A(n13472), .B(n[134]), .Z(n7898) );
  NAND U14654 ( .A(n8085), .B(n[134]), .Z(n13472) );
  NAND U14655 ( .A(n13473), .B(n[135]), .Z(n7893) );
  NAND U14656 ( .A(n8085), .B(n[135]), .Z(n13473) );
  NAND U14657 ( .A(n13474), .B(n[136]), .Z(n7888) );
  NAND U14658 ( .A(n8085), .B(n[136]), .Z(n13474) );
  NAND U14659 ( .A(n13475), .B(n[137]), .Z(n7883) );
  NAND U14660 ( .A(n8085), .B(n[137]), .Z(n13475) );
  NAND U14661 ( .A(n13476), .B(n[138]), .Z(n7878) );
  NAND U14662 ( .A(n8085), .B(n[138]), .Z(n13476) );
  NAND U14663 ( .A(n13477), .B(n[139]), .Z(n7873) );
  NAND U14664 ( .A(n8085), .B(n[139]), .Z(n13477) );
  NAND U14665 ( .A(n13478), .B(n[140]), .Z(n7863) );
  NAND U14666 ( .A(n8085), .B(n[140]), .Z(n13478) );
  NAND U14667 ( .A(n13479), .B(n[141]), .Z(n7858) );
  NAND U14668 ( .A(n8085), .B(n[141]), .Z(n13479) );
  NAND U14669 ( .A(n13480), .B(n[142]), .Z(n7853) );
  NAND U14670 ( .A(n8085), .B(n[142]), .Z(n13480) );
  NAND U14671 ( .A(n13481), .B(n[143]), .Z(n7848) );
  NAND U14672 ( .A(n8085), .B(n[143]), .Z(n13481) );
  NAND U14673 ( .A(n13482), .B(n[144]), .Z(n7843) );
  NAND U14674 ( .A(n8085), .B(n[144]), .Z(n13482) );
  NAND U14675 ( .A(n13483), .B(n[145]), .Z(n7838) );
  NAND U14676 ( .A(n8085), .B(n[145]), .Z(n13483) );
  NAND U14677 ( .A(n13484), .B(n[146]), .Z(n7833) );
  NAND U14678 ( .A(n8085), .B(n[146]), .Z(n13484) );
  NAND U14679 ( .A(n13485), .B(n[147]), .Z(n7828) );
  NAND U14680 ( .A(n8085), .B(n[147]), .Z(n13485) );
  NAND U14681 ( .A(n13486), .B(n[148]), .Z(n7823) );
  NAND U14682 ( .A(n8085), .B(n[148]), .Z(n13486) );
  NAND U14683 ( .A(n13487), .B(n[149]), .Z(n7818) );
  NAND U14684 ( .A(n8085), .B(n[149]), .Z(n13487) );
  NAND U14685 ( .A(n13488), .B(n[150]), .Z(n7808) );
  NAND U14686 ( .A(n8085), .B(n[150]), .Z(n13488) );
  NAND U14687 ( .A(n13489), .B(n[151]), .Z(n7803) );
  NAND U14688 ( .A(n8085), .B(n[151]), .Z(n13489) );
  NAND U14689 ( .A(n13490), .B(n[152]), .Z(n7798) );
  NAND U14690 ( .A(n8085), .B(n[152]), .Z(n13490) );
  NAND U14691 ( .A(n13491), .B(n[153]), .Z(n7793) );
  NAND U14692 ( .A(n8085), .B(n[153]), .Z(n13491) );
  NAND U14693 ( .A(n13492), .B(n[154]), .Z(n7788) );
  NAND U14694 ( .A(n8085), .B(n[154]), .Z(n13492) );
  NAND U14695 ( .A(n13493), .B(n[155]), .Z(n7783) );
  NAND U14696 ( .A(n8085), .B(n[155]), .Z(n13493) );
  NAND U14697 ( .A(n13494), .B(n[156]), .Z(n7778) );
  NAND U14698 ( .A(n8085), .B(n[156]), .Z(n13494) );
  NAND U14699 ( .A(n13495), .B(n[157]), .Z(n7773) );
  NAND U14700 ( .A(n8085), .B(n[157]), .Z(n13495) );
  NAND U14701 ( .A(n13496), .B(n[158]), .Z(n7768) );
  NAND U14702 ( .A(n8085), .B(n[158]), .Z(n13496) );
  NAND U14703 ( .A(n13497), .B(n[159]), .Z(n7763) );
  NAND U14704 ( .A(n8085), .B(n[159]), .Z(n13497) );
  NAND U14705 ( .A(n13498), .B(n[160]), .Z(n7753) );
  NAND U14706 ( .A(n8085), .B(n[160]), .Z(n13498) );
  NAND U14707 ( .A(n13499), .B(n[161]), .Z(n7748) );
  NAND U14708 ( .A(n8085), .B(n[161]), .Z(n13499) );
  NAND U14709 ( .A(n13500), .B(n[162]), .Z(n7743) );
  NAND U14710 ( .A(n8085), .B(n[162]), .Z(n13500) );
  NAND U14711 ( .A(n13501), .B(n[163]), .Z(n7738) );
  NAND U14712 ( .A(n8085), .B(n[163]), .Z(n13501) );
  NAND U14713 ( .A(n13502), .B(n[164]), .Z(n7733) );
  NAND U14714 ( .A(n8085), .B(n[164]), .Z(n13502) );
  NAND U14715 ( .A(n13503), .B(n[165]), .Z(n7728) );
  NAND U14716 ( .A(n8085), .B(n[165]), .Z(n13503) );
  NAND U14717 ( .A(n13504), .B(n[166]), .Z(n7723) );
  NAND U14718 ( .A(n8085), .B(n[166]), .Z(n13504) );
  NAND U14719 ( .A(n13505), .B(n[167]), .Z(n7718) );
  NAND U14720 ( .A(n8085), .B(n[167]), .Z(n13505) );
  NAND U14721 ( .A(n13506), .B(n[168]), .Z(n7713) );
  NAND U14722 ( .A(n8085), .B(n[168]), .Z(n13506) );
  NAND U14723 ( .A(n13507), .B(n[169]), .Z(n7708) );
  NAND U14724 ( .A(n8085), .B(n[169]), .Z(n13507) );
  NAND U14725 ( .A(n13508), .B(n[170]), .Z(n7698) );
  NAND U14726 ( .A(n8085), .B(n[170]), .Z(n13508) );
  NAND U14727 ( .A(n13509), .B(n[171]), .Z(n7693) );
  NAND U14728 ( .A(n8085), .B(n[171]), .Z(n13509) );
  NAND U14729 ( .A(n13510), .B(n[172]), .Z(n7688) );
  NAND U14730 ( .A(n8085), .B(n[172]), .Z(n13510) );
  NAND U14731 ( .A(n13511), .B(n[173]), .Z(n7683) );
  NAND U14732 ( .A(n8085), .B(n[173]), .Z(n13511) );
  NAND U14733 ( .A(n13512), .B(n[174]), .Z(n7678) );
  NAND U14734 ( .A(n8085), .B(n[174]), .Z(n13512) );
  NAND U14735 ( .A(n13513), .B(n[175]), .Z(n7673) );
  NAND U14736 ( .A(n8085), .B(n[175]), .Z(n13513) );
  NAND U14737 ( .A(n13514), .B(n[176]), .Z(n7668) );
  NAND U14738 ( .A(n8085), .B(n[176]), .Z(n13514) );
  NAND U14739 ( .A(n13515), .B(n[177]), .Z(n7663) );
  NAND U14740 ( .A(n8085), .B(n[177]), .Z(n13515) );
  NAND U14741 ( .A(n13516), .B(n[178]), .Z(n7658) );
  NAND U14742 ( .A(n8085), .B(n[178]), .Z(n13516) );
  NAND U14743 ( .A(n13517), .B(n[179]), .Z(n7653) );
  NAND U14744 ( .A(n8085), .B(n[179]), .Z(n13517) );
  NAND U14745 ( .A(n13518), .B(n[180]), .Z(n7643) );
  NAND U14746 ( .A(n8085), .B(n[180]), .Z(n13518) );
  NAND U14747 ( .A(n13519), .B(n[181]), .Z(n7638) );
  NAND U14748 ( .A(n8085), .B(n[181]), .Z(n13519) );
  NAND U14749 ( .A(n13520), .B(n[182]), .Z(n7633) );
  NAND U14750 ( .A(n8085), .B(n[182]), .Z(n13520) );
  NAND U14751 ( .A(n13521), .B(n[183]), .Z(n7628) );
  NAND U14752 ( .A(n8085), .B(n[183]), .Z(n13521) );
  NAND U14753 ( .A(n13522), .B(n[184]), .Z(n7623) );
  NAND U14754 ( .A(n8085), .B(n[184]), .Z(n13522) );
  NAND U14755 ( .A(n13523), .B(n[185]), .Z(n7618) );
  NAND U14756 ( .A(n8085), .B(n[185]), .Z(n13523) );
  NAND U14757 ( .A(n13524), .B(n[186]), .Z(n7613) );
  NAND U14758 ( .A(n8085), .B(n[186]), .Z(n13524) );
  NAND U14759 ( .A(n13525), .B(n[187]), .Z(n7608) );
  NAND U14760 ( .A(n8085), .B(n[187]), .Z(n13525) );
  NAND U14761 ( .A(n13526), .B(n[188]), .Z(n7603) );
  NAND U14762 ( .A(n8085), .B(n[188]), .Z(n13526) );
  NAND U14763 ( .A(n13527), .B(n[189]), .Z(n7598) );
  NAND U14764 ( .A(n8085), .B(n[189]), .Z(n13527) );
  NAND U14765 ( .A(n13528), .B(n[190]), .Z(n7588) );
  NAND U14766 ( .A(n8085), .B(n[190]), .Z(n13528) );
  NAND U14767 ( .A(n13529), .B(n[191]), .Z(n7583) );
  NAND U14768 ( .A(n8085), .B(n[191]), .Z(n13529) );
  NAND U14769 ( .A(n13530), .B(n[192]), .Z(n7578) );
  NAND U14770 ( .A(n8085), .B(n[192]), .Z(n13530) );
  NAND U14771 ( .A(n13531), .B(n[193]), .Z(n7573) );
  NAND U14772 ( .A(n8085), .B(n[193]), .Z(n13531) );
  NAND U14773 ( .A(n13532), .B(n[194]), .Z(n7568) );
  NAND U14774 ( .A(n8085), .B(n[194]), .Z(n13532) );
  NAND U14775 ( .A(n13533), .B(n[195]), .Z(n7563) );
  NAND U14776 ( .A(n8085), .B(n[195]), .Z(n13533) );
  NAND U14777 ( .A(n13534), .B(n[196]), .Z(n7558) );
  NAND U14778 ( .A(n8085), .B(n[196]), .Z(n13534) );
  NAND U14779 ( .A(n13535), .B(n[197]), .Z(n7553) );
  NAND U14780 ( .A(n8085), .B(n[197]), .Z(n13535) );
  NAND U14781 ( .A(n13536), .B(n[198]), .Z(n7548) );
  NAND U14782 ( .A(n8085), .B(n[198]), .Z(n13536) );
  NAND U14783 ( .A(n13537), .B(n[199]), .Z(n7543) );
  NAND U14784 ( .A(n8085), .B(n[199]), .Z(n13537) );
  NAND U14785 ( .A(n13538), .B(n[200]), .Z(n7528) );
  NAND U14786 ( .A(n8085), .B(n[200]), .Z(n13538) );
  NAND U14787 ( .A(n13539), .B(n[201]), .Z(n7523) );
  NAND U14788 ( .A(n8085), .B(n[201]), .Z(n13539) );
  NAND U14789 ( .A(n13540), .B(n[202]), .Z(n7518) );
  NAND U14790 ( .A(n8085), .B(n[202]), .Z(n13540) );
  NAND U14791 ( .A(n13541), .B(n[203]), .Z(n7513) );
  NAND U14792 ( .A(n8085), .B(n[203]), .Z(n13541) );
  NAND U14793 ( .A(n13542), .B(n[204]), .Z(n7508) );
  NAND U14794 ( .A(n8085), .B(n[204]), .Z(n13542) );
  NAND U14795 ( .A(n13543), .B(n[205]), .Z(n7503) );
  NAND U14796 ( .A(n8085), .B(n[205]), .Z(n13543) );
  NAND U14797 ( .A(n13544), .B(n[206]), .Z(n7498) );
  NAND U14798 ( .A(n8085), .B(n[206]), .Z(n13544) );
  NAND U14799 ( .A(n13545), .B(n[207]), .Z(n7493) );
  NAND U14800 ( .A(n8085), .B(n[207]), .Z(n13545) );
  NAND U14801 ( .A(n13546), .B(n[208]), .Z(n7488) );
  NAND U14802 ( .A(n8085), .B(n[208]), .Z(n13546) );
  NAND U14803 ( .A(n13547), .B(n[209]), .Z(n7483) );
  NAND U14804 ( .A(n8085), .B(n[209]), .Z(n13547) );
  NAND U14805 ( .A(n13548), .B(n[210]), .Z(n7473) );
  NAND U14806 ( .A(n8085), .B(n[210]), .Z(n13548) );
  NAND U14807 ( .A(n13549), .B(n[211]), .Z(n7468) );
  NAND U14808 ( .A(n8085), .B(n[211]), .Z(n13549) );
  NAND U14809 ( .A(n13550), .B(n[212]), .Z(n7463) );
  NAND U14810 ( .A(n8085), .B(n[212]), .Z(n13550) );
  NAND U14811 ( .A(n13551), .B(n[213]), .Z(n7458) );
  NAND U14812 ( .A(n8085), .B(n[213]), .Z(n13551) );
  NAND U14813 ( .A(n13552), .B(n[214]), .Z(n7453) );
  NAND U14814 ( .A(n8085), .B(n[214]), .Z(n13552) );
  NAND U14815 ( .A(n13553), .B(n[215]), .Z(n7448) );
  NAND U14816 ( .A(n8085), .B(n[215]), .Z(n13553) );
  NAND U14817 ( .A(n13554), .B(n[216]), .Z(n7443) );
  NAND U14818 ( .A(n8085), .B(n[216]), .Z(n13554) );
  NAND U14819 ( .A(n13555), .B(n[217]), .Z(n7438) );
  NAND U14820 ( .A(n8085), .B(n[217]), .Z(n13555) );
  NAND U14821 ( .A(n13556), .B(n[218]), .Z(n7433) );
  NAND U14822 ( .A(n8085), .B(n[218]), .Z(n13556) );
  NAND U14823 ( .A(n13557), .B(n[219]), .Z(n7428) );
  NAND U14824 ( .A(n8085), .B(n[219]), .Z(n13557) );
  NAND U14825 ( .A(n13558), .B(n[220]), .Z(n7418) );
  NAND U14826 ( .A(n8085), .B(n[220]), .Z(n13558) );
  NAND U14827 ( .A(n13559), .B(n[221]), .Z(n7413) );
  NAND U14828 ( .A(n8085), .B(n[221]), .Z(n13559) );
  NAND U14829 ( .A(n13560), .B(n[222]), .Z(n7408) );
  NAND U14830 ( .A(n8085), .B(n[222]), .Z(n13560) );
  NAND U14831 ( .A(n13561), .B(n[223]), .Z(n7403) );
  NAND U14832 ( .A(n8085), .B(n[223]), .Z(n13561) );
  NAND U14833 ( .A(n13562), .B(n[224]), .Z(n7398) );
  NAND U14834 ( .A(n8085), .B(n[224]), .Z(n13562) );
  NAND U14835 ( .A(n13563), .B(n[225]), .Z(n7393) );
  NAND U14836 ( .A(n8085), .B(n[225]), .Z(n13563) );
  NAND U14837 ( .A(n13564), .B(n[226]), .Z(n7388) );
  NAND U14838 ( .A(n8085), .B(n[226]), .Z(n13564) );
  NAND U14839 ( .A(n13565), .B(n[227]), .Z(n7383) );
  NAND U14840 ( .A(n8085), .B(n[227]), .Z(n13565) );
  NAND U14841 ( .A(n13566), .B(n[228]), .Z(n7378) );
  NAND U14842 ( .A(n8085), .B(n[228]), .Z(n13566) );
  NAND U14843 ( .A(n13567), .B(n[229]), .Z(n7373) );
  NAND U14844 ( .A(n8085), .B(n[229]), .Z(n13567) );
  NAND U14845 ( .A(n13568), .B(n[230]), .Z(n7363) );
  NAND U14846 ( .A(n8085), .B(n[230]), .Z(n13568) );
  NAND U14847 ( .A(n13569), .B(n[231]), .Z(n7358) );
  NAND U14848 ( .A(n8085), .B(n[231]), .Z(n13569) );
  NAND U14849 ( .A(n13570), .B(n[232]), .Z(n7353) );
  NAND U14850 ( .A(n8085), .B(n[232]), .Z(n13570) );
  NAND U14851 ( .A(n13571), .B(n[233]), .Z(n7348) );
  NAND U14852 ( .A(n8085), .B(n[233]), .Z(n13571) );
  NAND U14853 ( .A(n13572), .B(n[234]), .Z(n7343) );
  NAND U14854 ( .A(n8085), .B(n[234]), .Z(n13572) );
  NAND U14855 ( .A(n13573), .B(n[235]), .Z(n7338) );
  NAND U14856 ( .A(n8085), .B(n[235]), .Z(n13573) );
  NAND U14857 ( .A(n13574), .B(n[236]), .Z(n7333) );
  NAND U14858 ( .A(n8085), .B(n[236]), .Z(n13574) );
  NAND U14859 ( .A(n13575), .B(n[237]), .Z(n7328) );
  NAND U14860 ( .A(n8085), .B(n[237]), .Z(n13575) );
  NAND U14861 ( .A(n13576), .B(n[238]), .Z(n7323) );
  NAND U14862 ( .A(n8085), .B(n[238]), .Z(n13576) );
  NAND U14863 ( .A(n13577), .B(n[239]), .Z(n7318) );
  NAND U14864 ( .A(n8085), .B(n[239]), .Z(n13577) );
  NAND U14865 ( .A(n13578), .B(n[240]), .Z(n7308) );
  NAND U14866 ( .A(n8085), .B(n[240]), .Z(n13578) );
  NAND U14867 ( .A(n13579), .B(n[241]), .Z(n7303) );
  NAND U14868 ( .A(n8085), .B(n[241]), .Z(n13579) );
  NAND U14869 ( .A(n13580), .B(n[242]), .Z(n7298) );
  NAND U14870 ( .A(n8085), .B(n[242]), .Z(n13580) );
  NAND U14871 ( .A(n13581), .B(n[243]), .Z(n7293) );
  NAND U14872 ( .A(n8085), .B(n[243]), .Z(n13581) );
  NAND U14873 ( .A(n13582), .B(n[244]), .Z(n7288) );
  NAND U14874 ( .A(n8085), .B(n[244]), .Z(n13582) );
  NAND U14875 ( .A(n13583), .B(n[245]), .Z(n7283) );
  NAND U14876 ( .A(n8085), .B(n[245]), .Z(n13583) );
  NAND U14877 ( .A(n13584), .B(n[246]), .Z(n7278) );
  NAND U14878 ( .A(n8085), .B(n[246]), .Z(n13584) );
  NAND U14879 ( .A(n13585), .B(n[247]), .Z(n7273) );
  NAND U14880 ( .A(n8085), .B(n[247]), .Z(n13585) );
  NAND U14881 ( .A(n13586), .B(n[248]), .Z(n7268) );
  NAND U14882 ( .A(n8085), .B(n[248]), .Z(n13586) );
  NAND U14883 ( .A(n13587), .B(n[249]), .Z(n7263) );
  NAND U14884 ( .A(n8085), .B(n[249]), .Z(n13587) );
  NAND U14885 ( .A(n13588), .B(n[250]), .Z(n7253) );
  NAND U14886 ( .A(n8085), .B(n[250]), .Z(n13588) );
  NAND U14887 ( .A(n13589), .B(n[251]), .Z(n7248) );
  NAND U14888 ( .A(n8085), .B(n[251]), .Z(n13589) );
  NAND U14889 ( .A(n13590), .B(n[252]), .Z(n7243) );
  NAND U14890 ( .A(n8085), .B(n[252]), .Z(n13590) );
  NAND U14891 ( .A(n13591), .B(n[253]), .Z(n7238) );
  NAND U14892 ( .A(n8085), .B(n[253]), .Z(n13591) );
  NAND U14893 ( .A(n13592), .B(n[254]), .Z(n7233) );
  NAND U14894 ( .A(n8085), .B(n[254]), .Z(n13592) );
  NAND U14895 ( .A(n13593), .B(n[255]), .Z(n7228) );
  NAND U14896 ( .A(n8085), .B(n[255]), .Z(n13593) );
  NAND U14897 ( .A(n13594), .B(n[256]), .Z(n7223) );
  NAND U14898 ( .A(n8085), .B(n[256]), .Z(n13594) );
  NAND U14899 ( .A(n13595), .B(n[257]), .Z(n7218) );
  NAND U14900 ( .A(n8085), .B(n[257]), .Z(n13595) );
  NAND U14901 ( .A(n13596), .B(n[258]), .Z(n7213) );
  NAND U14902 ( .A(n8085), .B(n[258]), .Z(n13596) );
  NAND U14903 ( .A(n13597), .B(n[259]), .Z(n7208) );
  NAND U14904 ( .A(n8085), .B(n[259]), .Z(n13597) );
  NAND U14905 ( .A(n13598), .B(n[260]), .Z(n7198) );
  NAND U14906 ( .A(n8085), .B(n[260]), .Z(n13598) );
  NAND U14907 ( .A(n13599), .B(n[261]), .Z(n7193) );
  NAND U14908 ( .A(n8085), .B(n[261]), .Z(n13599) );
  NAND U14909 ( .A(n13600), .B(n[262]), .Z(n7188) );
  NAND U14910 ( .A(n8085), .B(n[262]), .Z(n13600) );
  NAND U14911 ( .A(n13601), .B(n[263]), .Z(n7183) );
  NAND U14912 ( .A(n8085), .B(n[263]), .Z(n13601) );
  NAND U14913 ( .A(n13602), .B(n[264]), .Z(n7178) );
  NAND U14914 ( .A(n8085), .B(n[264]), .Z(n13602) );
  NAND U14915 ( .A(n13603), .B(n[265]), .Z(n7173) );
  NAND U14916 ( .A(n8085), .B(n[265]), .Z(n13603) );
  NAND U14917 ( .A(n13604), .B(n[266]), .Z(n7168) );
  NAND U14918 ( .A(n8085), .B(n[266]), .Z(n13604) );
  NAND U14919 ( .A(n13605), .B(n[267]), .Z(n7163) );
  NAND U14920 ( .A(n8085), .B(n[267]), .Z(n13605) );
  NAND U14921 ( .A(n13606), .B(n[268]), .Z(n7158) );
  NAND U14922 ( .A(n8085), .B(n[268]), .Z(n13606) );
  NAND U14923 ( .A(n13607), .B(n[269]), .Z(n7153) );
  NAND U14924 ( .A(n8085), .B(n[269]), .Z(n13607) );
  NAND U14925 ( .A(n13608), .B(n[270]), .Z(n7143) );
  NAND U14926 ( .A(n8085), .B(n[270]), .Z(n13608) );
  NAND U14927 ( .A(n13609), .B(n[271]), .Z(n7138) );
  NAND U14928 ( .A(n8085), .B(n[271]), .Z(n13609) );
  NAND U14929 ( .A(n13610), .B(n[272]), .Z(n7133) );
  NAND U14930 ( .A(n8085), .B(n[272]), .Z(n13610) );
  NAND U14931 ( .A(n13611), .B(n[273]), .Z(n7128) );
  NAND U14932 ( .A(n8085), .B(n[273]), .Z(n13611) );
  NAND U14933 ( .A(n13612), .B(n[274]), .Z(n7123) );
  NAND U14934 ( .A(n8085), .B(n[274]), .Z(n13612) );
  NAND U14935 ( .A(n13613), .B(n[275]), .Z(n7118) );
  NAND U14936 ( .A(n8085), .B(n[275]), .Z(n13613) );
  NAND U14937 ( .A(n13614), .B(n[276]), .Z(n7113) );
  NAND U14938 ( .A(n8085), .B(n[276]), .Z(n13614) );
  NAND U14939 ( .A(n13615), .B(n[277]), .Z(n7108) );
  NAND U14940 ( .A(n8085), .B(n[277]), .Z(n13615) );
  NAND U14941 ( .A(n13616), .B(n[278]), .Z(n7103) );
  NAND U14942 ( .A(n8085), .B(n[278]), .Z(n13616) );
  NAND U14943 ( .A(n13617), .B(n[279]), .Z(n7098) );
  NAND U14944 ( .A(n8085), .B(n[279]), .Z(n13617) );
  NAND U14945 ( .A(n13618), .B(n[280]), .Z(n7088) );
  NAND U14946 ( .A(n8085), .B(n[280]), .Z(n13618) );
  NAND U14947 ( .A(n13619), .B(n[281]), .Z(n7083) );
  NAND U14948 ( .A(n8085), .B(n[281]), .Z(n13619) );
  NAND U14949 ( .A(n13620), .B(n[282]), .Z(n7078) );
  NAND U14950 ( .A(n8085), .B(n[282]), .Z(n13620) );
  NAND U14951 ( .A(n13621), .B(n[283]), .Z(n7073) );
  NAND U14952 ( .A(n8085), .B(n[283]), .Z(n13621) );
  NAND U14953 ( .A(n13622), .B(n[284]), .Z(n7068) );
  NAND U14954 ( .A(n8085), .B(n[284]), .Z(n13622) );
  NAND U14955 ( .A(n13623), .B(n[285]), .Z(n7063) );
  NAND U14956 ( .A(n8085), .B(n[285]), .Z(n13623) );
  NAND U14957 ( .A(n13624), .B(n[286]), .Z(n7058) );
  NAND U14958 ( .A(n8085), .B(n[286]), .Z(n13624) );
  NAND U14959 ( .A(n13625), .B(n[287]), .Z(n7053) );
  NAND U14960 ( .A(n8085), .B(n[287]), .Z(n13625) );
  NAND U14961 ( .A(n13626), .B(n[288]), .Z(n7048) );
  NAND U14962 ( .A(n8085), .B(n[288]), .Z(n13626) );
  NAND U14963 ( .A(n13627), .B(n[289]), .Z(n7043) );
  NAND U14964 ( .A(n8085), .B(n[289]), .Z(n13627) );
  NAND U14965 ( .A(n13628), .B(n[290]), .Z(n7033) );
  NAND U14966 ( .A(n8085), .B(n[290]), .Z(n13628) );
  NAND U14967 ( .A(n13629), .B(n[291]), .Z(n7028) );
  NAND U14968 ( .A(n8085), .B(n[291]), .Z(n13629) );
  NAND U14969 ( .A(n13630), .B(n[292]), .Z(n7023) );
  NAND U14970 ( .A(n8085), .B(n[292]), .Z(n13630) );
  NAND U14971 ( .A(n13631), .B(n[293]), .Z(n7018) );
  NAND U14972 ( .A(n8085), .B(n[293]), .Z(n13631) );
  NAND U14973 ( .A(n13632), .B(n[294]), .Z(n7013) );
  NAND U14974 ( .A(n8085), .B(n[294]), .Z(n13632) );
  NAND U14975 ( .A(n13633), .B(n[295]), .Z(n7008) );
  NAND U14976 ( .A(n8085), .B(n[295]), .Z(n13633) );
  NAND U14977 ( .A(n13634), .B(n[296]), .Z(n7003) );
  NAND U14978 ( .A(n8085), .B(n[296]), .Z(n13634) );
  NAND U14979 ( .A(n13635), .B(n[297]), .Z(n6998) );
  NAND U14980 ( .A(n8085), .B(n[297]), .Z(n13635) );
  NAND U14981 ( .A(n13636), .B(n[298]), .Z(n6993) );
  NAND U14982 ( .A(n8085), .B(n[298]), .Z(n13636) );
  NAND U14983 ( .A(n13637), .B(n[299]), .Z(n6988) );
  NAND U14984 ( .A(n8085), .B(n[299]), .Z(n13637) );
  NAND U14985 ( .A(n13638), .B(n[300]), .Z(n6973) );
  NAND U14986 ( .A(n8085), .B(n[300]), .Z(n13638) );
  NAND U14987 ( .A(n13639), .B(n[301]), .Z(n6968) );
  NAND U14988 ( .A(n8085), .B(n[301]), .Z(n13639) );
  NAND U14989 ( .A(n13640), .B(n[302]), .Z(n6963) );
  NAND U14990 ( .A(n8085), .B(n[302]), .Z(n13640) );
  NAND U14991 ( .A(n13641), .B(n[303]), .Z(n6958) );
  NAND U14992 ( .A(n8085), .B(n[303]), .Z(n13641) );
  NAND U14993 ( .A(n13642), .B(n[304]), .Z(n6953) );
  NAND U14994 ( .A(n8085), .B(n[304]), .Z(n13642) );
  NAND U14995 ( .A(n13643), .B(n[305]), .Z(n6948) );
  NAND U14996 ( .A(n8085), .B(n[305]), .Z(n13643) );
  NAND U14997 ( .A(n13644), .B(n[306]), .Z(n6943) );
  NAND U14998 ( .A(n8085), .B(n[306]), .Z(n13644) );
  NAND U14999 ( .A(n13645), .B(n[307]), .Z(n6938) );
  NAND U15000 ( .A(n8085), .B(n[307]), .Z(n13645) );
  NAND U15001 ( .A(n13646), .B(n[308]), .Z(n6933) );
  NAND U15002 ( .A(n8085), .B(n[308]), .Z(n13646) );
  NAND U15003 ( .A(n13647), .B(n[309]), .Z(n6928) );
  NAND U15004 ( .A(n8085), .B(n[309]), .Z(n13647) );
  NAND U15005 ( .A(n13648), .B(n[310]), .Z(n6918) );
  NAND U15006 ( .A(n8085), .B(n[310]), .Z(n13648) );
  NAND U15007 ( .A(n13649), .B(n[311]), .Z(n6913) );
  NAND U15008 ( .A(n8085), .B(n[311]), .Z(n13649) );
  NAND U15009 ( .A(n13650), .B(n[312]), .Z(n6908) );
  NAND U15010 ( .A(n8085), .B(n[312]), .Z(n13650) );
  NAND U15011 ( .A(n13651), .B(n[313]), .Z(n6903) );
  NAND U15012 ( .A(n8085), .B(n[313]), .Z(n13651) );
  NAND U15013 ( .A(n13652), .B(n[314]), .Z(n6898) );
  NAND U15014 ( .A(n8085), .B(n[314]), .Z(n13652) );
  NAND U15015 ( .A(n13653), .B(n[315]), .Z(n6893) );
  NAND U15016 ( .A(n8085), .B(n[315]), .Z(n13653) );
  NAND U15017 ( .A(n13654), .B(n[316]), .Z(n6888) );
  NAND U15018 ( .A(n8085), .B(n[316]), .Z(n13654) );
  NAND U15019 ( .A(n13655), .B(n[317]), .Z(n6883) );
  NAND U15020 ( .A(n8085), .B(n[317]), .Z(n13655) );
  NAND U15021 ( .A(n13656), .B(n[318]), .Z(n6878) );
  NAND U15022 ( .A(n8085), .B(n[318]), .Z(n13656) );
  NAND U15023 ( .A(n13657), .B(n[319]), .Z(n6873) );
  NAND U15024 ( .A(n8085), .B(n[319]), .Z(n13657) );
  NAND U15025 ( .A(n13658), .B(n[320]), .Z(n6863) );
  NAND U15026 ( .A(n8085), .B(n[320]), .Z(n13658) );
  NAND U15027 ( .A(n13659), .B(n[321]), .Z(n6858) );
  NAND U15028 ( .A(n8085), .B(n[321]), .Z(n13659) );
  NAND U15029 ( .A(n13660), .B(n[322]), .Z(n6853) );
  NAND U15030 ( .A(n8085), .B(n[322]), .Z(n13660) );
  NAND U15031 ( .A(n13661), .B(n[323]), .Z(n6848) );
  NAND U15032 ( .A(n8085), .B(n[323]), .Z(n13661) );
  NAND U15033 ( .A(n13662), .B(n[324]), .Z(n6843) );
  NAND U15034 ( .A(n8085), .B(n[324]), .Z(n13662) );
  NAND U15035 ( .A(n13663), .B(n[325]), .Z(n6838) );
  NAND U15036 ( .A(n8085), .B(n[325]), .Z(n13663) );
  NAND U15037 ( .A(n13664), .B(n[326]), .Z(n6833) );
  NAND U15038 ( .A(n8085), .B(n[326]), .Z(n13664) );
  NAND U15039 ( .A(n13665), .B(n[327]), .Z(n6828) );
  NAND U15040 ( .A(n8085), .B(n[327]), .Z(n13665) );
  NAND U15041 ( .A(n13666), .B(n[328]), .Z(n6823) );
  NAND U15042 ( .A(n8085), .B(n[328]), .Z(n13666) );
  NAND U15043 ( .A(n13667), .B(n[329]), .Z(n6818) );
  NAND U15044 ( .A(n8085), .B(n[329]), .Z(n13667) );
  NAND U15045 ( .A(n13668), .B(n[330]), .Z(n6808) );
  NAND U15046 ( .A(n8085), .B(n[330]), .Z(n13668) );
  NAND U15047 ( .A(n13669), .B(n[331]), .Z(n6803) );
  NAND U15048 ( .A(n8085), .B(n[331]), .Z(n13669) );
  NAND U15049 ( .A(n13670), .B(n[332]), .Z(n6798) );
  NAND U15050 ( .A(n8085), .B(n[332]), .Z(n13670) );
  NAND U15051 ( .A(n13671), .B(n[333]), .Z(n6793) );
  NAND U15052 ( .A(n8085), .B(n[333]), .Z(n13671) );
  NAND U15053 ( .A(n13672), .B(n[334]), .Z(n6788) );
  NAND U15054 ( .A(n8085), .B(n[334]), .Z(n13672) );
  NAND U15055 ( .A(n13673), .B(n[335]), .Z(n6783) );
  NAND U15056 ( .A(n8085), .B(n[335]), .Z(n13673) );
  NAND U15057 ( .A(n13674), .B(n[336]), .Z(n6778) );
  NAND U15058 ( .A(n8085), .B(n[336]), .Z(n13674) );
  NAND U15059 ( .A(n13675), .B(n[337]), .Z(n6773) );
  NAND U15060 ( .A(n8085), .B(n[337]), .Z(n13675) );
  NAND U15061 ( .A(n13676), .B(n[338]), .Z(n6768) );
  NAND U15062 ( .A(n8085), .B(n[338]), .Z(n13676) );
  NAND U15063 ( .A(n13677), .B(n[339]), .Z(n6763) );
  NAND U15064 ( .A(n8085), .B(n[339]), .Z(n13677) );
  NAND U15065 ( .A(n13678), .B(n[340]), .Z(n6753) );
  NAND U15066 ( .A(n8085), .B(n[340]), .Z(n13678) );
  NAND U15067 ( .A(n13679), .B(n[341]), .Z(n6748) );
  NAND U15068 ( .A(n8085), .B(n[341]), .Z(n13679) );
  NAND U15069 ( .A(n13680), .B(n[342]), .Z(n6743) );
  NAND U15070 ( .A(n8085), .B(n[342]), .Z(n13680) );
  NAND U15071 ( .A(n13681), .B(n[343]), .Z(n6738) );
  NAND U15072 ( .A(n8085), .B(n[343]), .Z(n13681) );
  NAND U15073 ( .A(n13682), .B(n[344]), .Z(n6733) );
  NAND U15074 ( .A(n8085), .B(n[344]), .Z(n13682) );
  NAND U15075 ( .A(n13683), .B(n[345]), .Z(n6728) );
  NAND U15076 ( .A(n8085), .B(n[345]), .Z(n13683) );
  NAND U15077 ( .A(n13684), .B(n[346]), .Z(n6723) );
  NAND U15078 ( .A(n8085), .B(n[346]), .Z(n13684) );
  NAND U15079 ( .A(n13685), .B(n[347]), .Z(n6718) );
  NAND U15080 ( .A(n8085), .B(n[347]), .Z(n13685) );
  NAND U15081 ( .A(n13686), .B(n[348]), .Z(n6713) );
  NAND U15082 ( .A(n8085), .B(n[348]), .Z(n13686) );
  NAND U15083 ( .A(n13687), .B(n[349]), .Z(n6708) );
  NAND U15084 ( .A(n8085), .B(n[349]), .Z(n13687) );
  NAND U15085 ( .A(n13688), .B(n[350]), .Z(n6698) );
  NAND U15086 ( .A(n8085), .B(n[350]), .Z(n13688) );
  NAND U15087 ( .A(n13689), .B(n[351]), .Z(n6693) );
  NAND U15088 ( .A(n8085), .B(n[351]), .Z(n13689) );
  NAND U15089 ( .A(n13690), .B(n[352]), .Z(n6688) );
  NAND U15090 ( .A(n8085), .B(n[352]), .Z(n13690) );
  NAND U15091 ( .A(n13691), .B(n[353]), .Z(n6683) );
  NAND U15092 ( .A(n8085), .B(n[353]), .Z(n13691) );
  NAND U15093 ( .A(n13692), .B(n[354]), .Z(n6678) );
  NAND U15094 ( .A(n8085), .B(n[354]), .Z(n13692) );
  NAND U15095 ( .A(n13693), .B(n[355]), .Z(n6673) );
  NAND U15096 ( .A(n8085), .B(n[355]), .Z(n13693) );
  NAND U15097 ( .A(n13694), .B(n[356]), .Z(n6668) );
  NAND U15098 ( .A(n8085), .B(n[356]), .Z(n13694) );
  NAND U15099 ( .A(n13695), .B(n[357]), .Z(n6663) );
  NAND U15100 ( .A(n8085), .B(n[357]), .Z(n13695) );
  NAND U15101 ( .A(n13696), .B(n[358]), .Z(n6658) );
  NAND U15102 ( .A(n8085), .B(n[358]), .Z(n13696) );
  NAND U15103 ( .A(n13697), .B(n[359]), .Z(n6653) );
  NAND U15104 ( .A(n8085), .B(n[359]), .Z(n13697) );
  NAND U15105 ( .A(n13698), .B(n[360]), .Z(n6643) );
  NAND U15106 ( .A(n8085), .B(n[360]), .Z(n13698) );
  NAND U15107 ( .A(n13699), .B(n[361]), .Z(n6638) );
  NAND U15108 ( .A(n8085), .B(n[361]), .Z(n13699) );
  NAND U15109 ( .A(n13700), .B(n[362]), .Z(n6633) );
  NAND U15110 ( .A(n8085), .B(n[362]), .Z(n13700) );
  NAND U15111 ( .A(n13701), .B(n[363]), .Z(n6628) );
  NAND U15112 ( .A(n8085), .B(n[363]), .Z(n13701) );
  NAND U15113 ( .A(n13702), .B(n[364]), .Z(n6623) );
  NAND U15114 ( .A(n8085), .B(n[364]), .Z(n13702) );
  NAND U15115 ( .A(n13703), .B(n[365]), .Z(n6618) );
  NAND U15116 ( .A(n8085), .B(n[365]), .Z(n13703) );
  NAND U15117 ( .A(n13704), .B(n[366]), .Z(n6613) );
  NAND U15118 ( .A(n8085), .B(n[366]), .Z(n13704) );
  NAND U15119 ( .A(n13705), .B(n[367]), .Z(n6608) );
  NAND U15120 ( .A(n8085), .B(n[367]), .Z(n13705) );
  NAND U15121 ( .A(n13706), .B(n[368]), .Z(n6603) );
  NAND U15122 ( .A(n8085), .B(n[368]), .Z(n13706) );
  NAND U15123 ( .A(n13707), .B(n[369]), .Z(n6598) );
  NAND U15124 ( .A(n8085), .B(n[369]), .Z(n13707) );
  NAND U15125 ( .A(n13708), .B(n[370]), .Z(n6588) );
  NAND U15126 ( .A(n8085), .B(n[370]), .Z(n13708) );
  NAND U15127 ( .A(n13709), .B(n[371]), .Z(n6583) );
  NAND U15128 ( .A(n8085), .B(n[371]), .Z(n13709) );
  NAND U15129 ( .A(n13710), .B(n[372]), .Z(n6578) );
  NAND U15130 ( .A(n8085), .B(n[372]), .Z(n13710) );
  NAND U15131 ( .A(n13711), .B(n[373]), .Z(n6573) );
  NAND U15132 ( .A(n8085), .B(n[373]), .Z(n13711) );
  NAND U15133 ( .A(n13712), .B(n[374]), .Z(n6568) );
  NAND U15134 ( .A(n8085), .B(n[374]), .Z(n13712) );
  NAND U15135 ( .A(n13713), .B(n[375]), .Z(n6563) );
  NAND U15136 ( .A(n8085), .B(n[375]), .Z(n13713) );
  NAND U15137 ( .A(n13714), .B(n[376]), .Z(n6558) );
  NAND U15138 ( .A(n8085), .B(n[376]), .Z(n13714) );
  NAND U15139 ( .A(n13715), .B(n[377]), .Z(n6553) );
  NAND U15140 ( .A(n8085), .B(n[377]), .Z(n13715) );
  NAND U15141 ( .A(n13716), .B(n[378]), .Z(n6548) );
  NAND U15142 ( .A(n8085), .B(n[378]), .Z(n13716) );
  NAND U15143 ( .A(n13717), .B(n[379]), .Z(n6543) );
  NAND U15144 ( .A(n8085), .B(n[379]), .Z(n13717) );
  NAND U15145 ( .A(n13718), .B(n[380]), .Z(n6533) );
  NAND U15146 ( .A(n8085), .B(n[380]), .Z(n13718) );
  NAND U15147 ( .A(n13719), .B(n[381]), .Z(n6528) );
  NAND U15148 ( .A(n8085), .B(n[381]), .Z(n13719) );
  NAND U15149 ( .A(n13720), .B(n[382]), .Z(n6523) );
  NAND U15150 ( .A(n8085), .B(n[382]), .Z(n13720) );
  NAND U15151 ( .A(n13721), .B(n[383]), .Z(n6518) );
  NAND U15152 ( .A(n8085), .B(n[383]), .Z(n13721) );
  NAND U15153 ( .A(n13722), .B(n[384]), .Z(n6513) );
  NAND U15154 ( .A(n8085), .B(n[384]), .Z(n13722) );
  NAND U15155 ( .A(n13723), .B(n[385]), .Z(n6508) );
  NAND U15156 ( .A(n8085), .B(n[385]), .Z(n13723) );
  NAND U15157 ( .A(n13724), .B(n[386]), .Z(n6503) );
  NAND U15158 ( .A(n8085), .B(n[386]), .Z(n13724) );
  NAND U15159 ( .A(n13725), .B(n[387]), .Z(n6498) );
  NAND U15160 ( .A(n8085), .B(n[387]), .Z(n13725) );
  NAND U15161 ( .A(n13726), .B(n[388]), .Z(n6493) );
  NAND U15162 ( .A(n8085), .B(n[388]), .Z(n13726) );
  NAND U15163 ( .A(n13727), .B(n[389]), .Z(n6488) );
  NAND U15164 ( .A(n8085), .B(n[389]), .Z(n13727) );
  NAND U15165 ( .A(n13728), .B(n[390]), .Z(n6478) );
  NAND U15166 ( .A(n8085), .B(n[390]), .Z(n13728) );
  NAND U15167 ( .A(n13729), .B(n[391]), .Z(n6473) );
  NAND U15168 ( .A(n8085), .B(n[391]), .Z(n13729) );
  NAND U15169 ( .A(n13730), .B(n[392]), .Z(n6468) );
  NAND U15170 ( .A(n8085), .B(n[392]), .Z(n13730) );
  NAND U15171 ( .A(n13731), .B(n[393]), .Z(n6463) );
  NAND U15172 ( .A(n8085), .B(n[393]), .Z(n13731) );
  NAND U15173 ( .A(n13732), .B(n[394]), .Z(n6458) );
  NAND U15174 ( .A(n8085), .B(n[394]), .Z(n13732) );
  NAND U15175 ( .A(n13733), .B(n[395]), .Z(n6453) );
  NAND U15176 ( .A(n8085), .B(n[395]), .Z(n13733) );
  NAND U15177 ( .A(n13734), .B(n[396]), .Z(n6448) );
  NAND U15178 ( .A(n8085), .B(n[396]), .Z(n13734) );
  NAND U15179 ( .A(n13735), .B(n[397]), .Z(n6443) );
  NAND U15180 ( .A(n8085), .B(n[397]), .Z(n13735) );
  NAND U15181 ( .A(n13736), .B(n[398]), .Z(n6438) );
  NAND U15182 ( .A(n8085), .B(n[398]), .Z(n13736) );
  NAND U15183 ( .A(n13737), .B(n[399]), .Z(n6433) );
  NAND U15184 ( .A(n8085), .B(n[399]), .Z(n13737) );
  NAND U15185 ( .A(n13738), .B(n[400]), .Z(n6418) );
  NAND U15186 ( .A(n8085), .B(n[400]), .Z(n13738) );
  NAND U15187 ( .A(n13739), .B(n[401]), .Z(n6413) );
  NAND U15188 ( .A(n8085), .B(n[401]), .Z(n13739) );
  NAND U15189 ( .A(n13740), .B(n[402]), .Z(n6408) );
  NAND U15190 ( .A(n8085), .B(n[402]), .Z(n13740) );
  NAND U15191 ( .A(n13741), .B(n[403]), .Z(n6403) );
  NAND U15192 ( .A(n8085), .B(n[403]), .Z(n13741) );
  NAND U15193 ( .A(n13742), .B(n[404]), .Z(n6398) );
  NAND U15194 ( .A(n8085), .B(n[404]), .Z(n13742) );
  NAND U15195 ( .A(n13743), .B(n[405]), .Z(n6393) );
  NAND U15196 ( .A(n8085), .B(n[405]), .Z(n13743) );
  NAND U15197 ( .A(n13744), .B(n[406]), .Z(n6388) );
  NAND U15198 ( .A(n8085), .B(n[406]), .Z(n13744) );
  NAND U15199 ( .A(n13745), .B(n[407]), .Z(n6383) );
  NAND U15200 ( .A(n8085), .B(n[407]), .Z(n13745) );
  NAND U15201 ( .A(n13746), .B(n[408]), .Z(n6378) );
  NAND U15202 ( .A(n8085), .B(n[408]), .Z(n13746) );
  NAND U15203 ( .A(n13747), .B(n[409]), .Z(n6373) );
  NAND U15204 ( .A(n8085), .B(n[409]), .Z(n13747) );
  NAND U15205 ( .A(n13748), .B(n[410]), .Z(n6363) );
  NAND U15206 ( .A(n8085), .B(n[410]), .Z(n13748) );
  NAND U15207 ( .A(n13749), .B(n[411]), .Z(n6358) );
  NAND U15208 ( .A(n8085), .B(n[411]), .Z(n13749) );
  NAND U15209 ( .A(n13750), .B(n[412]), .Z(n6353) );
  NAND U15210 ( .A(n8085), .B(n[412]), .Z(n13750) );
  NAND U15211 ( .A(n13751), .B(n[413]), .Z(n6348) );
  NAND U15212 ( .A(n8085), .B(n[413]), .Z(n13751) );
  NAND U15213 ( .A(n13752), .B(n[414]), .Z(n6343) );
  NAND U15214 ( .A(n8085), .B(n[414]), .Z(n13752) );
  NAND U15215 ( .A(n13753), .B(n[415]), .Z(n6338) );
  NAND U15216 ( .A(n8085), .B(n[415]), .Z(n13753) );
  NAND U15217 ( .A(n13754), .B(n[416]), .Z(n6333) );
  NAND U15218 ( .A(n8085), .B(n[416]), .Z(n13754) );
  NAND U15219 ( .A(n13755), .B(n[417]), .Z(n6328) );
  NAND U15220 ( .A(n8085), .B(n[417]), .Z(n13755) );
  NAND U15221 ( .A(n13756), .B(n[418]), .Z(n6323) );
  NAND U15222 ( .A(n8085), .B(n[418]), .Z(n13756) );
  NAND U15223 ( .A(n13757), .B(n[419]), .Z(n6318) );
  NAND U15224 ( .A(n8085), .B(n[419]), .Z(n13757) );
  NAND U15225 ( .A(n13758), .B(n[420]), .Z(n6308) );
  NAND U15226 ( .A(n8085), .B(n[420]), .Z(n13758) );
  NAND U15227 ( .A(n13759), .B(n[421]), .Z(n6303) );
  NAND U15228 ( .A(n8085), .B(n[421]), .Z(n13759) );
  NAND U15229 ( .A(n13760), .B(n[422]), .Z(n6298) );
  NAND U15230 ( .A(n8085), .B(n[422]), .Z(n13760) );
  NAND U15231 ( .A(n13761), .B(n[423]), .Z(n6293) );
  NAND U15232 ( .A(n8085), .B(n[423]), .Z(n13761) );
  NAND U15233 ( .A(n13762), .B(n[424]), .Z(n6288) );
  NAND U15234 ( .A(n8085), .B(n[424]), .Z(n13762) );
  NAND U15235 ( .A(n13763), .B(n[425]), .Z(n6283) );
  NAND U15236 ( .A(n8085), .B(n[425]), .Z(n13763) );
  NAND U15237 ( .A(n13764), .B(n[426]), .Z(n6278) );
  NAND U15238 ( .A(n8085), .B(n[426]), .Z(n13764) );
  NAND U15239 ( .A(n13765), .B(n[427]), .Z(n6273) );
  NAND U15240 ( .A(n8085), .B(n[427]), .Z(n13765) );
  NAND U15241 ( .A(n13766), .B(n[428]), .Z(n6268) );
  NAND U15242 ( .A(n8085), .B(n[428]), .Z(n13766) );
  NAND U15243 ( .A(n13767), .B(n[429]), .Z(n6263) );
  NAND U15244 ( .A(n8085), .B(n[429]), .Z(n13767) );
  NAND U15245 ( .A(n13768), .B(n[430]), .Z(n6253) );
  NAND U15246 ( .A(n8085), .B(n[430]), .Z(n13768) );
  NAND U15247 ( .A(n13769), .B(n[431]), .Z(n6248) );
  NAND U15248 ( .A(n8085), .B(n[431]), .Z(n13769) );
  NAND U15249 ( .A(n13770), .B(n[432]), .Z(n6243) );
  NAND U15250 ( .A(n8085), .B(n[432]), .Z(n13770) );
  NAND U15251 ( .A(n13771), .B(n[433]), .Z(n6238) );
  NAND U15252 ( .A(n8085), .B(n[433]), .Z(n13771) );
  NAND U15253 ( .A(n13772), .B(n[434]), .Z(n6233) );
  NAND U15254 ( .A(n8085), .B(n[434]), .Z(n13772) );
  NAND U15255 ( .A(n13773), .B(n[435]), .Z(n6228) );
  NAND U15256 ( .A(n8085), .B(n[435]), .Z(n13773) );
  NAND U15257 ( .A(n13774), .B(n[436]), .Z(n6223) );
  NAND U15258 ( .A(n8085), .B(n[436]), .Z(n13774) );
  NAND U15259 ( .A(n13775), .B(n[437]), .Z(n6218) );
  NAND U15260 ( .A(n8085), .B(n[437]), .Z(n13775) );
  NAND U15261 ( .A(n13776), .B(n[438]), .Z(n6213) );
  NAND U15262 ( .A(n8085), .B(n[438]), .Z(n13776) );
  NAND U15263 ( .A(n13777), .B(n[439]), .Z(n6208) );
  NAND U15264 ( .A(n8085), .B(n[439]), .Z(n13777) );
  NAND U15265 ( .A(n13778), .B(n[440]), .Z(n6198) );
  NAND U15266 ( .A(n8085), .B(n[440]), .Z(n13778) );
  NAND U15267 ( .A(n13779), .B(n[441]), .Z(n6193) );
  NAND U15268 ( .A(n8085), .B(n[441]), .Z(n13779) );
  NAND U15269 ( .A(n13780), .B(n[442]), .Z(n6188) );
  NAND U15270 ( .A(n8085), .B(n[442]), .Z(n13780) );
  NAND U15271 ( .A(n13781), .B(n[443]), .Z(n6183) );
  NAND U15272 ( .A(n8085), .B(n[443]), .Z(n13781) );
  NAND U15273 ( .A(n13782), .B(n[444]), .Z(n6178) );
  NAND U15274 ( .A(n8085), .B(n[444]), .Z(n13782) );
  NAND U15275 ( .A(n13783), .B(n[445]), .Z(n6173) );
  NAND U15276 ( .A(n8085), .B(n[445]), .Z(n13783) );
  NAND U15277 ( .A(n13784), .B(n[446]), .Z(n6168) );
  NAND U15278 ( .A(n8085), .B(n[446]), .Z(n13784) );
  NAND U15279 ( .A(n13785), .B(n[447]), .Z(n6163) );
  NAND U15280 ( .A(n8085), .B(n[447]), .Z(n13785) );
  NAND U15281 ( .A(n13786), .B(n[448]), .Z(n6158) );
  NAND U15282 ( .A(n8085), .B(n[448]), .Z(n13786) );
  NAND U15283 ( .A(n13787), .B(n[449]), .Z(n6153) );
  NAND U15284 ( .A(n8085), .B(n[449]), .Z(n13787) );
  NAND U15285 ( .A(n13788), .B(n[450]), .Z(n6143) );
  NAND U15286 ( .A(n8085), .B(n[450]), .Z(n13788) );
  NAND U15287 ( .A(n13789), .B(n[451]), .Z(n6138) );
  NAND U15288 ( .A(n8085), .B(n[451]), .Z(n13789) );
  NAND U15289 ( .A(n13790), .B(n[452]), .Z(n6133) );
  NAND U15290 ( .A(n8085), .B(n[452]), .Z(n13790) );
  NAND U15291 ( .A(n13791), .B(n[453]), .Z(n6128) );
  NAND U15292 ( .A(n8085), .B(n[453]), .Z(n13791) );
  NAND U15293 ( .A(n13792), .B(n[454]), .Z(n6123) );
  NAND U15294 ( .A(n8085), .B(n[454]), .Z(n13792) );
  NAND U15295 ( .A(n13793), .B(n[455]), .Z(n6118) );
  NAND U15296 ( .A(n8085), .B(n[455]), .Z(n13793) );
  NAND U15297 ( .A(n13794), .B(n[456]), .Z(n6113) );
  NAND U15298 ( .A(n8085), .B(n[456]), .Z(n13794) );
  NAND U15299 ( .A(n13795), .B(n[457]), .Z(n6108) );
  NAND U15300 ( .A(n8085), .B(n[457]), .Z(n13795) );
  NAND U15301 ( .A(n13796), .B(n[458]), .Z(n6103) );
  NAND U15302 ( .A(n8085), .B(n[458]), .Z(n13796) );
  NAND U15303 ( .A(n13797), .B(n[459]), .Z(n6098) );
  NAND U15304 ( .A(n8085), .B(n[459]), .Z(n13797) );
  NAND U15305 ( .A(n13798), .B(n[460]), .Z(n6088) );
  NAND U15306 ( .A(n8085), .B(n[460]), .Z(n13798) );
  NAND U15307 ( .A(n13799), .B(n[461]), .Z(n6083) );
  NAND U15308 ( .A(n8085), .B(n[461]), .Z(n13799) );
  NAND U15309 ( .A(n13800), .B(n[462]), .Z(n6078) );
  NAND U15310 ( .A(n8085), .B(n[462]), .Z(n13800) );
  NAND U15311 ( .A(n13801), .B(n[463]), .Z(n6073) );
  NAND U15312 ( .A(n8085), .B(n[463]), .Z(n13801) );
  NAND U15313 ( .A(n13802), .B(n[464]), .Z(n6068) );
  NAND U15314 ( .A(n8085), .B(n[464]), .Z(n13802) );
  NAND U15315 ( .A(n13803), .B(n[465]), .Z(n6063) );
  NAND U15316 ( .A(n8085), .B(n[465]), .Z(n13803) );
  NAND U15317 ( .A(n13804), .B(n[466]), .Z(n6058) );
  NAND U15318 ( .A(n8085), .B(n[466]), .Z(n13804) );
  NAND U15319 ( .A(n13805), .B(n[467]), .Z(n6053) );
  NAND U15320 ( .A(n8085), .B(n[467]), .Z(n13805) );
  NAND U15321 ( .A(n13806), .B(n[468]), .Z(n6048) );
  NAND U15322 ( .A(n8085), .B(n[468]), .Z(n13806) );
  NAND U15323 ( .A(n13807), .B(n[469]), .Z(n6043) );
  NAND U15324 ( .A(n8085), .B(n[469]), .Z(n13807) );
  NAND U15325 ( .A(n13808), .B(n[470]), .Z(n6033) );
  NAND U15326 ( .A(n8085), .B(n[470]), .Z(n13808) );
  NAND U15327 ( .A(n13809), .B(n[471]), .Z(n6028) );
  NAND U15328 ( .A(n8085), .B(n[471]), .Z(n13809) );
  NAND U15329 ( .A(n13810), .B(n[472]), .Z(n6023) );
  NAND U15330 ( .A(n8085), .B(n[472]), .Z(n13810) );
  NAND U15331 ( .A(n13811), .B(n[473]), .Z(n6018) );
  NAND U15332 ( .A(n8085), .B(n[473]), .Z(n13811) );
  NAND U15333 ( .A(n13812), .B(n[474]), .Z(n6013) );
  NAND U15334 ( .A(n8085), .B(n[474]), .Z(n13812) );
  NAND U15335 ( .A(n13813), .B(n[475]), .Z(n6008) );
  NAND U15336 ( .A(n8085), .B(n[475]), .Z(n13813) );
  NAND U15337 ( .A(n13814), .B(n[476]), .Z(n6003) );
  NAND U15338 ( .A(n8085), .B(n[476]), .Z(n13814) );
  NAND U15339 ( .A(n13815), .B(n[477]), .Z(n5998) );
  NAND U15340 ( .A(n8085), .B(n[477]), .Z(n13815) );
  NAND U15341 ( .A(n13816), .B(n[478]), .Z(n5993) );
  NAND U15342 ( .A(n8085), .B(n[478]), .Z(n13816) );
  NAND U15343 ( .A(n13817), .B(n[479]), .Z(n5988) );
  NAND U15344 ( .A(n8085), .B(n[479]), .Z(n13817) );
  NAND U15345 ( .A(n13818), .B(n[480]), .Z(n5978) );
  NAND U15346 ( .A(n8085), .B(n[480]), .Z(n13818) );
  NAND U15347 ( .A(n13819), .B(n[481]), .Z(n5973) );
  NAND U15348 ( .A(n8085), .B(n[481]), .Z(n13819) );
  NAND U15349 ( .A(n13820), .B(n[482]), .Z(n5968) );
  NAND U15350 ( .A(n8085), .B(n[482]), .Z(n13820) );
  NAND U15351 ( .A(n13821), .B(n[483]), .Z(n5963) );
  NAND U15352 ( .A(n8085), .B(n[483]), .Z(n13821) );
  NAND U15353 ( .A(n13822), .B(n[484]), .Z(n5958) );
  NAND U15354 ( .A(n8085), .B(n[484]), .Z(n13822) );
  NAND U15355 ( .A(n13823), .B(n[485]), .Z(n5953) );
  NAND U15356 ( .A(n8085), .B(n[485]), .Z(n13823) );
  NAND U15357 ( .A(n13824), .B(n[486]), .Z(n5948) );
  NAND U15358 ( .A(n8085), .B(n[486]), .Z(n13824) );
  NAND U15359 ( .A(n13825), .B(n[487]), .Z(n5943) );
  NAND U15360 ( .A(n8085), .B(n[487]), .Z(n13825) );
  NAND U15361 ( .A(n13826), .B(n[488]), .Z(n5938) );
  NAND U15362 ( .A(n8085), .B(n[488]), .Z(n13826) );
  NAND U15363 ( .A(n13827), .B(n[489]), .Z(n5933) );
  NAND U15364 ( .A(n8085), .B(n[489]), .Z(n13827) );
  NAND U15365 ( .A(n13828), .B(n[490]), .Z(n5923) );
  NAND U15366 ( .A(n8085), .B(n[490]), .Z(n13828) );
  NAND U15367 ( .A(n13829), .B(n[491]), .Z(n5918) );
  NAND U15368 ( .A(n8085), .B(n[491]), .Z(n13829) );
  NAND U15369 ( .A(n13830), .B(n[492]), .Z(n5913) );
  NAND U15370 ( .A(n8085), .B(n[492]), .Z(n13830) );
  NAND U15371 ( .A(n13831), .B(n[493]), .Z(n5908) );
  NAND U15372 ( .A(n8085), .B(n[493]), .Z(n13831) );
  NAND U15373 ( .A(n13832), .B(n[494]), .Z(n5903) );
  NAND U15374 ( .A(n8085), .B(n[494]), .Z(n13832) );
  NAND U15375 ( .A(n13833), .B(n[495]), .Z(n5898) );
  NAND U15376 ( .A(n8085), .B(n[495]), .Z(n13833) );
  NAND U15377 ( .A(n13834), .B(n[496]), .Z(n5893) );
  NAND U15378 ( .A(n8085), .B(n[496]), .Z(n13834) );
  NAND U15379 ( .A(n13835), .B(n[497]), .Z(n5888) );
  NAND U15380 ( .A(n8085), .B(n[497]), .Z(n13835) );
  NAND U15381 ( .A(n13836), .B(n[498]), .Z(n5883) );
  NAND U15382 ( .A(n8085), .B(n[498]), .Z(n13836) );
  NAND U15383 ( .A(n13837), .B(n[499]), .Z(n5878) );
  NAND U15384 ( .A(n8085), .B(n[499]), .Z(n13837) );
  NAND U15385 ( .A(n13838), .B(n[500]), .Z(n5863) );
  NAND U15386 ( .A(n8085), .B(n[500]), .Z(n13838) );
  NAND U15387 ( .A(n13839), .B(n[501]), .Z(n5858) );
  NAND U15388 ( .A(n8085), .B(n[501]), .Z(n13839) );
  NAND U15389 ( .A(n13840), .B(n[502]), .Z(n5853) );
  NAND U15390 ( .A(n8085), .B(n[502]), .Z(n13840) );
  NAND U15391 ( .A(n13841), .B(n[503]), .Z(n5848) );
  NAND U15392 ( .A(n8085), .B(n[503]), .Z(n13841) );
  NAND U15393 ( .A(n13842), .B(n[504]), .Z(n5843) );
  NAND U15394 ( .A(n8085), .B(n[504]), .Z(n13842) );
  NAND U15395 ( .A(n13843), .B(n[505]), .Z(n5838) );
  NAND U15396 ( .A(n8085), .B(n[505]), .Z(n13843) );
  NAND U15397 ( .A(n13844), .B(n[506]), .Z(n5833) );
  NAND U15398 ( .A(n8085), .B(n[506]), .Z(n13844) );
  NAND U15399 ( .A(n13845), .B(n[507]), .Z(n5828) );
  NAND U15400 ( .A(n8085), .B(n[507]), .Z(n13845) );
  NAND U15401 ( .A(n13846), .B(n[508]), .Z(n5823) );
  NAND U15402 ( .A(n8085), .B(n[508]), .Z(n13846) );
  NAND U15403 ( .A(n13847), .B(n[509]), .Z(n5818) );
  NAND U15404 ( .A(n8085), .B(n[509]), .Z(n13847) );
  NAND U15405 ( .A(n13848), .B(n[510]), .Z(n5808) );
  NAND U15406 ( .A(n8085), .B(n[510]), .Z(n13848) );
  NAND U15407 ( .A(n13849), .B(n[511]), .Z(n5803) );
  NAND U15408 ( .A(n8085), .B(n[511]), .Z(n13849) );
  NAND U15409 ( .A(n13850), .B(n[512]), .Z(n5798) );
  NAND U15410 ( .A(n8085), .B(n[512]), .Z(n13850) );
  NAND U15411 ( .A(n13851), .B(n[513]), .Z(n5793) );
  NAND U15412 ( .A(n8085), .B(n[513]), .Z(n13851) );
  NAND U15413 ( .A(n13852), .B(n[514]), .Z(n5788) );
  NAND U15414 ( .A(n8085), .B(n[514]), .Z(n13852) );
  NAND U15415 ( .A(n13853), .B(n[515]), .Z(n5783) );
  NAND U15416 ( .A(n8085), .B(n[515]), .Z(n13853) );
  NAND U15417 ( .A(n13854), .B(n[516]), .Z(n5778) );
  NAND U15418 ( .A(n8085), .B(n[516]), .Z(n13854) );
  NAND U15419 ( .A(n13855), .B(n[517]), .Z(n5773) );
  NAND U15420 ( .A(n8085), .B(n[517]), .Z(n13855) );
  NAND U15421 ( .A(n13856), .B(n[518]), .Z(n5768) );
  NAND U15422 ( .A(n8085), .B(n[518]), .Z(n13856) );
  NAND U15423 ( .A(n13857), .B(n[519]), .Z(n5763) );
  NAND U15424 ( .A(n8085), .B(n[519]), .Z(n13857) );
  NAND U15425 ( .A(n13858), .B(n[520]), .Z(n5753) );
  NAND U15426 ( .A(n8085), .B(n[520]), .Z(n13858) );
  NAND U15427 ( .A(n13859), .B(n[521]), .Z(n5748) );
  NAND U15428 ( .A(n8085), .B(n[521]), .Z(n13859) );
  NAND U15429 ( .A(n13860), .B(n[522]), .Z(n5743) );
  NAND U15430 ( .A(n8085), .B(n[522]), .Z(n13860) );
  NAND U15431 ( .A(n13861), .B(n[523]), .Z(n5738) );
  NAND U15432 ( .A(n8085), .B(n[523]), .Z(n13861) );
  NAND U15433 ( .A(n13862), .B(n[524]), .Z(n5733) );
  NAND U15434 ( .A(n8085), .B(n[524]), .Z(n13862) );
  NAND U15435 ( .A(n13863), .B(n[525]), .Z(n5728) );
  NAND U15436 ( .A(n8085), .B(n[525]), .Z(n13863) );
  NAND U15437 ( .A(n13864), .B(n[526]), .Z(n5723) );
  NAND U15438 ( .A(n8085), .B(n[526]), .Z(n13864) );
  NAND U15439 ( .A(n13865), .B(n[527]), .Z(n5718) );
  NAND U15440 ( .A(n8085), .B(n[527]), .Z(n13865) );
  NAND U15441 ( .A(n13866), .B(n[528]), .Z(n5713) );
  NAND U15442 ( .A(n8085), .B(n[528]), .Z(n13866) );
  NAND U15443 ( .A(n13867), .B(n[529]), .Z(n5708) );
  NAND U15444 ( .A(n8085), .B(n[529]), .Z(n13867) );
  NAND U15445 ( .A(n13868), .B(n[530]), .Z(n5698) );
  NAND U15446 ( .A(n8085), .B(n[530]), .Z(n13868) );
  NAND U15447 ( .A(n13869), .B(n[531]), .Z(n5693) );
  NAND U15448 ( .A(n8085), .B(n[531]), .Z(n13869) );
  NAND U15449 ( .A(n13870), .B(n[532]), .Z(n5688) );
  NAND U15450 ( .A(n8085), .B(n[532]), .Z(n13870) );
  NAND U15451 ( .A(n13871), .B(n[533]), .Z(n5683) );
  NAND U15452 ( .A(n8085), .B(n[533]), .Z(n13871) );
  NAND U15453 ( .A(n13872), .B(n[534]), .Z(n5678) );
  NAND U15454 ( .A(n8085), .B(n[534]), .Z(n13872) );
  NAND U15455 ( .A(n13873), .B(n[535]), .Z(n5673) );
  NAND U15456 ( .A(n8085), .B(n[535]), .Z(n13873) );
  NAND U15457 ( .A(n13874), .B(n[536]), .Z(n5668) );
  NAND U15458 ( .A(n8085), .B(n[536]), .Z(n13874) );
  NAND U15459 ( .A(n13875), .B(n[537]), .Z(n5663) );
  NAND U15460 ( .A(n8085), .B(n[537]), .Z(n13875) );
  NAND U15461 ( .A(n13876), .B(n[538]), .Z(n5658) );
  NAND U15462 ( .A(n8085), .B(n[538]), .Z(n13876) );
  NAND U15463 ( .A(n13877), .B(n[539]), .Z(n5653) );
  NAND U15464 ( .A(n8085), .B(n[539]), .Z(n13877) );
  NAND U15465 ( .A(n13878), .B(n[540]), .Z(n5643) );
  NAND U15466 ( .A(n8085), .B(n[540]), .Z(n13878) );
  NAND U15467 ( .A(n13879), .B(n[541]), .Z(n5638) );
  NAND U15468 ( .A(n8085), .B(n[541]), .Z(n13879) );
  NAND U15469 ( .A(n13880), .B(n[542]), .Z(n5633) );
  NAND U15470 ( .A(n8085), .B(n[542]), .Z(n13880) );
  NAND U15471 ( .A(n13881), .B(n[543]), .Z(n5628) );
  NAND U15472 ( .A(n8085), .B(n[543]), .Z(n13881) );
  NAND U15473 ( .A(n13882), .B(n[544]), .Z(n5623) );
  NAND U15474 ( .A(n8085), .B(n[544]), .Z(n13882) );
  NAND U15475 ( .A(n13883), .B(n[545]), .Z(n5618) );
  NAND U15476 ( .A(n8085), .B(n[545]), .Z(n13883) );
  NAND U15477 ( .A(n13884), .B(n[546]), .Z(n5613) );
  NAND U15478 ( .A(n8085), .B(n[546]), .Z(n13884) );
  NAND U15479 ( .A(n13885), .B(n[547]), .Z(n5608) );
  NAND U15480 ( .A(n8085), .B(n[547]), .Z(n13885) );
  NAND U15481 ( .A(n13886), .B(n[548]), .Z(n5603) );
  NAND U15482 ( .A(n8085), .B(n[548]), .Z(n13886) );
  NAND U15483 ( .A(n13887), .B(n[549]), .Z(n5598) );
  NAND U15484 ( .A(n8085), .B(n[549]), .Z(n13887) );
  NAND U15485 ( .A(n13888), .B(n[550]), .Z(n5588) );
  NAND U15486 ( .A(n8085), .B(n[550]), .Z(n13888) );
  NAND U15487 ( .A(n13889), .B(n[551]), .Z(n5583) );
  NAND U15488 ( .A(n8085), .B(n[551]), .Z(n13889) );
  NAND U15489 ( .A(n13890), .B(n[552]), .Z(n5578) );
  NAND U15490 ( .A(n8085), .B(n[552]), .Z(n13890) );
  NAND U15491 ( .A(n13891), .B(n[553]), .Z(n5573) );
  NAND U15492 ( .A(n8085), .B(n[553]), .Z(n13891) );
  NAND U15493 ( .A(n13892), .B(n[554]), .Z(n5568) );
  NAND U15494 ( .A(n8085), .B(n[554]), .Z(n13892) );
  NAND U15495 ( .A(n13893), .B(n[555]), .Z(n5563) );
  NAND U15496 ( .A(n8085), .B(n[555]), .Z(n13893) );
  NAND U15497 ( .A(n13894), .B(n[556]), .Z(n5558) );
  NAND U15498 ( .A(n8085), .B(n[556]), .Z(n13894) );
  NAND U15499 ( .A(n13895), .B(n[557]), .Z(n5553) );
  NAND U15500 ( .A(n8085), .B(n[557]), .Z(n13895) );
  NAND U15501 ( .A(n13896), .B(n[558]), .Z(n5548) );
  NAND U15502 ( .A(n8085), .B(n[558]), .Z(n13896) );
  NAND U15503 ( .A(n13897), .B(n[559]), .Z(n5543) );
  NAND U15504 ( .A(n8085), .B(n[559]), .Z(n13897) );
  NAND U15505 ( .A(n13898), .B(n[560]), .Z(n5533) );
  NAND U15506 ( .A(n8085), .B(n[560]), .Z(n13898) );
  NAND U15507 ( .A(n13899), .B(n[561]), .Z(n5528) );
  NAND U15508 ( .A(n8085), .B(n[561]), .Z(n13899) );
  NAND U15509 ( .A(n13900), .B(n[562]), .Z(n5523) );
  NAND U15510 ( .A(n8085), .B(n[562]), .Z(n13900) );
  NAND U15511 ( .A(n13901), .B(n[563]), .Z(n5518) );
  NAND U15512 ( .A(n8085), .B(n[563]), .Z(n13901) );
  NAND U15513 ( .A(n13902), .B(n[564]), .Z(n5513) );
  NAND U15514 ( .A(n8085), .B(n[564]), .Z(n13902) );
  NAND U15515 ( .A(n13903), .B(n[565]), .Z(n5508) );
  NAND U15516 ( .A(n8085), .B(n[565]), .Z(n13903) );
  NAND U15517 ( .A(n13904), .B(n[566]), .Z(n5503) );
  NAND U15518 ( .A(n8085), .B(n[566]), .Z(n13904) );
  NAND U15519 ( .A(n13905), .B(n[567]), .Z(n5498) );
  NAND U15520 ( .A(n8085), .B(n[567]), .Z(n13905) );
  NAND U15521 ( .A(n13906), .B(n[568]), .Z(n5493) );
  NAND U15522 ( .A(n8085), .B(n[568]), .Z(n13906) );
  NAND U15523 ( .A(n13907), .B(n[569]), .Z(n5488) );
  NAND U15524 ( .A(n8085), .B(n[569]), .Z(n13907) );
  NAND U15525 ( .A(n13908), .B(n[570]), .Z(n5478) );
  NAND U15526 ( .A(n8085), .B(n[570]), .Z(n13908) );
  NAND U15527 ( .A(n13909), .B(n[571]), .Z(n5473) );
  NAND U15528 ( .A(n8085), .B(n[571]), .Z(n13909) );
  NAND U15529 ( .A(n13910), .B(n[572]), .Z(n5468) );
  NAND U15530 ( .A(n8085), .B(n[572]), .Z(n13910) );
  NAND U15531 ( .A(n13911), .B(n[573]), .Z(n5463) );
  NAND U15532 ( .A(n8085), .B(n[573]), .Z(n13911) );
  NAND U15533 ( .A(n13912), .B(n[574]), .Z(n5458) );
  NAND U15534 ( .A(n8085), .B(n[574]), .Z(n13912) );
  NAND U15535 ( .A(n13913), .B(n[575]), .Z(n5453) );
  NAND U15536 ( .A(n8085), .B(n[575]), .Z(n13913) );
  NAND U15537 ( .A(n13914), .B(n[576]), .Z(n5448) );
  NAND U15538 ( .A(n8085), .B(n[576]), .Z(n13914) );
  NAND U15539 ( .A(n13915), .B(n[577]), .Z(n5443) );
  NAND U15540 ( .A(n8085), .B(n[577]), .Z(n13915) );
  NAND U15541 ( .A(n13916), .B(n[578]), .Z(n5438) );
  NAND U15542 ( .A(n8085), .B(n[578]), .Z(n13916) );
  NAND U15543 ( .A(n13917), .B(n[579]), .Z(n5433) );
  NAND U15544 ( .A(n8085), .B(n[579]), .Z(n13917) );
  NAND U15545 ( .A(n13918), .B(n[580]), .Z(n5423) );
  NAND U15546 ( .A(n8085), .B(n[580]), .Z(n13918) );
  NAND U15547 ( .A(n13919), .B(n[581]), .Z(n5418) );
  NAND U15548 ( .A(n8085), .B(n[581]), .Z(n13919) );
  NAND U15549 ( .A(n13920), .B(n[582]), .Z(n5413) );
  NAND U15550 ( .A(n8085), .B(n[582]), .Z(n13920) );
  NAND U15551 ( .A(n13921), .B(n[583]), .Z(n5408) );
  NAND U15552 ( .A(n8085), .B(n[583]), .Z(n13921) );
  NAND U15553 ( .A(n13922), .B(n[584]), .Z(n5403) );
  NAND U15554 ( .A(n8085), .B(n[584]), .Z(n13922) );
  NAND U15555 ( .A(n13923), .B(n[585]), .Z(n5398) );
  NAND U15556 ( .A(n8085), .B(n[585]), .Z(n13923) );
  NAND U15557 ( .A(n13924), .B(n[586]), .Z(n5393) );
  NAND U15558 ( .A(n8085), .B(n[586]), .Z(n13924) );
  NAND U15559 ( .A(n13925), .B(n[587]), .Z(n5388) );
  NAND U15560 ( .A(n8085), .B(n[587]), .Z(n13925) );
  NAND U15561 ( .A(n13926), .B(n[588]), .Z(n5383) );
  NAND U15562 ( .A(n8085), .B(n[588]), .Z(n13926) );
  NAND U15563 ( .A(n13927), .B(n[589]), .Z(n5378) );
  NAND U15564 ( .A(n8085), .B(n[589]), .Z(n13927) );
  NAND U15565 ( .A(n13928), .B(n[590]), .Z(n5368) );
  NAND U15566 ( .A(n8085), .B(n[590]), .Z(n13928) );
  NAND U15567 ( .A(n13929), .B(n[591]), .Z(n5363) );
  NAND U15568 ( .A(n8085), .B(n[591]), .Z(n13929) );
  NAND U15569 ( .A(n13930), .B(n[592]), .Z(n5358) );
  NAND U15570 ( .A(n8085), .B(n[592]), .Z(n13930) );
  NAND U15571 ( .A(n13931), .B(n[593]), .Z(n5353) );
  NAND U15572 ( .A(n8085), .B(n[593]), .Z(n13931) );
  NAND U15573 ( .A(n13932), .B(n[594]), .Z(n5348) );
  NAND U15574 ( .A(n8085), .B(n[594]), .Z(n13932) );
  NAND U15575 ( .A(n13933), .B(n[595]), .Z(n5343) );
  NAND U15576 ( .A(n8085), .B(n[595]), .Z(n13933) );
  NAND U15577 ( .A(n13934), .B(n[596]), .Z(n5338) );
  NAND U15578 ( .A(n8085), .B(n[596]), .Z(n13934) );
  NAND U15579 ( .A(n13935), .B(n[597]), .Z(n5333) );
  NAND U15580 ( .A(n8085), .B(n[597]), .Z(n13935) );
  NAND U15581 ( .A(n13936), .B(n[598]), .Z(n5328) );
  NAND U15582 ( .A(n8085), .B(n[598]), .Z(n13936) );
  NAND U15583 ( .A(n13937), .B(n[599]), .Z(n5323) );
  NAND U15584 ( .A(n8085), .B(n[599]), .Z(n13937) );
  NAND U15585 ( .A(n13938), .B(n[600]), .Z(n5308) );
  NAND U15586 ( .A(n8085), .B(n[600]), .Z(n13938) );
  NAND U15587 ( .A(n13939), .B(n[601]), .Z(n5303) );
  NAND U15588 ( .A(n8085), .B(n[601]), .Z(n13939) );
  NAND U15589 ( .A(n13940), .B(n[602]), .Z(n5298) );
  NAND U15590 ( .A(n8085), .B(n[602]), .Z(n13940) );
  NAND U15591 ( .A(n13941), .B(n[603]), .Z(n5293) );
  NAND U15592 ( .A(n8085), .B(n[603]), .Z(n13941) );
  NAND U15593 ( .A(n13942), .B(n[604]), .Z(n5288) );
  NAND U15594 ( .A(n8085), .B(n[604]), .Z(n13942) );
  NAND U15595 ( .A(n13943), .B(n[605]), .Z(n5283) );
  NAND U15596 ( .A(n8085), .B(n[605]), .Z(n13943) );
  NAND U15597 ( .A(n13944), .B(n[606]), .Z(n5278) );
  NAND U15598 ( .A(n8085), .B(n[606]), .Z(n13944) );
  NAND U15599 ( .A(n13945), .B(n[607]), .Z(n5273) );
  NAND U15600 ( .A(n8085), .B(n[607]), .Z(n13945) );
  NAND U15601 ( .A(n13946), .B(n[608]), .Z(n5268) );
  NAND U15602 ( .A(n8085), .B(n[608]), .Z(n13946) );
  NAND U15603 ( .A(n13947), .B(n[609]), .Z(n5263) );
  NAND U15604 ( .A(n8085), .B(n[609]), .Z(n13947) );
  NAND U15605 ( .A(n13948), .B(n[610]), .Z(n5253) );
  NAND U15606 ( .A(n8085), .B(n[610]), .Z(n13948) );
  NAND U15607 ( .A(n13949), .B(n[611]), .Z(n5248) );
  NAND U15608 ( .A(n8085), .B(n[611]), .Z(n13949) );
  NAND U15609 ( .A(n13950), .B(n[612]), .Z(n5243) );
  NAND U15610 ( .A(n8085), .B(n[612]), .Z(n13950) );
  NAND U15611 ( .A(n13951), .B(n[613]), .Z(n5238) );
  NAND U15612 ( .A(n8085), .B(n[613]), .Z(n13951) );
  NAND U15613 ( .A(n13952), .B(n[614]), .Z(n5233) );
  NAND U15614 ( .A(n8085), .B(n[614]), .Z(n13952) );
  NAND U15615 ( .A(n13953), .B(n[615]), .Z(n5228) );
  NAND U15616 ( .A(n8085), .B(n[615]), .Z(n13953) );
  NAND U15617 ( .A(n13954), .B(n[616]), .Z(n5223) );
  NAND U15618 ( .A(n8085), .B(n[616]), .Z(n13954) );
  NAND U15619 ( .A(n13955), .B(n[617]), .Z(n5218) );
  NAND U15620 ( .A(n8085), .B(n[617]), .Z(n13955) );
  NAND U15621 ( .A(n13956), .B(n[618]), .Z(n5213) );
  NAND U15622 ( .A(n8085), .B(n[618]), .Z(n13956) );
  NAND U15623 ( .A(n13957), .B(n[619]), .Z(n5208) );
  NAND U15624 ( .A(n8085), .B(n[619]), .Z(n13957) );
  NAND U15625 ( .A(n13958), .B(n[620]), .Z(n5198) );
  NAND U15626 ( .A(n8085), .B(n[620]), .Z(n13958) );
  NAND U15627 ( .A(n13959), .B(n[621]), .Z(n5193) );
  NAND U15628 ( .A(n8085), .B(n[621]), .Z(n13959) );
  NAND U15629 ( .A(n13960), .B(n[622]), .Z(n5188) );
  NAND U15630 ( .A(n8085), .B(n[622]), .Z(n13960) );
  NAND U15631 ( .A(n13961), .B(n[623]), .Z(n5183) );
  NAND U15632 ( .A(n8085), .B(n[623]), .Z(n13961) );
  NAND U15633 ( .A(n13962), .B(n[624]), .Z(n5178) );
  NAND U15634 ( .A(n8085), .B(n[624]), .Z(n13962) );
  NAND U15635 ( .A(n13963), .B(n[625]), .Z(n5173) );
  NAND U15636 ( .A(n8085), .B(n[625]), .Z(n13963) );
  NAND U15637 ( .A(n13964), .B(n[626]), .Z(n5168) );
  NAND U15638 ( .A(n8085), .B(n[626]), .Z(n13964) );
  NAND U15639 ( .A(n13965), .B(n[627]), .Z(n5163) );
  NAND U15640 ( .A(n8085), .B(n[627]), .Z(n13965) );
  NAND U15641 ( .A(n13966), .B(n[628]), .Z(n5158) );
  NAND U15642 ( .A(n8085), .B(n[628]), .Z(n13966) );
  NAND U15643 ( .A(n13967), .B(n[629]), .Z(n5153) );
  NAND U15644 ( .A(n8085), .B(n[629]), .Z(n13967) );
  NAND U15645 ( .A(n13968), .B(n[630]), .Z(n5143) );
  NAND U15646 ( .A(n8085), .B(n[630]), .Z(n13968) );
  NAND U15647 ( .A(n13969), .B(n[631]), .Z(n5138) );
  NAND U15648 ( .A(n8085), .B(n[631]), .Z(n13969) );
  NAND U15649 ( .A(n13970), .B(n[632]), .Z(n5133) );
  NAND U15650 ( .A(n8085), .B(n[632]), .Z(n13970) );
  NAND U15651 ( .A(n13971), .B(n[633]), .Z(n5128) );
  NAND U15652 ( .A(n8085), .B(n[633]), .Z(n13971) );
  NAND U15653 ( .A(n13972), .B(n[634]), .Z(n5123) );
  NAND U15654 ( .A(n8085), .B(n[634]), .Z(n13972) );
  NAND U15655 ( .A(n13973), .B(n[635]), .Z(n5118) );
  NAND U15656 ( .A(n8085), .B(n[635]), .Z(n13973) );
  NAND U15657 ( .A(n13974), .B(n[636]), .Z(n5113) );
  NAND U15658 ( .A(n8085), .B(n[636]), .Z(n13974) );
  NAND U15659 ( .A(n13975), .B(n[637]), .Z(n5108) );
  NAND U15660 ( .A(n8085), .B(n[637]), .Z(n13975) );
  NAND U15661 ( .A(n13976), .B(n[638]), .Z(n5103) );
  NAND U15662 ( .A(n8085), .B(n[638]), .Z(n13976) );
  NAND U15663 ( .A(n13977), .B(n[639]), .Z(n5098) );
  NAND U15664 ( .A(n8085), .B(n[639]), .Z(n13977) );
  NAND U15665 ( .A(n13978), .B(n[640]), .Z(n5088) );
  NAND U15666 ( .A(n8085), .B(n[640]), .Z(n13978) );
  NAND U15667 ( .A(n13979), .B(n[641]), .Z(n5083) );
  NAND U15668 ( .A(n8085), .B(n[641]), .Z(n13979) );
  NAND U15669 ( .A(n13980), .B(n[642]), .Z(n5078) );
  NAND U15670 ( .A(n8085), .B(n[642]), .Z(n13980) );
  NAND U15671 ( .A(n13981), .B(n[643]), .Z(n5073) );
  NAND U15672 ( .A(n8085), .B(n[643]), .Z(n13981) );
  NAND U15673 ( .A(n13982), .B(n[644]), .Z(n5068) );
  NAND U15674 ( .A(n8085), .B(n[644]), .Z(n13982) );
  NAND U15675 ( .A(n13983), .B(n[645]), .Z(n5063) );
  NAND U15676 ( .A(n8085), .B(n[645]), .Z(n13983) );
  NAND U15677 ( .A(n13984), .B(n[646]), .Z(n5058) );
  NAND U15678 ( .A(n8085), .B(n[646]), .Z(n13984) );
  NAND U15679 ( .A(n13985), .B(n[647]), .Z(n5053) );
  NAND U15680 ( .A(n8085), .B(n[647]), .Z(n13985) );
  NAND U15681 ( .A(n13986), .B(n[648]), .Z(n5048) );
  NAND U15682 ( .A(n8085), .B(n[648]), .Z(n13986) );
  NAND U15683 ( .A(n13987), .B(n[649]), .Z(n5043) );
  NAND U15684 ( .A(n8085), .B(n[649]), .Z(n13987) );
  NAND U15685 ( .A(n13988), .B(n[650]), .Z(n5033) );
  NAND U15686 ( .A(n8085), .B(n[650]), .Z(n13988) );
  NAND U15687 ( .A(n13989), .B(n[651]), .Z(n5028) );
  NAND U15688 ( .A(n8085), .B(n[651]), .Z(n13989) );
  NAND U15689 ( .A(n13990), .B(n[652]), .Z(n5023) );
  NAND U15690 ( .A(n8085), .B(n[652]), .Z(n13990) );
  NAND U15691 ( .A(n13991), .B(n[653]), .Z(n5018) );
  NAND U15692 ( .A(n8085), .B(n[653]), .Z(n13991) );
  NAND U15693 ( .A(n13992), .B(n[654]), .Z(n5013) );
  NAND U15694 ( .A(n8085), .B(n[654]), .Z(n13992) );
  NAND U15695 ( .A(n13993), .B(n[655]), .Z(n5008) );
  NAND U15696 ( .A(n8085), .B(n[655]), .Z(n13993) );
  NAND U15697 ( .A(n13994), .B(n[656]), .Z(n5003) );
  NAND U15698 ( .A(n8085), .B(n[656]), .Z(n13994) );
  NAND U15699 ( .A(n13995), .B(n[657]), .Z(n4998) );
  NAND U15700 ( .A(n8085), .B(n[657]), .Z(n13995) );
  NAND U15701 ( .A(n13996), .B(n[658]), .Z(n4993) );
  NAND U15702 ( .A(n8085), .B(n[658]), .Z(n13996) );
  NAND U15703 ( .A(n13997), .B(n[659]), .Z(n4988) );
  NAND U15704 ( .A(n8085), .B(n[659]), .Z(n13997) );
  NAND U15705 ( .A(n13998), .B(n[660]), .Z(n4978) );
  NAND U15706 ( .A(n8085), .B(n[660]), .Z(n13998) );
  NAND U15707 ( .A(n13999), .B(n[661]), .Z(n4973) );
  NAND U15708 ( .A(n8085), .B(n[661]), .Z(n13999) );
  NAND U15709 ( .A(n14000), .B(n[662]), .Z(n4968) );
  NAND U15710 ( .A(n8085), .B(n[662]), .Z(n14000) );
  NAND U15711 ( .A(n14001), .B(n[663]), .Z(n4963) );
  NAND U15712 ( .A(n8085), .B(n[663]), .Z(n14001) );
  NAND U15713 ( .A(n14002), .B(n[664]), .Z(n4958) );
  NAND U15714 ( .A(n8085), .B(n[664]), .Z(n14002) );
  NAND U15715 ( .A(n14003), .B(n[665]), .Z(n4953) );
  NAND U15716 ( .A(n8085), .B(n[665]), .Z(n14003) );
  NAND U15717 ( .A(n14004), .B(n[666]), .Z(n4948) );
  NAND U15718 ( .A(n8085), .B(n[666]), .Z(n14004) );
  NAND U15719 ( .A(n14005), .B(n[667]), .Z(n4943) );
  NAND U15720 ( .A(n8085), .B(n[667]), .Z(n14005) );
  NAND U15721 ( .A(n14006), .B(n[668]), .Z(n4938) );
  NAND U15722 ( .A(n8085), .B(n[668]), .Z(n14006) );
  NAND U15723 ( .A(n14007), .B(n[669]), .Z(n4933) );
  NAND U15724 ( .A(n8085), .B(n[669]), .Z(n14007) );
  NAND U15725 ( .A(n14008), .B(n[670]), .Z(n4923) );
  NAND U15726 ( .A(n8085), .B(n[670]), .Z(n14008) );
  NAND U15727 ( .A(n14009), .B(n[671]), .Z(n4918) );
  NAND U15728 ( .A(n8085), .B(n[671]), .Z(n14009) );
  NAND U15729 ( .A(n14010), .B(n[672]), .Z(n4913) );
  NAND U15730 ( .A(n8085), .B(n[672]), .Z(n14010) );
  NAND U15731 ( .A(n14011), .B(n[673]), .Z(n4908) );
  NAND U15732 ( .A(n8085), .B(n[673]), .Z(n14011) );
  NAND U15733 ( .A(n14012), .B(n[674]), .Z(n4903) );
  NAND U15734 ( .A(n8085), .B(n[674]), .Z(n14012) );
  NAND U15735 ( .A(n14013), .B(n[675]), .Z(n4898) );
  NAND U15736 ( .A(n8085), .B(n[675]), .Z(n14013) );
  NAND U15737 ( .A(n14014), .B(n[676]), .Z(n4893) );
  NAND U15738 ( .A(n8085), .B(n[676]), .Z(n14014) );
  NAND U15739 ( .A(n14015), .B(n[677]), .Z(n4888) );
  NAND U15740 ( .A(n8085), .B(n[677]), .Z(n14015) );
  NAND U15741 ( .A(n14016), .B(n[678]), .Z(n4883) );
  NAND U15742 ( .A(n8085), .B(n[678]), .Z(n14016) );
  NAND U15743 ( .A(n14017), .B(n[679]), .Z(n4878) );
  NAND U15744 ( .A(n8085), .B(n[679]), .Z(n14017) );
  NAND U15745 ( .A(n14018), .B(n[680]), .Z(n4868) );
  NAND U15746 ( .A(n8085), .B(n[680]), .Z(n14018) );
  NAND U15747 ( .A(n14019), .B(n[681]), .Z(n4863) );
  NAND U15748 ( .A(n8085), .B(n[681]), .Z(n14019) );
  NAND U15749 ( .A(n14020), .B(n[682]), .Z(n4858) );
  NAND U15750 ( .A(n8085), .B(n[682]), .Z(n14020) );
  NAND U15751 ( .A(n14021), .B(n[683]), .Z(n4853) );
  NAND U15752 ( .A(n8085), .B(n[683]), .Z(n14021) );
  NAND U15753 ( .A(n14022), .B(n[684]), .Z(n4848) );
  NAND U15754 ( .A(n8085), .B(n[684]), .Z(n14022) );
  NAND U15755 ( .A(n14023), .B(n[685]), .Z(n4843) );
  NAND U15756 ( .A(n8085), .B(n[685]), .Z(n14023) );
  NAND U15757 ( .A(n14024), .B(n[686]), .Z(n4838) );
  NAND U15758 ( .A(n8085), .B(n[686]), .Z(n14024) );
  NAND U15759 ( .A(n14025), .B(n[687]), .Z(n4833) );
  NAND U15760 ( .A(n8085), .B(n[687]), .Z(n14025) );
  NAND U15761 ( .A(n14026), .B(n[688]), .Z(n4828) );
  NAND U15762 ( .A(n8085), .B(n[688]), .Z(n14026) );
  NAND U15763 ( .A(n14027), .B(n[689]), .Z(n4823) );
  NAND U15764 ( .A(n8085), .B(n[689]), .Z(n14027) );
  NAND U15765 ( .A(n14028), .B(n[690]), .Z(n4813) );
  NAND U15766 ( .A(n8085), .B(n[690]), .Z(n14028) );
  NAND U15767 ( .A(n14029), .B(n[691]), .Z(n4808) );
  NAND U15768 ( .A(n8085), .B(n[691]), .Z(n14029) );
  NAND U15769 ( .A(n14030), .B(n[692]), .Z(n4803) );
  NAND U15770 ( .A(n8085), .B(n[692]), .Z(n14030) );
  NAND U15771 ( .A(n14031), .B(n[693]), .Z(n4798) );
  NAND U15772 ( .A(n8085), .B(n[693]), .Z(n14031) );
  NAND U15773 ( .A(n14032), .B(n[694]), .Z(n4793) );
  NAND U15774 ( .A(n8085), .B(n[694]), .Z(n14032) );
  NAND U15775 ( .A(n14033), .B(n[695]), .Z(n4788) );
  NAND U15776 ( .A(n8085), .B(n[695]), .Z(n14033) );
  NAND U15777 ( .A(n14034), .B(n[696]), .Z(n4783) );
  NAND U15778 ( .A(n8085), .B(n[696]), .Z(n14034) );
  NAND U15779 ( .A(n14035), .B(n[697]), .Z(n4778) );
  NAND U15780 ( .A(n8085), .B(n[697]), .Z(n14035) );
  NAND U15781 ( .A(n14036), .B(n[698]), .Z(n4773) );
  NAND U15782 ( .A(n8085), .B(n[698]), .Z(n14036) );
  NAND U15783 ( .A(n14037), .B(n[699]), .Z(n4768) );
  NAND U15784 ( .A(n8085), .B(n[699]), .Z(n14037) );
  NAND U15785 ( .A(n14038), .B(n[700]), .Z(n4753) );
  NAND U15786 ( .A(n8085), .B(n[700]), .Z(n14038) );
  NAND U15787 ( .A(n14039), .B(n[701]), .Z(n4748) );
  NAND U15788 ( .A(n8085), .B(n[701]), .Z(n14039) );
  NAND U15789 ( .A(n14040), .B(n[702]), .Z(n4743) );
  NAND U15790 ( .A(n8085), .B(n[702]), .Z(n14040) );
  NAND U15791 ( .A(n14041), .B(n[703]), .Z(n4738) );
  NAND U15792 ( .A(n8085), .B(n[703]), .Z(n14041) );
  NAND U15793 ( .A(n14042), .B(n[704]), .Z(n4733) );
  NAND U15794 ( .A(n8085), .B(n[704]), .Z(n14042) );
  NAND U15795 ( .A(n14043), .B(n[705]), .Z(n4728) );
  NAND U15796 ( .A(n8085), .B(n[705]), .Z(n14043) );
  NAND U15797 ( .A(n14044), .B(n[706]), .Z(n4723) );
  NAND U15798 ( .A(n8085), .B(n[706]), .Z(n14044) );
  NAND U15799 ( .A(n14045), .B(n[707]), .Z(n4718) );
  NAND U15800 ( .A(n8085), .B(n[707]), .Z(n14045) );
  NAND U15801 ( .A(n14046), .B(n[708]), .Z(n4713) );
  NAND U15802 ( .A(n8085), .B(n[708]), .Z(n14046) );
  NAND U15803 ( .A(n14047), .B(n[709]), .Z(n4708) );
  NAND U15804 ( .A(n8085), .B(n[709]), .Z(n14047) );
  NAND U15805 ( .A(n14048), .B(n[710]), .Z(n4698) );
  NAND U15806 ( .A(n8085), .B(n[710]), .Z(n14048) );
  NAND U15807 ( .A(n14049), .B(n[711]), .Z(n4693) );
  NAND U15808 ( .A(n8085), .B(n[711]), .Z(n14049) );
  NAND U15809 ( .A(n14050), .B(n[712]), .Z(n4688) );
  NAND U15810 ( .A(n8085), .B(n[712]), .Z(n14050) );
  NAND U15811 ( .A(n14051), .B(n[713]), .Z(n4683) );
  NAND U15812 ( .A(n8085), .B(n[713]), .Z(n14051) );
  NAND U15813 ( .A(n14052), .B(n[714]), .Z(n4678) );
  NAND U15814 ( .A(n8085), .B(n[714]), .Z(n14052) );
  NAND U15815 ( .A(n14053), .B(n[715]), .Z(n4673) );
  NAND U15816 ( .A(n8085), .B(n[715]), .Z(n14053) );
  NAND U15817 ( .A(n14054), .B(n[716]), .Z(n4668) );
  NAND U15818 ( .A(n8085), .B(n[716]), .Z(n14054) );
  NAND U15819 ( .A(n14055), .B(n[717]), .Z(n4663) );
  NAND U15820 ( .A(n8085), .B(n[717]), .Z(n14055) );
  NAND U15821 ( .A(n14056), .B(n[718]), .Z(n4658) );
  NAND U15822 ( .A(n8085), .B(n[718]), .Z(n14056) );
  NAND U15823 ( .A(n14057), .B(n[719]), .Z(n4653) );
  NAND U15824 ( .A(n8085), .B(n[719]), .Z(n14057) );
  NAND U15825 ( .A(n14058), .B(n[720]), .Z(n4643) );
  NAND U15826 ( .A(n8085), .B(n[720]), .Z(n14058) );
  NAND U15827 ( .A(n14059), .B(n[721]), .Z(n4638) );
  NAND U15828 ( .A(n8085), .B(n[721]), .Z(n14059) );
  NAND U15829 ( .A(n14060), .B(n[722]), .Z(n4633) );
  NAND U15830 ( .A(n8085), .B(n[722]), .Z(n14060) );
  NAND U15831 ( .A(n14061), .B(n[723]), .Z(n4628) );
  NAND U15832 ( .A(n8085), .B(n[723]), .Z(n14061) );
  NAND U15833 ( .A(n14062), .B(n[724]), .Z(n4623) );
  NAND U15834 ( .A(n8085), .B(n[724]), .Z(n14062) );
  NAND U15835 ( .A(n14063), .B(n[725]), .Z(n4618) );
  NAND U15836 ( .A(n8085), .B(n[725]), .Z(n14063) );
  NAND U15837 ( .A(n14064), .B(n[726]), .Z(n4613) );
  NAND U15838 ( .A(n8085), .B(n[726]), .Z(n14064) );
  NAND U15839 ( .A(n14065), .B(n[727]), .Z(n4608) );
  NAND U15840 ( .A(n8085), .B(n[727]), .Z(n14065) );
  NAND U15841 ( .A(n14066), .B(n[728]), .Z(n4603) );
  NAND U15842 ( .A(n8085), .B(n[728]), .Z(n14066) );
  NAND U15843 ( .A(n14067), .B(n[729]), .Z(n4598) );
  NAND U15844 ( .A(n8085), .B(n[729]), .Z(n14067) );
  NAND U15845 ( .A(n14068), .B(n[730]), .Z(n4588) );
  NAND U15846 ( .A(n8085), .B(n[730]), .Z(n14068) );
  NAND U15847 ( .A(n14069), .B(n[731]), .Z(n4583) );
  NAND U15848 ( .A(n8085), .B(n[731]), .Z(n14069) );
  NAND U15849 ( .A(n14070), .B(n[732]), .Z(n4578) );
  NAND U15850 ( .A(n8085), .B(n[732]), .Z(n14070) );
  NAND U15851 ( .A(n14071), .B(n[733]), .Z(n4573) );
  NAND U15852 ( .A(n8085), .B(n[733]), .Z(n14071) );
  NAND U15853 ( .A(n14072), .B(n[734]), .Z(n4568) );
  NAND U15854 ( .A(n8085), .B(n[734]), .Z(n14072) );
  NAND U15855 ( .A(n14073), .B(n[735]), .Z(n4563) );
  NAND U15856 ( .A(n8085), .B(n[735]), .Z(n14073) );
  NAND U15857 ( .A(n14074), .B(n[736]), .Z(n4558) );
  NAND U15858 ( .A(n8085), .B(n[736]), .Z(n14074) );
  NAND U15859 ( .A(n14075), .B(n[737]), .Z(n4553) );
  NAND U15860 ( .A(n8085), .B(n[737]), .Z(n14075) );
  NAND U15861 ( .A(n14076), .B(n[738]), .Z(n4548) );
  NAND U15862 ( .A(n8085), .B(n[738]), .Z(n14076) );
  NAND U15863 ( .A(n14077), .B(n[739]), .Z(n4543) );
  NAND U15864 ( .A(n8085), .B(n[739]), .Z(n14077) );
  NAND U15865 ( .A(n14078), .B(n[740]), .Z(n4533) );
  NAND U15866 ( .A(n8085), .B(n[740]), .Z(n14078) );
  NAND U15867 ( .A(n14079), .B(n[741]), .Z(n4528) );
  NAND U15868 ( .A(n8085), .B(n[741]), .Z(n14079) );
  NAND U15869 ( .A(n14080), .B(n[742]), .Z(n4523) );
  NAND U15870 ( .A(n8085), .B(n[742]), .Z(n14080) );
  NAND U15871 ( .A(n14081), .B(n[743]), .Z(n4518) );
  NAND U15872 ( .A(n8085), .B(n[743]), .Z(n14081) );
  NAND U15873 ( .A(n14082), .B(n[744]), .Z(n4513) );
  NAND U15874 ( .A(n8085), .B(n[744]), .Z(n14082) );
  NAND U15875 ( .A(n14083), .B(n[745]), .Z(n4508) );
  NAND U15876 ( .A(n8085), .B(n[745]), .Z(n14083) );
  NAND U15877 ( .A(n14084), .B(n[746]), .Z(n4503) );
  NAND U15878 ( .A(n8085), .B(n[746]), .Z(n14084) );
  NAND U15879 ( .A(n14085), .B(n[747]), .Z(n4498) );
  NAND U15880 ( .A(n8085), .B(n[747]), .Z(n14085) );
  NAND U15881 ( .A(n14086), .B(n[748]), .Z(n4493) );
  NAND U15882 ( .A(n8085), .B(n[748]), .Z(n14086) );
  NAND U15883 ( .A(n14087), .B(n[749]), .Z(n4488) );
  NAND U15884 ( .A(n8085), .B(n[749]), .Z(n14087) );
  NAND U15885 ( .A(n14088), .B(n[750]), .Z(n4478) );
  NAND U15886 ( .A(n8085), .B(n[750]), .Z(n14088) );
  NAND U15887 ( .A(n14089), .B(n[751]), .Z(n4473) );
  NAND U15888 ( .A(n8085), .B(n[751]), .Z(n14089) );
  NAND U15889 ( .A(n14090), .B(n[752]), .Z(n4468) );
  NAND U15890 ( .A(n8085), .B(n[752]), .Z(n14090) );
  NAND U15891 ( .A(n14091), .B(n[753]), .Z(n4463) );
  NAND U15892 ( .A(n8085), .B(n[753]), .Z(n14091) );
  NAND U15893 ( .A(n14092), .B(n[754]), .Z(n4458) );
  NAND U15894 ( .A(n8085), .B(n[754]), .Z(n14092) );
  NAND U15895 ( .A(n14093), .B(n[755]), .Z(n4453) );
  NAND U15896 ( .A(n8085), .B(n[755]), .Z(n14093) );
  NAND U15897 ( .A(n14094), .B(n[756]), .Z(n4448) );
  NAND U15898 ( .A(n8085), .B(n[756]), .Z(n14094) );
  NAND U15899 ( .A(n14095), .B(n[757]), .Z(n4443) );
  NAND U15900 ( .A(n8085), .B(n[757]), .Z(n14095) );
  NAND U15901 ( .A(n14096), .B(n[758]), .Z(n4438) );
  NAND U15902 ( .A(n8085), .B(n[758]), .Z(n14096) );
  NAND U15903 ( .A(n14097), .B(n[759]), .Z(n4433) );
  NAND U15904 ( .A(n8085), .B(n[759]), .Z(n14097) );
  NAND U15905 ( .A(n14098), .B(n[760]), .Z(n4423) );
  NAND U15906 ( .A(n8085), .B(n[760]), .Z(n14098) );
  NAND U15907 ( .A(n14099), .B(n[761]), .Z(n4418) );
  NAND U15908 ( .A(n8085), .B(n[761]), .Z(n14099) );
  NAND U15909 ( .A(n14100), .B(n[762]), .Z(n4413) );
  NAND U15910 ( .A(n8085), .B(n[762]), .Z(n14100) );
  NAND U15911 ( .A(n14101), .B(n[763]), .Z(n4408) );
  NAND U15912 ( .A(n8085), .B(n[763]), .Z(n14101) );
  NAND U15913 ( .A(n14102), .B(n[764]), .Z(n4403) );
  NAND U15914 ( .A(n8085), .B(n[764]), .Z(n14102) );
  NAND U15915 ( .A(n14103), .B(n[765]), .Z(n4398) );
  NAND U15916 ( .A(n8085), .B(n[765]), .Z(n14103) );
  NAND U15917 ( .A(n14104), .B(n[766]), .Z(n4393) );
  NAND U15918 ( .A(n8085), .B(n[766]), .Z(n14104) );
  NAND U15919 ( .A(n14105), .B(n[767]), .Z(n4388) );
  NAND U15920 ( .A(n8085), .B(n[767]), .Z(n14105) );
  NAND U15921 ( .A(n14106), .B(n[768]), .Z(n4383) );
  NAND U15922 ( .A(n8085), .B(n[768]), .Z(n14106) );
  NAND U15923 ( .A(n14107), .B(n[769]), .Z(n4378) );
  NAND U15924 ( .A(n8085), .B(n[769]), .Z(n14107) );
  NAND U15925 ( .A(n14108), .B(n[770]), .Z(n4368) );
  NAND U15926 ( .A(n8085), .B(n[770]), .Z(n14108) );
  NAND U15927 ( .A(n14109), .B(n[771]), .Z(n4363) );
  NAND U15928 ( .A(n8085), .B(n[771]), .Z(n14109) );
  NAND U15929 ( .A(n14110), .B(n[772]), .Z(n4358) );
  NAND U15930 ( .A(n8085), .B(n[772]), .Z(n14110) );
  NAND U15931 ( .A(n14111), .B(n[773]), .Z(n4353) );
  NAND U15932 ( .A(n8085), .B(n[773]), .Z(n14111) );
  NAND U15933 ( .A(n14112), .B(n[774]), .Z(n4348) );
  NAND U15934 ( .A(n8085), .B(n[774]), .Z(n14112) );
  NAND U15935 ( .A(n14113), .B(n[775]), .Z(n4343) );
  NAND U15936 ( .A(n8085), .B(n[775]), .Z(n14113) );
  NAND U15937 ( .A(n14114), .B(n[776]), .Z(n4338) );
  NAND U15938 ( .A(n8085), .B(n[776]), .Z(n14114) );
  NAND U15939 ( .A(n14115), .B(n[777]), .Z(n4333) );
  NAND U15940 ( .A(n8085), .B(n[777]), .Z(n14115) );
  NAND U15941 ( .A(n14116), .B(n[778]), .Z(n4328) );
  NAND U15942 ( .A(n8085), .B(n[778]), .Z(n14116) );
  NAND U15943 ( .A(n14117), .B(n[779]), .Z(n4323) );
  NAND U15944 ( .A(n8085), .B(n[779]), .Z(n14117) );
  NAND U15945 ( .A(n14118), .B(n[780]), .Z(n4313) );
  NAND U15946 ( .A(n8085), .B(n[780]), .Z(n14118) );
  NAND U15947 ( .A(n14119), .B(n[781]), .Z(n4308) );
  NAND U15948 ( .A(n8085), .B(n[781]), .Z(n14119) );
  NAND U15949 ( .A(n14120), .B(n[782]), .Z(n4303) );
  NAND U15950 ( .A(n8085), .B(n[782]), .Z(n14120) );
  NAND U15951 ( .A(n14121), .B(n[783]), .Z(n4298) );
  NAND U15952 ( .A(n8085), .B(n[783]), .Z(n14121) );
  NAND U15953 ( .A(n14122), .B(n[784]), .Z(n4293) );
  NAND U15954 ( .A(n8085), .B(n[784]), .Z(n14122) );
  NAND U15955 ( .A(n14123), .B(n[785]), .Z(n4288) );
  NAND U15956 ( .A(n8085), .B(n[785]), .Z(n14123) );
  NAND U15957 ( .A(n14124), .B(n[786]), .Z(n4283) );
  NAND U15958 ( .A(n8085), .B(n[786]), .Z(n14124) );
  NAND U15959 ( .A(n14125), .B(n[787]), .Z(n4278) );
  NAND U15960 ( .A(n8085), .B(n[787]), .Z(n14125) );
  NAND U15961 ( .A(n14126), .B(n[788]), .Z(n4273) );
  NAND U15962 ( .A(n8085), .B(n[788]), .Z(n14126) );
  NAND U15963 ( .A(n14127), .B(n[789]), .Z(n4268) );
  NAND U15964 ( .A(n8085), .B(n[789]), .Z(n14127) );
  NAND U15965 ( .A(n14128), .B(n[790]), .Z(n4258) );
  NAND U15966 ( .A(n8085), .B(n[790]), .Z(n14128) );
  NAND U15967 ( .A(n14129), .B(n[791]), .Z(n4253) );
  NAND U15968 ( .A(n8085), .B(n[791]), .Z(n14129) );
  NAND U15969 ( .A(n14130), .B(n[792]), .Z(n4248) );
  NAND U15970 ( .A(n8085), .B(n[792]), .Z(n14130) );
  NAND U15971 ( .A(n14131), .B(n[793]), .Z(n4243) );
  NAND U15972 ( .A(n8085), .B(n[793]), .Z(n14131) );
  NAND U15973 ( .A(n14132), .B(n[794]), .Z(n4238) );
  NAND U15974 ( .A(n8085), .B(n[794]), .Z(n14132) );
  NAND U15975 ( .A(n14133), .B(n[795]), .Z(n4233) );
  NAND U15976 ( .A(n8085), .B(n[795]), .Z(n14133) );
  NAND U15977 ( .A(n14134), .B(n[796]), .Z(n4228) );
  NAND U15978 ( .A(n8085), .B(n[796]), .Z(n14134) );
  NAND U15979 ( .A(n14135), .B(n[797]), .Z(n4223) );
  NAND U15980 ( .A(n8085), .B(n[797]), .Z(n14135) );
  NAND U15981 ( .A(n14136), .B(n[798]), .Z(n4218) );
  NAND U15982 ( .A(n8085), .B(n[798]), .Z(n14136) );
  NAND U15983 ( .A(n14137), .B(n[799]), .Z(n4213) );
  NAND U15984 ( .A(n8085), .B(n[799]), .Z(n14137) );
  NAND U15985 ( .A(n14138), .B(n[800]), .Z(n4198) );
  NAND U15986 ( .A(n8085), .B(n[800]), .Z(n14138) );
  NAND U15987 ( .A(n14139), .B(n[801]), .Z(n4193) );
  NAND U15988 ( .A(n8085), .B(n[801]), .Z(n14139) );
  NAND U15989 ( .A(n14140), .B(n[802]), .Z(n4188) );
  NAND U15990 ( .A(n8085), .B(n[802]), .Z(n14140) );
  NAND U15991 ( .A(n14141), .B(n[803]), .Z(n4183) );
  NAND U15992 ( .A(n8085), .B(n[803]), .Z(n14141) );
  NAND U15993 ( .A(n14142), .B(n[804]), .Z(n4178) );
  NAND U15994 ( .A(n8085), .B(n[804]), .Z(n14142) );
  NAND U15995 ( .A(n14143), .B(n[805]), .Z(n4173) );
  NAND U15996 ( .A(n8085), .B(n[805]), .Z(n14143) );
  NAND U15997 ( .A(n14144), .B(n[806]), .Z(n4168) );
  NAND U15998 ( .A(n8085), .B(n[806]), .Z(n14144) );
  NAND U15999 ( .A(n14145), .B(n[807]), .Z(n4163) );
  NAND U16000 ( .A(n8085), .B(n[807]), .Z(n14145) );
  NAND U16001 ( .A(n14146), .B(n[808]), .Z(n4158) );
  NAND U16002 ( .A(n8085), .B(n[808]), .Z(n14146) );
  NAND U16003 ( .A(n14147), .B(n[809]), .Z(n4153) );
  NAND U16004 ( .A(n8085), .B(n[809]), .Z(n14147) );
  NAND U16005 ( .A(n14148), .B(n[810]), .Z(n4143) );
  NAND U16006 ( .A(n8085), .B(n[810]), .Z(n14148) );
  NAND U16007 ( .A(n14149), .B(n[811]), .Z(n4138) );
  NAND U16008 ( .A(n8085), .B(n[811]), .Z(n14149) );
  NAND U16009 ( .A(n14150), .B(n[812]), .Z(n4133) );
  NAND U16010 ( .A(n8085), .B(n[812]), .Z(n14150) );
  NAND U16011 ( .A(n14151), .B(n[813]), .Z(n4128) );
  NAND U16012 ( .A(n8085), .B(n[813]), .Z(n14151) );
  NAND U16013 ( .A(n14152), .B(n[814]), .Z(n4123) );
  NAND U16014 ( .A(n8085), .B(n[814]), .Z(n14152) );
  NAND U16015 ( .A(n14153), .B(n[815]), .Z(n4118) );
  NAND U16016 ( .A(n8085), .B(n[815]), .Z(n14153) );
  NAND U16017 ( .A(n14154), .B(n[816]), .Z(n4113) );
  NAND U16018 ( .A(n8085), .B(n[816]), .Z(n14154) );
  NAND U16019 ( .A(n14155), .B(n[817]), .Z(n4108) );
  NAND U16020 ( .A(n8085), .B(n[817]), .Z(n14155) );
  NAND U16021 ( .A(n14156), .B(n[818]), .Z(n4103) );
  NAND U16022 ( .A(n8085), .B(n[818]), .Z(n14156) );
  NAND U16023 ( .A(n14157), .B(n[819]), .Z(n4098) );
  NAND U16024 ( .A(n8085), .B(n[819]), .Z(n14157) );
  NAND U16025 ( .A(n14158), .B(n[820]), .Z(n4088) );
  NAND U16026 ( .A(n8085), .B(n[820]), .Z(n14158) );
  NAND U16027 ( .A(n14159), .B(n[821]), .Z(n4083) );
  NAND U16028 ( .A(n8085), .B(n[821]), .Z(n14159) );
  NAND U16029 ( .A(n14160), .B(n[822]), .Z(n4078) );
  NAND U16030 ( .A(n8085), .B(n[822]), .Z(n14160) );
  NAND U16031 ( .A(n14161), .B(n[823]), .Z(n4073) );
  NAND U16032 ( .A(n8085), .B(n[823]), .Z(n14161) );
  NAND U16033 ( .A(n14162), .B(n[824]), .Z(n4068) );
  NAND U16034 ( .A(n8085), .B(n[824]), .Z(n14162) );
  NAND U16035 ( .A(n14163), .B(n[825]), .Z(n4063) );
  NAND U16036 ( .A(n8085), .B(n[825]), .Z(n14163) );
  NAND U16037 ( .A(n14164), .B(n[826]), .Z(n4058) );
  NAND U16038 ( .A(n8085), .B(n[826]), .Z(n14164) );
  NAND U16039 ( .A(n14165), .B(n[827]), .Z(n4053) );
  NAND U16040 ( .A(n8085), .B(n[827]), .Z(n14165) );
  NAND U16041 ( .A(n14166), .B(n[828]), .Z(n4048) );
  NAND U16042 ( .A(n8085), .B(n[828]), .Z(n14166) );
  NAND U16043 ( .A(n14167), .B(n[829]), .Z(n4043) );
  NAND U16044 ( .A(n8085), .B(n[829]), .Z(n14167) );
  NAND U16045 ( .A(n14168), .B(n[830]), .Z(n4033) );
  NAND U16046 ( .A(n8085), .B(n[830]), .Z(n14168) );
  NAND U16047 ( .A(n14169), .B(n[831]), .Z(n4028) );
  NAND U16048 ( .A(n8085), .B(n[831]), .Z(n14169) );
  NAND U16049 ( .A(n14170), .B(n[832]), .Z(n4023) );
  NAND U16050 ( .A(n8085), .B(n[832]), .Z(n14170) );
  NAND U16051 ( .A(n14171), .B(n[833]), .Z(n4018) );
  NAND U16052 ( .A(n8085), .B(n[833]), .Z(n14171) );
  NAND U16053 ( .A(n14172), .B(n[834]), .Z(n4013) );
  NAND U16054 ( .A(n8085), .B(n[834]), .Z(n14172) );
  NAND U16055 ( .A(n14173), .B(n[835]), .Z(n4008) );
  NAND U16056 ( .A(n8085), .B(n[835]), .Z(n14173) );
  NAND U16057 ( .A(n14174), .B(n[836]), .Z(n4003) );
  NAND U16058 ( .A(n8085), .B(n[836]), .Z(n14174) );
  NAND U16059 ( .A(n14175), .B(n[837]), .Z(n3998) );
  NAND U16060 ( .A(n8085), .B(n[837]), .Z(n14175) );
  NAND U16061 ( .A(n14176), .B(n[838]), .Z(n3993) );
  NAND U16062 ( .A(n8085), .B(n[838]), .Z(n14176) );
  NAND U16063 ( .A(n14177), .B(n[839]), .Z(n3988) );
  NAND U16064 ( .A(n8085), .B(n[839]), .Z(n14177) );
  NAND U16065 ( .A(n14178), .B(n[840]), .Z(n3978) );
  NAND U16066 ( .A(n8085), .B(n[840]), .Z(n14178) );
  NAND U16067 ( .A(n14179), .B(n[841]), .Z(n3973) );
  NAND U16068 ( .A(n8085), .B(n[841]), .Z(n14179) );
  NAND U16069 ( .A(n14180), .B(n[842]), .Z(n3968) );
  NAND U16070 ( .A(n8085), .B(n[842]), .Z(n14180) );
  NAND U16071 ( .A(n14181), .B(n[843]), .Z(n3963) );
  NAND U16072 ( .A(n8085), .B(n[843]), .Z(n14181) );
  NAND U16073 ( .A(n14182), .B(n[844]), .Z(n3958) );
  NAND U16074 ( .A(n8085), .B(n[844]), .Z(n14182) );
  NAND U16075 ( .A(n14183), .B(n[845]), .Z(n3953) );
  NAND U16076 ( .A(n8085), .B(n[845]), .Z(n14183) );
  NAND U16077 ( .A(n14184), .B(n[846]), .Z(n3948) );
  NAND U16078 ( .A(n8085), .B(n[846]), .Z(n14184) );
  NAND U16079 ( .A(n14185), .B(n[847]), .Z(n3943) );
  NAND U16080 ( .A(n8085), .B(n[847]), .Z(n14185) );
  NAND U16081 ( .A(n14186), .B(n[848]), .Z(n3938) );
  NAND U16082 ( .A(n8085), .B(n[848]), .Z(n14186) );
  NAND U16083 ( .A(n14187), .B(n[849]), .Z(n3933) );
  NAND U16084 ( .A(n8085), .B(n[849]), .Z(n14187) );
  NAND U16085 ( .A(n14188), .B(n[850]), .Z(n3923) );
  NAND U16086 ( .A(n8085), .B(n[850]), .Z(n14188) );
  NAND U16087 ( .A(n14189), .B(n[851]), .Z(n3918) );
  NAND U16088 ( .A(n8085), .B(n[851]), .Z(n14189) );
  NAND U16089 ( .A(n14190), .B(n[852]), .Z(n3913) );
  NAND U16090 ( .A(n8085), .B(n[852]), .Z(n14190) );
  NAND U16091 ( .A(n14191), .B(n[853]), .Z(n3908) );
  NAND U16092 ( .A(n8085), .B(n[853]), .Z(n14191) );
  NAND U16093 ( .A(n14192), .B(n[854]), .Z(n3903) );
  NAND U16094 ( .A(n8085), .B(n[854]), .Z(n14192) );
  NAND U16095 ( .A(n14193), .B(n[855]), .Z(n3898) );
  NAND U16096 ( .A(n8085), .B(n[855]), .Z(n14193) );
  NAND U16097 ( .A(n14194), .B(n[856]), .Z(n3893) );
  NAND U16098 ( .A(n8085), .B(n[856]), .Z(n14194) );
  NAND U16099 ( .A(n14195), .B(n[857]), .Z(n3888) );
  NAND U16100 ( .A(n8085), .B(n[857]), .Z(n14195) );
  NAND U16101 ( .A(n14196), .B(n[858]), .Z(n3883) );
  NAND U16102 ( .A(n8085), .B(n[858]), .Z(n14196) );
  NAND U16103 ( .A(n14197), .B(n[859]), .Z(n3878) );
  NAND U16104 ( .A(n8085), .B(n[859]), .Z(n14197) );
  NAND U16105 ( .A(n14198), .B(n[860]), .Z(n3868) );
  NAND U16106 ( .A(n8085), .B(n[860]), .Z(n14198) );
  NAND U16107 ( .A(n14199), .B(n[861]), .Z(n3863) );
  NAND U16108 ( .A(n8085), .B(n[861]), .Z(n14199) );
  NAND U16109 ( .A(n14200), .B(n[862]), .Z(n3858) );
  NAND U16110 ( .A(n8085), .B(n[862]), .Z(n14200) );
  NAND U16111 ( .A(n14201), .B(n[863]), .Z(n3853) );
  NAND U16112 ( .A(n8085), .B(n[863]), .Z(n14201) );
  NAND U16113 ( .A(n14202), .B(n[864]), .Z(n3848) );
  NAND U16114 ( .A(n8085), .B(n[864]), .Z(n14202) );
  NAND U16115 ( .A(n14203), .B(n[865]), .Z(n3843) );
  NAND U16116 ( .A(n8085), .B(n[865]), .Z(n14203) );
  NAND U16117 ( .A(n14204), .B(n[866]), .Z(n3838) );
  NAND U16118 ( .A(n8085), .B(n[866]), .Z(n14204) );
  NAND U16119 ( .A(n14205), .B(n[867]), .Z(n3833) );
  NAND U16120 ( .A(n8085), .B(n[867]), .Z(n14205) );
  NAND U16121 ( .A(n14206), .B(n[868]), .Z(n3828) );
  NAND U16122 ( .A(n8085), .B(n[868]), .Z(n14206) );
  NAND U16123 ( .A(n14207), .B(n[869]), .Z(n3823) );
  NAND U16124 ( .A(n8085), .B(n[869]), .Z(n14207) );
  NAND U16125 ( .A(n14208), .B(n[870]), .Z(n3813) );
  NAND U16126 ( .A(n8085), .B(n[870]), .Z(n14208) );
  NAND U16127 ( .A(n14209), .B(n[871]), .Z(n3808) );
  NAND U16128 ( .A(n8085), .B(n[871]), .Z(n14209) );
  NAND U16129 ( .A(n14210), .B(n[872]), .Z(n3803) );
  NAND U16130 ( .A(n8085), .B(n[872]), .Z(n14210) );
  NAND U16131 ( .A(n14211), .B(n[873]), .Z(n3798) );
  NAND U16132 ( .A(n8085), .B(n[873]), .Z(n14211) );
  NAND U16133 ( .A(n14212), .B(n[874]), .Z(n3793) );
  NAND U16134 ( .A(n8085), .B(n[874]), .Z(n14212) );
  NAND U16135 ( .A(n14213), .B(n[875]), .Z(n3788) );
  NAND U16136 ( .A(n8085), .B(n[875]), .Z(n14213) );
  NAND U16137 ( .A(n14214), .B(n[876]), .Z(n3783) );
  NAND U16138 ( .A(n8085), .B(n[876]), .Z(n14214) );
  NAND U16139 ( .A(n14215), .B(n[877]), .Z(n3778) );
  NAND U16140 ( .A(n8085), .B(n[877]), .Z(n14215) );
  NAND U16141 ( .A(n14216), .B(n[878]), .Z(n3773) );
  NAND U16142 ( .A(n8085), .B(n[878]), .Z(n14216) );
  NAND U16143 ( .A(n14217), .B(n[879]), .Z(n3768) );
  NAND U16144 ( .A(n8085), .B(n[879]), .Z(n14217) );
  NAND U16145 ( .A(n14218), .B(n[880]), .Z(n3758) );
  NAND U16146 ( .A(n8085), .B(n[880]), .Z(n14218) );
  NAND U16147 ( .A(n14219), .B(n[881]), .Z(n3753) );
  NAND U16148 ( .A(n8085), .B(n[881]), .Z(n14219) );
  NAND U16149 ( .A(n14220), .B(n[882]), .Z(n3748) );
  NAND U16150 ( .A(n8085), .B(n[882]), .Z(n14220) );
  NAND U16151 ( .A(n14221), .B(n[883]), .Z(n3743) );
  NAND U16152 ( .A(n8085), .B(n[883]), .Z(n14221) );
  NAND U16153 ( .A(n14222), .B(n[884]), .Z(n3738) );
  NAND U16154 ( .A(n8085), .B(n[884]), .Z(n14222) );
  NAND U16155 ( .A(n14223), .B(n[885]), .Z(n3733) );
  NAND U16156 ( .A(n8085), .B(n[885]), .Z(n14223) );
  NAND U16157 ( .A(n14224), .B(n[886]), .Z(n3728) );
  NAND U16158 ( .A(n8085), .B(n[886]), .Z(n14224) );
  NAND U16159 ( .A(n14225), .B(n[887]), .Z(n3723) );
  NAND U16160 ( .A(n8085), .B(n[887]), .Z(n14225) );
  NAND U16161 ( .A(n14226), .B(n[888]), .Z(n3718) );
  NAND U16162 ( .A(n8085), .B(n[888]), .Z(n14226) );
  NAND U16163 ( .A(n14227), .B(n[889]), .Z(n3713) );
  NAND U16164 ( .A(n8085), .B(n[889]), .Z(n14227) );
  NAND U16165 ( .A(n14228), .B(n[890]), .Z(n3703) );
  NAND U16166 ( .A(n8085), .B(n[890]), .Z(n14228) );
  NAND U16167 ( .A(n14229), .B(n[891]), .Z(n3698) );
  NAND U16168 ( .A(n8085), .B(n[891]), .Z(n14229) );
  NAND U16169 ( .A(n14230), .B(n[892]), .Z(n3693) );
  NAND U16170 ( .A(n8085), .B(n[892]), .Z(n14230) );
  NAND U16171 ( .A(n14231), .B(n[893]), .Z(n3688) );
  NAND U16172 ( .A(n8085), .B(n[893]), .Z(n14231) );
  NAND U16173 ( .A(n14232), .B(n[894]), .Z(n3683) );
  NAND U16174 ( .A(n8085), .B(n[894]), .Z(n14232) );
  NAND U16175 ( .A(n14233), .B(n[895]), .Z(n3678) );
  NAND U16176 ( .A(n8085), .B(n[895]), .Z(n14233) );
  NAND U16177 ( .A(n14234), .B(n[896]), .Z(n3673) );
  NAND U16178 ( .A(n8085), .B(n[896]), .Z(n14234) );
  NAND U16179 ( .A(n14235), .B(n[897]), .Z(n3668) );
  NAND U16180 ( .A(n8085), .B(n[897]), .Z(n14235) );
  NAND U16181 ( .A(n14236), .B(n[898]), .Z(n3663) );
  NAND U16182 ( .A(n8085), .B(n[898]), .Z(n14236) );
  NAND U16183 ( .A(n14237), .B(n[899]), .Z(n3658) );
  NAND U16184 ( .A(n8085), .B(n[899]), .Z(n14237) );
  NAND U16185 ( .A(n14238), .B(n[900]), .Z(n3643) );
  NAND U16186 ( .A(n8085), .B(n[900]), .Z(n14238) );
  NAND U16187 ( .A(n14239), .B(n[901]), .Z(n3638) );
  NAND U16188 ( .A(n8085), .B(n[901]), .Z(n14239) );
  NAND U16189 ( .A(n14240), .B(n[902]), .Z(n3633) );
  NAND U16190 ( .A(n8085), .B(n[902]), .Z(n14240) );
  NAND U16191 ( .A(n14241), .B(n[903]), .Z(n3628) );
  NAND U16192 ( .A(n8085), .B(n[903]), .Z(n14241) );
  NAND U16193 ( .A(n14242), .B(n[904]), .Z(n3623) );
  NAND U16194 ( .A(n8085), .B(n[904]), .Z(n14242) );
  NAND U16195 ( .A(n14243), .B(n[905]), .Z(n3618) );
  NAND U16196 ( .A(n8085), .B(n[905]), .Z(n14243) );
  NAND U16197 ( .A(n14244), .B(n[906]), .Z(n3613) );
  NAND U16198 ( .A(n8085), .B(n[906]), .Z(n14244) );
  NAND U16199 ( .A(n14245), .B(n[907]), .Z(n3608) );
  NAND U16200 ( .A(n8085), .B(n[907]), .Z(n14245) );
  NAND U16201 ( .A(n14246), .B(n[908]), .Z(n3603) );
  NAND U16202 ( .A(n8085), .B(n[908]), .Z(n14246) );
  NAND U16203 ( .A(n14247), .B(n[909]), .Z(n3598) );
  NAND U16204 ( .A(n8085), .B(n[909]), .Z(n14247) );
  NAND U16205 ( .A(n14248), .B(n[910]), .Z(n3588) );
  NAND U16206 ( .A(n8085), .B(n[910]), .Z(n14248) );
  NAND U16207 ( .A(n14249), .B(n[911]), .Z(n3583) );
  NAND U16208 ( .A(n8085), .B(n[911]), .Z(n14249) );
  NAND U16209 ( .A(n14250), .B(n[912]), .Z(n3578) );
  NAND U16210 ( .A(n8085), .B(n[912]), .Z(n14250) );
  NAND U16211 ( .A(n14251), .B(n[913]), .Z(n3573) );
  NAND U16212 ( .A(n8085), .B(n[913]), .Z(n14251) );
  NAND U16213 ( .A(n14252), .B(n[914]), .Z(n3568) );
  NAND U16214 ( .A(n8085), .B(n[914]), .Z(n14252) );
  NAND U16215 ( .A(n14253), .B(n[915]), .Z(n3563) );
  NAND U16216 ( .A(n8085), .B(n[915]), .Z(n14253) );
  NAND U16217 ( .A(n14254), .B(n[916]), .Z(n3558) );
  NAND U16218 ( .A(n8085), .B(n[916]), .Z(n14254) );
  NAND U16219 ( .A(n14255), .B(n[917]), .Z(n3553) );
  NAND U16220 ( .A(n8085), .B(n[917]), .Z(n14255) );
  NAND U16221 ( .A(n14256), .B(n[918]), .Z(n3548) );
  NAND U16222 ( .A(n8085), .B(n[918]), .Z(n14256) );
  NAND U16223 ( .A(n14257), .B(n[919]), .Z(n3543) );
  NAND U16224 ( .A(n8085), .B(n[919]), .Z(n14257) );
  NAND U16225 ( .A(n14258), .B(n[920]), .Z(n3533) );
  NAND U16226 ( .A(n8085), .B(n[920]), .Z(n14258) );
  NAND U16227 ( .A(n14259), .B(n[921]), .Z(n3528) );
  NAND U16228 ( .A(n8085), .B(n[921]), .Z(n14259) );
  NAND U16229 ( .A(n14260), .B(n[922]), .Z(n3523) );
  NAND U16230 ( .A(n8085), .B(n[922]), .Z(n14260) );
  NAND U16231 ( .A(n14261), .B(n[923]), .Z(n3518) );
  NAND U16232 ( .A(n8085), .B(n[923]), .Z(n14261) );
  NAND U16233 ( .A(n14262), .B(n[924]), .Z(n3513) );
  NAND U16234 ( .A(n8085), .B(n[924]), .Z(n14262) );
  NAND U16235 ( .A(n14263), .B(n[925]), .Z(n3508) );
  NAND U16236 ( .A(n8085), .B(n[925]), .Z(n14263) );
  NAND U16237 ( .A(n14264), .B(n[926]), .Z(n3503) );
  NAND U16238 ( .A(n8085), .B(n[926]), .Z(n14264) );
  NAND U16239 ( .A(n14265), .B(n[927]), .Z(n3498) );
  NAND U16240 ( .A(n8085), .B(n[927]), .Z(n14265) );
  NAND U16241 ( .A(n14266), .B(n[928]), .Z(n3493) );
  NAND U16242 ( .A(n8085), .B(n[928]), .Z(n14266) );
  NAND U16243 ( .A(n14267), .B(n[929]), .Z(n3488) );
  NAND U16244 ( .A(n8085), .B(n[929]), .Z(n14267) );
  NAND U16245 ( .A(n14268), .B(n[930]), .Z(n3478) );
  NAND U16246 ( .A(n8085), .B(n[930]), .Z(n14268) );
  NAND U16247 ( .A(n14269), .B(n[931]), .Z(n3473) );
  NAND U16248 ( .A(n8085), .B(n[931]), .Z(n14269) );
  NAND U16249 ( .A(n14270), .B(n[932]), .Z(n3468) );
  NAND U16250 ( .A(n8085), .B(n[932]), .Z(n14270) );
  NAND U16251 ( .A(n14271), .B(n[933]), .Z(n3463) );
  NAND U16252 ( .A(n8085), .B(n[933]), .Z(n14271) );
  NAND U16253 ( .A(n14272), .B(n[934]), .Z(n3458) );
  NAND U16254 ( .A(n8085), .B(n[934]), .Z(n14272) );
  NAND U16255 ( .A(n14273), .B(n[935]), .Z(n3453) );
  NAND U16256 ( .A(n8085), .B(n[935]), .Z(n14273) );
  NAND U16257 ( .A(n14274), .B(n[936]), .Z(n3448) );
  NAND U16258 ( .A(n8085), .B(n[936]), .Z(n14274) );
  NAND U16259 ( .A(n14275), .B(n[937]), .Z(n3443) );
  NAND U16260 ( .A(n8085), .B(n[937]), .Z(n14275) );
  NAND U16261 ( .A(n14276), .B(n[938]), .Z(n3438) );
  NAND U16262 ( .A(n8085), .B(n[938]), .Z(n14276) );
  NAND U16263 ( .A(n14277), .B(n[939]), .Z(n3433) );
  NAND U16264 ( .A(n8085), .B(n[939]), .Z(n14277) );
  NAND U16265 ( .A(n14278), .B(n[940]), .Z(n3423) );
  NAND U16266 ( .A(n8085), .B(n[940]), .Z(n14278) );
  NAND U16267 ( .A(n14279), .B(n[941]), .Z(n3418) );
  NAND U16268 ( .A(n8085), .B(n[941]), .Z(n14279) );
  NAND U16269 ( .A(n14280), .B(n[942]), .Z(n3413) );
  NAND U16270 ( .A(n8085), .B(n[942]), .Z(n14280) );
  NAND U16271 ( .A(n14281), .B(n[943]), .Z(n3408) );
  NAND U16272 ( .A(n8085), .B(n[943]), .Z(n14281) );
  NAND U16273 ( .A(n14282), .B(n[944]), .Z(n3403) );
  NAND U16274 ( .A(n8085), .B(n[944]), .Z(n14282) );
  NAND U16275 ( .A(n14283), .B(n[945]), .Z(n3398) );
  NAND U16276 ( .A(n8085), .B(n[945]), .Z(n14283) );
  NAND U16277 ( .A(n14284), .B(n[946]), .Z(n3393) );
  NAND U16278 ( .A(n8085), .B(n[946]), .Z(n14284) );
  NAND U16279 ( .A(n14285), .B(n[947]), .Z(n3388) );
  NAND U16280 ( .A(n8085), .B(n[947]), .Z(n14285) );
  NAND U16281 ( .A(n14286), .B(n[948]), .Z(n3383) );
  NAND U16282 ( .A(n8085), .B(n[948]), .Z(n14286) );
  NAND U16283 ( .A(n14287), .B(n[949]), .Z(n3378) );
  NAND U16284 ( .A(n8085), .B(n[949]), .Z(n14287) );
  NAND U16285 ( .A(n14288), .B(n[950]), .Z(n3368) );
  NAND U16286 ( .A(n8085), .B(n[950]), .Z(n14288) );
  NAND U16287 ( .A(n14289), .B(n[951]), .Z(n3363) );
  NAND U16288 ( .A(n8085), .B(n[951]), .Z(n14289) );
  NAND U16289 ( .A(n14290), .B(n[952]), .Z(n3358) );
  NAND U16290 ( .A(n8085), .B(n[952]), .Z(n14290) );
  NAND U16291 ( .A(n14291), .B(n[953]), .Z(n3353) );
  NAND U16292 ( .A(n8085), .B(n[953]), .Z(n14291) );
  NAND U16293 ( .A(n14292), .B(n[954]), .Z(n3348) );
  NAND U16294 ( .A(n8085), .B(n[954]), .Z(n14292) );
  NAND U16295 ( .A(n14293), .B(n[955]), .Z(n3343) );
  NAND U16296 ( .A(n8085), .B(n[955]), .Z(n14293) );
  NAND U16297 ( .A(n14294), .B(n[956]), .Z(n3338) );
  NAND U16298 ( .A(n8085), .B(n[956]), .Z(n14294) );
  NAND U16299 ( .A(n14295), .B(n[957]), .Z(n3333) );
  NAND U16300 ( .A(n8085), .B(n[957]), .Z(n14295) );
  NAND U16301 ( .A(n14296), .B(n[958]), .Z(n3328) );
  NAND U16302 ( .A(n8085), .B(n[958]), .Z(n14296) );
  NAND U16303 ( .A(n14297), .B(n[959]), .Z(n3323) );
  NAND U16304 ( .A(n8085), .B(n[959]), .Z(n14297) );
  NAND U16305 ( .A(n14298), .B(n[960]), .Z(n3313) );
  NAND U16306 ( .A(n8085), .B(n[960]), .Z(n14298) );
  NAND U16307 ( .A(n14299), .B(n[961]), .Z(n3308) );
  NAND U16308 ( .A(n8085), .B(n[961]), .Z(n14299) );
  NAND U16309 ( .A(n14300), .B(n[962]), .Z(n3303) );
  NAND U16310 ( .A(n8085), .B(n[962]), .Z(n14300) );
  NAND U16311 ( .A(n14301), .B(n[963]), .Z(n3298) );
  NAND U16312 ( .A(n8085), .B(n[963]), .Z(n14301) );
  NAND U16313 ( .A(n14302), .B(n[964]), .Z(n3293) );
  NAND U16314 ( .A(n8085), .B(n[964]), .Z(n14302) );
  NAND U16315 ( .A(n14303), .B(n[965]), .Z(n3288) );
  NAND U16316 ( .A(n8085), .B(n[965]), .Z(n14303) );
  NAND U16317 ( .A(n14304), .B(n[966]), .Z(n3283) );
  NAND U16318 ( .A(n8085), .B(n[966]), .Z(n14304) );
  NAND U16319 ( .A(n14305), .B(n[967]), .Z(n3278) );
  NAND U16320 ( .A(n8085), .B(n[967]), .Z(n14305) );
  NAND U16321 ( .A(n14306), .B(n[968]), .Z(n3273) );
  NAND U16322 ( .A(n8085), .B(n[968]), .Z(n14306) );
  NAND U16323 ( .A(n14307), .B(n[969]), .Z(n3268) );
  NAND U16324 ( .A(n8085), .B(n[969]), .Z(n14307) );
  NAND U16325 ( .A(n14308), .B(n[970]), .Z(n3258) );
  NAND U16326 ( .A(n8085), .B(n[970]), .Z(n14308) );
  NAND U16327 ( .A(n14309), .B(n[971]), .Z(n3253) );
  NAND U16328 ( .A(n8085), .B(n[971]), .Z(n14309) );
  NAND U16329 ( .A(n14310), .B(n[972]), .Z(n3248) );
  NAND U16330 ( .A(n8085), .B(n[972]), .Z(n14310) );
  NAND U16331 ( .A(n14311), .B(n[973]), .Z(n3243) );
  NAND U16332 ( .A(n8085), .B(n[973]), .Z(n14311) );
  NAND U16333 ( .A(n14312), .B(n[974]), .Z(n3238) );
  NAND U16334 ( .A(n8085), .B(n[974]), .Z(n14312) );
  NAND U16335 ( .A(n14313), .B(n[975]), .Z(n3233) );
  NAND U16336 ( .A(n8085), .B(n[975]), .Z(n14313) );
  NAND U16337 ( .A(n14314), .B(n[976]), .Z(n3228) );
  NAND U16338 ( .A(n8085), .B(n[976]), .Z(n14314) );
  NAND U16339 ( .A(n14315), .B(n[977]), .Z(n3223) );
  NAND U16340 ( .A(n8085), .B(n[977]), .Z(n14315) );
  NAND U16341 ( .A(n14316), .B(n[978]), .Z(n3218) );
  NAND U16342 ( .A(n8085), .B(n[978]), .Z(n14316) );
  NAND U16343 ( .A(n14317), .B(n[979]), .Z(n3213) );
  NAND U16344 ( .A(n8085), .B(n[979]), .Z(n14317) );
  NAND U16345 ( .A(n14318), .B(n[980]), .Z(n3203) );
  NAND U16346 ( .A(n8085), .B(n[980]), .Z(n14318) );
  NAND U16347 ( .A(n14319), .B(n[981]), .Z(n3198) );
  NAND U16348 ( .A(n8085), .B(n[981]), .Z(n14319) );
  NAND U16349 ( .A(n14320), .B(n[982]), .Z(n3193) );
  NAND U16350 ( .A(n8085), .B(n[982]), .Z(n14320) );
  NAND U16351 ( .A(n14321), .B(n[983]), .Z(n3188) );
  NAND U16352 ( .A(n8085), .B(n[983]), .Z(n14321) );
  NAND U16353 ( .A(n14322), .B(n[984]), .Z(n3183) );
  NAND U16354 ( .A(n8085), .B(n[984]), .Z(n14322) );
  NAND U16355 ( .A(n14323), .B(n[985]), .Z(n3178) );
  NAND U16356 ( .A(n8085), .B(n[985]), .Z(n14323) );
  NAND U16357 ( .A(n14324), .B(n[986]), .Z(n3173) );
  NAND U16358 ( .A(n8085), .B(n[986]), .Z(n14324) );
  NAND U16359 ( .A(n14325), .B(n[987]), .Z(n3168) );
  NAND U16360 ( .A(n8085), .B(n[987]), .Z(n14325) );
  NAND U16361 ( .A(n14326), .B(n[988]), .Z(n3163) );
  NAND U16362 ( .A(n8085), .B(n[988]), .Z(n14326) );
  NAND U16363 ( .A(n14327), .B(n[989]), .Z(n3158) );
  NAND U16364 ( .A(n8085), .B(n[989]), .Z(n14327) );
  NAND U16365 ( .A(n14328), .B(n[990]), .Z(n3148) );
  NAND U16366 ( .A(n8085), .B(n[990]), .Z(n14328) );
  NAND U16367 ( .A(n14329), .B(n[991]), .Z(n3143) );
  NAND U16368 ( .A(n8085), .B(n[991]), .Z(n14329) );
  NAND U16369 ( .A(n14330), .B(n[992]), .Z(n3138) );
  NAND U16370 ( .A(n8085), .B(n[992]), .Z(n14330) );
  NAND U16371 ( .A(n14331), .B(n[993]), .Z(n3133) );
  NAND U16372 ( .A(n8085), .B(n[993]), .Z(n14331) );
  NAND U16373 ( .A(n14332), .B(n[994]), .Z(n3128) );
  NAND U16374 ( .A(n8085), .B(n[994]), .Z(n14332) );
  NAND U16375 ( .A(n14333), .B(n[995]), .Z(n3123) );
  NAND U16376 ( .A(n8085), .B(n[995]), .Z(n14333) );
  NAND U16377 ( .A(n14334), .B(n[996]), .Z(n3118) );
  NAND U16378 ( .A(n8085), .B(n[996]), .Z(n14334) );
  NAND U16379 ( .A(n14335), .B(n[997]), .Z(n3113) );
  NAND U16380 ( .A(n8085), .B(n[997]), .Z(n14335) );
  NAND U16381 ( .A(n14336), .B(n[998]), .Z(n3108) );
  NAND U16382 ( .A(n8085), .B(n[998]), .Z(n14336) );
  NAND U16383 ( .A(n14337), .B(n[999]), .Z(n3103) );
  NAND U16384 ( .A(n8085), .B(n[999]), .Z(n14337) );
  NAND U16385 ( .A(n14338), .B(n[1000]), .Z(n8336) );
  NAND U16386 ( .A(n8085), .B(n[1000]), .Z(n14338) );
  XOR U16387 ( .A(n14339), .B(o[0]), .Z(creg_next[0]) );
  AND U16388 ( .A(n3090), .B(n14340), .Z(n14339) );
  XOR U16389 ( .A(c[0]), .B(o[0]), .Z(n14340) );
  XOR U16390 ( .A(n13338), .B(n13339), .Z(o[0]) );
  NAND U16391 ( .A(n14341), .B(n[0]), .Z(n13338) );
  NAND U16392 ( .A(n8085), .B(n[0]), .Z(n14341) );
  XNOR U16393 ( .A(n14342), .B(n14343), .Z(n8085) );
  ANDN U16394 ( .B(n14344), .A(n14345), .Z(n14342) );
  XOR U16395 ( .A(n14346), .B(n14347), .Z(n14344) );
  XNOR U16396 ( .A(n14348), .B(n14345), .Z(n14347) );
  IV U16397 ( .A(n14343), .Z(n14345) );
  XOR U16398 ( .A(n14349), .B(n14350), .Z(n14343) );
  ANDN U16399 ( .B(n14351), .A(n14352), .Z(n14349) );
  IV U16400 ( .A(n14350), .Z(n14352) );
  XNOR U16401 ( .A(n14350), .B(n1038), .Z(n14351) );
  XOR U16402 ( .A(n14353), .B(n14354), .Z(n14350) );
  AND U16403 ( .A(n14355), .B(n14356), .Z(n14353) );
  XOR U16404 ( .A(n14354), .B(n8078), .Z(n14356) );
  XNOR U16405 ( .A(n14357), .B(n14358), .Z(n8078) );
  XNOR U16406 ( .A(n[1023]), .B(n14359), .Z(n14355) );
  IV U16407 ( .A(n14354), .Z(n14359) );
  XOR U16408 ( .A(n14360), .B(n14361), .Z(n14354) );
  AND U16409 ( .A(n14362), .B(n14363), .Z(n14360) );
  XOR U16410 ( .A(n14361), .B(n8089), .Z(n14363) );
  XNOR U16411 ( .A(n14364), .B(n14365), .Z(n8089) );
  XNOR U16412 ( .A(n[1022]), .B(n14366), .Z(n14362) );
  IV U16413 ( .A(n14361), .Z(n14366) );
  XOR U16414 ( .A(n14367), .B(n14368), .Z(n14361) );
  AND U16415 ( .A(n14369), .B(n14370), .Z(n14367) );
  XOR U16416 ( .A(n14368), .B(n8100), .Z(n14370) );
  XNOR U16417 ( .A(n14371), .B(n14372), .Z(n8100) );
  XNOR U16418 ( .A(n[1021]), .B(n14373), .Z(n14369) );
  IV U16419 ( .A(n14368), .Z(n14373) );
  XOR U16420 ( .A(n14374), .B(n14375), .Z(n14368) );
  AND U16421 ( .A(n14376), .B(n14377), .Z(n14374) );
  XOR U16422 ( .A(n14375), .B(n8111), .Z(n14377) );
  XNOR U16423 ( .A(n14378), .B(n14379), .Z(n8111) );
  XNOR U16424 ( .A(n[1020]), .B(n14380), .Z(n14376) );
  IV U16425 ( .A(n14375), .Z(n14380) );
  XOR U16426 ( .A(n14381), .B(n14382), .Z(n14375) );
  AND U16427 ( .A(n14383), .B(n14384), .Z(n14381) );
  XOR U16428 ( .A(n14382), .B(n8127), .Z(n14384) );
  XNOR U16429 ( .A(n14385), .B(n14386), .Z(n8127) );
  XNOR U16430 ( .A(n[1019]), .B(n14387), .Z(n14383) );
  IV U16431 ( .A(n14382), .Z(n14387) );
  XOR U16432 ( .A(n14388), .B(n14389), .Z(n14382) );
  AND U16433 ( .A(n14390), .B(n14391), .Z(n14388) );
  XOR U16434 ( .A(n14389), .B(n8138), .Z(n14391) );
  XNOR U16435 ( .A(n14392), .B(n14393), .Z(n8138) );
  XNOR U16436 ( .A(n[1018]), .B(n14394), .Z(n14390) );
  IV U16437 ( .A(n14389), .Z(n14394) );
  XOR U16438 ( .A(n14395), .B(n14396), .Z(n14389) );
  AND U16439 ( .A(n14397), .B(n14398), .Z(n14395) );
  XOR U16440 ( .A(n14396), .B(n8149), .Z(n14398) );
  XNOR U16441 ( .A(n14399), .B(n14400), .Z(n8149) );
  XNOR U16442 ( .A(n[1017]), .B(n14401), .Z(n14397) );
  IV U16443 ( .A(n14396), .Z(n14401) );
  XOR U16444 ( .A(n14402), .B(n14403), .Z(n14396) );
  AND U16445 ( .A(n14404), .B(n14405), .Z(n14402) );
  XOR U16446 ( .A(n14403), .B(n8160), .Z(n14405) );
  XNOR U16447 ( .A(n14406), .B(n14407), .Z(n8160) );
  XNOR U16448 ( .A(n[1016]), .B(n14408), .Z(n14404) );
  IV U16449 ( .A(n14403), .Z(n14408) );
  XOR U16450 ( .A(n14409), .B(n14410), .Z(n14403) );
  AND U16451 ( .A(n14411), .B(n14412), .Z(n14409) );
  XOR U16452 ( .A(n14410), .B(n8171), .Z(n14412) );
  XNOR U16453 ( .A(n14413), .B(n14414), .Z(n8171) );
  XNOR U16454 ( .A(n[1015]), .B(n14415), .Z(n14411) );
  IV U16455 ( .A(n14410), .Z(n14415) );
  XOR U16456 ( .A(n14416), .B(n14417), .Z(n14410) );
  AND U16457 ( .A(n14418), .B(n14419), .Z(n14416) );
  XOR U16458 ( .A(n14417), .B(n8182), .Z(n14419) );
  XNOR U16459 ( .A(n14420), .B(n14421), .Z(n8182) );
  XNOR U16460 ( .A(n[1014]), .B(n14422), .Z(n14418) );
  IV U16461 ( .A(n14417), .Z(n14422) );
  XOR U16462 ( .A(n14423), .B(n14424), .Z(n14417) );
  AND U16463 ( .A(n14425), .B(n14426), .Z(n14423) );
  XOR U16464 ( .A(n14424), .B(n8193), .Z(n14426) );
  XNOR U16465 ( .A(n14427), .B(n14428), .Z(n8193) );
  XNOR U16466 ( .A(n[1013]), .B(n14429), .Z(n14425) );
  IV U16467 ( .A(n14424), .Z(n14429) );
  XOR U16468 ( .A(n14430), .B(n14431), .Z(n14424) );
  AND U16469 ( .A(n14432), .B(n14433), .Z(n14430) );
  XOR U16470 ( .A(n14431), .B(n8204), .Z(n14433) );
  XNOR U16471 ( .A(n14434), .B(n14435), .Z(n8204) );
  XNOR U16472 ( .A(n[1012]), .B(n14436), .Z(n14432) );
  IV U16473 ( .A(n14431), .Z(n14436) );
  XOR U16474 ( .A(n14437), .B(n14438), .Z(n14431) );
  AND U16475 ( .A(n14439), .B(n14440), .Z(n14437) );
  XOR U16476 ( .A(n14438), .B(n8215), .Z(n14440) );
  XNOR U16477 ( .A(n14441), .B(n14442), .Z(n8215) );
  XNOR U16478 ( .A(n[1011]), .B(n14443), .Z(n14439) );
  IV U16479 ( .A(n14438), .Z(n14443) );
  XOR U16480 ( .A(n14444), .B(n14445), .Z(n14438) );
  AND U16481 ( .A(n14446), .B(n14447), .Z(n14444) );
  XOR U16482 ( .A(n14445), .B(n8226), .Z(n14447) );
  XNOR U16483 ( .A(n14448), .B(n14449), .Z(n8226) );
  XNOR U16484 ( .A(n[1010]), .B(n14450), .Z(n14446) );
  IV U16485 ( .A(n14445), .Z(n14450) );
  XOR U16486 ( .A(n14451), .B(n14452), .Z(n14445) );
  AND U16487 ( .A(n14453), .B(n14454), .Z(n14451) );
  XOR U16488 ( .A(n14452), .B(n8242), .Z(n14454) );
  XNOR U16489 ( .A(n14455), .B(n14456), .Z(n8242) );
  XNOR U16490 ( .A(n[1009]), .B(n14457), .Z(n14453) );
  IV U16491 ( .A(n14452), .Z(n14457) );
  XOR U16492 ( .A(n14458), .B(n14459), .Z(n14452) );
  AND U16493 ( .A(n14460), .B(n14461), .Z(n14458) );
  XOR U16494 ( .A(n14459), .B(n8253), .Z(n14461) );
  XNOR U16495 ( .A(n14462), .B(n14463), .Z(n8253) );
  XNOR U16496 ( .A(n[1008]), .B(n14464), .Z(n14460) );
  IV U16497 ( .A(n14459), .Z(n14464) );
  XOR U16498 ( .A(n14465), .B(n14466), .Z(n14459) );
  AND U16499 ( .A(n14467), .B(n14468), .Z(n14465) );
  XOR U16500 ( .A(n14466), .B(n8264), .Z(n14468) );
  XNOR U16501 ( .A(n14469), .B(n14470), .Z(n8264) );
  XNOR U16502 ( .A(n[1007]), .B(n14471), .Z(n14467) );
  IV U16503 ( .A(n14466), .Z(n14471) );
  XOR U16504 ( .A(n14472), .B(n14473), .Z(n14466) );
  AND U16505 ( .A(n14474), .B(n14475), .Z(n14472) );
  XOR U16506 ( .A(n14473), .B(n8275), .Z(n14475) );
  XNOR U16507 ( .A(n14476), .B(n14477), .Z(n8275) );
  XNOR U16508 ( .A(n[1006]), .B(n14478), .Z(n14474) );
  IV U16509 ( .A(n14473), .Z(n14478) );
  XOR U16510 ( .A(n14479), .B(n14480), .Z(n14473) );
  AND U16511 ( .A(n14481), .B(n14482), .Z(n14479) );
  XOR U16512 ( .A(n14480), .B(n8286), .Z(n14482) );
  XNOR U16513 ( .A(n14483), .B(n14484), .Z(n8286) );
  XNOR U16514 ( .A(n[1005]), .B(n14485), .Z(n14481) );
  IV U16515 ( .A(n14480), .Z(n14485) );
  XOR U16516 ( .A(n14486), .B(n14487), .Z(n14480) );
  AND U16517 ( .A(n14488), .B(n14489), .Z(n14486) );
  XOR U16518 ( .A(n14487), .B(n8297), .Z(n14489) );
  XNOR U16519 ( .A(n14490), .B(n14491), .Z(n8297) );
  XNOR U16520 ( .A(n[1004]), .B(n14492), .Z(n14488) );
  IV U16521 ( .A(n14487), .Z(n14492) );
  XOR U16522 ( .A(n14493), .B(n14494), .Z(n14487) );
  AND U16523 ( .A(n14495), .B(n14496), .Z(n14493) );
  XOR U16524 ( .A(n14494), .B(n8308), .Z(n14496) );
  XNOR U16525 ( .A(n14497), .B(n14498), .Z(n8308) );
  XNOR U16526 ( .A(n[1003]), .B(n14499), .Z(n14495) );
  IV U16527 ( .A(n14494), .Z(n14499) );
  XOR U16528 ( .A(n14500), .B(n14501), .Z(n14494) );
  AND U16529 ( .A(n14502), .B(n14503), .Z(n14500) );
  XOR U16530 ( .A(n14501), .B(n8319), .Z(n14503) );
  XNOR U16531 ( .A(n14504), .B(n14505), .Z(n8319) );
  XNOR U16532 ( .A(n[1002]), .B(n14506), .Z(n14502) );
  IV U16533 ( .A(n14501), .Z(n14506) );
  XOR U16534 ( .A(n14507), .B(n14508), .Z(n14501) );
  AND U16535 ( .A(n14509), .B(n14510), .Z(n14507) );
  XOR U16536 ( .A(n14508), .B(n8330), .Z(n14510) );
  XNOR U16537 ( .A(n14511), .B(n14512), .Z(n8330) );
  XNOR U16538 ( .A(n[1001]), .B(n14513), .Z(n14509) );
  IV U16539 ( .A(n14508), .Z(n14513) );
  XOR U16540 ( .A(n14514), .B(n14515), .Z(n14508) );
  AND U16541 ( .A(n14516), .B(n14517), .Z(n14514) );
  XOR U16542 ( .A(n14515), .B(n8341), .Z(n14517) );
  XNOR U16543 ( .A(n14518), .B(n14519), .Z(n8341) );
  XNOR U16544 ( .A(n[1000]), .B(n14520), .Z(n14516) );
  IV U16545 ( .A(n14515), .Z(n14520) );
  XOR U16546 ( .A(n14521), .B(n14522), .Z(n14515) );
  AND U16547 ( .A(n14523), .B(n14524), .Z(n14521) );
  XOR U16548 ( .A(n14522), .B(n8346), .Z(n14524) );
  XNOR U16549 ( .A(n14525), .B(n14526), .Z(n8346) );
  XNOR U16550 ( .A(n[999]), .B(n14527), .Z(n14523) );
  IV U16551 ( .A(n14522), .Z(n14527) );
  XOR U16552 ( .A(n14528), .B(n14529), .Z(n14522) );
  AND U16553 ( .A(n14530), .B(n14531), .Z(n14528) );
  XOR U16554 ( .A(n14529), .B(n8351), .Z(n14531) );
  XNOR U16555 ( .A(n14532), .B(n14533), .Z(n8351) );
  XNOR U16556 ( .A(n[998]), .B(n14534), .Z(n14530) );
  IV U16557 ( .A(n14529), .Z(n14534) );
  XOR U16558 ( .A(n14535), .B(n14536), .Z(n14529) );
  AND U16559 ( .A(n14537), .B(n14538), .Z(n14535) );
  XOR U16560 ( .A(n14536), .B(n8356), .Z(n14538) );
  XNOR U16561 ( .A(n14539), .B(n14540), .Z(n8356) );
  XNOR U16562 ( .A(n[997]), .B(n14541), .Z(n14537) );
  IV U16563 ( .A(n14536), .Z(n14541) );
  XOR U16564 ( .A(n14542), .B(n14543), .Z(n14536) );
  AND U16565 ( .A(n14544), .B(n14545), .Z(n14542) );
  XOR U16566 ( .A(n14543), .B(n8361), .Z(n14545) );
  XNOR U16567 ( .A(n14546), .B(n14547), .Z(n8361) );
  XNOR U16568 ( .A(n[996]), .B(n14548), .Z(n14544) );
  IV U16569 ( .A(n14543), .Z(n14548) );
  XOR U16570 ( .A(n14549), .B(n14550), .Z(n14543) );
  AND U16571 ( .A(n14551), .B(n14552), .Z(n14549) );
  XOR U16572 ( .A(n14550), .B(n8366), .Z(n14552) );
  XNOR U16573 ( .A(n14553), .B(n14554), .Z(n8366) );
  XNOR U16574 ( .A(n[995]), .B(n14555), .Z(n14551) );
  IV U16575 ( .A(n14550), .Z(n14555) );
  XOR U16576 ( .A(n14556), .B(n14557), .Z(n14550) );
  AND U16577 ( .A(n14558), .B(n14559), .Z(n14556) );
  XOR U16578 ( .A(n14557), .B(n8371), .Z(n14559) );
  XNOR U16579 ( .A(n14560), .B(n14561), .Z(n8371) );
  XNOR U16580 ( .A(n[994]), .B(n14562), .Z(n14558) );
  IV U16581 ( .A(n14557), .Z(n14562) );
  XOR U16582 ( .A(n14563), .B(n14564), .Z(n14557) );
  AND U16583 ( .A(n14565), .B(n14566), .Z(n14563) );
  XOR U16584 ( .A(n14564), .B(n8376), .Z(n14566) );
  XNOR U16585 ( .A(n14567), .B(n14568), .Z(n8376) );
  XNOR U16586 ( .A(n[993]), .B(n14569), .Z(n14565) );
  IV U16587 ( .A(n14564), .Z(n14569) );
  XOR U16588 ( .A(n14570), .B(n14571), .Z(n14564) );
  AND U16589 ( .A(n14572), .B(n14573), .Z(n14570) );
  XOR U16590 ( .A(n14571), .B(n8381), .Z(n14573) );
  XNOR U16591 ( .A(n14574), .B(n14575), .Z(n8381) );
  XNOR U16592 ( .A(n[992]), .B(n14576), .Z(n14572) );
  IV U16593 ( .A(n14571), .Z(n14576) );
  XOR U16594 ( .A(n14577), .B(n14578), .Z(n14571) );
  AND U16595 ( .A(n14579), .B(n14580), .Z(n14577) );
  XOR U16596 ( .A(n14578), .B(n8386), .Z(n14580) );
  XNOR U16597 ( .A(n14581), .B(n14582), .Z(n8386) );
  XNOR U16598 ( .A(n[991]), .B(n14583), .Z(n14579) );
  IV U16599 ( .A(n14578), .Z(n14583) );
  XOR U16600 ( .A(n14584), .B(n14585), .Z(n14578) );
  AND U16601 ( .A(n14586), .B(n14587), .Z(n14584) );
  XOR U16602 ( .A(n14585), .B(n8391), .Z(n14587) );
  XNOR U16603 ( .A(n14588), .B(n14589), .Z(n8391) );
  XNOR U16604 ( .A(n[990]), .B(n14590), .Z(n14586) );
  IV U16605 ( .A(n14585), .Z(n14590) );
  XOR U16606 ( .A(n14591), .B(n14592), .Z(n14585) );
  AND U16607 ( .A(n14593), .B(n14594), .Z(n14591) );
  XOR U16608 ( .A(n14592), .B(n8396), .Z(n14594) );
  XNOR U16609 ( .A(n14595), .B(n14596), .Z(n8396) );
  XNOR U16610 ( .A(n[989]), .B(n14597), .Z(n14593) );
  IV U16611 ( .A(n14592), .Z(n14597) );
  XOR U16612 ( .A(n14598), .B(n14599), .Z(n14592) );
  AND U16613 ( .A(n14600), .B(n14601), .Z(n14598) );
  XOR U16614 ( .A(n14599), .B(n8401), .Z(n14601) );
  XNOR U16615 ( .A(n14602), .B(n14603), .Z(n8401) );
  XNOR U16616 ( .A(n[988]), .B(n14604), .Z(n14600) );
  IV U16617 ( .A(n14599), .Z(n14604) );
  XOR U16618 ( .A(n14605), .B(n14606), .Z(n14599) );
  AND U16619 ( .A(n14607), .B(n14608), .Z(n14605) );
  XOR U16620 ( .A(n14606), .B(n8406), .Z(n14608) );
  XNOR U16621 ( .A(n14609), .B(n14610), .Z(n8406) );
  XNOR U16622 ( .A(n[987]), .B(n14611), .Z(n14607) );
  IV U16623 ( .A(n14606), .Z(n14611) );
  XOR U16624 ( .A(n14612), .B(n14613), .Z(n14606) );
  AND U16625 ( .A(n14614), .B(n14615), .Z(n14612) );
  XOR U16626 ( .A(n14613), .B(n8411), .Z(n14615) );
  XNOR U16627 ( .A(n14616), .B(n14617), .Z(n8411) );
  XNOR U16628 ( .A(n[986]), .B(n14618), .Z(n14614) );
  IV U16629 ( .A(n14613), .Z(n14618) );
  XOR U16630 ( .A(n14619), .B(n14620), .Z(n14613) );
  AND U16631 ( .A(n14621), .B(n14622), .Z(n14619) );
  XOR U16632 ( .A(n14620), .B(n8416), .Z(n14622) );
  XNOR U16633 ( .A(n14623), .B(n14624), .Z(n8416) );
  XNOR U16634 ( .A(n[985]), .B(n14625), .Z(n14621) );
  IV U16635 ( .A(n14620), .Z(n14625) );
  XOR U16636 ( .A(n14626), .B(n14627), .Z(n14620) );
  AND U16637 ( .A(n14628), .B(n14629), .Z(n14626) );
  XOR U16638 ( .A(n14627), .B(n8421), .Z(n14629) );
  XNOR U16639 ( .A(n14630), .B(n14631), .Z(n8421) );
  XNOR U16640 ( .A(n[984]), .B(n14632), .Z(n14628) );
  IV U16641 ( .A(n14627), .Z(n14632) );
  XOR U16642 ( .A(n14633), .B(n14634), .Z(n14627) );
  AND U16643 ( .A(n14635), .B(n14636), .Z(n14633) );
  XOR U16644 ( .A(n14634), .B(n8426), .Z(n14636) );
  XNOR U16645 ( .A(n14637), .B(n14638), .Z(n8426) );
  XNOR U16646 ( .A(n[983]), .B(n14639), .Z(n14635) );
  IV U16647 ( .A(n14634), .Z(n14639) );
  XOR U16648 ( .A(n14640), .B(n14641), .Z(n14634) );
  AND U16649 ( .A(n14642), .B(n14643), .Z(n14640) );
  XOR U16650 ( .A(n14641), .B(n8431), .Z(n14643) );
  XNOR U16651 ( .A(n14644), .B(n14645), .Z(n8431) );
  XNOR U16652 ( .A(n[982]), .B(n14646), .Z(n14642) );
  IV U16653 ( .A(n14641), .Z(n14646) );
  XOR U16654 ( .A(n14647), .B(n14648), .Z(n14641) );
  AND U16655 ( .A(n14649), .B(n14650), .Z(n14647) );
  XOR U16656 ( .A(n14648), .B(n8436), .Z(n14650) );
  XNOR U16657 ( .A(n14651), .B(n14652), .Z(n8436) );
  XNOR U16658 ( .A(n[981]), .B(n14653), .Z(n14649) );
  IV U16659 ( .A(n14648), .Z(n14653) );
  XOR U16660 ( .A(n14654), .B(n14655), .Z(n14648) );
  AND U16661 ( .A(n14656), .B(n14657), .Z(n14654) );
  XOR U16662 ( .A(n14655), .B(n8441), .Z(n14657) );
  XNOR U16663 ( .A(n14658), .B(n14659), .Z(n8441) );
  XNOR U16664 ( .A(n[980]), .B(n14660), .Z(n14656) );
  IV U16665 ( .A(n14655), .Z(n14660) );
  XOR U16666 ( .A(n14661), .B(n14662), .Z(n14655) );
  AND U16667 ( .A(n14663), .B(n14664), .Z(n14661) );
  XOR U16668 ( .A(n14662), .B(n8446), .Z(n14664) );
  XNOR U16669 ( .A(n14665), .B(n14666), .Z(n8446) );
  XNOR U16670 ( .A(n[979]), .B(n14667), .Z(n14663) );
  IV U16671 ( .A(n14662), .Z(n14667) );
  XOR U16672 ( .A(n14668), .B(n14669), .Z(n14662) );
  AND U16673 ( .A(n14670), .B(n14671), .Z(n14668) );
  XOR U16674 ( .A(n14669), .B(n8451), .Z(n14671) );
  XNOR U16675 ( .A(n14672), .B(n14673), .Z(n8451) );
  XNOR U16676 ( .A(n[978]), .B(n14674), .Z(n14670) );
  IV U16677 ( .A(n14669), .Z(n14674) );
  XOR U16678 ( .A(n14675), .B(n14676), .Z(n14669) );
  AND U16679 ( .A(n14677), .B(n14678), .Z(n14675) );
  XOR U16680 ( .A(n14676), .B(n8456), .Z(n14678) );
  XNOR U16681 ( .A(n14679), .B(n14680), .Z(n8456) );
  XNOR U16682 ( .A(n[977]), .B(n14681), .Z(n14677) );
  IV U16683 ( .A(n14676), .Z(n14681) );
  XOR U16684 ( .A(n14682), .B(n14683), .Z(n14676) );
  AND U16685 ( .A(n14684), .B(n14685), .Z(n14682) );
  XOR U16686 ( .A(n14683), .B(n8461), .Z(n14685) );
  XNOR U16687 ( .A(n14686), .B(n14687), .Z(n8461) );
  XNOR U16688 ( .A(n[976]), .B(n14688), .Z(n14684) );
  IV U16689 ( .A(n14683), .Z(n14688) );
  XOR U16690 ( .A(n14689), .B(n14690), .Z(n14683) );
  AND U16691 ( .A(n14691), .B(n14692), .Z(n14689) );
  XOR U16692 ( .A(n14690), .B(n8466), .Z(n14692) );
  XNOR U16693 ( .A(n14693), .B(n14694), .Z(n8466) );
  XNOR U16694 ( .A(n[975]), .B(n14695), .Z(n14691) );
  IV U16695 ( .A(n14690), .Z(n14695) );
  XOR U16696 ( .A(n14696), .B(n14697), .Z(n14690) );
  AND U16697 ( .A(n14698), .B(n14699), .Z(n14696) );
  XOR U16698 ( .A(n14697), .B(n8471), .Z(n14699) );
  XNOR U16699 ( .A(n14700), .B(n14701), .Z(n8471) );
  XNOR U16700 ( .A(n[974]), .B(n14702), .Z(n14698) );
  IV U16701 ( .A(n14697), .Z(n14702) );
  XOR U16702 ( .A(n14703), .B(n14704), .Z(n14697) );
  AND U16703 ( .A(n14705), .B(n14706), .Z(n14703) );
  XOR U16704 ( .A(n14704), .B(n8476), .Z(n14706) );
  XNOR U16705 ( .A(n14707), .B(n14708), .Z(n8476) );
  XNOR U16706 ( .A(n[973]), .B(n14709), .Z(n14705) );
  IV U16707 ( .A(n14704), .Z(n14709) );
  XOR U16708 ( .A(n14710), .B(n14711), .Z(n14704) );
  AND U16709 ( .A(n14712), .B(n14713), .Z(n14710) );
  XOR U16710 ( .A(n14711), .B(n8481), .Z(n14713) );
  XNOR U16711 ( .A(n14714), .B(n14715), .Z(n8481) );
  XNOR U16712 ( .A(n[972]), .B(n14716), .Z(n14712) );
  IV U16713 ( .A(n14711), .Z(n14716) );
  XOR U16714 ( .A(n14717), .B(n14718), .Z(n14711) );
  AND U16715 ( .A(n14719), .B(n14720), .Z(n14717) );
  XOR U16716 ( .A(n14718), .B(n8486), .Z(n14720) );
  XNOR U16717 ( .A(n14721), .B(n14722), .Z(n8486) );
  XNOR U16718 ( .A(n[971]), .B(n14723), .Z(n14719) );
  IV U16719 ( .A(n14718), .Z(n14723) );
  XOR U16720 ( .A(n14724), .B(n14725), .Z(n14718) );
  AND U16721 ( .A(n14726), .B(n14727), .Z(n14724) );
  XOR U16722 ( .A(n14725), .B(n8491), .Z(n14727) );
  XNOR U16723 ( .A(n14728), .B(n14729), .Z(n8491) );
  XNOR U16724 ( .A(n[970]), .B(n14730), .Z(n14726) );
  IV U16725 ( .A(n14725), .Z(n14730) );
  XOR U16726 ( .A(n14731), .B(n14732), .Z(n14725) );
  AND U16727 ( .A(n14733), .B(n14734), .Z(n14731) );
  XOR U16728 ( .A(n14732), .B(n8496), .Z(n14734) );
  XNOR U16729 ( .A(n14735), .B(n14736), .Z(n8496) );
  XNOR U16730 ( .A(n[969]), .B(n14737), .Z(n14733) );
  IV U16731 ( .A(n14732), .Z(n14737) );
  XOR U16732 ( .A(n14738), .B(n14739), .Z(n14732) );
  AND U16733 ( .A(n14740), .B(n14741), .Z(n14738) );
  XOR U16734 ( .A(n14739), .B(n8501), .Z(n14741) );
  XNOR U16735 ( .A(n14742), .B(n14743), .Z(n8501) );
  XNOR U16736 ( .A(n[968]), .B(n14744), .Z(n14740) );
  IV U16737 ( .A(n14739), .Z(n14744) );
  XOR U16738 ( .A(n14745), .B(n14746), .Z(n14739) );
  AND U16739 ( .A(n14747), .B(n14748), .Z(n14745) );
  XOR U16740 ( .A(n14746), .B(n8506), .Z(n14748) );
  XNOR U16741 ( .A(n14749), .B(n14750), .Z(n8506) );
  XNOR U16742 ( .A(n[967]), .B(n14751), .Z(n14747) );
  IV U16743 ( .A(n14746), .Z(n14751) );
  XOR U16744 ( .A(n14752), .B(n14753), .Z(n14746) );
  AND U16745 ( .A(n14754), .B(n14755), .Z(n14752) );
  XOR U16746 ( .A(n14753), .B(n8511), .Z(n14755) );
  XNOR U16747 ( .A(n14756), .B(n14757), .Z(n8511) );
  XNOR U16748 ( .A(n[966]), .B(n14758), .Z(n14754) );
  IV U16749 ( .A(n14753), .Z(n14758) );
  XOR U16750 ( .A(n14759), .B(n14760), .Z(n14753) );
  AND U16751 ( .A(n14761), .B(n14762), .Z(n14759) );
  XOR U16752 ( .A(n14760), .B(n8516), .Z(n14762) );
  XNOR U16753 ( .A(n14763), .B(n14764), .Z(n8516) );
  XNOR U16754 ( .A(n[965]), .B(n14765), .Z(n14761) );
  IV U16755 ( .A(n14760), .Z(n14765) );
  XOR U16756 ( .A(n14766), .B(n14767), .Z(n14760) );
  AND U16757 ( .A(n14768), .B(n14769), .Z(n14766) );
  XOR U16758 ( .A(n14767), .B(n8521), .Z(n14769) );
  XNOR U16759 ( .A(n14770), .B(n14771), .Z(n8521) );
  XNOR U16760 ( .A(n[964]), .B(n14772), .Z(n14768) );
  IV U16761 ( .A(n14767), .Z(n14772) );
  XOR U16762 ( .A(n14773), .B(n14774), .Z(n14767) );
  AND U16763 ( .A(n14775), .B(n14776), .Z(n14773) );
  XOR U16764 ( .A(n14774), .B(n8526), .Z(n14776) );
  XNOR U16765 ( .A(n14777), .B(n14778), .Z(n8526) );
  XNOR U16766 ( .A(n[963]), .B(n14779), .Z(n14775) );
  IV U16767 ( .A(n14774), .Z(n14779) );
  XOR U16768 ( .A(n14780), .B(n14781), .Z(n14774) );
  AND U16769 ( .A(n14782), .B(n14783), .Z(n14780) );
  XOR U16770 ( .A(n14781), .B(n8531), .Z(n14783) );
  XNOR U16771 ( .A(n14784), .B(n14785), .Z(n8531) );
  XNOR U16772 ( .A(n[962]), .B(n14786), .Z(n14782) );
  IV U16773 ( .A(n14781), .Z(n14786) );
  XOR U16774 ( .A(n14787), .B(n14788), .Z(n14781) );
  AND U16775 ( .A(n14789), .B(n14790), .Z(n14787) );
  XOR U16776 ( .A(n14788), .B(n8536), .Z(n14790) );
  XNOR U16777 ( .A(n14791), .B(n14792), .Z(n8536) );
  XNOR U16778 ( .A(n[961]), .B(n14793), .Z(n14789) );
  IV U16779 ( .A(n14788), .Z(n14793) );
  XOR U16780 ( .A(n14794), .B(n14795), .Z(n14788) );
  AND U16781 ( .A(n14796), .B(n14797), .Z(n14794) );
  XOR U16782 ( .A(n14795), .B(n8541), .Z(n14797) );
  XNOR U16783 ( .A(n14798), .B(n14799), .Z(n8541) );
  XNOR U16784 ( .A(n[960]), .B(n14800), .Z(n14796) );
  IV U16785 ( .A(n14795), .Z(n14800) );
  XOR U16786 ( .A(n14801), .B(n14802), .Z(n14795) );
  AND U16787 ( .A(n14803), .B(n14804), .Z(n14801) );
  XOR U16788 ( .A(n14802), .B(n8546), .Z(n14804) );
  XNOR U16789 ( .A(n14805), .B(n14806), .Z(n8546) );
  XNOR U16790 ( .A(n[959]), .B(n14807), .Z(n14803) );
  IV U16791 ( .A(n14802), .Z(n14807) );
  XOR U16792 ( .A(n14808), .B(n14809), .Z(n14802) );
  AND U16793 ( .A(n14810), .B(n14811), .Z(n14808) );
  XOR U16794 ( .A(n14809), .B(n8551), .Z(n14811) );
  XNOR U16795 ( .A(n14812), .B(n14813), .Z(n8551) );
  XNOR U16796 ( .A(n[958]), .B(n14814), .Z(n14810) );
  IV U16797 ( .A(n14809), .Z(n14814) );
  XOR U16798 ( .A(n14815), .B(n14816), .Z(n14809) );
  AND U16799 ( .A(n14817), .B(n14818), .Z(n14815) );
  XOR U16800 ( .A(n14816), .B(n8556), .Z(n14818) );
  XNOR U16801 ( .A(n14819), .B(n14820), .Z(n8556) );
  XNOR U16802 ( .A(n[957]), .B(n14821), .Z(n14817) );
  IV U16803 ( .A(n14816), .Z(n14821) );
  XOR U16804 ( .A(n14822), .B(n14823), .Z(n14816) );
  AND U16805 ( .A(n14824), .B(n14825), .Z(n14822) );
  XOR U16806 ( .A(n14823), .B(n8561), .Z(n14825) );
  XNOR U16807 ( .A(n14826), .B(n14827), .Z(n8561) );
  XNOR U16808 ( .A(n[956]), .B(n14828), .Z(n14824) );
  IV U16809 ( .A(n14823), .Z(n14828) );
  XOR U16810 ( .A(n14829), .B(n14830), .Z(n14823) );
  AND U16811 ( .A(n14831), .B(n14832), .Z(n14829) );
  XOR U16812 ( .A(n14830), .B(n8566), .Z(n14832) );
  XNOR U16813 ( .A(n14833), .B(n14834), .Z(n8566) );
  XNOR U16814 ( .A(n[955]), .B(n14835), .Z(n14831) );
  IV U16815 ( .A(n14830), .Z(n14835) );
  XOR U16816 ( .A(n14836), .B(n14837), .Z(n14830) );
  AND U16817 ( .A(n14838), .B(n14839), .Z(n14836) );
  XOR U16818 ( .A(n14837), .B(n8571), .Z(n14839) );
  XNOR U16819 ( .A(n14840), .B(n14841), .Z(n8571) );
  XNOR U16820 ( .A(n[954]), .B(n14842), .Z(n14838) );
  IV U16821 ( .A(n14837), .Z(n14842) );
  XOR U16822 ( .A(n14843), .B(n14844), .Z(n14837) );
  AND U16823 ( .A(n14845), .B(n14846), .Z(n14843) );
  XOR U16824 ( .A(n14844), .B(n8576), .Z(n14846) );
  XNOR U16825 ( .A(n14847), .B(n14848), .Z(n8576) );
  XNOR U16826 ( .A(n[953]), .B(n14849), .Z(n14845) );
  IV U16827 ( .A(n14844), .Z(n14849) );
  XOR U16828 ( .A(n14850), .B(n14851), .Z(n14844) );
  AND U16829 ( .A(n14852), .B(n14853), .Z(n14850) );
  XOR U16830 ( .A(n14851), .B(n8581), .Z(n14853) );
  XNOR U16831 ( .A(n14854), .B(n14855), .Z(n8581) );
  XNOR U16832 ( .A(n[952]), .B(n14856), .Z(n14852) );
  IV U16833 ( .A(n14851), .Z(n14856) );
  XOR U16834 ( .A(n14857), .B(n14858), .Z(n14851) );
  AND U16835 ( .A(n14859), .B(n14860), .Z(n14857) );
  XOR U16836 ( .A(n14858), .B(n8586), .Z(n14860) );
  XNOR U16837 ( .A(n14861), .B(n14862), .Z(n8586) );
  XNOR U16838 ( .A(n[951]), .B(n14863), .Z(n14859) );
  IV U16839 ( .A(n14858), .Z(n14863) );
  XOR U16840 ( .A(n14864), .B(n14865), .Z(n14858) );
  AND U16841 ( .A(n14866), .B(n14867), .Z(n14864) );
  XOR U16842 ( .A(n14865), .B(n8591), .Z(n14867) );
  XNOR U16843 ( .A(n14868), .B(n14869), .Z(n8591) );
  XNOR U16844 ( .A(n[950]), .B(n14870), .Z(n14866) );
  IV U16845 ( .A(n14865), .Z(n14870) );
  XOR U16846 ( .A(n14871), .B(n14872), .Z(n14865) );
  AND U16847 ( .A(n14873), .B(n14874), .Z(n14871) );
  XOR U16848 ( .A(n14872), .B(n8596), .Z(n14874) );
  XNOR U16849 ( .A(n14875), .B(n14876), .Z(n8596) );
  XNOR U16850 ( .A(n[949]), .B(n14877), .Z(n14873) );
  IV U16851 ( .A(n14872), .Z(n14877) );
  XOR U16852 ( .A(n14878), .B(n14879), .Z(n14872) );
  AND U16853 ( .A(n14880), .B(n14881), .Z(n14878) );
  XOR U16854 ( .A(n14879), .B(n8601), .Z(n14881) );
  XNOR U16855 ( .A(n14882), .B(n14883), .Z(n8601) );
  XNOR U16856 ( .A(n[948]), .B(n14884), .Z(n14880) );
  IV U16857 ( .A(n14879), .Z(n14884) );
  XOR U16858 ( .A(n14885), .B(n14886), .Z(n14879) );
  AND U16859 ( .A(n14887), .B(n14888), .Z(n14885) );
  XOR U16860 ( .A(n14886), .B(n8606), .Z(n14888) );
  XNOR U16861 ( .A(n14889), .B(n14890), .Z(n8606) );
  XNOR U16862 ( .A(n[947]), .B(n14891), .Z(n14887) );
  IV U16863 ( .A(n14886), .Z(n14891) );
  XOR U16864 ( .A(n14892), .B(n14893), .Z(n14886) );
  AND U16865 ( .A(n14894), .B(n14895), .Z(n14892) );
  XOR U16866 ( .A(n14893), .B(n8611), .Z(n14895) );
  XNOR U16867 ( .A(n14896), .B(n14897), .Z(n8611) );
  XNOR U16868 ( .A(n[946]), .B(n14898), .Z(n14894) );
  IV U16869 ( .A(n14893), .Z(n14898) );
  XOR U16870 ( .A(n14899), .B(n14900), .Z(n14893) );
  AND U16871 ( .A(n14901), .B(n14902), .Z(n14899) );
  XOR U16872 ( .A(n14900), .B(n8616), .Z(n14902) );
  XNOR U16873 ( .A(n14903), .B(n14904), .Z(n8616) );
  XNOR U16874 ( .A(n[945]), .B(n14905), .Z(n14901) );
  IV U16875 ( .A(n14900), .Z(n14905) );
  XOR U16876 ( .A(n14906), .B(n14907), .Z(n14900) );
  AND U16877 ( .A(n14908), .B(n14909), .Z(n14906) );
  XOR U16878 ( .A(n14907), .B(n8621), .Z(n14909) );
  XNOR U16879 ( .A(n14910), .B(n14911), .Z(n8621) );
  XNOR U16880 ( .A(n[944]), .B(n14912), .Z(n14908) );
  IV U16881 ( .A(n14907), .Z(n14912) );
  XOR U16882 ( .A(n14913), .B(n14914), .Z(n14907) );
  AND U16883 ( .A(n14915), .B(n14916), .Z(n14913) );
  XOR U16884 ( .A(n14914), .B(n8626), .Z(n14916) );
  XNOR U16885 ( .A(n14917), .B(n14918), .Z(n8626) );
  XNOR U16886 ( .A(n[943]), .B(n14919), .Z(n14915) );
  IV U16887 ( .A(n14914), .Z(n14919) );
  XOR U16888 ( .A(n14920), .B(n14921), .Z(n14914) );
  AND U16889 ( .A(n14922), .B(n14923), .Z(n14920) );
  XOR U16890 ( .A(n14921), .B(n8631), .Z(n14923) );
  XNOR U16891 ( .A(n14924), .B(n14925), .Z(n8631) );
  XNOR U16892 ( .A(n[942]), .B(n14926), .Z(n14922) );
  IV U16893 ( .A(n14921), .Z(n14926) );
  XOR U16894 ( .A(n14927), .B(n14928), .Z(n14921) );
  AND U16895 ( .A(n14929), .B(n14930), .Z(n14927) );
  XOR U16896 ( .A(n14928), .B(n8636), .Z(n14930) );
  XNOR U16897 ( .A(n14931), .B(n14932), .Z(n8636) );
  XNOR U16898 ( .A(n[941]), .B(n14933), .Z(n14929) );
  IV U16899 ( .A(n14928), .Z(n14933) );
  XOR U16900 ( .A(n14934), .B(n14935), .Z(n14928) );
  AND U16901 ( .A(n14936), .B(n14937), .Z(n14934) );
  XOR U16902 ( .A(n14935), .B(n8641), .Z(n14937) );
  XNOR U16903 ( .A(n14938), .B(n14939), .Z(n8641) );
  XNOR U16904 ( .A(n[940]), .B(n14940), .Z(n14936) );
  IV U16905 ( .A(n14935), .Z(n14940) );
  XOR U16906 ( .A(n14941), .B(n14942), .Z(n14935) );
  AND U16907 ( .A(n14943), .B(n14944), .Z(n14941) );
  XOR U16908 ( .A(n14942), .B(n8646), .Z(n14944) );
  XNOR U16909 ( .A(n14945), .B(n14946), .Z(n8646) );
  XNOR U16910 ( .A(n[939]), .B(n14947), .Z(n14943) );
  IV U16911 ( .A(n14942), .Z(n14947) );
  XOR U16912 ( .A(n14948), .B(n14949), .Z(n14942) );
  AND U16913 ( .A(n14950), .B(n14951), .Z(n14948) );
  XOR U16914 ( .A(n14949), .B(n8651), .Z(n14951) );
  XNOR U16915 ( .A(n14952), .B(n14953), .Z(n8651) );
  XNOR U16916 ( .A(n[938]), .B(n14954), .Z(n14950) );
  IV U16917 ( .A(n14949), .Z(n14954) );
  XOR U16918 ( .A(n14955), .B(n14956), .Z(n14949) );
  AND U16919 ( .A(n14957), .B(n14958), .Z(n14955) );
  XOR U16920 ( .A(n14956), .B(n8656), .Z(n14958) );
  XNOR U16921 ( .A(n14959), .B(n14960), .Z(n8656) );
  XNOR U16922 ( .A(n[937]), .B(n14961), .Z(n14957) );
  IV U16923 ( .A(n14956), .Z(n14961) );
  XOR U16924 ( .A(n14962), .B(n14963), .Z(n14956) );
  AND U16925 ( .A(n14964), .B(n14965), .Z(n14962) );
  XOR U16926 ( .A(n14963), .B(n8661), .Z(n14965) );
  XNOR U16927 ( .A(n14966), .B(n14967), .Z(n8661) );
  XNOR U16928 ( .A(n[936]), .B(n14968), .Z(n14964) );
  IV U16929 ( .A(n14963), .Z(n14968) );
  XOR U16930 ( .A(n14969), .B(n14970), .Z(n14963) );
  AND U16931 ( .A(n14971), .B(n14972), .Z(n14969) );
  XOR U16932 ( .A(n14970), .B(n8666), .Z(n14972) );
  XNOR U16933 ( .A(n14973), .B(n14974), .Z(n8666) );
  XNOR U16934 ( .A(n[935]), .B(n14975), .Z(n14971) );
  IV U16935 ( .A(n14970), .Z(n14975) );
  XOR U16936 ( .A(n14976), .B(n14977), .Z(n14970) );
  AND U16937 ( .A(n14978), .B(n14979), .Z(n14976) );
  XOR U16938 ( .A(n14977), .B(n8671), .Z(n14979) );
  XNOR U16939 ( .A(n14980), .B(n14981), .Z(n8671) );
  XNOR U16940 ( .A(n[934]), .B(n14982), .Z(n14978) );
  IV U16941 ( .A(n14977), .Z(n14982) );
  XOR U16942 ( .A(n14983), .B(n14984), .Z(n14977) );
  AND U16943 ( .A(n14985), .B(n14986), .Z(n14983) );
  XOR U16944 ( .A(n14984), .B(n8676), .Z(n14986) );
  XNOR U16945 ( .A(n14987), .B(n14988), .Z(n8676) );
  XNOR U16946 ( .A(n[933]), .B(n14989), .Z(n14985) );
  IV U16947 ( .A(n14984), .Z(n14989) );
  XOR U16948 ( .A(n14990), .B(n14991), .Z(n14984) );
  AND U16949 ( .A(n14992), .B(n14993), .Z(n14990) );
  XOR U16950 ( .A(n14991), .B(n8681), .Z(n14993) );
  XNOR U16951 ( .A(n14994), .B(n14995), .Z(n8681) );
  XNOR U16952 ( .A(n[932]), .B(n14996), .Z(n14992) );
  IV U16953 ( .A(n14991), .Z(n14996) );
  XOR U16954 ( .A(n14997), .B(n14998), .Z(n14991) );
  AND U16955 ( .A(n14999), .B(n15000), .Z(n14997) );
  XOR U16956 ( .A(n14998), .B(n8686), .Z(n15000) );
  XNOR U16957 ( .A(n15001), .B(n15002), .Z(n8686) );
  XNOR U16958 ( .A(n[931]), .B(n15003), .Z(n14999) );
  IV U16959 ( .A(n14998), .Z(n15003) );
  XOR U16960 ( .A(n15004), .B(n15005), .Z(n14998) );
  AND U16961 ( .A(n15006), .B(n15007), .Z(n15004) );
  XOR U16962 ( .A(n15005), .B(n8691), .Z(n15007) );
  XNOR U16963 ( .A(n15008), .B(n15009), .Z(n8691) );
  XNOR U16964 ( .A(n[930]), .B(n15010), .Z(n15006) );
  IV U16965 ( .A(n15005), .Z(n15010) );
  XOR U16966 ( .A(n15011), .B(n15012), .Z(n15005) );
  AND U16967 ( .A(n15013), .B(n15014), .Z(n15011) );
  XOR U16968 ( .A(n15012), .B(n8696), .Z(n15014) );
  XNOR U16969 ( .A(n15015), .B(n15016), .Z(n8696) );
  XNOR U16970 ( .A(n[929]), .B(n15017), .Z(n15013) );
  IV U16971 ( .A(n15012), .Z(n15017) );
  XOR U16972 ( .A(n15018), .B(n15019), .Z(n15012) );
  AND U16973 ( .A(n15020), .B(n15021), .Z(n15018) );
  XOR U16974 ( .A(n15019), .B(n8701), .Z(n15021) );
  XNOR U16975 ( .A(n15022), .B(n15023), .Z(n8701) );
  XNOR U16976 ( .A(n[928]), .B(n15024), .Z(n15020) );
  IV U16977 ( .A(n15019), .Z(n15024) );
  XOR U16978 ( .A(n15025), .B(n15026), .Z(n15019) );
  AND U16979 ( .A(n15027), .B(n15028), .Z(n15025) );
  XOR U16980 ( .A(n15026), .B(n8706), .Z(n15028) );
  XNOR U16981 ( .A(n15029), .B(n15030), .Z(n8706) );
  XNOR U16982 ( .A(n[927]), .B(n15031), .Z(n15027) );
  IV U16983 ( .A(n15026), .Z(n15031) );
  XOR U16984 ( .A(n15032), .B(n15033), .Z(n15026) );
  AND U16985 ( .A(n15034), .B(n15035), .Z(n15032) );
  XOR U16986 ( .A(n15033), .B(n8711), .Z(n15035) );
  XNOR U16987 ( .A(n15036), .B(n15037), .Z(n8711) );
  XNOR U16988 ( .A(n[926]), .B(n15038), .Z(n15034) );
  IV U16989 ( .A(n15033), .Z(n15038) );
  XOR U16990 ( .A(n15039), .B(n15040), .Z(n15033) );
  AND U16991 ( .A(n15041), .B(n15042), .Z(n15039) );
  XOR U16992 ( .A(n15040), .B(n8716), .Z(n15042) );
  XNOR U16993 ( .A(n15043), .B(n15044), .Z(n8716) );
  XNOR U16994 ( .A(n[925]), .B(n15045), .Z(n15041) );
  IV U16995 ( .A(n15040), .Z(n15045) );
  XOR U16996 ( .A(n15046), .B(n15047), .Z(n15040) );
  AND U16997 ( .A(n15048), .B(n15049), .Z(n15046) );
  XOR U16998 ( .A(n15047), .B(n8721), .Z(n15049) );
  XNOR U16999 ( .A(n15050), .B(n15051), .Z(n8721) );
  XNOR U17000 ( .A(n[924]), .B(n15052), .Z(n15048) );
  IV U17001 ( .A(n15047), .Z(n15052) );
  XOR U17002 ( .A(n15053), .B(n15054), .Z(n15047) );
  AND U17003 ( .A(n15055), .B(n15056), .Z(n15053) );
  XOR U17004 ( .A(n15054), .B(n8726), .Z(n15056) );
  XNOR U17005 ( .A(n15057), .B(n15058), .Z(n8726) );
  XNOR U17006 ( .A(n[923]), .B(n15059), .Z(n15055) );
  IV U17007 ( .A(n15054), .Z(n15059) );
  XOR U17008 ( .A(n15060), .B(n15061), .Z(n15054) );
  AND U17009 ( .A(n15062), .B(n15063), .Z(n15060) );
  XOR U17010 ( .A(n15061), .B(n8731), .Z(n15063) );
  XNOR U17011 ( .A(n15064), .B(n15065), .Z(n8731) );
  XNOR U17012 ( .A(n[922]), .B(n15066), .Z(n15062) );
  IV U17013 ( .A(n15061), .Z(n15066) );
  XOR U17014 ( .A(n15067), .B(n15068), .Z(n15061) );
  AND U17015 ( .A(n15069), .B(n15070), .Z(n15067) );
  XOR U17016 ( .A(n15068), .B(n8736), .Z(n15070) );
  XNOR U17017 ( .A(n15071), .B(n15072), .Z(n8736) );
  XNOR U17018 ( .A(n[921]), .B(n15073), .Z(n15069) );
  IV U17019 ( .A(n15068), .Z(n15073) );
  XOR U17020 ( .A(n15074), .B(n15075), .Z(n15068) );
  AND U17021 ( .A(n15076), .B(n15077), .Z(n15074) );
  XOR U17022 ( .A(n15075), .B(n8741), .Z(n15077) );
  XNOR U17023 ( .A(n15078), .B(n15079), .Z(n8741) );
  XNOR U17024 ( .A(n[920]), .B(n15080), .Z(n15076) );
  IV U17025 ( .A(n15075), .Z(n15080) );
  XOR U17026 ( .A(n15081), .B(n15082), .Z(n15075) );
  AND U17027 ( .A(n15083), .B(n15084), .Z(n15081) );
  XOR U17028 ( .A(n15082), .B(n8746), .Z(n15084) );
  XNOR U17029 ( .A(n15085), .B(n15086), .Z(n8746) );
  XNOR U17030 ( .A(n[919]), .B(n15087), .Z(n15083) );
  IV U17031 ( .A(n15082), .Z(n15087) );
  XOR U17032 ( .A(n15088), .B(n15089), .Z(n15082) );
  AND U17033 ( .A(n15090), .B(n15091), .Z(n15088) );
  XOR U17034 ( .A(n15089), .B(n8751), .Z(n15091) );
  XNOR U17035 ( .A(n15092), .B(n15093), .Z(n8751) );
  XNOR U17036 ( .A(n[918]), .B(n15094), .Z(n15090) );
  IV U17037 ( .A(n15089), .Z(n15094) );
  XOR U17038 ( .A(n15095), .B(n15096), .Z(n15089) );
  AND U17039 ( .A(n15097), .B(n15098), .Z(n15095) );
  XOR U17040 ( .A(n15096), .B(n8756), .Z(n15098) );
  XNOR U17041 ( .A(n15099), .B(n15100), .Z(n8756) );
  XNOR U17042 ( .A(n[917]), .B(n15101), .Z(n15097) );
  IV U17043 ( .A(n15096), .Z(n15101) );
  XOR U17044 ( .A(n15102), .B(n15103), .Z(n15096) );
  AND U17045 ( .A(n15104), .B(n15105), .Z(n15102) );
  XOR U17046 ( .A(n15103), .B(n8761), .Z(n15105) );
  XNOR U17047 ( .A(n15106), .B(n15107), .Z(n8761) );
  XNOR U17048 ( .A(n[916]), .B(n15108), .Z(n15104) );
  IV U17049 ( .A(n15103), .Z(n15108) );
  XOR U17050 ( .A(n15109), .B(n15110), .Z(n15103) );
  AND U17051 ( .A(n15111), .B(n15112), .Z(n15109) );
  XOR U17052 ( .A(n15110), .B(n8766), .Z(n15112) );
  XNOR U17053 ( .A(n15113), .B(n15114), .Z(n8766) );
  XNOR U17054 ( .A(n[915]), .B(n15115), .Z(n15111) );
  IV U17055 ( .A(n15110), .Z(n15115) );
  XOR U17056 ( .A(n15116), .B(n15117), .Z(n15110) );
  AND U17057 ( .A(n15118), .B(n15119), .Z(n15116) );
  XOR U17058 ( .A(n15117), .B(n8771), .Z(n15119) );
  XNOR U17059 ( .A(n15120), .B(n15121), .Z(n8771) );
  XNOR U17060 ( .A(n[914]), .B(n15122), .Z(n15118) );
  IV U17061 ( .A(n15117), .Z(n15122) );
  XOR U17062 ( .A(n15123), .B(n15124), .Z(n15117) );
  AND U17063 ( .A(n15125), .B(n15126), .Z(n15123) );
  XOR U17064 ( .A(n15124), .B(n8776), .Z(n15126) );
  XNOR U17065 ( .A(n15127), .B(n15128), .Z(n8776) );
  XNOR U17066 ( .A(n[913]), .B(n15129), .Z(n15125) );
  IV U17067 ( .A(n15124), .Z(n15129) );
  XOR U17068 ( .A(n15130), .B(n15131), .Z(n15124) );
  AND U17069 ( .A(n15132), .B(n15133), .Z(n15130) );
  XOR U17070 ( .A(n15131), .B(n8781), .Z(n15133) );
  XNOR U17071 ( .A(n15134), .B(n15135), .Z(n8781) );
  XNOR U17072 ( .A(n[912]), .B(n15136), .Z(n15132) );
  IV U17073 ( .A(n15131), .Z(n15136) );
  XOR U17074 ( .A(n15137), .B(n15138), .Z(n15131) );
  AND U17075 ( .A(n15139), .B(n15140), .Z(n15137) );
  XOR U17076 ( .A(n15138), .B(n8786), .Z(n15140) );
  XNOR U17077 ( .A(n15141), .B(n15142), .Z(n8786) );
  XNOR U17078 ( .A(n[911]), .B(n15143), .Z(n15139) );
  IV U17079 ( .A(n15138), .Z(n15143) );
  XOR U17080 ( .A(n15144), .B(n15145), .Z(n15138) );
  AND U17081 ( .A(n15146), .B(n15147), .Z(n15144) );
  XOR U17082 ( .A(n15145), .B(n8791), .Z(n15147) );
  XNOR U17083 ( .A(n15148), .B(n15149), .Z(n8791) );
  XNOR U17084 ( .A(n[910]), .B(n15150), .Z(n15146) );
  IV U17085 ( .A(n15145), .Z(n15150) );
  XOR U17086 ( .A(n15151), .B(n15152), .Z(n15145) );
  AND U17087 ( .A(n15153), .B(n15154), .Z(n15151) );
  XOR U17088 ( .A(n15152), .B(n8796), .Z(n15154) );
  XNOR U17089 ( .A(n15155), .B(n15156), .Z(n8796) );
  XNOR U17090 ( .A(n[909]), .B(n15157), .Z(n15153) );
  IV U17091 ( .A(n15152), .Z(n15157) );
  XOR U17092 ( .A(n15158), .B(n15159), .Z(n15152) );
  AND U17093 ( .A(n15160), .B(n15161), .Z(n15158) );
  XOR U17094 ( .A(n15159), .B(n8801), .Z(n15161) );
  XNOR U17095 ( .A(n15162), .B(n15163), .Z(n8801) );
  XNOR U17096 ( .A(n[908]), .B(n15164), .Z(n15160) );
  IV U17097 ( .A(n15159), .Z(n15164) );
  XOR U17098 ( .A(n15165), .B(n15166), .Z(n15159) );
  AND U17099 ( .A(n15167), .B(n15168), .Z(n15165) );
  XOR U17100 ( .A(n15166), .B(n8806), .Z(n15168) );
  XNOR U17101 ( .A(n15169), .B(n15170), .Z(n8806) );
  XNOR U17102 ( .A(n[907]), .B(n15171), .Z(n15167) );
  IV U17103 ( .A(n15166), .Z(n15171) );
  XOR U17104 ( .A(n15172), .B(n15173), .Z(n15166) );
  AND U17105 ( .A(n15174), .B(n15175), .Z(n15172) );
  XOR U17106 ( .A(n15173), .B(n8811), .Z(n15175) );
  XNOR U17107 ( .A(n15176), .B(n15177), .Z(n8811) );
  XNOR U17108 ( .A(n[906]), .B(n15178), .Z(n15174) );
  IV U17109 ( .A(n15173), .Z(n15178) );
  XOR U17110 ( .A(n15179), .B(n15180), .Z(n15173) );
  AND U17111 ( .A(n15181), .B(n15182), .Z(n15179) );
  XOR U17112 ( .A(n15180), .B(n8816), .Z(n15182) );
  XNOR U17113 ( .A(n15183), .B(n15184), .Z(n8816) );
  XNOR U17114 ( .A(n[905]), .B(n15185), .Z(n15181) );
  IV U17115 ( .A(n15180), .Z(n15185) );
  XOR U17116 ( .A(n15186), .B(n15187), .Z(n15180) );
  AND U17117 ( .A(n15188), .B(n15189), .Z(n15186) );
  XOR U17118 ( .A(n15187), .B(n8821), .Z(n15189) );
  XNOR U17119 ( .A(n15190), .B(n15191), .Z(n8821) );
  XNOR U17120 ( .A(n[904]), .B(n15192), .Z(n15188) );
  IV U17121 ( .A(n15187), .Z(n15192) );
  XOR U17122 ( .A(n15193), .B(n15194), .Z(n15187) );
  AND U17123 ( .A(n15195), .B(n15196), .Z(n15193) );
  XOR U17124 ( .A(n15194), .B(n8826), .Z(n15196) );
  XNOR U17125 ( .A(n15197), .B(n15198), .Z(n8826) );
  XNOR U17126 ( .A(n[903]), .B(n15199), .Z(n15195) );
  IV U17127 ( .A(n15194), .Z(n15199) );
  XOR U17128 ( .A(n15200), .B(n15201), .Z(n15194) );
  AND U17129 ( .A(n15202), .B(n15203), .Z(n15200) );
  XOR U17130 ( .A(n15201), .B(n8831), .Z(n15203) );
  XNOR U17131 ( .A(n15204), .B(n15205), .Z(n8831) );
  XNOR U17132 ( .A(n[902]), .B(n15206), .Z(n15202) );
  IV U17133 ( .A(n15201), .Z(n15206) );
  XOR U17134 ( .A(n15207), .B(n15208), .Z(n15201) );
  AND U17135 ( .A(n15209), .B(n15210), .Z(n15207) );
  XOR U17136 ( .A(n15208), .B(n8836), .Z(n15210) );
  XNOR U17137 ( .A(n15211), .B(n15212), .Z(n8836) );
  XNOR U17138 ( .A(n[901]), .B(n15213), .Z(n15209) );
  IV U17139 ( .A(n15208), .Z(n15213) );
  XOR U17140 ( .A(n15214), .B(n15215), .Z(n15208) );
  AND U17141 ( .A(n15216), .B(n15217), .Z(n15214) );
  XOR U17142 ( .A(n15215), .B(n8841), .Z(n15217) );
  XNOR U17143 ( .A(n15218), .B(n15219), .Z(n8841) );
  XNOR U17144 ( .A(n[900]), .B(n15220), .Z(n15216) );
  IV U17145 ( .A(n15215), .Z(n15220) );
  XOR U17146 ( .A(n15221), .B(n15222), .Z(n15215) );
  AND U17147 ( .A(n15223), .B(n15224), .Z(n15221) );
  XOR U17148 ( .A(n15222), .B(n8846), .Z(n15224) );
  XNOR U17149 ( .A(n15225), .B(n15226), .Z(n8846) );
  XNOR U17150 ( .A(n[899]), .B(n15227), .Z(n15223) );
  IV U17151 ( .A(n15222), .Z(n15227) );
  XOR U17152 ( .A(n15228), .B(n15229), .Z(n15222) );
  AND U17153 ( .A(n15230), .B(n15231), .Z(n15228) );
  XOR U17154 ( .A(n15229), .B(n8851), .Z(n15231) );
  XNOR U17155 ( .A(n15232), .B(n15233), .Z(n8851) );
  XNOR U17156 ( .A(n[898]), .B(n15234), .Z(n15230) );
  IV U17157 ( .A(n15229), .Z(n15234) );
  XOR U17158 ( .A(n15235), .B(n15236), .Z(n15229) );
  AND U17159 ( .A(n15237), .B(n15238), .Z(n15235) );
  XOR U17160 ( .A(n15236), .B(n8856), .Z(n15238) );
  XNOR U17161 ( .A(n15239), .B(n15240), .Z(n8856) );
  XNOR U17162 ( .A(n[897]), .B(n15241), .Z(n15237) );
  IV U17163 ( .A(n15236), .Z(n15241) );
  XOR U17164 ( .A(n15242), .B(n15243), .Z(n15236) );
  AND U17165 ( .A(n15244), .B(n15245), .Z(n15242) );
  XOR U17166 ( .A(n15243), .B(n8861), .Z(n15245) );
  XNOR U17167 ( .A(n15246), .B(n15247), .Z(n8861) );
  XNOR U17168 ( .A(n[896]), .B(n15248), .Z(n15244) );
  IV U17169 ( .A(n15243), .Z(n15248) );
  XOR U17170 ( .A(n15249), .B(n15250), .Z(n15243) );
  AND U17171 ( .A(n15251), .B(n15252), .Z(n15249) );
  XOR U17172 ( .A(n15250), .B(n8866), .Z(n15252) );
  XNOR U17173 ( .A(n15253), .B(n15254), .Z(n8866) );
  XNOR U17174 ( .A(n[895]), .B(n15255), .Z(n15251) );
  IV U17175 ( .A(n15250), .Z(n15255) );
  XOR U17176 ( .A(n15256), .B(n15257), .Z(n15250) );
  AND U17177 ( .A(n15258), .B(n15259), .Z(n15256) );
  XOR U17178 ( .A(n15257), .B(n8871), .Z(n15259) );
  XNOR U17179 ( .A(n15260), .B(n15261), .Z(n8871) );
  XNOR U17180 ( .A(n[894]), .B(n15262), .Z(n15258) );
  IV U17181 ( .A(n15257), .Z(n15262) );
  XOR U17182 ( .A(n15263), .B(n15264), .Z(n15257) );
  AND U17183 ( .A(n15265), .B(n15266), .Z(n15263) );
  XOR U17184 ( .A(n15264), .B(n8876), .Z(n15266) );
  XNOR U17185 ( .A(n15267), .B(n15268), .Z(n8876) );
  XNOR U17186 ( .A(n[893]), .B(n15269), .Z(n15265) );
  IV U17187 ( .A(n15264), .Z(n15269) );
  XOR U17188 ( .A(n15270), .B(n15271), .Z(n15264) );
  AND U17189 ( .A(n15272), .B(n15273), .Z(n15270) );
  XOR U17190 ( .A(n15271), .B(n8881), .Z(n15273) );
  XNOR U17191 ( .A(n15274), .B(n15275), .Z(n8881) );
  XNOR U17192 ( .A(n[892]), .B(n15276), .Z(n15272) );
  IV U17193 ( .A(n15271), .Z(n15276) );
  XOR U17194 ( .A(n15277), .B(n15278), .Z(n15271) );
  AND U17195 ( .A(n15279), .B(n15280), .Z(n15277) );
  XOR U17196 ( .A(n15278), .B(n8886), .Z(n15280) );
  XNOR U17197 ( .A(n15281), .B(n15282), .Z(n8886) );
  XNOR U17198 ( .A(n[891]), .B(n15283), .Z(n15279) );
  IV U17199 ( .A(n15278), .Z(n15283) );
  XOR U17200 ( .A(n15284), .B(n15285), .Z(n15278) );
  AND U17201 ( .A(n15286), .B(n15287), .Z(n15284) );
  XOR U17202 ( .A(n15285), .B(n8891), .Z(n15287) );
  XNOR U17203 ( .A(n15288), .B(n15289), .Z(n8891) );
  XNOR U17204 ( .A(n[890]), .B(n15290), .Z(n15286) );
  IV U17205 ( .A(n15285), .Z(n15290) );
  XOR U17206 ( .A(n15291), .B(n15292), .Z(n15285) );
  AND U17207 ( .A(n15293), .B(n15294), .Z(n15291) );
  XOR U17208 ( .A(n15292), .B(n8896), .Z(n15294) );
  XNOR U17209 ( .A(n15295), .B(n15296), .Z(n8896) );
  XNOR U17210 ( .A(n[889]), .B(n15297), .Z(n15293) );
  IV U17211 ( .A(n15292), .Z(n15297) );
  XOR U17212 ( .A(n15298), .B(n15299), .Z(n15292) );
  AND U17213 ( .A(n15300), .B(n15301), .Z(n15298) );
  XOR U17214 ( .A(n15299), .B(n8901), .Z(n15301) );
  XNOR U17215 ( .A(n15302), .B(n15303), .Z(n8901) );
  XNOR U17216 ( .A(n[888]), .B(n15304), .Z(n15300) );
  IV U17217 ( .A(n15299), .Z(n15304) );
  XOR U17218 ( .A(n15305), .B(n15306), .Z(n15299) );
  AND U17219 ( .A(n15307), .B(n15308), .Z(n15305) );
  XOR U17220 ( .A(n15306), .B(n8906), .Z(n15308) );
  XNOR U17221 ( .A(n15309), .B(n15310), .Z(n8906) );
  XNOR U17222 ( .A(n[887]), .B(n15311), .Z(n15307) );
  IV U17223 ( .A(n15306), .Z(n15311) );
  XOR U17224 ( .A(n15312), .B(n15313), .Z(n15306) );
  AND U17225 ( .A(n15314), .B(n15315), .Z(n15312) );
  XOR U17226 ( .A(n15313), .B(n8911), .Z(n15315) );
  XNOR U17227 ( .A(n15316), .B(n15317), .Z(n8911) );
  XNOR U17228 ( .A(n[886]), .B(n15318), .Z(n15314) );
  IV U17229 ( .A(n15313), .Z(n15318) );
  XOR U17230 ( .A(n15319), .B(n15320), .Z(n15313) );
  AND U17231 ( .A(n15321), .B(n15322), .Z(n15319) );
  XOR U17232 ( .A(n15320), .B(n8916), .Z(n15322) );
  XNOR U17233 ( .A(n15323), .B(n15324), .Z(n8916) );
  XNOR U17234 ( .A(n[885]), .B(n15325), .Z(n15321) );
  IV U17235 ( .A(n15320), .Z(n15325) );
  XOR U17236 ( .A(n15326), .B(n15327), .Z(n15320) );
  AND U17237 ( .A(n15328), .B(n15329), .Z(n15326) );
  XOR U17238 ( .A(n15327), .B(n8921), .Z(n15329) );
  XNOR U17239 ( .A(n15330), .B(n15331), .Z(n8921) );
  XNOR U17240 ( .A(n[884]), .B(n15332), .Z(n15328) );
  IV U17241 ( .A(n15327), .Z(n15332) );
  XOR U17242 ( .A(n15333), .B(n15334), .Z(n15327) );
  AND U17243 ( .A(n15335), .B(n15336), .Z(n15333) );
  XOR U17244 ( .A(n15334), .B(n8926), .Z(n15336) );
  XNOR U17245 ( .A(n15337), .B(n15338), .Z(n8926) );
  XNOR U17246 ( .A(n[883]), .B(n15339), .Z(n15335) );
  IV U17247 ( .A(n15334), .Z(n15339) );
  XOR U17248 ( .A(n15340), .B(n15341), .Z(n15334) );
  AND U17249 ( .A(n15342), .B(n15343), .Z(n15340) );
  XOR U17250 ( .A(n15341), .B(n8931), .Z(n15343) );
  XNOR U17251 ( .A(n15344), .B(n15345), .Z(n8931) );
  XNOR U17252 ( .A(n[882]), .B(n15346), .Z(n15342) );
  IV U17253 ( .A(n15341), .Z(n15346) );
  XOR U17254 ( .A(n15347), .B(n15348), .Z(n15341) );
  AND U17255 ( .A(n15349), .B(n15350), .Z(n15347) );
  XOR U17256 ( .A(n15348), .B(n8936), .Z(n15350) );
  XNOR U17257 ( .A(n15351), .B(n15352), .Z(n8936) );
  XNOR U17258 ( .A(n[881]), .B(n15353), .Z(n15349) );
  IV U17259 ( .A(n15348), .Z(n15353) );
  XOR U17260 ( .A(n15354), .B(n15355), .Z(n15348) );
  AND U17261 ( .A(n15356), .B(n15357), .Z(n15354) );
  XOR U17262 ( .A(n15355), .B(n8941), .Z(n15357) );
  XNOR U17263 ( .A(n15358), .B(n15359), .Z(n8941) );
  XNOR U17264 ( .A(n[880]), .B(n15360), .Z(n15356) );
  IV U17265 ( .A(n15355), .Z(n15360) );
  XOR U17266 ( .A(n15361), .B(n15362), .Z(n15355) );
  AND U17267 ( .A(n15363), .B(n15364), .Z(n15361) );
  XOR U17268 ( .A(n15362), .B(n8946), .Z(n15364) );
  XNOR U17269 ( .A(n15365), .B(n15366), .Z(n8946) );
  XNOR U17270 ( .A(n[879]), .B(n15367), .Z(n15363) );
  IV U17271 ( .A(n15362), .Z(n15367) );
  XOR U17272 ( .A(n15368), .B(n15369), .Z(n15362) );
  AND U17273 ( .A(n15370), .B(n15371), .Z(n15368) );
  XOR U17274 ( .A(n15369), .B(n8951), .Z(n15371) );
  XNOR U17275 ( .A(n15372), .B(n15373), .Z(n8951) );
  XNOR U17276 ( .A(n[878]), .B(n15374), .Z(n15370) );
  IV U17277 ( .A(n15369), .Z(n15374) );
  XOR U17278 ( .A(n15375), .B(n15376), .Z(n15369) );
  AND U17279 ( .A(n15377), .B(n15378), .Z(n15375) );
  XOR U17280 ( .A(n15376), .B(n8956), .Z(n15378) );
  XNOR U17281 ( .A(n15379), .B(n15380), .Z(n8956) );
  XNOR U17282 ( .A(n[877]), .B(n15381), .Z(n15377) );
  IV U17283 ( .A(n15376), .Z(n15381) );
  XOR U17284 ( .A(n15382), .B(n15383), .Z(n15376) );
  AND U17285 ( .A(n15384), .B(n15385), .Z(n15382) );
  XOR U17286 ( .A(n15383), .B(n8961), .Z(n15385) );
  XNOR U17287 ( .A(n15386), .B(n15387), .Z(n8961) );
  XNOR U17288 ( .A(n[876]), .B(n15388), .Z(n15384) );
  IV U17289 ( .A(n15383), .Z(n15388) );
  XOR U17290 ( .A(n15389), .B(n15390), .Z(n15383) );
  AND U17291 ( .A(n15391), .B(n15392), .Z(n15389) );
  XOR U17292 ( .A(n15390), .B(n8966), .Z(n15392) );
  XNOR U17293 ( .A(n15393), .B(n15394), .Z(n8966) );
  XNOR U17294 ( .A(n[875]), .B(n15395), .Z(n15391) );
  IV U17295 ( .A(n15390), .Z(n15395) );
  XOR U17296 ( .A(n15396), .B(n15397), .Z(n15390) );
  AND U17297 ( .A(n15398), .B(n15399), .Z(n15396) );
  XOR U17298 ( .A(n15397), .B(n8971), .Z(n15399) );
  XNOR U17299 ( .A(n15400), .B(n15401), .Z(n8971) );
  XNOR U17300 ( .A(n[874]), .B(n15402), .Z(n15398) );
  IV U17301 ( .A(n15397), .Z(n15402) );
  XOR U17302 ( .A(n15403), .B(n15404), .Z(n15397) );
  AND U17303 ( .A(n15405), .B(n15406), .Z(n15403) );
  XOR U17304 ( .A(n15404), .B(n8976), .Z(n15406) );
  XNOR U17305 ( .A(n15407), .B(n15408), .Z(n8976) );
  XNOR U17306 ( .A(n[873]), .B(n15409), .Z(n15405) );
  IV U17307 ( .A(n15404), .Z(n15409) );
  XOR U17308 ( .A(n15410), .B(n15411), .Z(n15404) );
  AND U17309 ( .A(n15412), .B(n15413), .Z(n15410) );
  XOR U17310 ( .A(n15411), .B(n8981), .Z(n15413) );
  XNOR U17311 ( .A(n15414), .B(n15415), .Z(n8981) );
  XNOR U17312 ( .A(n[872]), .B(n15416), .Z(n15412) );
  IV U17313 ( .A(n15411), .Z(n15416) );
  XOR U17314 ( .A(n15417), .B(n15418), .Z(n15411) );
  AND U17315 ( .A(n15419), .B(n15420), .Z(n15417) );
  XOR U17316 ( .A(n15418), .B(n8986), .Z(n15420) );
  XNOR U17317 ( .A(n15421), .B(n15422), .Z(n8986) );
  XNOR U17318 ( .A(n[871]), .B(n15423), .Z(n15419) );
  IV U17319 ( .A(n15418), .Z(n15423) );
  XOR U17320 ( .A(n15424), .B(n15425), .Z(n15418) );
  AND U17321 ( .A(n15426), .B(n15427), .Z(n15424) );
  XOR U17322 ( .A(n15425), .B(n8991), .Z(n15427) );
  XNOR U17323 ( .A(n15428), .B(n15429), .Z(n8991) );
  XNOR U17324 ( .A(n[870]), .B(n15430), .Z(n15426) );
  IV U17325 ( .A(n15425), .Z(n15430) );
  XOR U17326 ( .A(n15431), .B(n15432), .Z(n15425) );
  AND U17327 ( .A(n15433), .B(n15434), .Z(n15431) );
  XOR U17328 ( .A(n15432), .B(n8996), .Z(n15434) );
  XNOR U17329 ( .A(n15435), .B(n15436), .Z(n8996) );
  XNOR U17330 ( .A(n[869]), .B(n15437), .Z(n15433) );
  IV U17331 ( .A(n15432), .Z(n15437) );
  XOR U17332 ( .A(n15438), .B(n15439), .Z(n15432) );
  AND U17333 ( .A(n15440), .B(n15441), .Z(n15438) );
  XOR U17334 ( .A(n15439), .B(n9001), .Z(n15441) );
  XNOR U17335 ( .A(n15442), .B(n15443), .Z(n9001) );
  XNOR U17336 ( .A(n[868]), .B(n15444), .Z(n15440) );
  IV U17337 ( .A(n15439), .Z(n15444) );
  XOR U17338 ( .A(n15445), .B(n15446), .Z(n15439) );
  AND U17339 ( .A(n15447), .B(n15448), .Z(n15445) );
  XOR U17340 ( .A(n15446), .B(n9006), .Z(n15448) );
  XNOR U17341 ( .A(n15449), .B(n15450), .Z(n9006) );
  XNOR U17342 ( .A(n[867]), .B(n15451), .Z(n15447) );
  IV U17343 ( .A(n15446), .Z(n15451) );
  XOR U17344 ( .A(n15452), .B(n15453), .Z(n15446) );
  AND U17345 ( .A(n15454), .B(n15455), .Z(n15452) );
  XOR U17346 ( .A(n15453), .B(n9011), .Z(n15455) );
  XNOR U17347 ( .A(n15456), .B(n15457), .Z(n9011) );
  XNOR U17348 ( .A(n[866]), .B(n15458), .Z(n15454) );
  IV U17349 ( .A(n15453), .Z(n15458) );
  XOR U17350 ( .A(n15459), .B(n15460), .Z(n15453) );
  AND U17351 ( .A(n15461), .B(n15462), .Z(n15459) );
  XOR U17352 ( .A(n15460), .B(n9016), .Z(n15462) );
  XNOR U17353 ( .A(n15463), .B(n15464), .Z(n9016) );
  XNOR U17354 ( .A(n[865]), .B(n15465), .Z(n15461) );
  IV U17355 ( .A(n15460), .Z(n15465) );
  XOR U17356 ( .A(n15466), .B(n15467), .Z(n15460) );
  AND U17357 ( .A(n15468), .B(n15469), .Z(n15466) );
  XOR U17358 ( .A(n15467), .B(n9021), .Z(n15469) );
  XNOR U17359 ( .A(n15470), .B(n15471), .Z(n9021) );
  XNOR U17360 ( .A(n[864]), .B(n15472), .Z(n15468) );
  IV U17361 ( .A(n15467), .Z(n15472) );
  XOR U17362 ( .A(n15473), .B(n15474), .Z(n15467) );
  AND U17363 ( .A(n15475), .B(n15476), .Z(n15473) );
  XOR U17364 ( .A(n15474), .B(n9026), .Z(n15476) );
  XNOR U17365 ( .A(n15477), .B(n15478), .Z(n9026) );
  XNOR U17366 ( .A(n[863]), .B(n15479), .Z(n15475) );
  IV U17367 ( .A(n15474), .Z(n15479) );
  XOR U17368 ( .A(n15480), .B(n15481), .Z(n15474) );
  AND U17369 ( .A(n15482), .B(n15483), .Z(n15480) );
  XOR U17370 ( .A(n15481), .B(n9031), .Z(n15483) );
  XNOR U17371 ( .A(n15484), .B(n15485), .Z(n9031) );
  XNOR U17372 ( .A(n[862]), .B(n15486), .Z(n15482) );
  IV U17373 ( .A(n15481), .Z(n15486) );
  XOR U17374 ( .A(n15487), .B(n15488), .Z(n15481) );
  AND U17375 ( .A(n15489), .B(n15490), .Z(n15487) );
  XOR U17376 ( .A(n15488), .B(n9036), .Z(n15490) );
  XNOR U17377 ( .A(n15491), .B(n15492), .Z(n9036) );
  XNOR U17378 ( .A(n[861]), .B(n15493), .Z(n15489) );
  IV U17379 ( .A(n15488), .Z(n15493) );
  XOR U17380 ( .A(n15494), .B(n15495), .Z(n15488) );
  AND U17381 ( .A(n15496), .B(n15497), .Z(n15494) );
  XOR U17382 ( .A(n15495), .B(n9041), .Z(n15497) );
  XNOR U17383 ( .A(n15498), .B(n15499), .Z(n9041) );
  XNOR U17384 ( .A(n[860]), .B(n15500), .Z(n15496) );
  IV U17385 ( .A(n15495), .Z(n15500) );
  XOR U17386 ( .A(n15501), .B(n15502), .Z(n15495) );
  AND U17387 ( .A(n15503), .B(n15504), .Z(n15501) );
  XOR U17388 ( .A(n15502), .B(n9046), .Z(n15504) );
  XNOR U17389 ( .A(n15505), .B(n15506), .Z(n9046) );
  XNOR U17390 ( .A(n[859]), .B(n15507), .Z(n15503) );
  IV U17391 ( .A(n15502), .Z(n15507) );
  XOR U17392 ( .A(n15508), .B(n15509), .Z(n15502) );
  AND U17393 ( .A(n15510), .B(n15511), .Z(n15508) );
  XOR U17394 ( .A(n15509), .B(n9051), .Z(n15511) );
  XNOR U17395 ( .A(n15512), .B(n15513), .Z(n9051) );
  XNOR U17396 ( .A(n[858]), .B(n15514), .Z(n15510) );
  IV U17397 ( .A(n15509), .Z(n15514) );
  XOR U17398 ( .A(n15515), .B(n15516), .Z(n15509) );
  AND U17399 ( .A(n15517), .B(n15518), .Z(n15515) );
  XOR U17400 ( .A(n15516), .B(n9056), .Z(n15518) );
  XNOR U17401 ( .A(n15519), .B(n15520), .Z(n9056) );
  XNOR U17402 ( .A(n[857]), .B(n15521), .Z(n15517) );
  IV U17403 ( .A(n15516), .Z(n15521) );
  XOR U17404 ( .A(n15522), .B(n15523), .Z(n15516) );
  AND U17405 ( .A(n15524), .B(n15525), .Z(n15522) );
  XOR U17406 ( .A(n15523), .B(n9061), .Z(n15525) );
  XNOR U17407 ( .A(n15526), .B(n15527), .Z(n9061) );
  XNOR U17408 ( .A(n[856]), .B(n15528), .Z(n15524) );
  IV U17409 ( .A(n15523), .Z(n15528) );
  XOR U17410 ( .A(n15529), .B(n15530), .Z(n15523) );
  AND U17411 ( .A(n15531), .B(n15532), .Z(n15529) );
  XOR U17412 ( .A(n15530), .B(n9066), .Z(n15532) );
  XNOR U17413 ( .A(n15533), .B(n15534), .Z(n9066) );
  XNOR U17414 ( .A(n[855]), .B(n15535), .Z(n15531) );
  IV U17415 ( .A(n15530), .Z(n15535) );
  XOR U17416 ( .A(n15536), .B(n15537), .Z(n15530) );
  AND U17417 ( .A(n15538), .B(n15539), .Z(n15536) );
  XOR U17418 ( .A(n15537), .B(n9071), .Z(n15539) );
  XNOR U17419 ( .A(n15540), .B(n15541), .Z(n9071) );
  XNOR U17420 ( .A(n[854]), .B(n15542), .Z(n15538) );
  IV U17421 ( .A(n15537), .Z(n15542) );
  XOR U17422 ( .A(n15543), .B(n15544), .Z(n15537) );
  AND U17423 ( .A(n15545), .B(n15546), .Z(n15543) );
  XOR U17424 ( .A(n15544), .B(n9076), .Z(n15546) );
  XNOR U17425 ( .A(n15547), .B(n15548), .Z(n9076) );
  XNOR U17426 ( .A(n[853]), .B(n15549), .Z(n15545) );
  IV U17427 ( .A(n15544), .Z(n15549) );
  XOR U17428 ( .A(n15550), .B(n15551), .Z(n15544) );
  AND U17429 ( .A(n15552), .B(n15553), .Z(n15550) );
  XOR U17430 ( .A(n15551), .B(n9081), .Z(n15553) );
  XNOR U17431 ( .A(n15554), .B(n15555), .Z(n9081) );
  XNOR U17432 ( .A(n[852]), .B(n15556), .Z(n15552) );
  IV U17433 ( .A(n15551), .Z(n15556) );
  XOR U17434 ( .A(n15557), .B(n15558), .Z(n15551) );
  AND U17435 ( .A(n15559), .B(n15560), .Z(n15557) );
  XOR U17436 ( .A(n15558), .B(n9086), .Z(n15560) );
  XNOR U17437 ( .A(n15561), .B(n15562), .Z(n9086) );
  XNOR U17438 ( .A(n[851]), .B(n15563), .Z(n15559) );
  IV U17439 ( .A(n15558), .Z(n15563) );
  XOR U17440 ( .A(n15564), .B(n15565), .Z(n15558) );
  AND U17441 ( .A(n15566), .B(n15567), .Z(n15564) );
  XOR U17442 ( .A(n15565), .B(n9091), .Z(n15567) );
  XNOR U17443 ( .A(n15568), .B(n15569), .Z(n9091) );
  XNOR U17444 ( .A(n[850]), .B(n15570), .Z(n15566) );
  IV U17445 ( .A(n15565), .Z(n15570) );
  XOR U17446 ( .A(n15571), .B(n15572), .Z(n15565) );
  AND U17447 ( .A(n15573), .B(n15574), .Z(n15571) );
  XOR U17448 ( .A(n15572), .B(n9096), .Z(n15574) );
  XNOR U17449 ( .A(n15575), .B(n15576), .Z(n9096) );
  XNOR U17450 ( .A(n[849]), .B(n15577), .Z(n15573) );
  IV U17451 ( .A(n15572), .Z(n15577) );
  XOR U17452 ( .A(n15578), .B(n15579), .Z(n15572) );
  AND U17453 ( .A(n15580), .B(n15581), .Z(n15578) );
  XOR U17454 ( .A(n15579), .B(n9101), .Z(n15581) );
  XNOR U17455 ( .A(n15582), .B(n15583), .Z(n9101) );
  XNOR U17456 ( .A(n[848]), .B(n15584), .Z(n15580) );
  IV U17457 ( .A(n15579), .Z(n15584) );
  XOR U17458 ( .A(n15585), .B(n15586), .Z(n15579) );
  AND U17459 ( .A(n15587), .B(n15588), .Z(n15585) );
  XOR U17460 ( .A(n15586), .B(n9106), .Z(n15588) );
  XNOR U17461 ( .A(n15589), .B(n15590), .Z(n9106) );
  XNOR U17462 ( .A(n[847]), .B(n15591), .Z(n15587) );
  IV U17463 ( .A(n15586), .Z(n15591) );
  XOR U17464 ( .A(n15592), .B(n15593), .Z(n15586) );
  AND U17465 ( .A(n15594), .B(n15595), .Z(n15592) );
  XOR U17466 ( .A(n15593), .B(n9111), .Z(n15595) );
  XNOR U17467 ( .A(n15596), .B(n15597), .Z(n9111) );
  XNOR U17468 ( .A(n[846]), .B(n15598), .Z(n15594) );
  IV U17469 ( .A(n15593), .Z(n15598) );
  XOR U17470 ( .A(n15599), .B(n15600), .Z(n15593) );
  AND U17471 ( .A(n15601), .B(n15602), .Z(n15599) );
  XOR U17472 ( .A(n15600), .B(n9116), .Z(n15602) );
  XNOR U17473 ( .A(n15603), .B(n15604), .Z(n9116) );
  XNOR U17474 ( .A(n[845]), .B(n15605), .Z(n15601) );
  IV U17475 ( .A(n15600), .Z(n15605) );
  XOR U17476 ( .A(n15606), .B(n15607), .Z(n15600) );
  AND U17477 ( .A(n15608), .B(n15609), .Z(n15606) );
  XOR U17478 ( .A(n15607), .B(n9121), .Z(n15609) );
  XNOR U17479 ( .A(n15610), .B(n15611), .Z(n9121) );
  XNOR U17480 ( .A(n[844]), .B(n15612), .Z(n15608) );
  IV U17481 ( .A(n15607), .Z(n15612) );
  XOR U17482 ( .A(n15613), .B(n15614), .Z(n15607) );
  AND U17483 ( .A(n15615), .B(n15616), .Z(n15613) );
  XOR U17484 ( .A(n15614), .B(n9126), .Z(n15616) );
  XNOR U17485 ( .A(n15617), .B(n15618), .Z(n9126) );
  XNOR U17486 ( .A(n[843]), .B(n15619), .Z(n15615) );
  IV U17487 ( .A(n15614), .Z(n15619) );
  XOR U17488 ( .A(n15620), .B(n15621), .Z(n15614) );
  AND U17489 ( .A(n15622), .B(n15623), .Z(n15620) );
  XOR U17490 ( .A(n15621), .B(n9131), .Z(n15623) );
  XNOR U17491 ( .A(n15624), .B(n15625), .Z(n9131) );
  XNOR U17492 ( .A(n[842]), .B(n15626), .Z(n15622) );
  IV U17493 ( .A(n15621), .Z(n15626) );
  XOR U17494 ( .A(n15627), .B(n15628), .Z(n15621) );
  AND U17495 ( .A(n15629), .B(n15630), .Z(n15627) );
  XOR U17496 ( .A(n15628), .B(n9136), .Z(n15630) );
  XNOR U17497 ( .A(n15631), .B(n15632), .Z(n9136) );
  XNOR U17498 ( .A(n[841]), .B(n15633), .Z(n15629) );
  IV U17499 ( .A(n15628), .Z(n15633) );
  XOR U17500 ( .A(n15634), .B(n15635), .Z(n15628) );
  AND U17501 ( .A(n15636), .B(n15637), .Z(n15634) );
  XOR U17502 ( .A(n15635), .B(n9141), .Z(n15637) );
  XNOR U17503 ( .A(n15638), .B(n15639), .Z(n9141) );
  XNOR U17504 ( .A(n[840]), .B(n15640), .Z(n15636) );
  IV U17505 ( .A(n15635), .Z(n15640) );
  XOR U17506 ( .A(n15641), .B(n15642), .Z(n15635) );
  AND U17507 ( .A(n15643), .B(n15644), .Z(n15641) );
  XOR U17508 ( .A(n15642), .B(n9146), .Z(n15644) );
  XNOR U17509 ( .A(n15645), .B(n15646), .Z(n9146) );
  XNOR U17510 ( .A(n[839]), .B(n15647), .Z(n15643) );
  IV U17511 ( .A(n15642), .Z(n15647) );
  XOR U17512 ( .A(n15648), .B(n15649), .Z(n15642) );
  AND U17513 ( .A(n15650), .B(n15651), .Z(n15648) );
  XOR U17514 ( .A(n15649), .B(n9151), .Z(n15651) );
  XNOR U17515 ( .A(n15652), .B(n15653), .Z(n9151) );
  XNOR U17516 ( .A(n[838]), .B(n15654), .Z(n15650) );
  IV U17517 ( .A(n15649), .Z(n15654) );
  XOR U17518 ( .A(n15655), .B(n15656), .Z(n15649) );
  AND U17519 ( .A(n15657), .B(n15658), .Z(n15655) );
  XOR U17520 ( .A(n15656), .B(n9156), .Z(n15658) );
  XNOR U17521 ( .A(n15659), .B(n15660), .Z(n9156) );
  XNOR U17522 ( .A(n[837]), .B(n15661), .Z(n15657) );
  IV U17523 ( .A(n15656), .Z(n15661) );
  XOR U17524 ( .A(n15662), .B(n15663), .Z(n15656) );
  AND U17525 ( .A(n15664), .B(n15665), .Z(n15662) );
  XOR U17526 ( .A(n15663), .B(n9161), .Z(n15665) );
  XNOR U17527 ( .A(n15666), .B(n15667), .Z(n9161) );
  XNOR U17528 ( .A(n[836]), .B(n15668), .Z(n15664) );
  IV U17529 ( .A(n15663), .Z(n15668) );
  XOR U17530 ( .A(n15669), .B(n15670), .Z(n15663) );
  AND U17531 ( .A(n15671), .B(n15672), .Z(n15669) );
  XOR U17532 ( .A(n15670), .B(n9166), .Z(n15672) );
  XNOR U17533 ( .A(n15673), .B(n15674), .Z(n9166) );
  XNOR U17534 ( .A(n[835]), .B(n15675), .Z(n15671) );
  IV U17535 ( .A(n15670), .Z(n15675) );
  XOR U17536 ( .A(n15676), .B(n15677), .Z(n15670) );
  AND U17537 ( .A(n15678), .B(n15679), .Z(n15676) );
  XOR U17538 ( .A(n15677), .B(n9171), .Z(n15679) );
  XNOR U17539 ( .A(n15680), .B(n15681), .Z(n9171) );
  XNOR U17540 ( .A(n[834]), .B(n15682), .Z(n15678) );
  IV U17541 ( .A(n15677), .Z(n15682) );
  XOR U17542 ( .A(n15683), .B(n15684), .Z(n15677) );
  AND U17543 ( .A(n15685), .B(n15686), .Z(n15683) );
  XOR U17544 ( .A(n15684), .B(n9176), .Z(n15686) );
  XNOR U17545 ( .A(n15687), .B(n15688), .Z(n9176) );
  XNOR U17546 ( .A(n[833]), .B(n15689), .Z(n15685) );
  IV U17547 ( .A(n15684), .Z(n15689) );
  XOR U17548 ( .A(n15690), .B(n15691), .Z(n15684) );
  AND U17549 ( .A(n15692), .B(n15693), .Z(n15690) );
  XOR U17550 ( .A(n15691), .B(n9181), .Z(n15693) );
  XNOR U17551 ( .A(n15694), .B(n15695), .Z(n9181) );
  XNOR U17552 ( .A(n[832]), .B(n15696), .Z(n15692) );
  IV U17553 ( .A(n15691), .Z(n15696) );
  XOR U17554 ( .A(n15697), .B(n15698), .Z(n15691) );
  AND U17555 ( .A(n15699), .B(n15700), .Z(n15697) );
  XOR U17556 ( .A(n15698), .B(n9186), .Z(n15700) );
  XNOR U17557 ( .A(n15701), .B(n15702), .Z(n9186) );
  XNOR U17558 ( .A(n[831]), .B(n15703), .Z(n15699) );
  IV U17559 ( .A(n15698), .Z(n15703) );
  XOR U17560 ( .A(n15704), .B(n15705), .Z(n15698) );
  AND U17561 ( .A(n15706), .B(n15707), .Z(n15704) );
  XOR U17562 ( .A(n15705), .B(n9191), .Z(n15707) );
  XNOR U17563 ( .A(n15708), .B(n15709), .Z(n9191) );
  XNOR U17564 ( .A(n[830]), .B(n15710), .Z(n15706) );
  IV U17565 ( .A(n15705), .Z(n15710) );
  XOR U17566 ( .A(n15711), .B(n15712), .Z(n15705) );
  AND U17567 ( .A(n15713), .B(n15714), .Z(n15711) );
  XOR U17568 ( .A(n15712), .B(n9196), .Z(n15714) );
  XNOR U17569 ( .A(n15715), .B(n15716), .Z(n9196) );
  XNOR U17570 ( .A(n[829]), .B(n15717), .Z(n15713) );
  IV U17571 ( .A(n15712), .Z(n15717) );
  XOR U17572 ( .A(n15718), .B(n15719), .Z(n15712) );
  AND U17573 ( .A(n15720), .B(n15721), .Z(n15718) );
  XOR U17574 ( .A(n15719), .B(n9201), .Z(n15721) );
  XNOR U17575 ( .A(n15722), .B(n15723), .Z(n9201) );
  XNOR U17576 ( .A(n[828]), .B(n15724), .Z(n15720) );
  IV U17577 ( .A(n15719), .Z(n15724) );
  XOR U17578 ( .A(n15725), .B(n15726), .Z(n15719) );
  AND U17579 ( .A(n15727), .B(n15728), .Z(n15725) );
  XOR U17580 ( .A(n15726), .B(n9206), .Z(n15728) );
  XNOR U17581 ( .A(n15729), .B(n15730), .Z(n9206) );
  XNOR U17582 ( .A(n[827]), .B(n15731), .Z(n15727) );
  IV U17583 ( .A(n15726), .Z(n15731) );
  XOR U17584 ( .A(n15732), .B(n15733), .Z(n15726) );
  AND U17585 ( .A(n15734), .B(n15735), .Z(n15732) );
  XOR U17586 ( .A(n15733), .B(n9211), .Z(n15735) );
  XNOR U17587 ( .A(n15736), .B(n15737), .Z(n9211) );
  XNOR U17588 ( .A(n[826]), .B(n15738), .Z(n15734) );
  IV U17589 ( .A(n15733), .Z(n15738) );
  XOR U17590 ( .A(n15739), .B(n15740), .Z(n15733) );
  AND U17591 ( .A(n15741), .B(n15742), .Z(n15739) );
  XOR U17592 ( .A(n15740), .B(n9216), .Z(n15742) );
  XNOR U17593 ( .A(n15743), .B(n15744), .Z(n9216) );
  XNOR U17594 ( .A(n[825]), .B(n15745), .Z(n15741) );
  IV U17595 ( .A(n15740), .Z(n15745) );
  XOR U17596 ( .A(n15746), .B(n15747), .Z(n15740) );
  AND U17597 ( .A(n15748), .B(n15749), .Z(n15746) );
  XOR U17598 ( .A(n15747), .B(n9221), .Z(n15749) );
  XNOR U17599 ( .A(n15750), .B(n15751), .Z(n9221) );
  XNOR U17600 ( .A(n[824]), .B(n15752), .Z(n15748) );
  IV U17601 ( .A(n15747), .Z(n15752) );
  XOR U17602 ( .A(n15753), .B(n15754), .Z(n15747) );
  AND U17603 ( .A(n15755), .B(n15756), .Z(n15753) );
  XOR U17604 ( .A(n15754), .B(n9226), .Z(n15756) );
  XNOR U17605 ( .A(n15757), .B(n15758), .Z(n9226) );
  XNOR U17606 ( .A(n[823]), .B(n15759), .Z(n15755) );
  IV U17607 ( .A(n15754), .Z(n15759) );
  XOR U17608 ( .A(n15760), .B(n15761), .Z(n15754) );
  AND U17609 ( .A(n15762), .B(n15763), .Z(n15760) );
  XOR U17610 ( .A(n15761), .B(n9231), .Z(n15763) );
  XNOR U17611 ( .A(n15764), .B(n15765), .Z(n9231) );
  XNOR U17612 ( .A(n[822]), .B(n15766), .Z(n15762) );
  IV U17613 ( .A(n15761), .Z(n15766) );
  XOR U17614 ( .A(n15767), .B(n15768), .Z(n15761) );
  AND U17615 ( .A(n15769), .B(n15770), .Z(n15767) );
  XOR U17616 ( .A(n15768), .B(n9236), .Z(n15770) );
  XNOR U17617 ( .A(n15771), .B(n15772), .Z(n9236) );
  XNOR U17618 ( .A(n[821]), .B(n15773), .Z(n15769) );
  IV U17619 ( .A(n15768), .Z(n15773) );
  XOR U17620 ( .A(n15774), .B(n15775), .Z(n15768) );
  AND U17621 ( .A(n15776), .B(n15777), .Z(n15774) );
  XOR U17622 ( .A(n15775), .B(n9241), .Z(n15777) );
  XNOR U17623 ( .A(n15778), .B(n15779), .Z(n9241) );
  XNOR U17624 ( .A(n[820]), .B(n15780), .Z(n15776) );
  IV U17625 ( .A(n15775), .Z(n15780) );
  XOR U17626 ( .A(n15781), .B(n15782), .Z(n15775) );
  AND U17627 ( .A(n15783), .B(n15784), .Z(n15781) );
  XOR U17628 ( .A(n15782), .B(n9246), .Z(n15784) );
  XNOR U17629 ( .A(n15785), .B(n15786), .Z(n9246) );
  XNOR U17630 ( .A(n[819]), .B(n15787), .Z(n15783) );
  IV U17631 ( .A(n15782), .Z(n15787) );
  XOR U17632 ( .A(n15788), .B(n15789), .Z(n15782) );
  AND U17633 ( .A(n15790), .B(n15791), .Z(n15788) );
  XOR U17634 ( .A(n15789), .B(n9251), .Z(n15791) );
  XNOR U17635 ( .A(n15792), .B(n15793), .Z(n9251) );
  XNOR U17636 ( .A(n[818]), .B(n15794), .Z(n15790) );
  IV U17637 ( .A(n15789), .Z(n15794) );
  XOR U17638 ( .A(n15795), .B(n15796), .Z(n15789) );
  AND U17639 ( .A(n15797), .B(n15798), .Z(n15795) );
  XOR U17640 ( .A(n15796), .B(n9256), .Z(n15798) );
  XNOR U17641 ( .A(n15799), .B(n15800), .Z(n9256) );
  XNOR U17642 ( .A(n[817]), .B(n15801), .Z(n15797) );
  IV U17643 ( .A(n15796), .Z(n15801) );
  XOR U17644 ( .A(n15802), .B(n15803), .Z(n15796) );
  AND U17645 ( .A(n15804), .B(n15805), .Z(n15802) );
  XOR U17646 ( .A(n15803), .B(n9261), .Z(n15805) );
  XNOR U17647 ( .A(n15806), .B(n15807), .Z(n9261) );
  XNOR U17648 ( .A(n[816]), .B(n15808), .Z(n15804) );
  IV U17649 ( .A(n15803), .Z(n15808) );
  XOR U17650 ( .A(n15809), .B(n15810), .Z(n15803) );
  AND U17651 ( .A(n15811), .B(n15812), .Z(n15809) );
  XOR U17652 ( .A(n15810), .B(n9266), .Z(n15812) );
  XNOR U17653 ( .A(n15813), .B(n15814), .Z(n9266) );
  XNOR U17654 ( .A(n[815]), .B(n15815), .Z(n15811) );
  IV U17655 ( .A(n15810), .Z(n15815) );
  XOR U17656 ( .A(n15816), .B(n15817), .Z(n15810) );
  AND U17657 ( .A(n15818), .B(n15819), .Z(n15816) );
  XOR U17658 ( .A(n15817), .B(n9271), .Z(n15819) );
  XNOR U17659 ( .A(n15820), .B(n15821), .Z(n9271) );
  XNOR U17660 ( .A(n[814]), .B(n15822), .Z(n15818) );
  IV U17661 ( .A(n15817), .Z(n15822) );
  XOR U17662 ( .A(n15823), .B(n15824), .Z(n15817) );
  AND U17663 ( .A(n15825), .B(n15826), .Z(n15823) );
  XOR U17664 ( .A(n15824), .B(n9276), .Z(n15826) );
  XNOR U17665 ( .A(n15827), .B(n15828), .Z(n9276) );
  XNOR U17666 ( .A(n[813]), .B(n15829), .Z(n15825) );
  IV U17667 ( .A(n15824), .Z(n15829) );
  XOR U17668 ( .A(n15830), .B(n15831), .Z(n15824) );
  AND U17669 ( .A(n15832), .B(n15833), .Z(n15830) );
  XOR U17670 ( .A(n15831), .B(n9281), .Z(n15833) );
  XNOR U17671 ( .A(n15834), .B(n15835), .Z(n9281) );
  XNOR U17672 ( .A(n[812]), .B(n15836), .Z(n15832) );
  IV U17673 ( .A(n15831), .Z(n15836) );
  XOR U17674 ( .A(n15837), .B(n15838), .Z(n15831) );
  AND U17675 ( .A(n15839), .B(n15840), .Z(n15837) );
  XOR U17676 ( .A(n15838), .B(n9286), .Z(n15840) );
  XNOR U17677 ( .A(n15841), .B(n15842), .Z(n9286) );
  XNOR U17678 ( .A(n[811]), .B(n15843), .Z(n15839) );
  IV U17679 ( .A(n15838), .Z(n15843) );
  XOR U17680 ( .A(n15844), .B(n15845), .Z(n15838) );
  AND U17681 ( .A(n15846), .B(n15847), .Z(n15844) );
  XOR U17682 ( .A(n15845), .B(n9291), .Z(n15847) );
  XNOR U17683 ( .A(n15848), .B(n15849), .Z(n9291) );
  XNOR U17684 ( .A(n[810]), .B(n15850), .Z(n15846) );
  IV U17685 ( .A(n15845), .Z(n15850) );
  XOR U17686 ( .A(n15851), .B(n15852), .Z(n15845) );
  AND U17687 ( .A(n15853), .B(n15854), .Z(n15851) );
  XOR U17688 ( .A(n15852), .B(n9296), .Z(n15854) );
  XNOR U17689 ( .A(n15855), .B(n15856), .Z(n9296) );
  XNOR U17690 ( .A(n[809]), .B(n15857), .Z(n15853) );
  IV U17691 ( .A(n15852), .Z(n15857) );
  XOR U17692 ( .A(n15858), .B(n15859), .Z(n15852) );
  AND U17693 ( .A(n15860), .B(n15861), .Z(n15858) );
  XOR U17694 ( .A(n15859), .B(n9301), .Z(n15861) );
  XNOR U17695 ( .A(n15862), .B(n15863), .Z(n9301) );
  XNOR U17696 ( .A(n[808]), .B(n15864), .Z(n15860) );
  IV U17697 ( .A(n15859), .Z(n15864) );
  XOR U17698 ( .A(n15865), .B(n15866), .Z(n15859) );
  AND U17699 ( .A(n15867), .B(n15868), .Z(n15865) );
  XOR U17700 ( .A(n15866), .B(n9306), .Z(n15868) );
  XNOR U17701 ( .A(n15869), .B(n15870), .Z(n9306) );
  XNOR U17702 ( .A(n[807]), .B(n15871), .Z(n15867) );
  IV U17703 ( .A(n15866), .Z(n15871) );
  XOR U17704 ( .A(n15872), .B(n15873), .Z(n15866) );
  AND U17705 ( .A(n15874), .B(n15875), .Z(n15872) );
  XOR U17706 ( .A(n15873), .B(n9311), .Z(n15875) );
  XNOR U17707 ( .A(n15876), .B(n15877), .Z(n9311) );
  XNOR U17708 ( .A(n[806]), .B(n15878), .Z(n15874) );
  IV U17709 ( .A(n15873), .Z(n15878) );
  XOR U17710 ( .A(n15879), .B(n15880), .Z(n15873) );
  AND U17711 ( .A(n15881), .B(n15882), .Z(n15879) );
  XOR U17712 ( .A(n15880), .B(n9316), .Z(n15882) );
  XNOR U17713 ( .A(n15883), .B(n15884), .Z(n9316) );
  XNOR U17714 ( .A(n[805]), .B(n15885), .Z(n15881) );
  IV U17715 ( .A(n15880), .Z(n15885) );
  XOR U17716 ( .A(n15886), .B(n15887), .Z(n15880) );
  AND U17717 ( .A(n15888), .B(n15889), .Z(n15886) );
  XOR U17718 ( .A(n15887), .B(n9321), .Z(n15889) );
  XNOR U17719 ( .A(n15890), .B(n15891), .Z(n9321) );
  XNOR U17720 ( .A(n[804]), .B(n15892), .Z(n15888) );
  IV U17721 ( .A(n15887), .Z(n15892) );
  XOR U17722 ( .A(n15893), .B(n15894), .Z(n15887) );
  AND U17723 ( .A(n15895), .B(n15896), .Z(n15893) );
  XOR U17724 ( .A(n15894), .B(n9326), .Z(n15896) );
  XNOR U17725 ( .A(n15897), .B(n15898), .Z(n9326) );
  XNOR U17726 ( .A(n[803]), .B(n15899), .Z(n15895) );
  IV U17727 ( .A(n15894), .Z(n15899) );
  XOR U17728 ( .A(n15900), .B(n15901), .Z(n15894) );
  AND U17729 ( .A(n15902), .B(n15903), .Z(n15900) );
  XOR U17730 ( .A(n15901), .B(n9331), .Z(n15903) );
  XNOR U17731 ( .A(n15904), .B(n15905), .Z(n9331) );
  XNOR U17732 ( .A(n[802]), .B(n15906), .Z(n15902) );
  IV U17733 ( .A(n15901), .Z(n15906) );
  XOR U17734 ( .A(n15907), .B(n15908), .Z(n15901) );
  AND U17735 ( .A(n15909), .B(n15910), .Z(n15907) );
  XOR U17736 ( .A(n15908), .B(n9336), .Z(n15910) );
  XNOR U17737 ( .A(n15911), .B(n15912), .Z(n9336) );
  XNOR U17738 ( .A(n[801]), .B(n15913), .Z(n15909) );
  IV U17739 ( .A(n15908), .Z(n15913) );
  XOR U17740 ( .A(n15914), .B(n15915), .Z(n15908) );
  AND U17741 ( .A(n15916), .B(n15917), .Z(n15914) );
  XOR U17742 ( .A(n15915), .B(n9341), .Z(n15917) );
  XNOR U17743 ( .A(n15918), .B(n15919), .Z(n9341) );
  XNOR U17744 ( .A(n[800]), .B(n15920), .Z(n15916) );
  IV U17745 ( .A(n15915), .Z(n15920) );
  XOR U17746 ( .A(n15921), .B(n15922), .Z(n15915) );
  AND U17747 ( .A(n15923), .B(n15924), .Z(n15921) );
  XOR U17748 ( .A(n15922), .B(n9346), .Z(n15924) );
  XNOR U17749 ( .A(n15925), .B(n15926), .Z(n9346) );
  XNOR U17750 ( .A(n[799]), .B(n15927), .Z(n15923) );
  IV U17751 ( .A(n15922), .Z(n15927) );
  XOR U17752 ( .A(n15928), .B(n15929), .Z(n15922) );
  AND U17753 ( .A(n15930), .B(n15931), .Z(n15928) );
  XOR U17754 ( .A(n15929), .B(n9351), .Z(n15931) );
  XNOR U17755 ( .A(n15932), .B(n15933), .Z(n9351) );
  XNOR U17756 ( .A(n[798]), .B(n15934), .Z(n15930) );
  IV U17757 ( .A(n15929), .Z(n15934) );
  XOR U17758 ( .A(n15935), .B(n15936), .Z(n15929) );
  AND U17759 ( .A(n15937), .B(n15938), .Z(n15935) );
  XOR U17760 ( .A(n15936), .B(n9356), .Z(n15938) );
  XNOR U17761 ( .A(n15939), .B(n15940), .Z(n9356) );
  XNOR U17762 ( .A(n[797]), .B(n15941), .Z(n15937) );
  IV U17763 ( .A(n15936), .Z(n15941) );
  XOR U17764 ( .A(n15942), .B(n15943), .Z(n15936) );
  AND U17765 ( .A(n15944), .B(n15945), .Z(n15942) );
  XOR U17766 ( .A(n15943), .B(n9361), .Z(n15945) );
  XNOR U17767 ( .A(n15946), .B(n15947), .Z(n9361) );
  XNOR U17768 ( .A(n[796]), .B(n15948), .Z(n15944) );
  IV U17769 ( .A(n15943), .Z(n15948) );
  XOR U17770 ( .A(n15949), .B(n15950), .Z(n15943) );
  AND U17771 ( .A(n15951), .B(n15952), .Z(n15949) );
  XOR U17772 ( .A(n15950), .B(n9366), .Z(n15952) );
  XNOR U17773 ( .A(n15953), .B(n15954), .Z(n9366) );
  XNOR U17774 ( .A(n[795]), .B(n15955), .Z(n15951) );
  IV U17775 ( .A(n15950), .Z(n15955) );
  XOR U17776 ( .A(n15956), .B(n15957), .Z(n15950) );
  AND U17777 ( .A(n15958), .B(n15959), .Z(n15956) );
  XOR U17778 ( .A(n15957), .B(n9371), .Z(n15959) );
  XNOR U17779 ( .A(n15960), .B(n15961), .Z(n9371) );
  XNOR U17780 ( .A(n[794]), .B(n15962), .Z(n15958) );
  IV U17781 ( .A(n15957), .Z(n15962) );
  XOR U17782 ( .A(n15963), .B(n15964), .Z(n15957) );
  AND U17783 ( .A(n15965), .B(n15966), .Z(n15963) );
  XOR U17784 ( .A(n15964), .B(n9376), .Z(n15966) );
  XNOR U17785 ( .A(n15967), .B(n15968), .Z(n9376) );
  XNOR U17786 ( .A(n[793]), .B(n15969), .Z(n15965) );
  IV U17787 ( .A(n15964), .Z(n15969) );
  XOR U17788 ( .A(n15970), .B(n15971), .Z(n15964) );
  AND U17789 ( .A(n15972), .B(n15973), .Z(n15970) );
  XOR U17790 ( .A(n15971), .B(n9381), .Z(n15973) );
  XNOR U17791 ( .A(n15974), .B(n15975), .Z(n9381) );
  XNOR U17792 ( .A(n[792]), .B(n15976), .Z(n15972) );
  IV U17793 ( .A(n15971), .Z(n15976) );
  XOR U17794 ( .A(n15977), .B(n15978), .Z(n15971) );
  AND U17795 ( .A(n15979), .B(n15980), .Z(n15977) );
  XOR U17796 ( .A(n15978), .B(n9386), .Z(n15980) );
  XNOR U17797 ( .A(n15981), .B(n15982), .Z(n9386) );
  XNOR U17798 ( .A(n[791]), .B(n15983), .Z(n15979) );
  IV U17799 ( .A(n15978), .Z(n15983) );
  XOR U17800 ( .A(n15984), .B(n15985), .Z(n15978) );
  AND U17801 ( .A(n15986), .B(n15987), .Z(n15984) );
  XOR U17802 ( .A(n15985), .B(n9391), .Z(n15987) );
  XNOR U17803 ( .A(n15988), .B(n15989), .Z(n9391) );
  XNOR U17804 ( .A(n[790]), .B(n15990), .Z(n15986) );
  IV U17805 ( .A(n15985), .Z(n15990) );
  XOR U17806 ( .A(n15991), .B(n15992), .Z(n15985) );
  AND U17807 ( .A(n15993), .B(n15994), .Z(n15991) );
  XOR U17808 ( .A(n15992), .B(n9396), .Z(n15994) );
  XNOR U17809 ( .A(n15995), .B(n15996), .Z(n9396) );
  XNOR U17810 ( .A(n[789]), .B(n15997), .Z(n15993) );
  IV U17811 ( .A(n15992), .Z(n15997) );
  XOR U17812 ( .A(n15998), .B(n15999), .Z(n15992) );
  AND U17813 ( .A(n16000), .B(n16001), .Z(n15998) );
  XOR U17814 ( .A(n15999), .B(n9401), .Z(n16001) );
  XNOR U17815 ( .A(n16002), .B(n16003), .Z(n9401) );
  XNOR U17816 ( .A(n[788]), .B(n16004), .Z(n16000) );
  IV U17817 ( .A(n15999), .Z(n16004) );
  XOR U17818 ( .A(n16005), .B(n16006), .Z(n15999) );
  AND U17819 ( .A(n16007), .B(n16008), .Z(n16005) );
  XOR U17820 ( .A(n16006), .B(n9406), .Z(n16008) );
  XNOR U17821 ( .A(n16009), .B(n16010), .Z(n9406) );
  XNOR U17822 ( .A(n[787]), .B(n16011), .Z(n16007) );
  IV U17823 ( .A(n16006), .Z(n16011) );
  XOR U17824 ( .A(n16012), .B(n16013), .Z(n16006) );
  AND U17825 ( .A(n16014), .B(n16015), .Z(n16012) );
  XOR U17826 ( .A(n16013), .B(n9411), .Z(n16015) );
  XNOR U17827 ( .A(n16016), .B(n16017), .Z(n9411) );
  XNOR U17828 ( .A(n[786]), .B(n16018), .Z(n16014) );
  IV U17829 ( .A(n16013), .Z(n16018) );
  XOR U17830 ( .A(n16019), .B(n16020), .Z(n16013) );
  AND U17831 ( .A(n16021), .B(n16022), .Z(n16019) );
  XOR U17832 ( .A(n16020), .B(n9416), .Z(n16022) );
  XNOR U17833 ( .A(n16023), .B(n16024), .Z(n9416) );
  XNOR U17834 ( .A(n[785]), .B(n16025), .Z(n16021) );
  IV U17835 ( .A(n16020), .Z(n16025) );
  XOR U17836 ( .A(n16026), .B(n16027), .Z(n16020) );
  AND U17837 ( .A(n16028), .B(n16029), .Z(n16026) );
  XOR U17838 ( .A(n16027), .B(n9421), .Z(n16029) );
  XNOR U17839 ( .A(n16030), .B(n16031), .Z(n9421) );
  XNOR U17840 ( .A(n[784]), .B(n16032), .Z(n16028) );
  IV U17841 ( .A(n16027), .Z(n16032) );
  XOR U17842 ( .A(n16033), .B(n16034), .Z(n16027) );
  AND U17843 ( .A(n16035), .B(n16036), .Z(n16033) );
  XOR U17844 ( .A(n16034), .B(n9426), .Z(n16036) );
  XNOR U17845 ( .A(n16037), .B(n16038), .Z(n9426) );
  XNOR U17846 ( .A(n[783]), .B(n16039), .Z(n16035) );
  IV U17847 ( .A(n16034), .Z(n16039) );
  XOR U17848 ( .A(n16040), .B(n16041), .Z(n16034) );
  AND U17849 ( .A(n16042), .B(n16043), .Z(n16040) );
  XOR U17850 ( .A(n16041), .B(n9431), .Z(n16043) );
  XNOR U17851 ( .A(n16044), .B(n16045), .Z(n9431) );
  XNOR U17852 ( .A(n[782]), .B(n16046), .Z(n16042) );
  IV U17853 ( .A(n16041), .Z(n16046) );
  XOR U17854 ( .A(n16047), .B(n16048), .Z(n16041) );
  AND U17855 ( .A(n16049), .B(n16050), .Z(n16047) );
  XOR U17856 ( .A(n16048), .B(n9436), .Z(n16050) );
  XNOR U17857 ( .A(n16051), .B(n16052), .Z(n9436) );
  XNOR U17858 ( .A(n[781]), .B(n16053), .Z(n16049) );
  IV U17859 ( .A(n16048), .Z(n16053) );
  XOR U17860 ( .A(n16054), .B(n16055), .Z(n16048) );
  AND U17861 ( .A(n16056), .B(n16057), .Z(n16054) );
  XOR U17862 ( .A(n16055), .B(n9441), .Z(n16057) );
  XNOR U17863 ( .A(n16058), .B(n16059), .Z(n9441) );
  XNOR U17864 ( .A(n[780]), .B(n16060), .Z(n16056) );
  IV U17865 ( .A(n16055), .Z(n16060) );
  XOR U17866 ( .A(n16061), .B(n16062), .Z(n16055) );
  AND U17867 ( .A(n16063), .B(n16064), .Z(n16061) );
  XOR U17868 ( .A(n16062), .B(n9446), .Z(n16064) );
  XNOR U17869 ( .A(n16065), .B(n16066), .Z(n9446) );
  XNOR U17870 ( .A(n[779]), .B(n16067), .Z(n16063) );
  IV U17871 ( .A(n16062), .Z(n16067) );
  XOR U17872 ( .A(n16068), .B(n16069), .Z(n16062) );
  AND U17873 ( .A(n16070), .B(n16071), .Z(n16068) );
  XOR U17874 ( .A(n16069), .B(n9451), .Z(n16071) );
  XNOR U17875 ( .A(n16072), .B(n16073), .Z(n9451) );
  XNOR U17876 ( .A(n[778]), .B(n16074), .Z(n16070) );
  IV U17877 ( .A(n16069), .Z(n16074) );
  XOR U17878 ( .A(n16075), .B(n16076), .Z(n16069) );
  AND U17879 ( .A(n16077), .B(n16078), .Z(n16075) );
  XOR U17880 ( .A(n16076), .B(n9456), .Z(n16078) );
  XNOR U17881 ( .A(n16079), .B(n16080), .Z(n9456) );
  XNOR U17882 ( .A(n[777]), .B(n16081), .Z(n16077) );
  IV U17883 ( .A(n16076), .Z(n16081) );
  XOR U17884 ( .A(n16082), .B(n16083), .Z(n16076) );
  AND U17885 ( .A(n16084), .B(n16085), .Z(n16082) );
  XOR U17886 ( .A(n16083), .B(n9461), .Z(n16085) );
  XNOR U17887 ( .A(n16086), .B(n16087), .Z(n9461) );
  XNOR U17888 ( .A(n[776]), .B(n16088), .Z(n16084) );
  IV U17889 ( .A(n16083), .Z(n16088) );
  XOR U17890 ( .A(n16089), .B(n16090), .Z(n16083) );
  AND U17891 ( .A(n16091), .B(n16092), .Z(n16089) );
  XOR U17892 ( .A(n16090), .B(n9466), .Z(n16092) );
  XNOR U17893 ( .A(n16093), .B(n16094), .Z(n9466) );
  XNOR U17894 ( .A(n[775]), .B(n16095), .Z(n16091) );
  IV U17895 ( .A(n16090), .Z(n16095) );
  XOR U17896 ( .A(n16096), .B(n16097), .Z(n16090) );
  AND U17897 ( .A(n16098), .B(n16099), .Z(n16096) );
  XOR U17898 ( .A(n16097), .B(n9471), .Z(n16099) );
  XNOR U17899 ( .A(n16100), .B(n16101), .Z(n9471) );
  XNOR U17900 ( .A(n[774]), .B(n16102), .Z(n16098) );
  IV U17901 ( .A(n16097), .Z(n16102) );
  XOR U17902 ( .A(n16103), .B(n16104), .Z(n16097) );
  AND U17903 ( .A(n16105), .B(n16106), .Z(n16103) );
  XOR U17904 ( .A(n16104), .B(n9476), .Z(n16106) );
  XNOR U17905 ( .A(n16107), .B(n16108), .Z(n9476) );
  XNOR U17906 ( .A(n[773]), .B(n16109), .Z(n16105) );
  IV U17907 ( .A(n16104), .Z(n16109) );
  XOR U17908 ( .A(n16110), .B(n16111), .Z(n16104) );
  AND U17909 ( .A(n16112), .B(n16113), .Z(n16110) );
  XOR U17910 ( .A(n16111), .B(n9481), .Z(n16113) );
  XNOR U17911 ( .A(n16114), .B(n16115), .Z(n9481) );
  XNOR U17912 ( .A(n[772]), .B(n16116), .Z(n16112) );
  IV U17913 ( .A(n16111), .Z(n16116) );
  XOR U17914 ( .A(n16117), .B(n16118), .Z(n16111) );
  AND U17915 ( .A(n16119), .B(n16120), .Z(n16117) );
  XOR U17916 ( .A(n16118), .B(n9486), .Z(n16120) );
  XNOR U17917 ( .A(n16121), .B(n16122), .Z(n9486) );
  XNOR U17918 ( .A(n[771]), .B(n16123), .Z(n16119) );
  IV U17919 ( .A(n16118), .Z(n16123) );
  XOR U17920 ( .A(n16124), .B(n16125), .Z(n16118) );
  AND U17921 ( .A(n16126), .B(n16127), .Z(n16124) );
  XOR U17922 ( .A(n16125), .B(n9491), .Z(n16127) );
  XNOR U17923 ( .A(n16128), .B(n16129), .Z(n9491) );
  XNOR U17924 ( .A(n[770]), .B(n16130), .Z(n16126) );
  IV U17925 ( .A(n16125), .Z(n16130) );
  XOR U17926 ( .A(n16131), .B(n16132), .Z(n16125) );
  AND U17927 ( .A(n16133), .B(n16134), .Z(n16131) );
  XOR U17928 ( .A(n16132), .B(n9496), .Z(n16134) );
  XNOR U17929 ( .A(n16135), .B(n16136), .Z(n9496) );
  XNOR U17930 ( .A(n[769]), .B(n16137), .Z(n16133) );
  IV U17931 ( .A(n16132), .Z(n16137) );
  XOR U17932 ( .A(n16138), .B(n16139), .Z(n16132) );
  AND U17933 ( .A(n16140), .B(n16141), .Z(n16138) );
  XOR U17934 ( .A(n16139), .B(n9501), .Z(n16141) );
  XNOR U17935 ( .A(n16142), .B(n16143), .Z(n9501) );
  XNOR U17936 ( .A(n[768]), .B(n16144), .Z(n16140) );
  IV U17937 ( .A(n16139), .Z(n16144) );
  XOR U17938 ( .A(n16145), .B(n16146), .Z(n16139) );
  AND U17939 ( .A(n16147), .B(n16148), .Z(n16145) );
  XOR U17940 ( .A(n16146), .B(n9506), .Z(n16148) );
  XNOR U17941 ( .A(n16149), .B(n16150), .Z(n9506) );
  XNOR U17942 ( .A(n[767]), .B(n16151), .Z(n16147) );
  IV U17943 ( .A(n16146), .Z(n16151) );
  XOR U17944 ( .A(n16152), .B(n16153), .Z(n16146) );
  AND U17945 ( .A(n16154), .B(n16155), .Z(n16152) );
  XOR U17946 ( .A(n16153), .B(n9511), .Z(n16155) );
  XNOR U17947 ( .A(n16156), .B(n16157), .Z(n9511) );
  XNOR U17948 ( .A(n[766]), .B(n16158), .Z(n16154) );
  IV U17949 ( .A(n16153), .Z(n16158) );
  XOR U17950 ( .A(n16159), .B(n16160), .Z(n16153) );
  AND U17951 ( .A(n16161), .B(n16162), .Z(n16159) );
  XOR U17952 ( .A(n16160), .B(n9516), .Z(n16162) );
  XNOR U17953 ( .A(n16163), .B(n16164), .Z(n9516) );
  XNOR U17954 ( .A(n[765]), .B(n16165), .Z(n16161) );
  IV U17955 ( .A(n16160), .Z(n16165) );
  XOR U17956 ( .A(n16166), .B(n16167), .Z(n16160) );
  AND U17957 ( .A(n16168), .B(n16169), .Z(n16166) );
  XOR U17958 ( .A(n16167), .B(n9521), .Z(n16169) );
  XNOR U17959 ( .A(n16170), .B(n16171), .Z(n9521) );
  XNOR U17960 ( .A(n[764]), .B(n16172), .Z(n16168) );
  IV U17961 ( .A(n16167), .Z(n16172) );
  XOR U17962 ( .A(n16173), .B(n16174), .Z(n16167) );
  AND U17963 ( .A(n16175), .B(n16176), .Z(n16173) );
  XOR U17964 ( .A(n16174), .B(n9526), .Z(n16176) );
  XNOR U17965 ( .A(n16177), .B(n16178), .Z(n9526) );
  XNOR U17966 ( .A(n[763]), .B(n16179), .Z(n16175) );
  IV U17967 ( .A(n16174), .Z(n16179) );
  XOR U17968 ( .A(n16180), .B(n16181), .Z(n16174) );
  AND U17969 ( .A(n16182), .B(n16183), .Z(n16180) );
  XOR U17970 ( .A(n16181), .B(n9531), .Z(n16183) );
  XNOR U17971 ( .A(n16184), .B(n16185), .Z(n9531) );
  XNOR U17972 ( .A(n[762]), .B(n16186), .Z(n16182) );
  IV U17973 ( .A(n16181), .Z(n16186) );
  XOR U17974 ( .A(n16187), .B(n16188), .Z(n16181) );
  AND U17975 ( .A(n16189), .B(n16190), .Z(n16187) );
  XOR U17976 ( .A(n16188), .B(n9536), .Z(n16190) );
  XNOR U17977 ( .A(n16191), .B(n16192), .Z(n9536) );
  XNOR U17978 ( .A(n[761]), .B(n16193), .Z(n16189) );
  IV U17979 ( .A(n16188), .Z(n16193) );
  XOR U17980 ( .A(n16194), .B(n16195), .Z(n16188) );
  AND U17981 ( .A(n16196), .B(n16197), .Z(n16194) );
  XOR U17982 ( .A(n16195), .B(n9541), .Z(n16197) );
  XNOR U17983 ( .A(n16198), .B(n16199), .Z(n9541) );
  XNOR U17984 ( .A(n[760]), .B(n16200), .Z(n16196) );
  IV U17985 ( .A(n16195), .Z(n16200) );
  XOR U17986 ( .A(n16201), .B(n16202), .Z(n16195) );
  AND U17987 ( .A(n16203), .B(n16204), .Z(n16201) );
  XOR U17988 ( .A(n16202), .B(n9546), .Z(n16204) );
  XNOR U17989 ( .A(n16205), .B(n16206), .Z(n9546) );
  XNOR U17990 ( .A(n[759]), .B(n16207), .Z(n16203) );
  IV U17991 ( .A(n16202), .Z(n16207) );
  XOR U17992 ( .A(n16208), .B(n16209), .Z(n16202) );
  AND U17993 ( .A(n16210), .B(n16211), .Z(n16208) );
  XOR U17994 ( .A(n16209), .B(n9551), .Z(n16211) );
  XNOR U17995 ( .A(n16212), .B(n16213), .Z(n9551) );
  XNOR U17996 ( .A(n[758]), .B(n16214), .Z(n16210) );
  IV U17997 ( .A(n16209), .Z(n16214) );
  XOR U17998 ( .A(n16215), .B(n16216), .Z(n16209) );
  AND U17999 ( .A(n16217), .B(n16218), .Z(n16215) );
  XOR U18000 ( .A(n16216), .B(n9556), .Z(n16218) );
  XNOR U18001 ( .A(n16219), .B(n16220), .Z(n9556) );
  XNOR U18002 ( .A(n[757]), .B(n16221), .Z(n16217) );
  IV U18003 ( .A(n16216), .Z(n16221) );
  XOR U18004 ( .A(n16222), .B(n16223), .Z(n16216) );
  AND U18005 ( .A(n16224), .B(n16225), .Z(n16222) );
  XOR U18006 ( .A(n16223), .B(n9561), .Z(n16225) );
  XNOR U18007 ( .A(n16226), .B(n16227), .Z(n9561) );
  XNOR U18008 ( .A(n[756]), .B(n16228), .Z(n16224) );
  IV U18009 ( .A(n16223), .Z(n16228) );
  XOR U18010 ( .A(n16229), .B(n16230), .Z(n16223) );
  AND U18011 ( .A(n16231), .B(n16232), .Z(n16229) );
  XOR U18012 ( .A(n16230), .B(n9566), .Z(n16232) );
  XNOR U18013 ( .A(n16233), .B(n16234), .Z(n9566) );
  XNOR U18014 ( .A(n[755]), .B(n16235), .Z(n16231) );
  IV U18015 ( .A(n16230), .Z(n16235) );
  XOR U18016 ( .A(n16236), .B(n16237), .Z(n16230) );
  AND U18017 ( .A(n16238), .B(n16239), .Z(n16236) );
  XOR U18018 ( .A(n16237), .B(n9571), .Z(n16239) );
  XNOR U18019 ( .A(n16240), .B(n16241), .Z(n9571) );
  XNOR U18020 ( .A(n[754]), .B(n16242), .Z(n16238) );
  IV U18021 ( .A(n16237), .Z(n16242) );
  XOR U18022 ( .A(n16243), .B(n16244), .Z(n16237) );
  AND U18023 ( .A(n16245), .B(n16246), .Z(n16243) );
  XOR U18024 ( .A(n16244), .B(n9576), .Z(n16246) );
  XNOR U18025 ( .A(n16247), .B(n16248), .Z(n9576) );
  XNOR U18026 ( .A(n[753]), .B(n16249), .Z(n16245) );
  IV U18027 ( .A(n16244), .Z(n16249) );
  XOR U18028 ( .A(n16250), .B(n16251), .Z(n16244) );
  AND U18029 ( .A(n16252), .B(n16253), .Z(n16250) );
  XOR U18030 ( .A(n16251), .B(n9581), .Z(n16253) );
  XNOR U18031 ( .A(n16254), .B(n16255), .Z(n9581) );
  XNOR U18032 ( .A(n[752]), .B(n16256), .Z(n16252) );
  IV U18033 ( .A(n16251), .Z(n16256) );
  XOR U18034 ( .A(n16257), .B(n16258), .Z(n16251) );
  AND U18035 ( .A(n16259), .B(n16260), .Z(n16257) );
  XOR U18036 ( .A(n16258), .B(n9586), .Z(n16260) );
  XNOR U18037 ( .A(n16261), .B(n16262), .Z(n9586) );
  XNOR U18038 ( .A(n[751]), .B(n16263), .Z(n16259) );
  IV U18039 ( .A(n16258), .Z(n16263) );
  XOR U18040 ( .A(n16264), .B(n16265), .Z(n16258) );
  AND U18041 ( .A(n16266), .B(n16267), .Z(n16264) );
  XOR U18042 ( .A(n16265), .B(n9591), .Z(n16267) );
  XNOR U18043 ( .A(n16268), .B(n16269), .Z(n9591) );
  XNOR U18044 ( .A(n[750]), .B(n16270), .Z(n16266) );
  IV U18045 ( .A(n16265), .Z(n16270) );
  XOR U18046 ( .A(n16271), .B(n16272), .Z(n16265) );
  AND U18047 ( .A(n16273), .B(n16274), .Z(n16271) );
  XOR U18048 ( .A(n16272), .B(n9596), .Z(n16274) );
  XNOR U18049 ( .A(n16275), .B(n16276), .Z(n9596) );
  XNOR U18050 ( .A(n[749]), .B(n16277), .Z(n16273) );
  IV U18051 ( .A(n16272), .Z(n16277) );
  XOR U18052 ( .A(n16278), .B(n16279), .Z(n16272) );
  AND U18053 ( .A(n16280), .B(n16281), .Z(n16278) );
  XOR U18054 ( .A(n16279), .B(n9601), .Z(n16281) );
  XNOR U18055 ( .A(n16282), .B(n16283), .Z(n9601) );
  XNOR U18056 ( .A(n[748]), .B(n16284), .Z(n16280) );
  IV U18057 ( .A(n16279), .Z(n16284) );
  XOR U18058 ( .A(n16285), .B(n16286), .Z(n16279) );
  AND U18059 ( .A(n16287), .B(n16288), .Z(n16285) );
  XOR U18060 ( .A(n16286), .B(n9606), .Z(n16288) );
  XNOR U18061 ( .A(n16289), .B(n16290), .Z(n9606) );
  XNOR U18062 ( .A(n[747]), .B(n16291), .Z(n16287) );
  IV U18063 ( .A(n16286), .Z(n16291) );
  XOR U18064 ( .A(n16292), .B(n16293), .Z(n16286) );
  AND U18065 ( .A(n16294), .B(n16295), .Z(n16292) );
  XOR U18066 ( .A(n16293), .B(n9611), .Z(n16295) );
  XNOR U18067 ( .A(n16296), .B(n16297), .Z(n9611) );
  XNOR U18068 ( .A(n[746]), .B(n16298), .Z(n16294) );
  IV U18069 ( .A(n16293), .Z(n16298) );
  XOR U18070 ( .A(n16299), .B(n16300), .Z(n16293) );
  AND U18071 ( .A(n16301), .B(n16302), .Z(n16299) );
  XOR U18072 ( .A(n16300), .B(n9616), .Z(n16302) );
  XNOR U18073 ( .A(n16303), .B(n16304), .Z(n9616) );
  XNOR U18074 ( .A(n[745]), .B(n16305), .Z(n16301) );
  IV U18075 ( .A(n16300), .Z(n16305) );
  XOR U18076 ( .A(n16306), .B(n16307), .Z(n16300) );
  AND U18077 ( .A(n16308), .B(n16309), .Z(n16306) );
  XOR U18078 ( .A(n16307), .B(n9621), .Z(n16309) );
  XNOR U18079 ( .A(n16310), .B(n16311), .Z(n9621) );
  XNOR U18080 ( .A(n[744]), .B(n16312), .Z(n16308) );
  IV U18081 ( .A(n16307), .Z(n16312) );
  XOR U18082 ( .A(n16313), .B(n16314), .Z(n16307) );
  AND U18083 ( .A(n16315), .B(n16316), .Z(n16313) );
  XOR U18084 ( .A(n16314), .B(n9626), .Z(n16316) );
  XNOR U18085 ( .A(n16317), .B(n16318), .Z(n9626) );
  XNOR U18086 ( .A(n[743]), .B(n16319), .Z(n16315) );
  IV U18087 ( .A(n16314), .Z(n16319) );
  XOR U18088 ( .A(n16320), .B(n16321), .Z(n16314) );
  AND U18089 ( .A(n16322), .B(n16323), .Z(n16320) );
  XOR U18090 ( .A(n16321), .B(n9631), .Z(n16323) );
  XNOR U18091 ( .A(n16324), .B(n16325), .Z(n9631) );
  XNOR U18092 ( .A(n[742]), .B(n16326), .Z(n16322) );
  IV U18093 ( .A(n16321), .Z(n16326) );
  XOR U18094 ( .A(n16327), .B(n16328), .Z(n16321) );
  AND U18095 ( .A(n16329), .B(n16330), .Z(n16327) );
  XOR U18096 ( .A(n16328), .B(n9636), .Z(n16330) );
  XNOR U18097 ( .A(n16331), .B(n16332), .Z(n9636) );
  XNOR U18098 ( .A(n[741]), .B(n16333), .Z(n16329) );
  IV U18099 ( .A(n16328), .Z(n16333) );
  XOR U18100 ( .A(n16334), .B(n16335), .Z(n16328) );
  AND U18101 ( .A(n16336), .B(n16337), .Z(n16334) );
  XOR U18102 ( .A(n16335), .B(n9641), .Z(n16337) );
  XNOR U18103 ( .A(n16338), .B(n16339), .Z(n9641) );
  XNOR U18104 ( .A(n[740]), .B(n16340), .Z(n16336) );
  IV U18105 ( .A(n16335), .Z(n16340) );
  XOR U18106 ( .A(n16341), .B(n16342), .Z(n16335) );
  AND U18107 ( .A(n16343), .B(n16344), .Z(n16341) );
  XOR U18108 ( .A(n16342), .B(n9646), .Z(n16344) );
  XNOR U18109 ( .A(n16345), .B(n16346), .Z(n9646) );
  XNOR U18110 ( .A(n[739]), .B(n16347), .Z(n16343) );
  IV U18111 ( .A(n16342), .Z(n16347) );
  XOR U18112 ( .A(n16348), .B(n16349), .Z(n16342) );
  AND U18113 ( .A(n16350), .B(n16351), .Z(n16348) );
  XOR U18114 ( .A(n16349), .B(n9651), .Z(n16351) );
  XNOR U18115 ( .A(n16352), .B(n16353), .Z(n9651) );
  XNOR U18116 ( .A(n[738]), .B(n16354), .Z(n16350) );
  IV U18117 ( .A(n16349), .Z(n16354) );
  XOR U18118 ( .A(n16355), .B(n16356), .Z(n16349) );
  AND U18119 ( .A(n16357), .B(n16358), .Z(n16355) );
  XOR U18120 ( .A(n16356), .B(n9656), .Z(n16358) );
  XNOR U18121 ( .A(n16359), .B(n16360), .Z(n9656) );
  XNOR U18122 ( .A(n[737]), .B(n16361), .Z(n16357) );
  IV U18123 ( .A(n16356), .Z(n16361) );
  XOR U18124 ( .A(n16362), .B(n16363), .Z(n16356) );
  AND U18125 ( .A(n16364), .B(n16365), .Z(n16362) );
  XOR U18126 ( .A(n16363), .B(n9661), .Z(n16365) );
  XNOR U18127 ( .A(n16366), .B(n16367), .Z(n9661) );
  XNOR U18128 ( .A(n[736]), .B(n16368), .Z(n16364) );
  IV U18129 ( .A(n16363), .Z(n16368) );
  XOR U18130 ( .A(n16369), .B(n16370), .Z(n16363) );
  AND U18131 ( .A(n16371), .B(n16372), .Z(n16369) );
  XOR U18132 ( .A(n16370), .B(n9666), .Z(n16372) );
  XNOR U18133 ( .A(n16373), .B(n16374), .Z(n9666) );
  XNOR U18134 ( .A(n[735]), .B(n16375), .Z(n16371) );
  IV U18135 ( .A(n16370), .Z(n16375) );
  XOR U18136 ( .A(n16376), .B(n16377), .Z(n16370) );
  AND U18137 ( .A(n16378), .B(n16379), .Z(n16376) );
  XOR U18138 ( .A(n16377), .B(n9671), .Z(n16379) );
  XNOR U18139 ( .A(n16380), .B(n16381), .Z(n9671) );
  XNOR U18140 ( .A(n[734]), .B(n16382), .Z(n16378) );
  IV U18141 ( .A(n16377), .Z(n16382) );
  XOR U18142 ( .A(n16383), .B(n16384), .Z(n16377) );
  AND U18143 ( .A(n16385), .B(n16386), .Z(n16383) );
  XOR U18144 ( .A(n16384), .B(n9676), .Z(n16386) );
  XNOR U18145 ( .A(n16387), .B(n16388), .Z(n9676) );
  XNOR U18146 ( .A(n[733]), .B(n16389), .Z(n16385) );
  IV U18147 ( .A(n16384), .Z(n16389) );
  XOR U18148 ( .A(n16390), .B(n16391), .Z(n16384) );
  AND U18149 ( .A(n16392), .B(n16393), .Z(n16390) );
  XOR U18150 ( .A(n16391), .B(n9681), .Z(n16393) );
  XNOR U18151 ( .A(n16394), .B(n16395), .Z(n9681) );
  XNOR U18152 ( .A(n[732]), .B(n16396), .Z(n16392) );
  IV U18153 ( .A(n16391), .Z(n16396) );
  XOR U18154 ( .A(n16397), .B(n16398), .Z(n16391) );
  AND U18155 ( .A(n16399), .B(n16400), .Z(n16397) );
  XOR U18156 ( .A(n16398), .B(n9686), .Z(n16400) );
  XNOR U18157 ( .A(n16401), .B(n16402), .Z(n9686) );
  XNOR U18158 ( .A(n[731]), .B(n16403), .Z(n16399) );
  IV U18159 ( .A(n16398), .Z(n16403) );
  XOR U18160 ( .A(n16404), .B(n16405), .Z(n16398) );
  AND U18161 ( .A(n16406), .B(n16407), .Z(n16404) );
  XOR U18162 ( .A(n16405), .B(n9691), .Z(n16407) );
  XNOR U18163 ( .A(n16408), .B(n16409), .Z(n9691) );
  XNOR U18164 ( .A(n[730]), .B(n16410), .Z(n16406) );
  IV U18165 ( .A(n16405), .Z(n16410) );
  XOR U18166 ( .A(n16411), .B(n16412), .Z(n16405) );
  AND U18167 ( .A(n16413), .B(n16414), .Z(n16411) );
  XOR U18168 ( .A(n16412), .B(n9696), .Z(n16414) );
  XNOR U18169 ( .A(n16415), .B(n16416), .Z(n9696) );
  XNOR U18170 ( .A(n[729]), .B(n16417), .Z(n16413) );
  IV U18171 ( .A(n16412), .Z(n16417) );
  XOR U18172 ( .A(n16418), .B(n16419), .Z(n16412) );
  AND U18173 ( .A(n16420), .B(n16421), .Z(n16418) );
  XOR U18174 ( .A(n16419), .B(n9701), .Z(n16421) );
  XNOR U18175 ( .A(n16422), .B(n16423), .Z(n9701) );
  XNOR U18176 ( .A(n[728]), .B(n16424), .Z(n16420) );
  IV U18177 ( .A(n16419), .Z(n16424) );
  XOR U18178 ( .A(n16425), .B(n16426), .Z(n16419) );
  AND U18179 ( .A(n16427), .B(n16428), .Z(n16425) );
  XOR U18180 ( .A(n16426), .B(n9706), .Z(n16428) );
  XNOR U18181 ( .A(n16429), .B(n16430), .Z(n9706) );
  XNOR U18182 ( .A(n[727]), .B(n16431), .Z(n16427) );
  IV U18183 ( .A(n16426), .Z(n16431) );
  XOR U18184 ( .A(n16432), .B(n16433), .Z(n16426) );
  AND U18185 ( .A(n16434), .B(n16435), .Z(n16432) );
  XOR U18186 ( .A(n16433), .B(n9711), .Z(n16435) );
  XNOR U18187 ( .A(n16436), .B(n16437), .Z(n9711) );
  XNOR U18188 ( .A(n[726]), .B(n16438), .Z(n16434) );
  IV U18189 ( .A(n16433), .Z(n16438) );
  XOR U18190 ( .A(n16439), .B(n16440), .Z(n16433) );
  AND U18191 ( .A(n16441), .B(n16442), .Z(n16439) );
  XOR U18192 ( .A(n16440), .B(n9716), .Z(n16442) );
  XNOR U18193 ( .A(n16443), .B(n16444), .Z(n9716) );
  XNOR U18194 ( .A(n[725]), .B(n16445), .Z(n16441) );
  IV U18195 ( .A(n16440), .Z(n16445) );
  XOR U18196 ( .A(n16446), .B(n16447), .Z(n16440) );
  AND U18197 ( .A(n16448), .B(n16449), .Z(n16446) );
  XOR U18198 ( .A(n16447), .B(n9721), .Z(n16449) );
  XNOR U18199 ( .A(n16450), .B(n16451), .Z(n9721) );
  XNOR U18200 ( .A(n[724]), .B(n16452), .Z(n16448) );
  IV U18201 ( .A(n16447), .Z(n16452) );
  XOR U18202 ( .A(n16453), .B(n16454), .Z(n16447) );
  AND U18203 ( .A(n16455), .B(n16456), .Z(n16453) );
  XOR U18204 ( .A(n16454), .B(n9726), .Z(n16456) );
  XNOR U18205 ( .A(n16457), .B(n16458), .Z(n9726) );
  XNOR U18206 ( .A(n[723]), .B(n16459), .Z(n16455) );
  IV U18207 ( .A(n16454), .Z(n16459) );
  XOR U18208 ( .A(n16460), .B(n16461), .Z(n16454) );
  AND U18209 ( .A(n16462), .B(n16463), .Z(n16460) );
  XOR U18210 ( .A(n16461), .B(n9731), .Z(n16463) );
  XNOR U18211 ( .A(n16464), .B(n16465), .Z(n9731) );
  XNOR U18212 ( .A(n[722]), .B(n16466), .Z(n16462) );
  IV U18213 ( .A(n16461), .Z(n16466) );
  XOR U18214 ( .A(n16467), .B(n16468), .Z(n16461) );
  AND U18215 ( .A(n16469), .B(n16470), .Z(n16467) );
  XOR U18216 ( .A(n16468), .B(n9736), .Z(n16470) );
  XNOR U18217 ( .A(n16471), .B(n16472), .Z(n9736) );
  XNOR U18218 ( .A(n[721]), .B(n16473), .Z(n16469) );
  IV U18219 ( .A(n16468), .Z(n16473) );
  XOR U18220 ( .A(n16474), .B(n16475), .Z(n16468) );
  AND U18221 ( .A(n16476), .B(n16477), .Z(n16474) );
  XOR U18222 ( .A(n16475), .B(n9741), .Z(n16477) );
  XNOR U18223 ( .A(n16478), .B(n16479), .Z(n9741) );
  XNOR U18224 ( .A(n[720]), .B(n16480), .Z(n16476) );
  IV U18225 ( .A(n16475), .Z(n16480) );
  XOR U18226 ( .A(n16481), .B(n16482), .Z(n16475) );
  AND U18227 ( .A(n16483), .B(n16484), .Z(n16481) );
  XOR U18228 ( .A(n16482), .B(n9746), .Z(n16484) );
  XNOR U18229 ( .A(n16485), .B(n16486), .Z(n9746) );
  XNOR U18230 ( .A(n[719]), .B(n16487), .Z(n16483) );
  IV U18231 ( .A(n16482), .Z(n16487) );
  XOR U18232 ( .A(n16488), .B(n16489), .Z(n16482) );
  AND U18233 ( .A(n16490), .B(n16491), .Z(n16488) );
  XOR U18234 ( .A(n16489), .B(n9751), .Z(n16491) );
  XNOR U18235 ( .A(n16492), .B(n16493), .Z(n9751) );
  XNOR U18236 ( .A(n[718]), .B(n16494), .Z(n16490) );
  IV U18237 ( .A(n16489), .Z(n16494) );
  XOR U18238 ( .A(n16495), .B(n16496), .Z(n16489) );
  AND U18239 ( .A(n16497), .B(n16498), .Z(n16495) );
  XOR U18240 ( .A(n16496), .B(n9756), .Z(n16498) );
  XNOR U18241 ( .A(n16499), .B(n16500), .Z(n9756) );
  XNOR U18242 ( .A(n[717]), .B(n16501), .Z(n16497) );
  IV U18243 ( .A(n16496), .Z(n16501) );
  XOR U18244 ( .A(n16502), .B(n16503), .Z(n16496) );
  AND U18245 ( .A(n16504), .B(n16505), .Z(n16502) );
  XOR U18246 ( .A(n16503), .B(n9761), .Z(n16505) );
  XNOR U18247 ( .A(n16506), .B(n16507), .Z(n9761) );
  XNOR U18248 ( .A(n[716]), .B(n16508), .Z(n16504) );
  IV U18249 ( .A(n16503), .Z(n16508) );
  XOR U18250 ( .A(n16509), .B(n16510), .Z(n16503) );
  AND U18251 ( .A(n16511), .B(n16512), .Z(n16509) );
  XOR U18252 ( .A(n16510), .B(n9766), .Z(n16512) );
  XNOR U18253 ( .A(n16513), .B(n16514), .Z(n9766) );
  XNOR U18254 ( .A(n[715]), .B(n16515), .Z(n16511) );
  IV U18255 ( .A(n16510), .Z(n16515) );
  XOR U18256 ( .A(n16516), .B(n16517), .Z(n16510) );
  AND U18257 ( .A(n16518), .B(n16519), .Z(n16516) );
  XOR U18258 ( .A(n16517), .B(n9771), .Z(n16519) );
  XNOR U18259 ( .A(n16520), .B(n16521), .Z(n9771) );
  XNOR U18260 ( .A(n[714]), .B(n16522), .Z(n16518) );
  IV U18261 ( .A(n16517), .Z(n16522) );
  XOR U18262 ( .A(n16523), .B(n16524), .Z(n16517) );
  AND U18263 ( .A(n16525), .B(n16526), .Z(n16523) );
  XOR U18264 ( .A(n16524), .B(n9776), .Z(n16526) );
  XNOR U18265 ( .A(n16527), .B(n16528), .Z(n9776) );
  XNOR U18266 ( .A(n[713]), .B(n16529), .Z(n16525) );
  IV U18267 ( .A(n16524), .Z(n16529) );
  XOR U18268 ( .A(n16530), .B(n16531), .Z(n16524) );
  AND U18269 ( .A(n16532), .B(n16533), .Z(n16530) );
  XOR U18270 ( .A(n16531), .B(n9781), .Z(n16533) );
  XNOR U18271 ( .A(n16534), .B(n16535), .Z(n9781) );
  XNOR U18272 ( .A(n[712]), .B(n16536), .Z(n16532) );
  IV U18273 ( .A(n16531), .Z(n16536) );
  XOR U18274 ( .A(n16537), .B(n16538), .Z(n16531) );
  AND U18275 ( .A(n16539), .B(n16540), .Z(n16537) );
  XOR U18276 ( .A(n16538), .B(n9786), .Z(n16540) );
  XNOR U18277 ( .A(n16541), .B(n16542), .Z(n9786) );
  XNOR U18278 ( .A(n[711]), .B(n16543), .Z(n16539) );
  IV U18279 ( .A(n16538), .Z(n16543) );
  XOR U18280 ( .A(n16544), .B(n16545), .Z(n16538) );
  AND U18281 ( .A(n16546), .B(n16547), .Z(n16544) );
  XOR U18282 ( .A(n16545), .B(n9791), .Z(n16547) );
  XNOR U18283 ( .A(n16548), .B(n16549), .Z(n9791) );
  XNOR U18284 ( .A(n[710]), .B(n16550), .Z(n16546) );
  IV U18285 ( .A(n16545), .Z(n16550) );
  XOR U18286 ( .A(n16551), .B(n16552), .Z(n16545) );
  AND U18287 ( .A(n16553), .B(n16554), .Z(n16551) );
  XOR U18288 ( .A(n16552), .B(n9796), .Z(n16554) );
  XNOR U18289 ( .A(n16555), .B(n16556), .Z(n9796) );
  XNOR U18290 ( .A(n[709]), .B(n16557), .Z(n16553) );
  IV U18291 ( .A(n16552), .Z(n16557) );
  XOR U18292 ( .A(n16558), .B(n16559), .Z(n16552) );
  AND U18293 ( .A(n16560), .B(n16561), .Z(n16558) );
  XOR U18294 ( .A(n16559), .B(n9801), .Z(n16561) );
  XNOR U18295 ( .A(n16562), .B(n16563), .Z(n9801) );
  XNOR U18296 ( .A(n[708]), .B(n16564), .Z(n16560) );
  IV U18297 ( .A(n16559), .Z(n16564) );
  XOR U18298 ( .A(n16565), .B(n16566), .Z(n16559) );
  AND U18299 ( .A(n16567), .B(n16568), .Z(n16565) );
  XOR U18300 ( .A(n16566), .B(n9806), .Z(n16568) );
  XNOR U18301 ( .A(n16569), .B(n16570), .Z(n9806) );
  XNOR U18302 ( .A(n[707]), .B(n16571), .Z(n16567) );
  IV U18303 ( .A(n16566), .Z(n16571) );
  XOR U18304 ( .A(n16572), .B(n16573), .Z(n16566) );
  AND U18305 ( .A(n16574), .B(n16575), .Z(n16572) );
  XOR U18306 ( .A(n16573), .B(n9811), .Z(n16575) );
  XNOR U18307 ( .A(n16576), .B(n16577), .Z(n9811) );
  XNOR U18308 ( .A(n[706]), .B(n16578), .Z(n16574) );
  IV U18309 ( .A(n16573), .Z(n16578) );
  XOR U18310 ( .A(n16579), .B(n16580), .Z(n16573) );
  AND U18311 ( .A(n16581), .B(n16582), .Z(n16579) );
  XOR U18312 ( .A(n16580), .B(n9816), .Z(n16582) );
  XNOR U18313 ( .A(n16583), .B(n16584), .Z(n9816) );
  XNOR U18314 ( .A(n[705]), .B(n16585), .Z(n16581) );
  IV U18315 ( .A(n16580), .Z(n16585) );
  XOR U18316 ( .A(n16586), .B(n16587), .Z(n16580) );
  AND U18317 ( .A(n16588), .B(n16589), .Z(n16586) );
  XOR U18318 ( .A(n16587), .B(n9821), .Z(n16589) );
  XNOR U18319 ( .A(n16590), .B(n16591), .Z(n9821) );
  XNOR U18320 ( .A(n[704]), .B(n16592), .Z(n16588) );
  IV U18321 ( .A(n16587), .Z(n16592) );
  XOR U18322 ( .A(n16593), .B(n16594), .Z(n16587) );
  AND U18323 ( .A(n16595), .B(n16596), .Z(n16593) );
  XOR U18324 ( .A(n16594), .B(n9826), .Z(n16596) );
  XNOR U18325 ( .A(n16597), .B(n16598), .Z(n9826) );
  XNOR U18326 ( .A(n[703]), .B(n16599), .Z(n16595) );
  IV U18327 ( .A(n16594), .Z(n16599) );
  XOR U18328 ( .A(n16600), .B(n16601), .Z(n16594) );
  AND U18329 ( .A(n16602), .B(n16603), .Z(n16600) );
  XOR U18330 ( .A(n16601), .B(n9831), .Z(n16603) );
  XNOR U18331 ( .A(n16604), .B(n16605), .Z(n9831) );
  XNOR U18332 ( .A(n[702]), .B(n16606), .Z(n16602) );
  IV U18333 ( .A(n16601), .Z(n16606) );
  XOR U18334 ( .A(n16607), .B(n16608), .Z(n16601) );
  AND U18335 ( .A(n16609), .B(n16610), .Z(n16607) );
  XOR U18336 ( .A(n16608), .B(n9836), .Z(n16610) );
  XNOR U18337 ( .A(n16611), .B(n16612), .Z(n9836) );
  XNOR U18338 ( .A(n[701]), .B(n16613), .Z(n16609) );
  IV U18339 ( .A(n16608), .Z(n16613) );
  XOR U18340 ( .A(n16614), .B(n16615), .Z(n16608) );
  AND U18341 ( .A(n16616), .B(n16617), .Z(n16614) );
  XOR U18342 ( .A(n16615), .B(n9841), .Z(n16617) );
  XNOR U18343 ( .A(n16618), .B(n16619), .Z(n9841) );
  XNOR U18344 ( .A(n[700]), .B(n16620), .Z(n16616) );
  IV U18345 ( .A(n16615), .Z(n16620) );
  XOR U18346 ( .A(n16621), .B(n16622), .Z(n16615) );
  AND U18347 ( .A(n16623), .B(n16624), .Z(n16621) );
  XOR U18348 ( .A(n16622), .B(n9846), .Z(n16624) );
  XNOR U18349 ( .A(n16625), .B(n16626), .Z(n9846) );
  XNOR U18350 ( .A(n[699]), .B(n16627), .Z(n16623) );
  IV U18351 ( .A(n16622), .Z(n16627) );
  XOR U18352 ( .A(n16628), .B(n16629), .Z(n16622) );
  AND U18353 ( .A(n16630), .B(n16631), .Z(n16628) );
  XOR U18354 ( .A(n16629), .B(n9851), .Z(n16631) );
  XNOR U18355 ( .A(n16632), .B(n16633), .Z(n9851) );
  XNOR U18356 ( .A(n[698]), .B(n16634), .Z(n16630) );
  IV U18357 ( .A(n16629), .Z(n16634) );
  XOR U18358 ( .A(n16635), .B(n16636), .Z(n16629) );
  AND U18359 ( .A(n16637), .B(n16638), .Z(n16635) );
  XOR U18360 ( .A(n16636), .B(n9856), .Z(n16638) );
  XNOR U18361 ( .A(n16639), .B(n16640), .Z(n9856) );
  XNOR U18362 ( .A(n[697]), .B(n16641), .Z(n16637) );
  IV U18363 ( .A(n16636), .Z(n16641) );
  XOR U18364 ( .A(n16642), .B(n16643), .Z(n16636) );
  AND U18365 ( .A(n16644), .B(n16645), .Z(n16642) );
  XOR U18366 ( .A(n16643), .B(n9861), .Z(n16645) );
  XNOR U18367 ( .A(n16646), .B(n16647), .Z(n9861) );
  XNOR U18368 ( .A(n[696]), .B(n16648), .Z(n16644) );
  IV U18369 ( .A(n16643), .Z(n16648) );
  XOR U18370 ( .A(n16649), .B(n16650), .Z(n16643) );
  AND U18371 ( .A(n16651), .B(n16652), .Z(n16649) );
  XOR U18372 ( .A(n16650), .B(n9866), .Z(n16652) );
  XNOR U18373 ( .A(n16653), .B(n16654), .Z(n9866) );
  XNOR U18374 ( .A(n[695]), .B(n16655), .Z(n16651) );
  IV U18375 ( .A(n16650), .Z(n16655) );
  XOR U18376 ( .A(n16656), .B(n16657), .Z(n16650) );
  AND U18377 ( .A(n16658), .B(n16659), .Z(n16656) );
  XOR U18378 ( .A(n16657), .B(n9871), .Z(n16659) );
  XNOR U18379 ( .A(n16660), .B(n16661), .Z(n9871) );
  XNOR U18380 ( .A(n[694]), .B(n16662), .Z(n16658) );
  IV U18381 ( .A(n16657), .Z(n16662) );
  XOR U18382 ( .A(n16663), .B(n16664), .Z(n16657) );
  AND U18383 ( .A(n16665), .B(n16666), .Z(n16663) );
  XOR U18384 ( .A(n16664), .B(n9876), .Z(n16666) );
  XNOR U18385 ( .A(n16667), .B(n16668), .Z(n9876) );
  XNOR U18386 ( .A(n[693]), .B(n16669), .Z(n16665) );
  IV U18387 ( .A(n16664), .Z(n16669) );
  XOR U18388 ( .A(n16670), .B(n16671), .Z(n16664) );
  AND U18389 ( .A(n16672), .B(n16673), .Z(n16670) );
  XOR U18390 ( .A(n16671), .B(n9881), .Z(n16673) );
  XNOR U18391 ( .A(n16674), .B(n16675), .Z(n9881) );
  XNOR U18392 ( .A(n[692]), .B(n16676), .Z(n16672) );
  IV U18393 ( .A(n16671), .Z(n16676) );
  XOR U18394 ( .A(n16677), .B(n16678), .Z(n16671) );
  AND U18395 ( .A(n16679), .B(n16680), .Z(n16677) );
  XOR U18396 ( .A(n16678), .B(n9886), .Z(n16680) );
  XNOR U18397 ( .A(n16681), .B(n16682), .Z(n9886) );
  XNOR U18398 ( .A(n[691]), .B(n16683), .Z(n16679) );
  IV U18399 ( .A(n16678), .Z(n16683) );
  XOR U18400 ( .A(n16684), .B(n16685), .Z(n16678) );
  AND U18401 ( .A(n16686), .B(n16687), .Z(n16684) );
  XOR U18402 ( .A(n16685), .B(n9891), .Z(n16687) );
  XNOR U18403 ( .A(n16688), .B(n16689), .Z(n9891) );
  XNOR U18404 ( .A(n[690]), .B(n16690), .Z(n16686) );
  IV U18405 ( .A(n16685), .Z(n16690) );
  XOR U18406 ( .A(n16691), .B(n16692), .Z(n16685) );
  AND U18407 ( .A(n16693), .B(n16694), .Z(n16691) );
  XOR U18408 ( .A(n16692), .B(n9896), .Z(n16694) );
  XNOR U18409 ( .A(n16695), .B(n16696), .Z(n9896) );
  XNOR U18410 ( .A(n[689]), .B(n16697), .Z(n16693) );
  IV U18411 ( .A(n16692), .Z(n16697) );
  XOR U18412 ( .A(n16698), .B(n16699), .Z(n16692) );
  AND U18413 ( .A(n16700), .B(n16701), .Z(n16698) );
  XOR U18414 ( .A(n16699), .B(n9901), .Z(n16701) );
  XNOR U18415 ( .A(n16702), .B(n16703), .Z(n9901) );
  XNOR U18416 ( .A(n[688]), .B(n16704), .Z(n16700) );
  IV U18417 ( .A(n16699), .Z(n16704) );
  XOR U18418 ( .A(n16705), .B(n16706), .Z(n16699) );
  AND U18419 ( .A(n16707), .B(n16708), .Z(n16705) );
  XOR U18420 ( .A(n16706), .B(n9906), .Z(n16708) );
  XNOR U18421 ( .A(n16709), .B(n16710), .Z(n9906) );
  XNOR U18422 ( .A(n[687]), .B(n16711), .Z(n16707) );
  IV U18423 ( .A(n16706), .Z(n16711) );
  XOR U18424 ( .A(n16712), .B(n16713), .Z(n16706) );
  AND U18425 ( .A(n16714), .B(n16715), .Z(n16712) );
  XOR U18426 ( .A(n16713), .B(n9911), .Z(n16715) );
  XNOR U18427 ( .A(n16716), .B(n16717), .Z(n9911) );
  XNOR U18428 ( .A(n[686]), .B(n16718), .Z(n16714) );
  IV U18429 ( .A(n16713), .Z(n16718) );
  XOR U18430 ( .A(n16719), .B(n16720), .Z(n16713) );
  AND U18431 ( .A(n16721), .B(n16722), .Z(n16719) );
  XOR U18432 ( .A(n16720), .B(n9916), .Z(n16722) );
  XNOR U18433 ( .A(n16723), .B(n16724), .Z(n9916) );
  XNOR U18434 ( .A(n[685]), .B(n16725), .Z(n16721) );
  IV U18435 ( .A(n16720), .Z(n16725) );
  XOR U18436 ( .A(n16726), .B(n16727), .Z(n16720) );
  AND U18437 ( .A(n16728), .B(n16729), .Z(n16726) );
  XOR U18438 ( .A(n16727), .B(n9921), .Z(n16729) );
  XNOR U18439 ( .A(n16730), .B(n16731), .Z(n9921) );
  XNOR U18440 ( .A(n[684]), .B(n16732), .Z(n16728) );
  IV U18441 ( .A(n16727), .Z(n16732) );
  XOR U18442 ( .A(n16733), .B(n16734), .Z(n16727) );
  AND U18443 ( .A(n16735), .B(n16736), .Z(n16733) );
  XOR U18444 ( .A(n16734), .B(n9926), .Z(n16736) );
  XNOR U18445 ( .A(n16737), .B(n16738), .Z(n9926) );
  XNOR U18446 ( .A(n[683]), .B(n16739), .Z(n16735) );
  IV U18447 ( .A(n16734), .Z(n16739) );
  XOR U18448 ( .A(n16740), .B(n16741), .Z(n16734) );
  AND U18449 ( .A(n16742), .B(n16743), .Z(n16740) );
  XOR U18450 ( .A(n16741), .B(n9931), .Z(n16743) );
  XNOR U18451 ( .A(n16744), .B(n16745), .Z(n9931) );
  XNOR U18452 ( .A(n[682]), .B(n16746), .Z(n16742) );
  IV U18453 ( .A(n16741), .Z(n16746) );
  XOR U18454 ( .A(n16747), .B(n16748), .Z(n16741) );
  AND U18455 ( .A(n16749), .B(n16750), .Z(n16747) );
  XOR U18456 ( .A(n16748), .B(n9936), .Z(n16750) );
  XNOR U18457 ( .A(n16751), .B(n16752), .Z(n9936) );
  XNOR U18458 ( .A(n[681]), .B(n16753), .Z(n16749) );
  IV U18459 ( .A(n16748), .Z(n16753) );
  XOR U18460 ( .A(n16754), .B(n16755), .Z(n16748) );
  AND U18461 ( .A(n16756), .B(n16757), .Z(n16754) );
  XOR U18462 ( .A(n16755), .B(n9941), .Z(n16757) );
  XNOR U18463 ( .A(n16758), .B(n16759), .Z(n9941) );
  XNOR U18464 ( .A(n[680]), .B(n16760), .Z(n16756) );
  IV U18465 ( .A(n16755), .Z(n16760) );
  XOR U18466 ( .A(n16761), .B(n16762), .Z(n16755) );
  AND U18467 ( .A(n16763), .B(n16764), .Z(n16761) );
  XOR U18468 ( .A(n16762), .B(n9946), .Z(n16764) );
  XNOR U18469 ( .A(n16765), .B(n16766), .Z(n9946) );
  XNOR U18470 ( .A(n[679]), .B(n16767), .Z(n16763) );
  IV U18471 ( .A(n16762), .Z(n16767) );
  XOR U18472 ( .A(n16768), .B(n16769), .Z(n16762) );
  AND U18473 ( .A(n16770), .B(n16771), .Z(n16768) );
  XOR U18474 ( .A(n16769), .B(n9951), .Z(n16771) );
  XNOR U18475 ( .A(n16772), .B(n16773), .Z(n9951) );
  XNOR U18476 ( .A(n[678]), .B(n16774), .Z(n16770) );
  IV U18477 ( .A(n16769), .Z(n16774) );
  XOR U18478 ( .A(n16775), .B(n16776), .Z(n16769) );
  AND U18479 ( .A(n16777), .B(n16778), .Z(n16775) );
  XOR U18480 ( .A(n16776), .B(n9956), .Z(n16778) );
  XNOR U18481 ( .A(n16779), .B(n16780), .Z(n9956) );
  XNOR U18482 ( .A(n[677]), .B(n16781), .Z(n16777) );
  IV U18483 ( .A(n16776), .Z(n16781) );
  XOR U18484 ( .A(n16782), .B(n16783), .Z(n16776) );
  AND U18485 ( .A(n16784), .B(n16785), .Z(n16782) );
  XOR U18486 ( .A(n16783), .B(n9961), .Z(n16785) );
  XNOR U18487 ( .A(n16786), .B(n16787), .Z(n9961) );
  XNOR U18488 ( .A(n[676]), .B(n16788), .Z(n16784) );
  IV U18489 ( .A(n16783), .Z(n16788) );
  XOR U18490 ( .A(n16789), .B(n16790), .Z(n16783) );
  AND U18491 ( .A(n16791), .B(n16792), .Z(n16789) );
  XOR U18492 ( .A(n16790), .B(n9966), .Z(n16792) );
  XNOR U18493 ( .A(n16793), .B(n16794), .Z(n9966) );
  XNOR U18494 ( .A(n[675]), .B(n16795), .Z(n16791) );
  IV U18495 ( .A(n16790), .Z(n16795) );
  XOR U18496 ( .A(n16796), .B(n16797), .Z(n16790) );
  AND U18497 ( .A(n16798), .B(n16799), .Z(n16796) );
  XOR U18498 ( .A(n16797), .B(n9971), .Z(n16799) );
  XNOR U18499 ( .A(n16800), .B(n16801), .Z(n9971) );
  XNOR U18500 ( .A(n[674]), .B(n16802), .Z(n16798) );
  IV U18501 ( .A(n16797), .Z(n16802) );
  XOR U18502 ( .A(n16803), .B(n16804), .Z(n16797) );
  AND U18503 ( .A(n16805), .B(n16806), .Z(n16803) );
  XOR U18504 ( .A(n16804), .B(n9976), .Z(n16806) );
  XNOR U18505 ( .A(n16807), .B(n16808), .Z(n9976) );
  XNOR U18506 ( .A(n[673]), .B(n16809), .Z(n16805) );
  IV U18507 ( .A(n16804), .Z(n16809) );
  XOR U18508 ( .A(n16810), .B(n16811), .Z(n16804) );
  AND U18509 ( .A(n16812), .B(n16813), .Z(n16810) );
  XOR U18510 ( .A(n16811), .B(n9981), .Z(n16813) );
  XNOR U18511 ( .A(n16814), .B(n16815), .Z(n9981) );
  XNOR U18512 ( .A(n[672]), .B(n16816), .Z(n16812) );
  IV U18513 ( .A(n16811), .Z(n16816) );
  XOR U18514 ( .A(n16817), .B(n16818), .Z(n16811) );
  AND U18515 ( .A(n16819), .B(n16820), .Z(n16817) );
  XOR U18516 ( .A(n16818), .B(n9986), .Z(n16820) );
  XNOR U18517 ( .A(n16821), .B(n16822), .Z(n9986) );
  XNOR U18518 ( .A(n[671]), .B(n16823), .Z(n16819) );
  IV U18519 ( .A(n16818), .Z(n16823) );
  XOR U18520 ( .A(n16824), .B(n16825), .Z(n16818) );
  AND U18521 ( .A(n16826), .B(n16827), .Z(n16824) );
  XOR U18522 ( .A(n16825), .B(n9991), .Z(n16827) );
  XNOR U18523 ( .A(n16828), .B(n16829), .Z(n9991) );
  XNOR U18524 ( .A(n[670]), .B(n16830), .Z(n16826) );
  IV U18525 ( .A(n16825), .Z(n16830) );
  XOR U18526 ( .A(n16831), .B(n16832), .Z(n16825) );
  AND U18527 ( .A(n16833), .B(n16834), .Z(n16831) );
  XOR U18528 ( .A(n16832), .B(n9996), .Z(n16834) );
  XNOR U18529 ( .A(n16835), .B(n16836), .Z(n9996) );
  XNOR U18530 ( .A(n[669]), .B(n16837), .Z(n16833) );
  IV U18531 ( .A(n16832), .Z(n16837) );
  XOR U18532 ( .A(n16838), .B(n16839), .Z(n16832) );
  AND U18533 ( .A(n16840), .B(n16841), .Z(n16838) );
  XOR U18534 ( .A(n16839), .B(n10001), .Z(n16841) );
  XNOR U18535 ( .A(n16842), .B(n16843), .Z(n10001) );
  XNOR U18536 ( .A(n[668]), .B(n16844), .Z(n16840) );
  IV U18537 ( .A(n16839), .Z(n16844) );
  XOR U18538 ( .A(n16845), .B(n16846), .Z(n16839) );
  AND U18539 ( .A(n16847), .B(n16848), .Z(n16845) );
  XOR U18540 ( .A(n16846), .B(n10006), .Z(n16848) );
  XNOR U18541 ( .A(n16849), .B(n16850), .Z(n10006) );
  XNOR U18542 ( .A(n[667]), .B(n16851), .Z(n16847) );
  IV U18543 ( .A(n16846), .Z(n16851) );
  XOR U18544 ( .A(n16852), .B(n16853), .Z(n16846) );
  AND U18545 ( .A(n16854), .B(n16855), .Z(n16852) );
  XOR U18546 ( .A(n16853), .B(n10011), .Z(n16855) );
  XNOR U18547 ( .A(n16856), .B(n16857), .Z(n10011) );
  XNOR U18548 ( .A(n[666]), .B(n16858), .Z(n16854) );
  IV U18549 ( .A(n16853), .Z(n16858) );
  XOR U18550 ( .A(n16859), .B(n16860), .Z(n16853) );
  AND U18551 ( .A(n16861), .B(n16862), .Z(n16859) );
  XOR U18552 ( .A(n16860), .B(n10016), .Z(n16862) );
  XNOR U18553 ( .A(n16863), .B(n16864), .Z(n10016) );
  XNOR U18554 ( .A(n[665]), .B(n16865), .Z(n16861) );
  IV U18555 ( .A(n16860), .Z(n16865) );
  XOR U18556 ( .A(n16866), .B(n16867), .Z(n16860) );
  AND U18557 ( .A(n16868), .B(n16869), .Z(n16866) );
  XOR U18558 ( .A(n16867), .B(n10021), .Z(n16869) );
  XNOR U18559 ( .A(n16870), .B(n16871), .Z(n10021) );
  XNOR U18560 ( .A(n[664]), .B(n16872), .Z(n16868) );
  IV U18561 ( .A(n16867), .Z(n16872) );
  XOR U18562 ( .A(n16873), .B(n16874), .Z(n16867) );
  AND U18563 ( .A(n16875), .B(n16876), .Z(n16873) );
  XOR U18564 ( .A(n16874), .B(n10026), .Z(n16876) );
  XNOR U18565 ( .A(n16877), .B(n16878), .Z(n10026) );
  XNOR U18566 ( .A(n[663]), .B(n16879), .Z(n16875) );
  IV U18567 ( .A(n16874), .Z(n16879) );
  XOR U18568 ( .A(n16880), .B(n16881), .Z(n16874) );
  AND U18569 ( .A(n16882), .B(n16883), .Z(n16880) );
  XOR U18570 ( .A(n16881), .B(n10031), .Z(n16883) );
  XNOR U18571 ( .A(n16884), .B(n16885), .Z(n10031) );
  XNOR U18572 ( .A(n[662]), .B(n16886), .Z(n16882) );
  IV U18573 ( .A(n16881), .Z(n16886) );
  XOR U18574 ( .A(n16887), .B(n16888), .Z(n16881) );
  AND U18575 ( .A(n16889), .B(n16890), .Z(n16887) );
  XOR U18576 ( .A(n16888), .B(n10036), .Z(n16890) );
  XNOR U18577 ( .A(n16891), .B(n16892), .Z(n10036) );
  XNOR U18578 ( .A(n[661]), .B(n16893), .Z(n16889) );
  IV U18579 ( .A(n16888), .Z(n16893) );
  XOR U18580 ( .A(n16894), .B(n16895), .Z(n16888) );
  AND U18581 ( .A(n16896), .B(n16897), .Z(n16894) );
  XOR U18582 ( .A(n16895), .B(n10041), .Z(n16897) );
  XNOR U18583 ( .A(n16898), .B(n16899), .Z(n10041) );
  XNOR U18584 ( .A(n[660]), .B(n16900), .Z(n16896) );
  IV U18585 ( .A(n16895), .Z(n16900) );
  XOR U18586 ( .A(n16901), .B(n16902), .Z(n16895) );
  AND U18587 ( .A(n16903), .B(n16904), .Z(n16901) );
  XOR U18588 ( .A(n16902), .B(n10046), .Z(n16904) );
  XNOR U18589 ( .A(n16905), .B(n16906), .Z(n10046) );
  XNOR U18590 ( .A(n[659]), .B(n16907), .Z(n16903) );
  IV U18591 ( .A(n16902), .Z(n16907) );
  XOR U18592 ( .A(n16908), .B(n16909), .Z(n16902) );
  AND U18593 ( .A(n16910), .B(n16911), .Z(n16908) );
  XOR U18594 ( .A(n16909), .B(n10051), .Z(n16911) );
  XNOR U18595 ( .A(n16912), .B(n16913), .Z(n10051) );
  XNOR U18596 ( .A(n[658]), .B(n16914), .Z(n16910) );
  IV U18597 ( .A(n16909), .Z(n16914) );
  XOR U18598 ( .A(n16915), .B(n16916), .Z(n16909) );
  AND U18599 ( .A(n16917), .B(n16918), .Z(n16915) );
  XOR U18600 ( .A(n16916), .B(n10056), .Z(n16918) );
  XNOR U18601 ( .A(n16919), .B(n16920), .Z(n10056) );
  XNOR U18602 ( .A(n[657]), .B(n16921), .Z(n16917) );
  IV U18603 ( .A(n16916), .Z(n16921) );
  XOR U18604 ( .A(n16922), .B(n16923), .Z(n16916) );
  AND U18605 ( .A(n16924), .B(n16925), .Z(n16922) );
  XOR U18606 ( .A(n16923), .B(n10061), .Z(n16925) );
  XNOR U18607 ( .A(n16926), .B(n16927), .Z(n10061) );
  XNOR U18608 ( .A(n[656]), .B(n16928), .Z(n16924) );
  IV U18609 ( .A(n16923), .Z(n16928) );
  XOR U18610 ( .A(n16929), .B(n16930), .Z(n16923) );
  AND U18611 ( .A(n16931), .B(n16932), .Z(n16929) );
  XOR U18612 ( .A(n16930), .B(n10066), .Z(n16932) );
  XNOR U18613 ( .A(n16933), .B(n16934), .Z(n10066) );
  XNOR U18614 ( .A(n[655]), .B(n16935), .Z(n16931) );
  IV U18615 ( .A(n16930), .Z(n16935) );
  XOR U18616 ( .A(n16936), .B(n16937), .Z(n16930) );
  AND U18617 ( .A(n16938), .B(n16939), .Z(n16936) );
  XOR U18618 ( .A(n16937), .B(n10071), .Z(n16939) );
  XNOR U18619 ( .A(n16940), .B(n16941), .Z(n10071) );
  XNOR U18620 ( .A(n[654]), .B(n16942), .Z(n16938) );
  IV U18621 ( .A(n16937), .Z(n16942) );
  XOR U18622 ( .A(n16943), .B(n16944), .Z(n16937) );
  AND U18623 ( .A(n16945), .B(n16946), .Z(n16943) );
  XOR U18624 ( .A(n16944), .B(n10076), .Z(n16946) );
  XNOR U18625 ( .A(n16947), .B(n16948), .Z(n10076) );
  XNOR U18626 ( .A(n[653]), .B(n16949), .Z(n16945) );
  IV U18627 ( .A(n16944), .Z(n16949) );
  XOR U18628 ( .A(n16950), .B(n16951), .Z(n16944) );
  AND U18629 ( .A(n16952), .B(n16953), .Z(n16950) );
  XOR U18630 ( .A(n16951), .B(n10081), .Z(n16953) );
  XNOR U18631 ( .A(n16954), .B(n16955), .Z(n10081) );
  XNOR U18632 ( .A(n[652]), .B(n16956), .Z(n16952) );
  IV U18633 ( .A(n16951), .Z(n16956) );
  XOR U18634 ( .A(n16957), .B(n16958), .Z(n16951) );
  AND U18635 ( .A(n16959), .B(n16960), .Z(n16957) );
  XOR U18636 ( .A(n16958), .B(n10086), .Z(n16960) );
  XNOR U18637 ( .A(n16961), .B(n16962), .Z(n10086) );
  XNOR U18638 ( .A(n[651]), .B(n16963), .Z(n16959) );
  IV U18639 ( .A(n16958), .Z(n16963) );
  XOR U18640 ( .A(n16964), .B(n16965), .Z(n16958) );
  AND U18641 ( .A(n16966), .B(n16967), .Z(n16964) );
  XOR U18642 ( .A(n16965), .B(n10091), .Z(n16967) );
  XNOR U18643 ( .A(n16968), .B(n16969), .Z(n10091) );
  XNOR U18644 ( .A(n[650]), .B(n16970), .Z(n16966) );
  IV U18645 ( .A(n16965), .Z(n16970) );
  XOR U18646 ( .A(n16971), .B(n16972), .Z(n16965) );
  AND U18647 ( .A(n16973), .B(n16974), .Z(n16971) );
  XOR U18648 ( .A(n16972), .B(n10096), .Z(n16974) );
  XNOR U18649 ( .A(n16975), .B(n16976), .Z(n10096) );
  XNOR U18650 ( .A(n[649]), .B(n16977), .Z(n16973) );
  IV U18651 ( .A(n16972), .Z(n16977) );
  XOR U18652 ( .A(n16978), .B(n16979), .Z(n16972) );
  AND U18653 ( .A(n16980), .B(n16981), .Z(n16978) );
  XOR U18654 ( .A(n16979), .B(n10101), .Z(n16981) );
  XNOR U18655 ( .A(n16982), .B(n16983), .Z(n10101) );
  XNOR U18656 ( .A(n[648]), .B(n16984), .Z(n16980) );
  IV U18657 ( .A(n16979), .Z(n16984) );
  XOR U18658 ( .A(n16985), .B(n16986), .Z(n16979) );
  AND U18659 ( .A(n16987), .B(n16988), .Z(n16985) );
  XOR U18660 ( .A(n16986), .B(n10106), .Z(n16988) );
  XNOR U18661 ( .A(n16989), .B(n16990), .Z(n10106) );
  XNOR U18662 ( .A(n[647]), .B(n16991), .Z(n16987) );
  IV U18663 ( .A(n16986), .Z(n16991) );
  XOR U18664 ( .A(n16992), .B(n16993), .Z(n16986) );
  AND U18665 ( .A(n16994), .B(n16995), .Z(n16992) );
  XOR U18666 ( .A(n16993), .B(n10111), .Z(n16995) );
  XNOR U18667 ( .A(n16996), .B(n16997), .Z(n10111) );
  XNOR U18668 ( .A(n[646]), .B(n16998), .Z(n16994) );
  IV U18669 ( .A(n16993), .Z(n16998) );
  XOR U18670 ( .A(n16999), .B(n17000), .Z(n16993) );
  AND U18671 ( .A(n17001), .B(n17002), .Z(n16999) );
  XOR U18672 ( .A(n17000), .B(n10116), .Z(n17002) );
  XNOR U18673 ( .A(n17003), .B(n17004), .Z(n10116) );
  XNOR U18674 ( .A(n[645]), .B(n17005), .Z(n17001) );
  IV U18675 ( .A(n17000), .Z(n17005) );
  XOR U18676 ( .A(n17006), .B(n17007), .Z(n17000) );
  AND U18677 ( .A(n17008), .B(n17009), .Z(n17006) );
  XOR U18678 ( .A(n17007), .B(n10121), .Z(n17009) );
  XNOR U18679 ( .A(n17010), .B(n17011), .Z(n10121) );
  XNOR U18680 ( .A(n[644]), .B(n17012), .Z(n17008) );
  IV U18681 ( .A(n17007), .Z(n17012) );
  XOR U18682 ( .A(n17013), .B(n17014), .Z(n17007) );
  AND U18683 ( .A(n17015), .B(n17016), .Z(n17013) );
  XOR U18684 ( .A(n17014), .B(n10126), .Z(n17016) );
  XNOR U18685 ( .A(n17017), .B(n17018), .Z(n10126) );
  XNOR U18686 ( .A(n[643]), .B(n17019), .Z(n17015) );
  IV U18687 ( .A(n17014), .Z(n17019) );
  XOR U18688 ( .A(n17020), .B(n17021), .Z(n17014) );
  AND U18689 ( .A(n17022), .B(n17023), .Z(n17020) );
  XOR U18690 ( .A(n17021), .B(n10131), .Z(n17023) );
  XNOR U18691 ( .A(n17024), .B(n17025), .Z(n10131) );
  XNOR U18692 ( .A(n[642]), .B(n17026), .Z(n17022) );
  IV U18693 ( .A(n17021), .Z(n17026) );
  XOR U18694 ( .A(n17027), .B(n17028), .Z(n17021) );
  AND U18695 ( .A(n17029), .B(n17030), .Z(n17027) );
  XOR U18696 ( .A(n17028), .B(n10136), .Z(n17030) );
  XNOR U18697 ( .A(n17031), .B(n17032), .Z(n10136) );
  XNOR U18698 ( .A(n[641]), .B(n17033), .Z(n17029) );
  IV U18699 ( .A(n17028), .Z(n17033) );
  XOR U18700 ( .A(n17034), .B(n17035), .Z(n17028) );
  AND U18701 ( .A(n17036), .B(n17037), .Z(n17034) );
  XOR U18702 ( .A(n17035), .B(n10141), .Z(n17037) );
  XNOR U18703 ( .A(n17038), .B(n17039), .Z(n10141) );
  XNOR U18704 ( .A(n[640]), .B(n17040), .Z(n17036) );
  IV U18705 ( .A(n17035), .Z(n17040) );
  XOR U18706 ( .A(n17041), .B(n17042), .Z(n17035) );
  AND U18707 ( .A(n17043), .B(n17044), .Z(n17041) );
  XOR U18708 ( .A(n17042), .B(n10146), .Z(n17044) );
  XNOR U18709 ( .A(n17045), .B(n17046), .Z(n10146) );
  XNOR U18710 ( .A(n[639]), .B(n17047), .Z(n17043) );
  IV U18711 ( .A(n17042), .Z(n17047) );
  XOR U18712 ( .A(n17048), .B(n17049), .Z(n17042) );
  AND U18713 ( .A(n17050), .B(n17051), .Z(n17048) );
  XOR U18714 ( .A(n17049), .B(n10151), .Z(n17051) );
  XNOR U18715 ( .A(n17052), .B(n17053), .Z(n10151) );
  XNOR U18716 ( .A(n[638]), .B(n17054), .Z(n17050) );
  IV U18717 ( .A(n17049), .Z(n17054) );
  XOR U18718 ( .A(n17055), .B(n17056), .Z(n17049) );
  AND U18719 ( .A(n17057), .B(n17058), .Z(n17055) );
  XOR U18720 ( .A(n17056), .B(n10156), .Z(n17058) );
  XNOR U18721 ( .A(n17059), .B(n17060), .Z(n10156) );
  XNOR U18722 ( .A(n[637]), .B(n17061), .Z(n17057) );
  IV U18723 ( .A(n17056), .Z(n17061) );
  XOR U18724 ( .A(n17062), .B(n17063), .Z(n17056) );
  AND U18725 ( .A(n17064), .B(n17065), .Z(n17062) );
  XOR U18726 ( .A(n17063), .B(n10161), .Z(n17065) );
  XNOR U18727 ( .A(n17066), .B(n17067), .Z(n10161) );
  XNOR U18728 ( .A(n[636]), .B(n17068), .Z(n17064) );
  IV U18729 ( .A(n17063), .Z(n17068) );
  XOR U18730 ( .A(n17069), .B(n17070), .Z(n17063) );
  AND U18731 ( .A(n17071), .B(n17072), .Z(n17069) );
  XOR U18732 ( .A(n17070), .B(n10166), .Z(n17072) );
  XNOR U18733 ( .A(n17073), .B(n17074), .Z(n10166) );
  XNOR U18734 ( .A(n[635]), .B(n17075), .Z(n17071) );
  IV U18735 ( .A(n17070), .Z(n17075) );
  XOR U18736 ( .A(n17076), .B(n17077), .Z(n17070) );
  AND U18737 ( .A(n17078), .B(n17079), .Z(n17076) );
  XOR U18738 ( .A(n17077), .B(n10171), .Z(n17079) );
  XNOR U18739 ( .A(n17080), .B(n17081), .Z(n10171) );
  XNOR U18740 ( .A(n[634]), .B(n17082), .Z(n17078) );
  IV U18741 ( .A(n17077), .Z(n17082) );
  XOR U18742 ( .A(n17083), .B(n17084), .Z(n17077) );
  AND U18743 ( .A(n17085), .B(n17086), .Z(n17083) );
  XOR U18744 ( .A(n17084), .B(n10176), .Z(n17086) );
  XNOR U18745 ( .A(n17087), .B(n17088), .Z(n10176) );
  XNOR U18746 ( .A(n[633]), .B(n17089), .Z(n17085) );
  IV U18747 ( .A(n17084), .Z(n17089) );
  XOR U18748 ( .A(n17090), .B(n17091), .Z(n17084) );
  AND U18749 ( .A(n17092), .B(n17093), .Z(n17090) );
  XOR U18750 ( .A(n17091), .B(n10181), .Z(n17093) );
  XNOR U18751 ( .A(n17094), .B(n17095), .Z(n10181) );
  XNOR U18752 ( .A(n[632]), .B(n17096), .Z(n17092) );
  IV U18753 ( .A(n17091), .Z(n17096) );
  XOR U18754 ( .A(n17097), .B(n17098), .Z(n17091) );
  AND U18755 ( .A(n17099), .B(n17100), .Z(n17097) );
  XOR U18756 ( .A(n17098), .B(n10186), .Z(n17100) );
  XNOR U18757 ( .A(n17101), .B(n17102), .Z(n10186) );
  XNOR U18758 ( .A(n[631]), .B(n17103), .Z(n17099) );
  IV U18759 ( .A(n17098), .Z(n17103) );
  XOR U18760 ( .A(n17104), .B(n17105), .Z(n17098) );
  AND U18761 ( .A(n17106), .B(n17107), .Z(n17104) );
  XOR U18762 ( .A(n17105), .B(n10191), .Z(n17107) );
  XNOR U18763 ( .A(n17108), .B(n17109), .Z(n10191) );
  XNOR U18764 ( .A(n[630]), .B(n17110), .Z(n17106) );
  IV U18765 ( .A(n17105), .Z(n17110) );
  XOR U18766 ( .A(n17111), .B(n17112), .Z(n17105) );
  AND U18767 ( .A(n17113), .B(n17114), .Z(n17111) );
  XOR U18768 ( .A(n17112), .B(n10196), .Z(n17114) );
  XNOR U18769 ( .A(n17115), .B(n17116), .Z(n10196) );
  XNOR U18770 ( .A(n[629]), .B(n17117), .Z(n17113) );
  IV U18771 ( .A(n17112), .Z(n17117) );
  XOR U18772 ( .A(n17118), .B(n17119), .Z(n17112) );
  AND U18773 ( .A(n17120), .B(n17121), .Z(n17118) );
  XOR U18774 ( .A(n17119), .B(n10201), .Z(n17121) );
  XNOR U18775 ( .A(n17122), .B(n17123), .Z(n10201) );
  XNOR U18776 ( .A(n[628]), .B(n17124), .Z(n17120) );
  IV U18777 ( .A(n17119), .Z(n17124) );
  XOR U18778 ( .A(n17125), .B(n17126), .Z(n17119) );
  AND U18779 ( .A(n17127), .B(n17128), .Z(n17125) );
  XOR U18780 ( .A(n17126), .B(n10206), .Z(n17128) );
  XNOR U18781 ( .A(n17129), .B(n17130), .Z(n10206) );
  XNOR U18782 ( .A(n[627]), .B(n17131), .Z(n17127) );
  IV U18783 ( .A(n17126), .Z(n17131) );
  XOR U18784 ( .A(n17132), .B(n17133), .Z(n17126) );
  AND U18785 ( .A(n17134), .B(n17135), .Z(n17132) );
  XOR U18786 ( .A(n17133), .B(n10211), .Z(n17135) );
  XNOR U18787 ( .A(n17136), .B(n17137), .Z(n10211) );
  XNOR U18788 ( .A(n[626]), .B(n17138), .Z(n17134) );
  IV U18789 ( .A(n17133), .Z(n17138) );
  XOR U18790 ( .A(n17139), .B(n17140), .Z(n17133) );
  AND U18791 ( .A(n17141), .B(n17142), .Z(n17139) );
  XOR U18792 ( .A(n17140), .B(n10216), .Z(n17142) );
  XNOR U18793 ( .A(n17143), .B(n17144), .Z(n10216) );
  XNOR U18794 ( .A(n[625]), .B(n17145), .Z(n17141) );
  IV U18795 ( .A(n17140), .Z(n17145) );
  XOR U18796 ( .A(n17146), .B(n17147), .Z(n17140) );
  AND U18797 ( .A(n17148), .B(n17149), .Z(n17146) );
  XOR U18798 ( .A(n17147), .B(n10221), .Z(n17149) );
  XNOR U18799 ( .A(n17150), .B(n17151), .Z(n10221) );
  XNOR U18800 ( .A(n[624]), .B(n17152), .Z(n17148) );
  IV U18801 ( .A(n17147), .Z(n17152) );
  XOR U18802 ( .A(n17153), .B(n17154), .Z(n17147) );
  AND U18803 ( .A(n17155), .B(n17156), .Z(n17153) );
  XOR U18804 ( .A(n17154), .B(n10226), .Z(n17156) );
  XNOR U18805 ( .A(n17157), .B(n17158), .Z(n10226) );
  XNOR U18806 ( .A(n[623]), .B(n17159), .Z(n17155) );
  IV U18807 ( .A(n17154), .Z(n17159) );
  XOR U18808 ( .A(n17160), .B(n17161), .Z(n17154) );
  AND U18809 ( .A(n17162), .B(n17163), .Z(n17160) );
  XOR U18810 ( .A(n17161), .B(n10231), .Z(n17163) );
  XNOR U18811 ( .A(n17164), .B(n17165), .Z(n10231) );
  XNOR U18812 ( .A(n[622]), .B(n17166), .Z(n17162) );
  IV U18813 ( .A(n17161), .Z(n17166) );
  XOR U18814 ( .A(n17167), .B(n17168), .Z(n17161) );
  AND U18815 ( .A(n17169), .B(n17170), .Z(n17167) );
  XOR U18816 ( .A(n17168), .B(n10236), .Z(n17170) );
  XNOR U18817 ( .A(n17171), .B(n17172), .Z(n10236) );
  XNOR U18818 ( .A(n[621]), .B(n17173), .Z(n17169) );
  IV U18819 ( .A(n17168), .Z(n17173) );
  XOR U18820 ( .A(n17174), .B(n17175), .Z(n17168) );
  AND U18821 ( .A(n17176), .B(n17177), .Z(n17174) );
  XOR U18822 ( .A(n17175), .B(n10241), .Z(n17177) );
  XNOR U18823 ( .A(n17178), .B(n17179), .Z(n10241) );
  XNOR U18824 ( .A(n[620]), .B(n17180), .Z(n17176) );
  IV U18825 ( .A(n17175), .Z(n17180) );
  XOR U18826 ( .A(n17181), .B(n17182), .Z(n17175) );
  AND U18827 ( .A(n17183), .B(n17184), .Z(n17181) );
  XOR U18828 ( .A(n17182), .B(n10246), .Z(n17184) );
  XNOR U18829 ( .A(n17185), .B(n17186), .Z(n10246) );
  XNOR U18830 ( .A(n[619]), .B(n17187), .Z(n17183) );
  IV U18831 ( .A(n17182), .Z(n17187) );
  XOR U18832 ( .A(n17188), .B(n17189), .Z(n17182) );
  AND U18833 ( .A(n17190), .B(n17191), .Z(n17188) );
  XOR U18834 ( .A(n17189), .B(n10251), .Z(n17191) );
  XNOR U18835 ( .A(n17192), .B(n17193), .Z(n10251) );
  XNOR U18836 ( .A(n[618]), .B(n17194), .Z(n17190) );
  IV U18837 ( .A(n17189), .Z(n17194) );
  XOR U18838 ( .A(n17195), .B(n17196), .Z(n17189) );
  AND U18839 ( .A(n17197), .B(n17198), .Z(n17195) );
  XOR U18840 ( .A(n17196), .B(n10256), .Z(n17198) );
  XNOR U18841 ( .A(n17199), .B(n17200), .Z(n10256) );
  XNOR U18842 ( .A(n[617]), .B(n17201), .Z(n17197) );
  IV U18843 ( .A(n17196), .Z(n17201) );
  XOR U18844 ( .A(n17202), .B(n17203), .Z(n17196) );
  AND U18845 ( .A(n17204), .B(n17205), .Z(n17202) );
  XOR U18846 ( .A(n17203), .B(n10261), .Z(n17205) );
  XNOR U18847 ( .A(n17206), .B(n17207), .Z(n10261) );
  XNOR U18848 ( .A(n[616]), .B(n17208), .Z(n17204) );
  IV U18849 ( .A(n17203), .Z(n17208) );
  XOR U18850 ( .A(n17209), .B(n17210), .Z(n17203) );
  AND U18851 ( .A(n17211), .B(n17212), .Z(n17209) );
  XOR U18852 ( .A(n17210), .B(n10266), .Z(n17212) );
  XNOR U18853 ( .A(n17213), .B(n17214), .Z(n10266) );
  XNOR U18854 ( .A(n[615]), .B(n17215), .Z(n17211) );
  IV U18855 ( .A(n17210), .Z(n17215) );
  XOR U18856 ( .A(n17216), .B(n17217), .Z(n17210) );
  AND U18857 ( .A(n17218), .B(n17219), .Z(n17216) );
  XOR U18858 ( .A(n17217), .B(n10271), .Z(n17219) );
  XNOR U18859 ( .A(n17220), .B(n17221), .Z(n10271) );
  XNOR U18860 ( .A(n[614]), .B(n17222), .Z(n17218) );
  IV U18861 ( .A(n17217), .Z(n17222) );
  XOR U18862 ( .A(n17223), .B(n17224), .Z(n17217) );
  AND U18863 ( .A(n17225), .B(n17226), .Z(n17223) );
  XOR U18864 ( .A(n17224), .B(n10276), .Z(n17226) );
  XNOR U18865 ( .A(n17227), .B(n17228), .Z(n10276) );
  XNOR U18866 ( .A(n[613]), .B(n17229), .Z(n17225) );
  IV U18867 ( .A(n17224), .Z(n17229) );
  XOR U18868 ( .A(n17230), .B(n17231), .Z(n17224) );
  AND U18869 ( .A(n17232), .B(n17233), .Z(n17230) );
  XOR U18870 ( .A(n17231), .B(n10281), .Z(n17233) );
  XNOR U18871 ( .A(n17234), .B(n17235), .Z(n10281) );
  XNOR U18872 ( .A(n[612]), .B(n17236), .Z(n17232) );
  IV U18873 ( .A(n17231), .Z(n17236) );
  XOR U18874 ( .A(n17237), .B(n17238), .Z(n17231) );
  AND U18875 ( .A(n17239), .B(n17240), .Z(n17237) );
  XOR U18876 ( .A(n17238), .B(n10286), .Z(n17240) );
  XNOR U18877 ( .A(n17241), .B(n17242), .Z(n10286) );
  XNOR U18878 ( .A(n[611]), .B(n17243), .Z(n17239) );
  IV U18879 ( .A(n17238), .Z(n17243) );
  XOR U18880 ( .A(n17244), .B(n17245), .Z(n17238) );
  AND U18881 ( .A(n17246), .B(n17247), .Z(n17244) );
  XOR U18882 ( .A(n17245), .B(n10291), .Z(n17247) );
  XNOR U18883 ( .A(n17248), .B(n17249), .Z(n10291) );
  XNOR U18884 ( .A(n[610]), .B(n17250), .Z(n17246) );
  IV U18885 ( .A(n17245), .Z(n17250) );
  XOR U18886 ( .A(n17251), .B(n17252), .Z(n17245) );
  AND U18887 ( .A(n17253), .B(n17254), .Z(n17251) );
  XOR U18888 ( .A(n17252), .B(n10296), .Z(n17254) );
  XNOR U18889 ( .A(n17255), .B(n17256), .Z(n10296) );
  XNOR U18890 ( .A(n[609]), .B(n17257), .Z(n17253) );
  IV U18891 ( .A(n17252), .Z(n17257) );
  XOR U18892 ( .A(n17258), .B(n17259), .Z(n17252) );
  AND U18893 ( .A(n17260), .B(n17261), .Z(n17258) );
  XOR U18894 ( .A(n17259), .B(n10301), .Z(n17261) );
  XNOR U18895 ( .A(n17262), .B(n17263), .Z(n10301) );
  XNOR U18896 ( .A(n[608]), .B(n17264), .Z(n17260) );
  IV U18897 ( .A(n17259), .Z(n17264) );
  XOR U18898 ( .A(n17265), .B(n17266), .Z(n17259) );
  AND U18899 ( .A(n17267), .B(n17268), .Z(n17265) );
  XOR U18900 ( .A(n17266), .B(n10306), .Z(n17268) );
  XNOR U18901 ( .A(n17269), .B(n17270), .Z(n10306) );
  XNOR U18902 ( .A(n[607]), .B(n17271), .Z(n17267) );
  IV U18903 ( .A(n17266), .Z(n17271) );
  XOR U18904 ( .A(n17272), .B(n17273), .Z(n17266) );
  AND U18905 ( .A(n17274), .B(n17275), .Z(n17272) );
  XOR U18906 ( .A(n17273), .B(n10311), .Z(n17275) );
  XNOR U18907 ( .A(n17276), .B(n17277), .Z(n10311) );
  XNOR U18908 ( .A(n[606]), .B(n17278), .Z(n17274) );
  IV U18909 ( .A(n17273), .Z(n17278) );
  XOR U18910 ( .A(n17279), .B(n17280), .Z(n17273) );
  AND U18911 ( .A(n17281), .B(n17282), .Z(n17279) );
  XOR U18912 ( .A(n17280), .B(n10316), .Z(n17282) );
  XNOR U18913 ( .A(n17283), .B(n17284), .Z(n10316) );
  XNOR U18914 ( .A(n[605]), .B(n17285), .Z(n17281) );
  IV U18915 ( .A(n17280), .Z(n17285) );
  XOR U18916 ( .A(n17286), .B(n17287), .Z(n17280) );
  AND U18917 ( .A(n17288), .B(n17289), .Z(n17286) );
  XOR U18918 ( .A(n17287), .B(n10321), .Z(n17289) );
  XNOR U18919 ( .A(n17290), .B(n17291), .Z(n10321) );
  XNOR U18920 ( .A(n[604]), .B(n17292), .Z(n17288) );
  IV U18921 ( .A(n17287), .Z(n17292) );
  XOR U18922 ( .A(n17293), .B(n17294), .Z(n17287) );
  AND U18923 ( .A(n17295), .B(n17296), .Z(n17293) );
  XOR U18924 ( .A(n17294), .B(n10326), .Z(n17296) );
  XNOR U18925 ( .A(n17297), .B(n17298), .Z(n10326) );
  XNOR U18926 ( .A(n[603]), .B(n17299), .Z(n17295) );
  IV U18927 ( .A(n17294), .Z(n17299) );
  XOR U18928 ( .A(n17300), .B(n17301), .Z(n17294) );
  AND U18929 ( .A(n17302), .B(n17303), .Z(n17300) );
  XOR U18930 ( .A(n17301), .B(n10331), .Z(n17303) );
  XNOR U18931 ( .A(n17304), .B(n17305), .Z(n10331) );
  XNOR U18932 ( .A(n[602]), .B(n17306), .Z(n17302) );
  IV U18933 ( .A(n17301), .Z(n17306) );
  XOR U18934 ( .A(n17307), .B(n17308), .Z(n17301) );
  AND U18935 ( .A(n17309), .B(n17310), .Z(n17307) );
  XOR U18936 ( .A(n17308), .B(n10336), .Z(n17310) );
  XNOR U18937 ( .A(n17311), .B(n17312), .Z(n10336) );
  XNOR U18938 ( .A(n[601]), .B(n17313), .Z(n17309) );
  IV U18939 ( .A(n17308), .Z(n17313) );
  XOR U18940 ( .A(n17314), .B(n17315), .Z(n17308) );
  AND U18941 ( .A(n17316), .B(n17317), .Z(n17314) );
  XOR U18942 ( .A(n17315), .B(n10341), .Z(n17317) );
  XNOR U18943 ( .A(n17318), .B(n17319), .Z(n10341) );
  XNOR U18944 ( .A(n[600]), .B(n17320), .Z(n17316) );
  IV U18945 ( .A(n17315), .Z(n17320) );
  XOR U18946 ( .A(n17321), .B(n17322), .Z(n17315) );
  AND U18947 ( .A(n17323), .B(n17324), .Z(n17321) );
  XOR U18948 ( .A(n17322), .B(n10346), .Z(n17324) );
  XNOR U18949 ( .A(n17325), .B(n17326), .Z(n10346) );
  XNOR U18950 ( .A(n[599]), .B(n17327), .Z(n17323) );
  IV U18951 ( .A(n17322), .Z(n17327) );
  XOR U18952 ( .A(n17328), .B(n17329), .Z(n17322) );
  AND U18953 ( .A(n17330), .B(n17331), .Z(n17328) );
  XOR U18954 ( .A(n17329), .B(n10351), .Z(n17331) );
  XNOR U18955 ( .A(n17332), .B(n17333), .Z(n10351) );
  XNOR U18956 ( .A(n[598]), .B(n17334), .Z(n17330) );
  IV U18957 ( .A(n17329), .Z(n17334) );
  XOR U18958 ( .A(n17335), .B(n17336), .Z(n17329) );
  AND U18959 ( .A(n17337), .B(n17338), .Z(n17335) );
  XOR U18960 ( .A(n17336), .B(n10356), .Z(n17338) );
  XNOR U18961 ( .A(n17339), .B(n17340), .Z(n10356) );
  XNOR U18962 ( .A(n[597]), .B(n17341), .Z(n17337) );
  IV U18963 ( .A(n17336), .Z(n17341) );
  XOR U18964 ( .A(n17342), .B(n17343), .Z(n17336) );
  AND U18965 ( .A(n17344), .B(n17345), .Z(n17342) );
  XOR U18966 ( .A(n17343), .B(n10361), .Z(n17345) );
  XNOR U18967 ( .A(n17346), .B(n17347), .Z(n10361) );
  XNOR U18968 ( .A(n[596]), .B(n17348), .Z(n17344) );
  IV U18969 ( .A(n17343), .Z(n17348) );
  XOR U18970 ( .A(n17349), .B(n17350), .Z(n17343) );
  AND U18971 ( .A(n17351), .B(n17352), .Z(n17349) );
  XOR U18972 ( .A(n17350), .B(n10366), .Z(n17352) );
  XNOR U18973 ( .A(n17353), .B(n17354), .Z(n10366) );
  XNOR U18974 ( .A(n[595]), .B(n17355), .Z(n17351) );
  IV U18975 ( .A(n17350), .Z(n17355) );
  XOR U18976 ( .A(n17356), .B(n17357), .Z(n17350) );
  AND U18977 ( .A(n17358), .B(n17359), .Z(n17356) );
  XOR U18978 ( .A(n17357), .B(n10371), .Z(n17359) );
  XNOR U18979 ( .A(n17360), .B(n17361), .Z(n10371) );
  XNOR U18980 ( .A(n[594]), .B(n17362), .Z(n17358) );
  IV U18981 ( .A(n17357), .Z(n17362) );
  XOR U18982 ( .A(n17363), .B(n17364), .Z(n17357) );
  AND U18983 ( .A(n17365), .B(n17366), .Z(n17363) );
  XOR U18984 ( .A(n17364), .B(n10376), .Z(n17366) );
  XNOR U18985 ( .A(n17367), .B(n17368), .Z(n10376) );
  XNOR U18986 ( .A(n[593]), .B(n17369), .Z(n17365) );
  IV U18987 ( .A(n17364), .Z(n17369) );
  XOR U18988 ( .A(n17370), .B(n17371), .Z(n17364) );
  AND U18989 ( .A(n17372), .B(n17373), .Z(n17370) );
  XOR U18990 ( .A(n17371), .B(n10381), .Z(n17373) );
  XNOR U18991 ( .A(n17374), .B(n17375), .Z(n10381) );
  XNOR U18992 ( .A(n[592]), .B(n17376), .Z(n17372) );
  IV U18993 ( .A(n17371), .Z(n17376) );
  XOR U18994 ( .A(n17377), .B(n17378), .Z(n17371) );
  AND U18995 ( .A(n17379), .B(n17380), .Z(n17377) );
  XOR U18996 ( .A(n17378), .B(n10386), .Z(n17380) );
  XNOR U18997 ( .A(n17381), .B(n17382), .Z(n10386) );
  XNOR U18998 ( .A(n[591]), .B(n17383), .Z(n17379) );
  IV U18999 ( .A(n17378), .Z(n17383) );
  XOR U19000 ( .A(n17384), .B(n17385), .Z(n17378) );
  AND U19001 ( .A(n17386), .B(n17387), .Z(n17384) );
  XOR U19002 ( .A(n17385), .B(n10391), .Z(n17387) );
  XNOR U19003 ( .A(n17388), .B(n17389), .Z(n10391) );
  XNOR U19004 ( .A(n[590]), .B(n17390), .Z(n17386) );
  IV U19005 ( .A(n17385), .Z(n17390) );
  XOR U19006 ( .A(n17391), .B(n17392), .Z(n17385) );
  AND U19007 ( .A(n17393), .B(n17394), .Z(n17391) );
  XOR U19008 ( .A(n17392), .B(n10396), .Z(n17394) );
  XNOR U19009 ( .A(n17395), .B(n17396), .Z(n10396) );
  XNOR U19010 ( .A(n[589]), .B(n17397), .Z(n17393) );
  IV U19011 ( .A(n17392), .Z(n17397) );
  XOR U19012 ( .A(n17398), .B(n17399), .Z(n17392) );
  AND U19013 ( .A(n17400), .B(n17401), .Z(n17398) );
  XOR U19014 ( .A(n17399), .B(n10401), .Z(n17401) );
  XNOR U19015 ( .A(n17402), .B(n17403), .Z(n10401) );
  XNOR U19016 ( .A(n[588]), .B(n17404), .Z(n17400) );
  IV U19017 ( .A(n17399), .Z(n17404) );
  XOR U19018 ( .A(n17405), .B(n17406), .Z(n17399) );
  AND U19019 ( .A(n17407), .B(n17408), .Z(n17405) );
  XOR U19020 ( .A(n17406), .B(n10406), .Z(n17408) );
  XNOR U19021 ( .A(n17409), .B(n17410), .Z(n10406) );
  XNOR U19022 ( .A(n[587]), .B(n17411), .Z(n17407) );
  IV U19023 ( .A(n17406), .Z(n17411) );
  XOR U19024 ( .A(n17412), .B(n17413), .Z(n17406) );
  AND U19025 ( .A(n17414), .B(n17415), .Z(n17412) );
  XOR U19026 ( .A(n17413), .B(n10411), .Z(n17415) );
  XNOR U19027 ( .A(n17416), .B(n17417), .Z(n10411) );
  XNOR U19028 ( .A(n[586]), .B(n17418), .Z(n17414) );
  IV U19029 ( .A(n17413), .Z(n17418) );
  XOR U19030 ( .A(n17419), .B(n17420), .Z(n17413) );
  AND U19031 ( .A(n17421), .B(n17422), .Z(n17419) );
  XOR U19032 ( .A(n17420), .B(n10416), .Z(n17422) );
  XNOR U19033 ( .A(n17423), .B(n17424), .Z(n10416) );
  XNOR U19034 ( .A(n[585]), .B(n17425), .Z(n17421) );
  IV U19035 ( .A(n17420), .Z(n17425) );
  XOR U19036 ( .A(n17426), .B(n17427), .Z(n17420) );
  AND U19037 ( .A(n17428), .B(n17429), .Z(n17426) );
  XOR U19038 ( .A(n17427), .B(n10421), .Z(n17429) );
  XNOR U19039 ( .A(n17430), .B(n17431), .Z(n10421) );
  XNOR U19040 ( .A(n[584]), .B(n17432), .Z(n17428) );
  IV U19041 ( .A(n17427), .Z(n17432) );
  XOR U19042 ( .A(n17433), .B(n17434), .Z(n17427) );
  AND U19043 ( .A(n17435), .B(n17436), .Z(n17433) );
  XOR U19044 ( .A(n17434), .B(n10426), .Z(n17436) );
  XNOR U19045 ( .A(n17437), .B(n17438), .Z(n10426) );
  XNOR U19046 ( .A(n[583]), .B(n17439), .Z(n17435) );
  IV U19047 ( .A(n17434), .Z(n17439) );
  XOR U19048 ( .A(n17440), .B(n17441), .Z(n17434) );
  AND U19049 ( .A(n17442), .B(n17443), .Z(n17440) );
  XOR U19050 ( .A(n17441), .B(n10431), .Z(n17443) );
  XNOR U19051 ( .A(n17444), .B(n17445), .Z(n10431) );
  XNOR U19052 ( .A(n[582]), .B(n17446), .Z(n17442) );
  IV U19053 ( .A(n17441), .Z(n17446) );
  XOR U19054 ( .A(n17447), .B(n17448), .Z(n17441) );
  AND U19055 ( .A(n17449), .B(n17450), .Z(n17447) );
  XOR U19056 ( .A(n17448), .B(n10436), .Z(n17450) );
  XNOR U19057 ( .A(n17451), .B(n17452), .Z(n10436) );
  XNOR U19058 ( .A(n[581]), .B(n17453), .Z(n17449) );
  IV U19059 ( .A(n17448), .Z(n17453) );
  XOR U19060 ( .A(n17454), .B(n17455), .Z(n17448) );
  AND U19061 ( .A(n17456), .B(n17457), .Z(n17454) );
  XOR U19062 ( .A(n17455), .B(n10441), .Z(n17457) );
  XNOR U19063 ( .A(n17458), .B(n17459), .Z(n10441) );
  XNOR U19064 ( .A(n[580]), .B(n17460), .Z(n17456) );
  IV U19065 ( .A(n17455), .Z(n17460) );
  XOR U19066 ( .A(n17461), .B(n17462), .Z(n17455) );
  AND U19067 ( .A(n17463), .B(n17464), .Z(n17461) );
  XOR U19068 ( .A(n17462), .B(n10446), .Z(n17464) );
  XNOR U19069 ( .A(n17465), .B(n17466), .Z(n10446) );
  XNOR U19070 ( .A(n[579]), .B(n17467), .Z(n17463) );
  IV U19071 ( .A(n17462), .Z(n17467) );
  XOR U19072 ( .A(n17468), .B(n17469), .Z(n17462) );
  AND U19073 ( .A(n17470), .B(n17471), .Z(n17468) );
  XOR U19074 ( .A(n17469), .B(n10451), .Z(n17471) );
  XNOR U19075 ( .A(n17472), .B(n17473), .Z(n10451) );
  XNOR U19076 ( .A(n[578]), .B(n17474), .Z(n17470) );
  IV U19077 ( .A(n17469), .Z(n17474) );
  XOR U19078 ( .A(n17475), .B(n17476), .Z(n17469) );
  AND U19079 ( .A(n17477), .B(n17478), .Z(n17475) );
  XOR U19080 ( .A(n17476), .B(n10456), .Z(n17478) );
  XNOR U19081 ( .A(n17479), .B(n17480), .Z(n10456) );
  XNOR U19082 ( .A(n[577]), .B(n17481), .Z(n17477) );
  IV U19083 ( .A(n17476), .Z(n17481) );
  XOR U19084 ( .A(n17482), .B(n17483), .Z(n17476) );
  AND U19085 ( .A(n17484), .B(n17485), .Z(n17482) );
  XOR U19086 ( .A(n17483), .B(n10461), .Z(n17485) );
  XNOR U19087 ( .A(n17486), .B(n17487), .Z(n10461) );
  XNOR U19088 ( .A(n[576]), .B(n17488), .Z(n17484) );
  IV U19089 ( .A(n17483), .Z(n17488) );
  XOR U19090 ( .A(n17489), .B(n17490), .Z(n17483) );
  AND U19091 ( .A(n17491), .B(n17492), .Z(n17489) );
  XOR U19092 ( .A(n17490), .B(n10466), .Z(n17492) );
  XNOR U19093 ( .A(n17493), .B(n17494), .Z(n10466) );
  XNOR U19094 ( .A(n[575]), .B(n17495), .Z(n17491) );
  IV U19095 ( .A(n17490), .Z(n17495) );
  XOR U19096 ( .A(n17496), .B(n17497), .Z(n17490) );
  AND U19097 ( .A(n17498), .B(n17499), .Z(n17496) );
  XOR U19098 ( .A(n17497), .B(n10471), .Z(n17499) );
  XNOR U19099 ( .A(n17500), .B(n17501), .Z(n10471) );
  XNOR U19100 ( .A(n[574]), .B(n17502), .Z(n17498) );
  IV U19101 ( .A(n17497), .Z(n17502) );
  XOR U19102 ( .A(n17503), .B(n17504), .Z(n17497) );
  AND U19103 ( .A(n17505), .B(n17506), .Z(n17503) );
  XOR U19104 ( .A(n17504), .B(n10476), .Z(n17506) );
  XNOR U19105 ( .A(n17507), .B(n17508), .Z(n10476) );
  XNOR U19106 ( .A(n[573]), .B(n17509), .Z(n17505) );
  IV U19107 ( .A(n17504), .Z(n17509) );
  XOR U19108 ( .A(n17510), .B(n17511), .Z(n17504) );
  AND U19109 ( .A(n17512), .B(n17513), .Z(n17510) );
  XOR U19110 ( .A(n17511), .B(n10481), .Z(n17513) );
  XNOR U19111 ( .A(n17514), .B(n17515), .Z(n10481) );
  XNOR U19112 ( .A(n[572]), .B(n17516), .Z(n17512) );
  IV U19113 ( .A(n17511), .Z(n17516) );
  XOR U19114 ( .A(n17517), .B(n17518), .Z(n17511) );
  AND U19115 ( .A(n17519), .B(n17520), .Z(n17517) );
  XOR U19116 ( .A(n17518), .B(n10486), .Z(n17520) );
  XNOR U19117 ( .A(n17521), .B(n17522), .Z(n10486) );
  XNOR U19118 ( .A(n[571]), .B(n17523), .Z(n17519) );
  IV U19119 ( .A(n17518), .Z(n17523) );
  XOR U19120 ( .A(n17524), .B(n17525), .Z(n17518) );
  AND U19121 ( .A(n17526), .B(n17527), .Z(n17524) );
  XOR U19122 ( .A(n17525), .B(n10491), .Z(n17527) );
  XNOR U19123 ( .A(n17528), .B(n17529), .Z(n10491) );
  XNOR U19124 ( .A(n[570]), .B(n17530), .Z(n17526) );
  IV U19125 ( .A(n17525), .Z(n17530) );
  XOR U19126 ( .A(n17531), .B(n17532), .Z(n17525) );
  AND U19127 ( .A(n17533), .B(n17534), .Z(n17531) );
  XOR U19128 ( .A(n17532), .B(n10496), .Z(n17534) );
  XNOR U19129 ( .A(n17535), .B(n17536), .Z(n10496) );
  XNOR U19130 ( .A(n[569]), .B(n17537), .Z(n17533) );
  IV U19131 ( .A(n17532), .Z(n17537) );
  XOR U19132 ( .A(n17538), .B(n17539), .Z(n17532) );
  AND U19133 ( .A(n17540), .B(n17541), .Z(n17538) );
  XOR U19134 ( .A(n17539), .B(n10501), .Z(n17541) );
  XNOR U19135 ( .A(n17542), .B(n17543), .Z(n10501) );
  XNOR U19136 ( .A(n[568]), .B(n17544), .Z(n17540) );
  IV U19137 ( .A(n17539), .Z(n17544) );
  XOR U19138 ( .A(n17545), .B(n17546), .Z(n17539) );
  AND U19139 ( .A(n17547), .B(n17548), .Z(n17545) );
  XOR U19140 ( .A(n17546), .B(n10506), .Z(n17548) );
  XNOR U19141 ( .A(n17549), .B(n17550), .Z(n10506) );
  XNOR U19142 ( .A(n[567]), .B(n17551), .Z(n17547) );
  IV U19143 ( .A(n17546), .Z(n17551) );
  XOR U19144 ( .A(n17552), .B(n17553), .Z(n17546) );
  AND U19145 ( .A(n17554), .B(n17555), .Z(n17552) );
  XOR U19146 ( .A(n17553), .B(n10511), .Z(n17555) );
  XNOR U19147 ( .A(n17556), .B(n17557), .Z(n10511) );
  XNOR U19148 ( .A(n[566]), .B(n17558), .Z(n17554) );
  IV U19149 ( .A(n17553), .Z(n17558) );
  XOR U19150 ( .A(n17559), .B(n17560), .Z(n17553) );
  AND U19151 ( .A(n17561), .B(n17562), .Z(n17559) );
  XOR U19152 ( .A(n17560), .B(n10516), .Z(n17562) );
  XNOR U19153 ( .A(n17563), .B(n17564), .Z(n10516) );
  XNOR U19154 ( .A(n[565]), .B(n17565), .Z(n17561) );
  IV U19155 ( .A(n17560), .Z(n17565) );
  XOR U19156 ( .A(n17566), .B(n17567), .Z(n17560) );
  AND U19157 ( .A(n17568), .B(n17569), .Z(n17566) );
  XOR U19158 ( .A(n17567), .B(n10521), .Z(n17569) );
  XNOR U19159 ( .A(n17570), .B(n17571), .Z(n10521) );
  XNOR U19160 ( .A(n[564]), .B(n17572), .Z(n17568) );
  IV U19161 ( .A(n17567), .Z(n17572) );
  XOR U19162 ( .A(n17573), .B(n17574), .Z(n17567) );
  AND U19163 ( .A(n17575), .B(n17576), .Z(n17573) );
  XOR U19164 ( .A(n17574), .B(n10526), .Z(n17576) );
  XNOR U19165 ( .A(n17577), .B(n17578), .Z(n10526) );
  XNOR U19166 ( .A(n[563]), .B(n17579), .Z(n17575) );
  IV U19167 ( .A(n17574), .Z(n17579) );
  XOR U19168 ( .A(n17580), .B(n17581), .Z(n17574) );
  AND U19169 ( .A(n17582), .B(n17583), .Z(n17580) );
  XOR U19170 ( .A(n17581), .B(n10531), .Z(n17583) );
  XNOR U19171 ( .A(n17584), .B(n17585), .Z(n10531) );
  XNOR U19172 ( .A(n[562]), .B(n17586), .Z(n17582) );
  IV U19173 ( .A(n17581), .Z(n17586) );
  XOR U19174 ( .A(n17587), .B(n17588), .Z(n17581) );
  AND U19175 ( .A(n17589), .B(n17590), .Z(n17587) );
  XOR U19176 ( .A(n17588), .B(n10536), .Z(n17590) );
  XNOR U19177 ( .A(n17591), .B(n17592), .Z(n10536) );
  XNOR U19178 ( .A(n[561]), .B(n17593), .Z(n17589) );
  IV U19179 ( .A(n17588), .Z(n17593) );
  XOR U19180 ( .A(n17594), .B(n17595), .Z(n17588) );
  AND U19181 ( .A(n17596), .B(n17597), .Z(n17594) );
  XOR U19182 ( .A(n17595), .B(n10541), .Z(n17597) );
  XNOR U19183 ( .A(n17598), .B(n17599), .Z(n10541) );
  XNOR U19184 ( .A(n[560]), .B(n17600), .Z(n17596) );
  IV U19185 ( .A(n17595), .Z(n17600) );
  XOR U19186 ( .A(n17601), .B(n17602), .Z(n17595) );
  AND U19187 ( .A(n17603), .B(n17604), .Z(n17601) );
  XOR U19188 ( .A(n17602), .B(n10546), .Z(n17604) );
  XNOR U19189 ( .A(n17605), .B(n17606), .Z(n10546) );
  XNOR U19190 ( .A(n[559]), .B(n17607), .Z(n17603) );
  IV U19191 ( .A(n17602), .Z(n17607) );
  XOR U19192 ( .A(n17608), .B(n17609), .Z(n17602) );
  AND U19193 ( .A(n17610), .B(n17611), .Z(n17608) );
  XOR U19194 ( .A(n17609), .B(n10551), .Z(n17611) );
  XNOR U19195 ( .A(n17612), .B(n17613), .Z(n10551) );
  XNOR U19196 ( .A(n[558]), .B(n17614), .Z(n17610) );
  IV U19197 ( .A(n17609), .Z(n17614) );
  XOR U19198 ( .A(n17615), .B(n17616), .Z(n17609) );
  AND U19199 ( .A(n17617), .B(n17618), .Z(n17615) );
  XOR U19200 ( .A(n17616), .B(n10556), .Z(n17618) );
  XNOR U19201 ( .A(n17619), .B(n17620), .Z(n10556) );
  XNOR U19202 ( .A(n[557]), .B(n17621), .Z(n17617) );
  IV U19203 ( .A(n17616), .Z(n17621) );
  XOR U19204 ( .A(n17622), .B(n17623), .Z(n17616) );
  AND U19205 ( .A(n17624), .B(n17625), .Z(n17622) );
  XOR U19206 ( .A(n17623), .B(n10561), .Z(n17625) );
  XNOR U19207 ( .A(n17626), .B(n17627), .Z(n10561) );
  XNOR U19208 ( .A(n[556]), .B(n17628), .Z(n17624) );
  IV U19209 ( .A(n17623), .Z(n17628) );
  XOR U19210 ( .A(n17629), .B(n17630), .Z(n17623) );
  AND U19211 ( .A(n17631), .B(n17632), .Z(n17629) );
  XOR U19212 ( .A(n17630), .B(n10566), .Z(n17632) );
  XNOR U19213 ( .A(n17633), .B(n17634), .Z(n10566) );
  XNOR U19214 ( .A(n[555]), .B(n17635), .Z(n17631) );
  IV U19215 ( .A(n17630), .Z(n17635) );
  XOR U19216 ( .A(n17636), .B(n17637), .Z(n17630) );
  AND U19217 ( .A(n17638), .B(n17639), .Z(n17636) );
  XOR U19218 ( .A(n17637), .B(n10571), .Z(n17639) );
  XNOR U19219 ( .A(n17640), .B(n17641), .Z(n10571) );
  XNOR U19220 ( .A(n[554]), .B(n17642), .Z(n17638) );
  IV U19221 ( .A(n17637), .Z(n17642) );
  XOR U19222 ( .A(n17643), .B(n17644), .Z(n17637) );
  AND U19223 ( .A(n17645), .B(n17646), .Z(n17643) );
  XOR U19224 ( .A(n17644), .B(n10576), .Z(n17646) );
  XNOR U19225 ( .A(n17647), .B(n17648), .Z(n10576) );
  XNOR U19226 ( .A(n[553]), .B(n17649), .Z(n17645) );
  IV U19227 ( .A(n17644), .Z(n17649) );
  XOR U19228 ( .A(n17650), .B(n17651), .Z(n17644) );
  AND U19229 ( .A(n17652), .B(n17653), .Z(n17650) );
  XOR U19230 ( .A(n17651), .B(n10581), .Z(n17653) );
  XNOR U19231 ( .A(n17654), .B(n17655), .Z(n10581) );
  XNOR U19232 ( .A(n[552]), .B(n17656), .Z(n17652) );
  IV U19233 ( .A(n17651), .Z(n17656) );
  XOR U19234 ( .A(n17657), .B(n17658), .Z(n17651) );
  AND U19235 ( .A(n17659), .B(n17660), .Z(n17657) );
  XOR U19236 ( .A(n17658), .B(n10586), .Z(n17660) );
  XNOR U19237 ( .A(n17661), .B(n17662), .Z(n10586) );
  XNOR U19238 ( .A(n[551]), .B(n17663), .Z(n17659) );
  IV U19239 ( .A(n17658), .Z(n17663) );
  XOR U19240 ( .A(n17664), .B(n17665), .Z(n17658) );
  AND U19241 ( .A(n17666), .B(n17667), .Z(n17664) );
  XOR U19242 ( .A(n17665), .B(n10591), .Z(n17667) );
  XNOR U19243 ( .A(n17668), .B(n17669), .Z(n10591) );
  XNOR U19244 ( .A(n[550]), .B(n17670), .Z(n17666) );
  IV U19245 ( .A(n17665), .Z(n17670) );
  XOR U19246 ( .A(n17671), .B(n17672), .Z(n17665) );
  AND U19247 ( .A(n17673), .B(n17674), .Z(n17671) );
  XOR U19248 ( .A(n17672), .B(n10596), .Z(n17674) );
  XNOR U19249 ( .A(n17675), .B(n17676), .Z(n10596) );
  XNOR U19250 ( .A(n[549]), .B(n17677), .Z(n17673) );
  IV U19251 ( .A(n17672), .Z(n17677) );
  XOR U19252 ( .A(n17678), .B(n17679), .Z(n17672) );
  AND U19253 ( .A(n17680), .B(n17681), .Z(n17678) );
  XOR U19254 ( .A(n17679), .B(n10601), .Z(n17681) );
  XNOR U19255 ( .A(n17682), .B(n17683), .Z(n10601) );
  XNOR U19256 ( .A(n[548]), .B(n17684), .Z(n17680) );
  IV U19257 ( .A(n17679), .Z(n17684) );
  XOR U19258 ( .A(n17685), .B(n17686), .Z(n17679) );
  AND U19259 ( .A(n17687), .B(n17688), .Z(n17685) );
  XOR U19260 ( .A(n17686), .B(n10606), .Z(n17688) );
  XNOR U19261 ( .A(n17689), .B(n17690), .Z(n10606) );
  XNOR U19262 ( .A(n[547]), .B(n17691), .Z(n17687) );
  IV U19263 ( .A(n17686), .Z(n17691) );
  XOR U19264 ( .A(n17692), .B(n17693), .Z(n17686) );
  AND U19265 ( .A(n17694), .B(n17695), .Z(n17692) );
  XOR U19266 ( .A(n17693), .B(n10611), .Z(n17695) );
  XNOR U19267 ( .A(n17696), .B(n17697), .Z(n10611) );
  XNOR U19268 ( .A(n[546]), .B(n17698), .Z(n17694) );
  IV U19269 ( .A(n17693), .Z(n17698) );
  XOR U19270 ( .A(n17699), .B(n17700), .Z(n17693) );
  AND U19271 ( .A(n17701), .B(n17702), .Z(n17699) );
  XOR U19272 ( .A(n17700), .B(n10616), .Z(n17702) );
  XNOR U19273 ( .A(n17703), .B(n17704), .Z(n10616) );
  XNOR U19274 ( .A(n[545]), .B(n17705), .Z(n17701) );
  IV U19275 ( .A(n17700), .Z(n17705) );
  XOR U19276 ( .A(n17706), .B(n17707), .Z(n17700) );
  AND U19277 ( .A(n17708), .B(n17709), .Z(n17706) );
  XOR U19278 ( .A(n17707), .B(n10621), .Z(n17709) );
  XNOR U19279 ( .A(n17710), .B(n17711), .Z(n10621) );
  XNOR U19280 ( .A(n[544]), .B(n17712), .Z(n17708) );
  IV U19281 ( .A(n17707), .Z(n17712) );
  XOR U19282 ( .A(n17713), .B(n17714), .Z(n17707) );
  AND U19283 ( .A(n17715), .B(n17716), .Z(n17713) );
  XOR U19284 ( .A(n17714), .B(n10626), .Z(n17716) );
  XNOR U19285 ( .A(n17717), .B(n17718), .Z(n10626) );
  XNOR U19286 ( .A(n[543]), .B(n17719), .Z(n17715) );
  IV U19287 ( .A(n17714), .Z(n17719) );
  XOR U19288 ( .A(n17720), .B(n17721), .Z(n17714) );
  AND U19289 ( .A(n17722), .B(n17723), .Z(n17720) );
  XOR U19290 ( .A(n17721), .B(n10631), .Z(n17723) );
  XNOR U19291 ( .A(n17724), .B(n17725), .Z(n10631) );
  XNOR U19292 ( .A(n[542]), .B(n17726), .Z(n17722) );
  IV U19293 ( .A(n17721), .Z(n17726) );
  XOR U19294 ( .A(n17727), .B(n17728), .Z(n17721) );
  AND U19295 ( .A(n17729), .B(n17730), .Z(n17727) );
  XOR U19296 ( .A(n17728), .B(n10636), .Z(n17730) );
  XNOR U19297 ( .A(n17731), .B(n17732), .Z(n10636) );
  XNOR U19298 ( .A(n[541]), .B(n17733), .Z(n17729) );
  IV U19299 ( .A(n17728), .Z(n17733) );
  XOR U19300 ( .A(n17734), .B(n17735), .Z(n17728) );
  AND U19301 ( .A(n17736), .B(n17737), .Z(n17734) );
  XOR U19302 ( .A(n17735), .B(n10641), .Z(n17737) );
  XNOR U19303 ( .A(n17738), .B(n17739), .Z(n10641) );
  XNOR U19304 ( .A(n[540]), .B(n17740), .Z(n17736) );
  IV U19305 ( .A(n17735), .Z(n17740) );
  XOR U19306 ( .A(n17741), .B(n17742), .Z(n17735) );
  AND U19307 ( .A(n17743), .B(n17744), .Z(n17741) );
  XOR U19308 ( .A(n17742), .B(n10646), .Z(n17744) );
  XNOR U19309 ( .A(n17745), .B(n17746), .Z(n10646) );
  XNOR U19310 ( .A(n[539]), .B(n17747), .Z(n17743) );
  IV U19311 ( .A(n17742), .Z(n17747) );
  XOR U19312 ( .A(n17748), .B(n17749), .Z(n17742) );
  AND U19313 ( .A(n17750), .B(n17751), .Z(n17748) );
  XOR U19314 ( .A(n17749), .B(n10651), .Z(n17751) );
  XNOR U19315 ( .A(n17752), .B(n17753), .Z(n10651) );
  XNOR U19316 ( .A(n[538]), .B(n17754), .Z(n17750) );
  IV U19317 ( .A(n17749), .Z(n17754) );
  XOR U19318 ( .A(n17755), .B(n17756), .Z(n17749) );
  AND U19319 ( .A(n17757), .B(n17758), .Z(n17755) );
  XOR U19320 ( .A(n17756), .B(n10656), .Z(n17758) );
  XNOR U19321 ( .A(n17759), .B(n17760), .Z(n10656) );
  XNOR U19322 ( .A(n[537]), .B(n17761), .Z(n17757) );
  IV U19323 ( .A(n17756), .Z(n17761) );
  XOR U19324 ( .A(n17762), .B(n17763), .Z(n17756) );
  AND U19325 ( .A(n17764), .B(n17765), .Z(n17762) );
  XOR U19326 ( .A(n17763), .B(n10661), .Z(n17765) );
  XNOR U19327 ( .A(n17766), .B(n17767), .Z(n10661) );
  XNOR U19328 ( .A(n[536]), .B(n17768), .Z(n17764) );
  IV U19329 ( .A(n17763), .Z(n17768) );
  XOR U19330 ( .A(n17769), .B(n17770), .Z(n17763) );
  AND U19331 ( .A(n17771), .B(n17772), .Z(n17769) );
  XOR U19332 ( .A(n17770), .B(n10666), .Z(n17772) );
  XNOR U19333 ( .A(n17773), .B(n17774), .Z(n10666) );
  XNOR U19334 ( .A(n[535]), .B(n17775), .Z(n17771) );
  IV U19335 ( .A(n17770), .Z(n17775) );
  XOR U19336 ( .A(n17776), .B(n17777), .Z(n17770) );
  AND U19337 ( .A(n17778), .B(n17779), .Z(n17776) );
  XOR U19338 ( .A(n17777), .B(n10671), .Z(n17779) );
  XNOR U19339 ( .A(n17780), .B(n17781), .Z(n10671) );
  XNOR U19340 ( .A(n[534]), .B(n17782), .Z(n17778) );
  IV U19341 ( .A(n17777), .Z(n17782) );
  XOR U19342 ( .A(n17783), .B(n17784), .Z(n17777) );
  AND U19343 ( .A(n17785), .B(n17786), .Z(n17783) );
  XOR U19344 ( .A(n17784), .B(n10676), .Z(n17786) );
  XNOR U19345 ( .A(n17787), .B(n17788), .Z(n10676) );
  XNOR U19346 ( .A(n[533]), .B(n17789), .Z(n17785) );
  IV U19347 ( .A(n17784), .Z(n17789) );
  XOR U19348 ( .A(n17790), .B(n17791), .Z(n17784) );
  AND U19349 ( .A(n17792), .B(n17793), .Z(n17790) );
  XOR U19350 ( .A(n17791), .B(n10681), .Z(n17793) );
  XNOR U19351 ( .A(n17794), .B(n17795), .Z(n10681) );
  XNOR U19352 ( .A(n[532]), .B(n17796), .Z(n17792) );
  IV U19353 ( .A(n17791), .Z(n17796) );
  XOR U19354 ( .A(n17797), .B(n17798), .Z(n17791) );
  AND U19355 ( .A(n17799), .B(n17800), .Z(n17797) );
  XOR U19356 ( .A(n17798), .B(n10686), .Z(n17800) );
  XNOR U19357 ( .A(n17801), .B(n17802), .Z(n10686) );
  XNOR U19358 ( .A(n[531]), .B(n17803), .Z(n17799) );
  IV U19359 ( .A(n17798), .Z(n17803) );
  XOR U19360 ( .A(n17804), .B(n17805), .Z(n17798) );
  AND U19361 ( .A(n17806), .B(n17807), .Z(n17804) );
  XOR U19362 ( .A(n17805), .B(n10691), .Z(n17807) );
  XNOR U19363 ( .A(n17808), .B(n17809), .Z(n10691) );
  XNOR U19364 ( .A(n[530]), .B(n17810), .Z(n17806) );
  IV U19365 ( .A(n17805), .Z(n17810) );
  XOR U19366 ( .A(n17811), .B(n17812), .Z(n17805) );
  AND U19367 ( .A(n17813), .B(n17814), .Z(n17811) );
  XOR U19368 ( .A(n17812), .B(n10696), .Z(n17814) );
  XNOR U19369 ( .A(n17815), .B(n17816), .Z(n10696) );
  XNOR U19370 ( .A(n[529]), .B(n17817), .Z(n17813) );
  IV U19371 ( .A(n17812), .Z(n17817) );
  XOR U19372 ( .A(n17818), .B(n17819), .Z(n17812) );
  AND U19373 ( .A(n17820), .B(n17821), .Z(n17818) );
  XOR U19374 ( .A(n17819), .B(n10701), .Z(n17821) );
  XNOR U19375 ( .A(n17822), .B(n17823), .Z(n10701) );
  XNOR U19376 ( .A(n[528]), .B(n17824), .Z(n17820) );
  IV U19377 ( .A(n17819), .Z(n17824) );
  XOR U19378 ( .A(n17825), .B(n17826), .Z(n17819) );
  AND U19379 ( .A(n17827), .B(n17828), .Z(n17825) );
  XOR U19380 ( .A(n17826), .B(n10706), .Z(n17828) );
  XNOR U19381 ( .A(n17829), .B(n17830), .Z(n10706) );
  XNOR U19382 ( .A(n[527]), .B(n17831), .Z(n17827) );
  IV U19383 ( .A(n17826), .Z(n17831) );
  XOR U19384 ( .A(n17832), .B(n17833), .Z(n17826) );
  AND U19385 ( .A(n17834), .B(n17835), .Z(n17832) );
  XOR U19386 ( .A(n17833), .B(n10711), .Z(n17835) );
  XNOR U19387 ( .A(n17836), .B(n17837), .Z(n10711) );
  XNOR U19388 ( .A(n[526]), .B(n17838), .Z(n17834) );
  IV U19389 ( .A(n17833), .Z(n17838) );
  XOR U19390 ( .A(n17839), .B(n17840), .Z(n17833) );
  AND U19391 ( .A(n17841), .B(n17842), .Z(n17839) );
  XOR U19392 ( .A(n17840), .B(n10716), .Z(n17842) );
  XNOR U19393 ( .A(n17843), .B(n17844), .Z(n10716) );
  XNOR U19394 ( .A(n[525]), .B(n17845), .Z(n17841) );
  IV U19395 ( .A(n17840), .Z(n17845) );
  XOR U19396 ( .A(n17846), .B(n17847), .Z(n17840) );
  AND U19397 ( .A(n17848), .B(n17849), .Z(n17846) );
  XOR U19398 ( .A(n17847), .B(n10721), .Z(n17849) );
  XNOR U19399 ( .A(n17850), .B(n17851), .Z(n10721) );
  XNOR U19400 ( .A(n[524]), .B(n17852), .Z(n17848) );
  IV U19401 ( .A(n17847), .Z(n17852) );
  XOR U19402 ( .A(n17853), .B(n17854), .Z(n17847) );
  AND U19403 ( .A(n17855), .B(n17856), .Z(n17853) );
  XOR U19404 ( .A(n17854), .B(n10726), .Z(n17856) );
  XNOR U19405 ( .A(n17857), .B(n17858), .Z(n10726) );
  XNOR U19406 ( .A(n[523]), .B(n17859), .Z(n17855) );
  IV U19407 ( .A(n17854), .Z(n17859) );
  XOR U19408 ( .A(n17860), .B(n17861), .Z(n17854) );
  AND U19409 ( .A(n17862), .B(n17863), .Z(n17860) );
  XOR U19410 ( .A(n17861), .B(n10731), .Z(n17863) );
  XNOR U19411 ( .A(n17864), .B(n17865), .Z(n10731) );
  XNOR U19412 ( .A(n[522]), .B(n17866), .Z(n17862) );
  IV U19413 ( .A(n17861), .Z(n17866) );
  XOR U19414 ( .A(n17867), .B(n17868), .Z(n17861) );
  AND U19415 ( .A(n17869), .B(n17870), .Z(n17867) );
  XOR U19416 ( .A(n17868), .B(n10736), .Z(n17870) );
  XNOR U19417 ( .A(n17871), .B(n17872), .Z(n10736) );
  XNOR U19418 ( .A(n[521]), .B(n17873), .Z(n17869) );
  IV U19419 ( .A(n17868), .Z(n17873) );
  XOR U19420 ( .A(n17874), .B(n17875), .Z(n17868) );
  AND U19421 ( .A(n17876), .B(n17877), .Z(n17874) );
  XOR U19422 ( .A(n17875), .B(n10741), .Z(n17877) );
  XNOR U19423 ( .A(n17878), .B(n17879), .Z(n10741) );
  XNOR U19424 ( .A(n[520]), .B(n17880), .Z(n17876) );
  IV U19425 ( .A(n17875), .Z(n17880) );
  XOR U19426 ( .A(n17881), .B(n17882), .Z(n17875) );
  AND U19427 ( .A(n17883), .B(n17884), .Z(n17881) );
  XOR U19428 ( .A(n17882), .B(n10746), .Z(n17884) );
  XNOR U19429 ( .A(n17885), .B(n17886), .Z(n10746) );
  XNOR U19430 ( .A(n[519]), .B(n17887), .Z(n17883) );
  IV U19431 ( .A(n17882), .Z(n17887) );
  XOR U19432 ( .A(n17888), .B(n17889), .Z(n17882) );
  AND U19433 ( .A(n17890), .B(n17891), .Z(n17888) );
  XOR U19434 ( .A(n17889), .B(n10751), .Z(n17891) );
  XNOR U19435 ( .A(n17892), .B(n17893), .Z(n10751) );
  XNOR U19436 ( .A(n[518]), .B(n17894), .Z(n17890) );
  IV U19437 ( .A(n17889), .Z(n17894) );
  XOR U19438 ( .A(n17895), .B(n17896), .Z(n17889) );
  AND U19439 ( .A(n17897), .B(n17898), .Z(n17895) );
  XOR U19440 ( .A(n17896), .B(n10756), .Z(n17898) );
  XNOR U19441 ( .A(n17899), .B(n17900), .Z(n10756) );
  XNOR U19442 ( .A(n[517]), .B(n17901), .Z(n17897) );
  IV U19443 ( .A(n17896), .Z(n17901) );
  XOR U19444 ( .A(n17902), .B(n17903), .Z(n17896) );
  AND U19445 ( .A(n17904), .B(n17905), .Z(n17902) );
  XOR U19446 ( .A(n17903), .B(n10761), .Z(n17905) );
  XNOR U19447 ( .A(n17906), .B(n17907), .Z(n10761) );
  XNOR U19448 ( .A(n[516]), .B(n17908), .Z(n17904) );
  IV U19449 ( .A(n17903), .Z(n17908) );
  XOR U19450 ( .A(n17909), .B(n17910), .Z(n17903) );
  AND U19451 ( .A(n17911), .B(n17912), .Z(n17909) );
  XOR U19452 ( .A(n17910), .B(n10766), .Z(n17912) );
  XNOR U19453 ( .A(n17913), .B(n17914), .Z(n10766) );
  XNOR U19454 ( .A(n[515]), .B(n17915), .Z(n17911) );
  IV U19455 ( .A(n17910), .Z(n17915) );
  XOR U19456 ( .A(n17916), .B(n17917), .Z(n17910) );
  AND U19457 ( .A(n17918), .B(n17919), .Z(n17916) );
  XOR U19458 ( .A(n17917), .B(n10771), .Z(n17919) );
  XNOR U19459 ( .A(n17920), .B(n17921), .Z(n10771) );
  XNOR U19460 ( .A(n[514]), .B(n17922), .Z(n17918) );
  IV U19461 ( .A(n17917), .Z(n17922) );
  XOR U19462 ( .A(n17923), .B(n17924), .Z(n17917) );
  AND U19463 ( .A(n17925), .B(n17926), .Z(n17923) );
  XOR U19464 ( .A(n17924), .B(n10776), .Z(n17926) );
  XNOR U19465 ( .A(n17927), .B(n17928), .Z(n10776) );
  XNOR U19466 ( .A(n[513]), .B(n17929), .Z(n17925) );
  IV U19467 ( .A(n17924), .Z(n17929) );
  XOR U19468 ( .A(n17930), .B(n17931), .Z(n17924) );
  AND U19469 ( .A(n17932), .B(n17933), .Z(n17930) );
  XOR U19470 ( .A(n17931), .B(n10781), .Z(n17933) );
  XNOR U19471 ( .A(n17934), .B(n17935), .Z(n10781) );
  XNOR U19472 ( .A(n[512]), .B(n17936), .Z(n17932) );
  IV U19473 ( .A(n17931), .Z(n17936) );
  XOR U19474 ( .A(n17937), .B(n17938), .Z(n17931) );
  AND U19475 ( .A(n17939), .B(n17940), .Z(n17937) );
  XOR U19476 ( .A(n17938), .B(n10786), .Z(n17940) );
  XNOR U19477 ( .A(n17941), .B(n17942), .Z(n10786) );
  XNOR U19478 ( .A(n[511]), .B(n17943), .Z(n17939) );
  IV U19479 ( .A(n17938), .Z(n17943) );
  XOR U19480 ( .A(n17944), .B(n17945), .Z(n17938) );
  AND U19481 ( .A(n17946), .B(n17947), .Z(n17944) );
  XOR U19482 ( .A(n17945), .B(n10791), .Z(n17947) );
  XNOR U19483 ( .A(n17948), .B(n17949), .Z(n10791) );
  XNOR U19484 ( .A(n[510]), .B(n17950), .Z(n17946) );
  IV U19485 ( .A(n17945), .Z(n17950) );
  XOR U19486 ( .A(n17951), .B(n17952), .Z(n17945) );
  AND U19487 ( .A(n17953), .B(n17954), .Z(n17951) );
  XOR U19488 ( .A(n17952), .B(n10796), .Z(n17954) );
  XNOR U19489 ( .A(n17955), .B(n17956), .Z(n10796) );
  XNOR U19490 ( .A(n[509]), .B(n17957), .Z(n17953) );
  IV U19491 ( .A(n17952), .Z(n17957) );
  XOR U19492 ( .A(n17958), .B(n17959), .Z(n17952) );
  AND U19493 ( .A(n17960), .B(n17961), .Z(n17958) );
  XOR U19494 ( .A(n17959), .B(n10801), .Z(n17961) );
  XNOR U19495 ( .A(n17962), .B(n17963), .Z(n10801) );
  XNOR U19496 ( .A(n[508]), .B(n17964), .Z(n17960) );
  IV U19497 ( .A(n17959), .Z(n17964) );
  XOR U19498 ( .A(n17965), .B(n17966), .Z(n17959) );
  AND U19499 ( .A(n17967), .B(n17968), .Z(n17965) );
  XOR U19500 ( .A(n17966), .B(n10806), .Z(n17968) );
  XNOR U19501 ( .A(n17969), .B(n17970), .Z(n10806) );
  XNOR U19502 ( .A(n[507]), .B(n17971), .Z(n17967) );
  IV U19503 ( .A(n17966), .Z(n17971) );
  XOR U19504 ( .A(n17972), .B(n17973), .Z(n17966) );
  AND U19505 ( .A(n17974), .B(n17975), .Z(n17972) );
  XOR U19506 ( .A(n17973), .B(n10811), .Z(n17975) );
  XNOR U19507 ( .A(n17976), .B(n17977), .Z(n10811) );
  XNOR U19508 ( .A(n[506]), .B(n17978), .Z(n17974) );
  IV U19509 ( .A(n17973), .Z(n17978) );
  XOR U19510 ( .A(n17979), .B(n17980), .Z(n17973) );
  AND U19511 ( .A(n17981), .B(n17982), .Z(n17979) );
  XOR U19512 ( .A(n17980), .B(n10816), .Z(n17982) );
  XNOR U19513 ( .A(n17983), .B(n17984), .Z(n10816) );
  XNOR U19514 ( .A(n[505]), .B(n17985), .Z(n17981) );
  IV U19515 ( .A(n17980), .Z(n17985) );
  XOR U19516 ( .A(n17986), .B(n17987), .Z(n17980) );
  AND U19517 ( .A(n17988), .B(n17989), .Z(n17986) );
  XOR U19518 ( .A(n17987), .B(n10821), .Z(n17989) );
  XNOR U19519 ( .A(n17990), .B(n17991), .Z(n10821) );
  XNOR U19520 ( .A(n[504]), .B(n17992), .Z(n17988) );
  IV U19521 ( .A(n17987), .Z(n17992) );
  XOR U19522 ( .A(n17993), .B(n17994), .Z(n17987) );
  AND U19523 ( .A(n17995), .B(n17996), .Z(n17993) );
  XOR U19524 ( .A(n17994), .B(n10826), .Z(n17996) );
  XNOR U19525 ( .A(n17997), .B(n17998), .Z(n10826) );
  XNOR U19526 ( .A(n[503]), .B(n17999), .Z(n17995) );
  IV U19527 ( .A(n17994), .Z(n17999) );
  XOR U19528 ( .A(n18000), .B(n18001), .Z(n17994) );
  AND U19529 ( .A(n18002), .B(n18003), .Z(n18000) );
  XOR U19530 ( .A(n18001), .B(n10831), .Z(n18003) );
  XNOR U19531 ( .A(n18004), .B(n18005), .Z(n10831) );
  XNOR U19532 ( .A(n[502]), .B(n18006), .Z(n18002) );
  IV U19533 ( .A(n18001), .Z(n18006) );
  XOR U19534 ( .A(n18007), .B(n18008), .Z(n18001) );
  AND U19535 ( .A(n18009), .B(n18010), .Z(n18007) );
  XOR U19536 ( .A(n18008), .B(n10836), .Z(n18010) );
  XNOR U19537 ( .A(n18011), .B(n18012), .Z(n10836) );
  XNOR U19538 ( .A(n[501]), .B(n18013), .Z(n18009) );
  IV U19539 ( .A(n18008), .Z(n18013) );
  XOR U19540 ( .A(n18014), .B(n18015), .Z(n18008) );
  AND U19541 ( .A(n18016), .B(n18017), .Z(n18014) );
  XOR U19542 ( .A(n18015), .B(n10841), .Z(n18017) );
  XNOR U19543 ( .A(n18018), .B(n18019), .Z(n10841) );
  XNOR U19544 ( .A(n[500]), .B(n18020), .Z(n18016) );
  IV U19545 ( .A(n18015), .Z(n18020) );
  XOR U19546 ( .A(n18021), .B(n18022), .Z(n18015) );
  AND U19547 ( .A(n18023), .B(n18024), .Z(n18021) );
  XOR U19548 ( .A(n18022), .B(n10846), .Z(n18024) );
  XNOR U19549 ( .A(n18025), .B(n18026), .Z(n10846) );
  XNOR U19550 ( .A(n[499]), .B(n18027), .Z(n18023) );
  IV U19551 ( .A(n18022), .Z(n18027) );
  XOR U19552 ( .A(n18028), .B(n18029), .Z(n18022) );
  AND U19553 ( .A(n18030), .B(n18031), .Z(n18028) );
  XOR U19554 ( .A(n18029), .B(n10851), .Z(n18031) );
  XNOR U19555 ( .A(n18032), .B(n18033), .Z(n10851) );
  XNOR U19556 ( .A(n[498]), .B(n18034), .Z(n18030) );
  IV U19557 ( .A(n18029), .Z(n18034) );
  XOR U19558 ( .A(n18035), .B(n18036), .Z(n18029) );
  AND U19559 ( .A(n18037), .B(n18038), .Z(n18035) );
  XOR U19560 ( .A(n18036), .B(n10856), .Z(n18038) );
  XNOR U19561 ( .A(n18039), .B(n18040), .Z(n10856) );
  XNOR U19562 ( .A(n[497]), .B(n18041), .Z(n18037) );
  IV U19563 ( .A(n18036), .Z(n18041) );
  XOR U19564 ( .A(n18042), .B(n18043), .Z(n18036) );
  AND U19565 ( .A(n18044), .B(n18045), .Z(n18042) );
  XOR U19566 ( .A(n18043), .B(n10861), .Z(n18045) );
  XNOR U19567 ( .A(n18046), .B(n18047), .Z(n10861) );
  XNOR U19568 ( .A(n[496]), .B(n18048), .Z(n18044) );
  IV U19569 ( .A(n18043), .Z(n18048) );
  XOR U19570 ( .A(n18049), .B(n18050), .Z(n18043) );
  AND U19571 ( .A(n18051), .B(n18052), .Z(n18049) );
  XOR U19572 ( .A(n18050), .B(n10866), .Z(n18052) );
  XNOR U19573 ( .A(n18053), .B(n18054), .Z(n10866) );
  XNOR U19574 ( .A(n[495]), .B(n18055), .Z(n18051) );
  IV U19575 ( .A(n18050), .Z(n18055) );
  XOR U19576 ( .A(n18056), .B(n18057), .Z(n18050) );
  AND U19577 ( .A(n18058), .B(n18059), .Z(n18056) );
  XOR U19578 ( .A(n18057), .B(n10871), .Z(n18059) );
  XNOR U19579 ( .A(n18060), .B(n18061), .Z(n10871) );
  XNOR U19580 ( .A(n[494]), .B(n18062), .Z(n18058) );
  IV U19581 ( .A(n18057), .Z(n18062) );
  XOR U19582 ( .A(n18063), .B(n18064), .Z(n18057) );
  AND U19583 ( .A(n18065), .B(n18066), .Z(n18063) );
  XOR U19584 ( .A(n18064), .B(n10876), .Z(n18066) );
  XNOR U19585 ( .A(n18067), .B(n18068), .Z(n10876) );
  XNOR U19586 ( .A(n[493]), .B(n18069), .Z(n18065) );
  IV U19587 ( .A(n18064), .Z(n18069) );
  XOR U19588 ( .A(n18070), .B(n18071), .Z(n18064) );
  AND U19589 ( .A(n18072), .B(n18073), .Z(n18070) );
  XOR U19590 ( .A(n18071), .B(n10881), .Z(n18073) );
  XNOR U19591 ( .A(n18074), .B(n18075), .Z(n10881) );
  XNOR U19592 ( .A(n[492]), .B(n18076), .Z(n18072) );
  IV U19593 ( .A(n18071), .Z(n18076) );
  XOR U19594 ( .A(n18077), .B(n18078), .Z(n18071) );
  AND U19595 ( .A(n18079), .B(n18080), .Z(n18077) );
  XOR U19596 ( .A(n18078), .B(n10886), .Z(n18080) );
  XNOR U19597 ( .A(n18081), .B(n18082), .Z(n10886) );
  XNOR U19598 ( .A(n[491]), .B(n18083), .Z(n18079) );
  IV U19599 ( .A(n18078), .Z(n18083) );
  XOR U19600 ( .A(n18084), .B(n18085), .Z(n18078) );
  AND U19601 ( .A(n18086), .B(n18087), .Z(n18084) );
  XOR U19602 ( .A(n18085), .B(n10891), .Z(n18087) );
  XNOR U19603 ( .A(n18088), .B(n18089), .Z(n10891) );
  XNOR U19604 ( .A(n[490]), .B(n18090), .Z(n18086) );
  IV U19605 ( .A(n18085), .Z(n18090) );
  XOR U19606 ( .A(n18091), .B(n18092), .Z(n18085) );
  AND U19607 ( .A(n18093), .B(n18094), .Z(n18091) );
  XOR U19608 ( .A(n18092), .B(n10896), .Z(n18094) );
  XNOR U19609 ( .A(n18095), .B(n18096), .Z(n10896) );
  XNOR U19610 ( .A(n[489]), .B(n18097), .Z(n18093) );
  IV U19611 ( .A(n18092), .Z(n18097) );
  XOR U19612 ( .A(n18098), .B(n18099), .Z(n18092) );
  AND U19613 ( .A(n18100), .B(n18101), .Z(n18098) );
  XOR U19614 ( .A(n18099), .B(n10901), .Z(n18101) );
  XNOR U19615 ( .A(n18102), .B(n18103), .Z(n10901) );
  XNOR U19616 ( .A(n[488]), .B(n18104), .Z(n18100) );
  IV U19617 ( .A(n18099), .Z(n18104) );
  XOR U19618 ( .A(n18105), .B(n18106), .Z(n18099) );
  AND U19619 ( .A(n18107), .B(n18108), .Z(n18105) );
  XOR U19620 ( .A(n18106), .B(n10906), .Z(n18108) );
  XNOR U19621 ( .A(n18109), .B(n18110), .Z(n10906) );
  XNOR U19622 ( .A(n[487]), .B(n18111), .Z(n18107) );
  IV U19623 ( .A(n18106), .Z(n18111) );
  XOR U19624 ( .A(n18112), .B(n18113), .Z(n18106) );
  AND U19625 ( .A(n18114), .B(n18115), .Z(n18112) );
  XOR U19626 ( .A(n18113), .B(n10911), .Z(n18115) );
  XNOR U19627 ( .A(n18116), .B(n18117), .Z(n10911) );
  XNOR U19628 ( .A(n[486]), .B(n18118), .Z(n18114) );
  IV U19629 ( .A(n18113), .Z(n18118) );
  XOR U19630 ( .A(n18119), .B(n18120), .Z(n18113) );
  AND U19631 ( .A(n18121), .B(n18122), .Z(n18119) );
  XOR U19632 ( .A(n18120), .B(n10916), .Z(n18122) );
  XNOR U19633 ( .A(n18123), .B(n18124), .Z(n10916) );
  XNOR U19634 ( .A(n[485]), .B(n18125), .Z(n18121) );
  IV U19635 ( .A(n18120), .Z(n18125) );
  XOR U19636 ( .A(n18126), .B(n18127), .Z(n18120) );
  AND U19637 ( .A(n18128), .B(n18129), .Z(n18126) );
  XOR U19638 ( .A(n18127), .B(n10921), .Z(n18129) );
  XNOR U19639 ( .A(n18130), .B(n18131), .Z(n10921) );
  XNOR U19640 ( .A(n[484]), .B(n18132), .Z(n18128) );
  IV U19641 ( .A(n18127), .Z(n18132) );
  XOR U19642 ( .A(n18133), .B(n18134), .Z(n18127) );
  AND U19643 ( .A(n18135), .B(n18136), .Z(n18133) );
  XOR U19644 ( .A(n18134), .B(n10926), .Z(n18136) );
  XNOR U19645 ( .A(n18137), .B(n18138), .Z(n10926) );
  XNOR U19646 ( .A(n[483]), .B(n18139), .Z(n18135) );
  IV U19647 ( .A(n18134), .Z(n18139) );
  XOR U19648 ( .A(n18140), .B(n18141), .Z(n18134) );
  AND U19649 ( .A(n18142), .B(n18143), .Z(n18140) );
  XOR U19650 ( .A(n18141), .B(n10931), .Z(n18143) );
  XNOR U19651 ( .A(n18144), .B(n18145), .Z(n10931) );
  XNOR U19652 ( .A(n[482]), .B(n18146), .Z(n18142) );
  IV U19653 ( .A(n18141), .Z(n18146) );
  XOR U19654 ( .A(n18147), .B(n18148), .Z(n18141) );
  AND U19655 ( .A(n18149), .B(n18150), .Z(n18147) );
  XOR U19656 ( .A(n18148), .B(n10936), .Z(n18150) );
  XNOR U19657 ( .A(n18151), .B(n18152), .Z(n10936) );
  XNOR U19658 ( .A(n[481]), .B(n18153), .Z(n18149) );
  IV U19659 ( .A(n18148), .Z(n18153) );
  XOR U19660 ( .A(n18154), .B(n18155), .Z(n18148) );
  AND U19661 ( .A(n18156), .B(n18157), .Z(n18154) );
  XOR U19662 ( .A(n18155), .B(n10941), .Z(n18157) );
  XNOR U19663 ( .A(n18158), .B(n18159), .Z(n10941) );
  XNOR U19664 ( .A(n[480]), .B(n18160), .Z(n18156) );
  IV U19665 ( .A(n18155), .Z(n18160) );
  XOR U19666 ( .A(n18161), .B(n18162), .Z(n18155) );
  AND U19667 ( .A(n18163), .B(n18164), .Z(n18161) );
  XOR U19668 ( .A(n18162), .B(n10946), .Z(n18164) );
  XNOR U19669 ( .A(n18165), .B(n18166), .Z(n10946) );
  XNOR U19670 ( .A(n[479]), .B(n18167), .Z(n18163) );
  IV U19671 ( .A(n18162), .Z(n18167) );
  XOR U19672 ( .A(n18168), .B(n18169), .Z(n18162) );
  AND U19673 ( .A(n18170), .B(n18171), .Z(n18168) );
  XOR U19674 ( .A(n18169), .B(n10951), .Z(n18171) );
  XNOR U19675 ( .A(n18172), .B(n18173), .Z(n10951) );
  XNOR U19676 ( .A(n[478]), .B(n18174), .Z(n18170) );
  IV U19677 ( .A(n18169), .Z(n18174) );
  XOR U19678 ( .A(n18175), .B(n18176), .Z(n18169) );
  AND U19679 ( .A(n18177), .B(n18178), .Z(n18175) );
  XOR U19680 ( .A(n18176), .B(n10956), .Z(n18178) );
  XNOR U19681 ( .A(n18179), .B(n18180), .Z(n10956) );
  XNOR U19682 ( .A(n[477]), .B(n18181), .Z(n18177) );
  IV U19683 ( .A(n18176), .Z(n18181) );
  XOR U19684 ( .A(n18182), .B(n18183), .Z(n18176) );
  AND U19685 ( .A(n18184), .B(n18185), .Z(n18182) );
  XOR U19686 ( .A(n18183), .B(n10961), .Z(n18185) );
  XNOR U19687 ( .A(n18186), .B(n18187), .Z(n10961) );
  XNOR U19688 ( .A(n[476]), .B(n18188), .Z(n18184) );
  IV U19689 ( .A(n18183), .Z(n18188) );
  XOR U19690 ( .A(n18189), .B(n18190), .Z(n18183) );
  AND U19691 ( .A(n18191), .B(n18192), .Z(n18189) );
  XOR U19692 ( .A(n18190), .B(n10966), .Z(n18192) );
  XNOR U19693 ( .A(n18193), .B(n18194), .Z(n10966) );
  XNOR U19694 ( .A(n[475]), .B(n18195), .Z(n18191) );
  IV U19695 ( .A(n18190), .Z(n18195) );
  XOR U19696 ( .A(n18196), .B(n18197), .Z(n18190) );
  AND U19697 ( .A(n18198), .B(n18199), .Z(n18196) );
  XOR U19698 ( .A(n18197), .B(n10971), .Z(n18199) );
  XNOR U19699 ( .A(n18200), .B(n18201), .Z(n10971) );
  XNOR U19700 ( .A(n[474]), .B(n18202), .Z(n18198) );
  IV U19701 ( .A(n18197), .Z(n18202) );
  XOR U19702 ( .A(n18203), .B(n18204), .Z(n18197) );
  AND U19703 ( .A(n18205), .B(n18206), .Z(n18203) );
  XOR U19704 ( .A(n18204), .B(n10976), .Z(n18206) );
  XNOR U19705 ( .A(n18207), .B(n18208), .Z(n10976) );
  XNOR U19706 ( .A(n[473]), .B(n18209), .Z(n18205) );
  IV U19707 ( .A(n18204), .Z(n18209) );
  XOR U19708 ( .A(n18210), .B(n18211), .Z(n18204) );
  AND U19709 ( .A(n18212), .B(n18213), .Z(n18210) );
  XOR U19710 ( .A(n18211), .B(n10981), .Z(n18213) );
  XNOR U19711 ( .A(n18214), .B(n18215), .Z(n10981) );
  XNOR U19712 ( .A(n[472]), .B(n18216), .Z(n18212) );
  IV U19713 ( .A(n18211), .Z(n18216) );
  XOR U19714 ( .A(n18217), .B(n18218), .Z(n18211) );
  AND U19715 ( .A(n18219), .B(n18220), .Z(n18217) );
  XOR U19716 ( .A(n18218), .B(n10986), .Z(n18220) );
  XNOR U19717 ( .A(n18221), .B(n18222), .Z(n10986) );
  XNOR U19718 ( .A(n[471]), .B(n18223), .Z(n18219) );
  IV U19719 ( .A(n18218), .Z(n18223) );
  XOR U19720 ( .A(n18224), .B(n18225), .Z(n18218) );
  AND U19721 ( .A(n18226), .B(n18227), .Z(n18224) );
  XOR U19722 ( .A(n18225), .B(n10991), .Z(n18227) );
  XNOR U19723 ( .A(n18228), .B(n18229), .Z(n10991) );
  XNOR U19724 ( .A(n[470]), .B(n18230), .Z(n18226) );
  IV U19725 ( .A(n18225), .Z(n18230) );
  XOR U19726 ( .A(n18231), .B(n18232), .Z(n18225) );
  AND U19727 ( .A(n18233), .B(n18234), .Z(n18231) );
  XOR U19728 ( .A(n18232), .B(n10996), .Z(n18234) );
  XNOR U19729 ( .A(n18235), .B(n18236), .Z(n10996) );
  XNOR U19730 ( .A(n[469]), .B(n18237), .Z(n18233) );
  IV U19731 ( .A(n18232), .Z(n18237) );
  XOR U19732 ( .A(n18238), .B(n18239), .Z(n18232) );
  AND U19733 ( .A(n18240), .B(n18241), .Z(n18238) );
  XOR U19734 ( .A(n18239), .B(n11001), .Z(n18241) );
  XNOR U19735 ( .A(n18242), .B(n18243), .Z(n11001) );
  XNOR U19736 ( .A(n[468]), .B(n18244), .Z(n18240) );
  IV U19737 ( .A(n18239), .Z(n18244) );
  XOR U19738 ( .A(n18245), .B(n18246), .Z(n18239) );
  AND U19739 ( .A(n18247), .B(n18248), .Z(n18245) );
  XOR U19740 ( .A(n18246), .B(n11006), .Z(n18248) );
  XNOR U19741 ( .A(n18249), .B(n18250), .Z(n11006) );
  XNOR U19742 ( .A(n[467]), .B(n18251), .Z(n18247) );
  IV U19743 ( .A(n18246), .Z(n18251) );
  XOR U19744 ( .A(n18252), .B(n18253), .Z(n18246) );
  AND U19745 ( .A(n18254), .B(n18255), .Z(n18252) );
  XOR U19746 ( .A(n18253), .B(n11011), .Z(n18255) );
  XNOR U19747 ( .A(n18256), .B(n18257), .Z(n11011) );
  XNOR U19748 ( .A(n[466]), .B(n18258), .Z(n18254) );
  IV U19749 ( .A(n18253), .Z(n18258) );
  XOR U19750 ( .A(n18259), .B(n18260), .Z(n18253) );
  AND U19751 ( .A(n18261), .B(n18262), .Z(n18259) );
  XOR U19752 ( .A(n18260), .B(n11016), .Z(n18262) );
  XNOR U19753 ( .A(n18263), .B(n18264), .Z(n11016) );
  XNOR U19754 ( .A(n[465]), .B(n18265), .Z(n18261) );
  IV U19755 ( .A(n18260), .Z(n18265) );
  XOR U19756 ( .A(n18266), .B(n18267), .Z(n18260) );
  AND U19757 ( .A(n18268), .B(n18269), .Z(n18266) );
  XOR U19758 ( .A(n18267), .B(n11021), .Z(n18269) );
  XNOR U19759 ( .A(n18270), .B(n18271), .Z(n11021) );
  XNOR U19760 ( .A(n[464]), .B(n18272), .Z(n18268) );
  IV U19761 ( .A(n18267), .Z(n18272) );
  XOR U19762 ( .A(n18273), .B(n18274), .Z(n18267) );
  AND U19763 ( .A(n18275), .B(n18276), .Z(n18273) );
  XOR U19764 ( .A(n18274), .B(n11026), .Z(n18276) );
  XNOR U19765 ( .A(n18277), .B(n18278), .Z(n11026) );
  XNOR U19766 ( .A(n[463]), .B(n18279), .Z(n18275) );
  IV U19767 ( .A(n18274), .Z(n18279) );
  XOR U19768 ( .A(n18280), .B(n18281), .Z(n18274) );
  AND U19769 ( .A(n18282), .B(n18283), .Z(n18280) );
  XOR U19770 ( .A(n18281), .B(n11031), .Z(n18283) );
  XNOR U19771 ( .A(n18284), .B(n18285), .Z(n11031) );
  XNOR U19772 ( .A(n[462]), .B(n18286), .Z(n18282) );
  IV U19773 ( .A(n18281), .Z(n18286) );
  XOR U19774 ( .A(n18287), .B(n18288), .Z(n18281) );
  AND U19775 ( .A(n18289), .B(n18290), .Z(n18287) );
  XOR U19776 ( .A(n18288), .B(n11036), .Z(n18290) );
  XNOR U19777 ( .A(n18291), .B(n18292), .Z(n11036) );
  XNOR U19778 ( .A(n[461]), .B(n18293), .Z(n18289) );
  IV U19779 ( .A(n18288), .Z(n18293) );
  XOR U19780 ( .A(n18294), .B(n18295), .Z(n18288) );
  AND U19781 ( .A(n18296), .B(n18297), .Z(n18294) );
  XOR U19782 ( .A(n18295), .B(n11041), .Z(n18297) );
  XNOR U19783 ( .A(n18298), .B(n18299), .Z(n11041) );
  XNOR U19784 ( .A(n[460]), .B(n18300), .Z(n18296) );
  IV U19785 ( .A(n18295), .Z(n18300) );
  XOR U19786 ( .A(n18301), .B(n18302), .Z(n18295) );
  AND U19787 ( .A(n18303), .B(n18304), .Z(n18301) );
  XOR U19788 ( .A(n18302), .B(n11046), .Z(n18304) );
  XNOR U19789 ( .A(n18305), .B(n18306), .Z(n11046) );
  XNOR U19790 ( .A(n[459]), .B(n18307), .Z(n18303) );
  IV U19791 ( .A(n18302), .Z(n18307) );
  XOR U19792 ( .A(n18308), .B(n18309), .Z(n18302) );
  AND U19793 ( .A(n18310), .B(n18311), .Z(n18308) );
  XOR U19794 ( .A(n18309), .B(n11051), .Z(n18311) );
  XNOR U19795 ( .A(n18312), .B(n18313), .Z(n11051) );
  XNOR U19796 ( .A(n[458]), .B(n18314), .Z(n18310) );
  IV U19797 ( .A(n18309), .Z(n18314) );
  XOR U19798 ( .A(n18315), .B(n18316), .Z(n18309) );
  AND U19799 ( .A(n18317), .B(n18318), .Z(n18315) );
  XOR U19800 ( .A(n18316), .B(n11056), .Z(n18318) );
  XNOR U19801 ( .A(n18319), .B(n18320), .Z(n11056) );
  XNOR U19802 ( .A(n[457]), .B(n18321), .Z(n18317) );
  IV U19803 ( .A(n18316), .Z(n18321) );
  XOR U19804 ( .A(n18322), .B(n18323), .Z(n18316) );
  AND U19805 ( .A(n18324), .B(n18325), .Z(n18322) );
  XOR U19806 ( .A(n18323), .B(n11061), .Z(n18325) );
  XNOR U19807 ( .A(n18326), .B(n18327), .Z(n11061) );
  XNOR U19808 ( .A(n[456]), .B(n18328), .Z(n18324) );
  IV U19809 ( .A(n18323), .Z(n18328) );
  XOR U19810 ( .A(n18329), .B(n18330), .Z(n18323) );
  AND U19811 ( .A(n18331), .B(n18332), .Z(n18329) );
  XOR U19812 ( .A(n18330), .B(n11066), .Z(n18332) );
  XNOR U19813 ( .A(n18333), .B(n18334), .Z(n11066) );
  XNOR U19814 ( .A(n[455]), .B(n18335), .Z(n18331) );
  IV U19815 ( .A(n18330), .Z(n18335) );
  XOR U19816 ( .A(n18336), .B(n18337), .Z(n18330) );
  AND U19817 ( .A(n18338), .B(n18339), .Z(n18336) );
  XOR U19818 ( .A(n18337), .B(n11071), .Z(n18339) );
  XNOR U19819 ( .A(n18340), .B(n18341), .Z(n11071) );
  XNOR U19820 ( .A(n[454]), .B(n18342), .Z(n18338) );
  IV U19821 ( .A(n18337), .Z(n18342) );
  XOR U19822 ( .A(n18343), .B(n18344), .Z(n18337) );
  AND U19823 ( .A(n18345), .B(n18346), .Z(n18343) );
  XOR U19824 ( .A(n18344), .B(n11076), .Z(n18346) );
  XNOR U19825 ( .A(n18347), .B(n18348), .Z(n11076) );
  XNOR U19826 ( .A(n[453]), .B(n18349), .Z(n18345) );
  IV U19827 ( .A(n18344), .Z(n18349) );
  XOR U19828 ( .A(n18350), .B(n18351), .Z(n18344) );
  AND U19829 ( .A(n18352), .B(n18353), .Z(n18350) );
  XOR U19830 ( .A(n18351), .B(n11081), .Z(n18353) );
  XNOR U19831 ( .A(n18354), .B(n18355), .Z(n11081) );
  XNOR U19832 ( .A(n[452]), .B(n18356), .Z(n18352) );
  IV U19833 ( .A(n18351), .Z(n18356) );
  XOR U19834 ( .A(n18357), .B(n18358), .Z(n18351) );
  AND U19835 ( .A(n18359), .B(n18360), .Z(n18357) );
  XOR U19836 ( .A(n18358), .B(n11086), .Z(n18360) );
  XNOR U19837 ( .A(n18361), .B(n18362), .Z(n11086) );
  XNOR U19838 ( .A(n[451]), .B(n18363), .Z(n18359) );
  IV U19839 ( .A(n18358), .Z(n18363) );
  XOR U19840 ( .A(n18364), .B(n18365), .Z(n18358) );
  AND U19841 ( .A(n18366), .B(n18367), .Z(n18364) );
  XOR U19842 ( .A(n18365), .B(n11091), .Z(n18367) );
  XNOR U19843 ( .A(n18368), .B(n18369), .Z(n11091) );
  XNOR U19844 ( .A(n[450]), .B(n18370), .Z(n18366) );
  IV U19845 ( .A(n18365), .Z(n18370) );
  XOR U19846 ( .A(n18371), .B(n18372), .Z(n18365) );
  AND U19847 ( .A(n18373), .B(n18374), .Z(n18371) );
  XOR U19848 ( .A(n18372), .B(n11096), .Z(n18374) );
  XNOR U19849 ( .A(n18375), .B(n18376), .Z(n11096) );
  XNOR U19850 ( .A(n[449]), .B(n18377), .Z(n18373) );
  IV U19851 ( .A(n18372), .Z(n18377) );
  XOR U19852 ( .A(n18378), .B(n18379), .Z(n18372) );
  AND U19853 ( .A(n18380), .B(n18381), .Z(n18378) );
  XOR U19854 ( .A(n18379), .B(n11101), .Z(n18381) );
  XNOR U19855 ( .A(n18382), .B(n18383), .Z(n11101) );
  XNOR U19856 ( .A(n[448]), .B(n18384), .Z(n18380) );
  IV U19857 ( .A(n18379), .Z(n18384) );
  XOR U19858 ( .A(n18385), .B(n18386), .Z(n18379) );
  AND U19859 ( .A(n18387), .B(n18388), .Z(n18385) );
  XOR U19860 ( .A(n18386), .B(n11106), .Z(n18388) );
  XNOR U19861 ( .A(n18389), .B(n18390), .Z(n11106) );
  XNOR U19862 ( .A(n[447]), .B(n18391), .Z(n18387) );
  IV U19863 ( .A(n18386), .Z(n18391) );
  XOR U19864 ( .A(n18392), .B(n18393), .Z(n18386) );
  AND U19865 ( .A(n18394), .B(n18395), .Z(n18392) );
  XOR U19866 ( .A(n18393), .B(n11111), .Z(n18395) );
  XNOR U19867 ( .A(n18396), .B(n18397), .Z(n11111) );
  XNOR U19868 ( .A(n[446]), .B(n18398), .Z(n18394) );
  IV U19869 ( .A(n18393), .Z(n18398) );
  XOR U19870 ( .A(n18399), .B(n18400), .Z(n18393) );
  AND U19871 ( .A(n18401), .B(n18402), .Z(n18399) );
  XOR U19872 ( .A(n18400), .B(n11116), .Z(n18402) );
  XNOR U19873 ( .A(n18403), .B(n18404), .Z(n11116) );
  XNOR U19874 ( .A(n[445]), .B(n18405), .Z(n18401) );
  IV U19875 ( .A(n18400), .Z(n18405) );
  XOR U19876 ( .A(n18406), .B(n18407), .Z(n18400) );
  AND U19877 ( .A(n18408), .B(n18409), .Z(n18406) );
  XOR U19878 ( .A(n18407), .B(n11121), .Z(n18409) );
  XNOR U19879 ( .A(n18410), .B(n18411), .Z(n11121) );
  XNOR U19880 ( .A(n[444]), .B(n18412), .Z(n18408) );
  IV U19881 ( .A(n18407), .Z(n18412) );
  XOR U19882 ( .A(n18413), .B(n18414), .Z(n18407) );
  AND U19883 ( .A(n18415), .B(n18416), .Z(n18413) );
  XOR U19884 ( .A(n18414), .B(n11126), .Z(n18416) );
  XNOR U19885 ( .A(n18417), .B(n18418), .Z(n11126) );
  XNOR U19886 ( .A(n[443]), .B(n18419), .Z(n18415) );
  IV U19887 ( .A(n18414), .Z(n18419) );
  XOR U19888 ( .A(n18420), .B(n18421), .Z(n18414) );
  AND U19889 ( .A(n18422), .B(n18423), .Z(n18420) );
  XOR U19890 ( .A(n18421), .B(n11131), .Z(n18423) );
  XNOR U19891 ( .A(n18424), .B(n18425), .Z(n11131) );
  XNOR U19892 ( .A(n[442]), .B(n18426), .Z(n18422) );
  IV U19893 ( .A(n18421), .Z(n18426) );
  XOR U19894 ( .A(n18427), .B(n18428), .Z(n18421) );
  AND U19895 ( .A(n18429), .B(n18430), .Z(n18427) );
  XOR U19896 ( .A(n18428), .B(n11136), .Z(n18430) );
  XNOR U19897 ( .A(n18431), .B(n18432), .Z(n11136) );
  XNOR U19898 ( .A(n[441]), .B(n18433), .Z(n18429) );
  IV U19899 ( .A(n18428), .Z(n18433) );
  XOR U19900 ( .A(n18434), .B(n18435), .Z(n18428) );
  AND U19901 ( .A(n18436), .B(n18437), .Z(n18434) );
  XOR U19902 ( .A(n18435), .B(n11141), .Z(n18437) );
  XNOR U19903 ( .A(n18438), .B(n18439), .Z(n11141) );
  XNOR U19904 ( .A(n[440]), .B(n18440), .Z(n18436) );
  IV U19905 ( .A(n18435), .Z(n18440) );
  XOR U19906 ( .A(n18441), .B(n18442), .Z(n18435) );
  AND U19907 ( .A(n18443), .B(n18444), .Z(n18441) );
  XOR U19908 ( .A(n18442), .B(n11146), .Z(n18444) );
  XNOR U19909 ( .A(n18445), .B(n18446), .Z(n11146) );
  XNOR U19910 ( .A(n[439]), .B(n18447), .Z(n18443) );
  IV U19911 ( .A(n18442), .Z(n18447) );
  XOR U19912 ( .A(n18448), .B(n18449), .Z(n18442) );
  AND U19913 ( .A(n18450), .B(n18451), .Z(n18448) );
  XOR U19914 ( .A(n18449), .B(n11151), .Z(n18451) );
  XNOR U19915 ( .A(n18452), .B(n18453), .Z(n11151) );
  XNOR U19916 ( .A(n[438]), .B(n18454), .Z(n18450) );
  IV U19917 ( .A(n18449), .Z(n18454) );
  XOR U19918 ( .A(n18455), .B(n18456), .Z(n18449) );
  AND U19919 ( .A(n18457), .B(n18458), .Z(n18455) );
  XOR U19920 ( .A(n18456), .B(n11156), .Z(n18458) );
  XNOR U19921 ( .A(n18459), .B(n18460), .Z(n11156) );
  XNOR U19922 ( .A(n[437]), .B(n18461), .Z(n18457) );
  IV U19923 ( .A(n18456), .Z(n18461) );
  XOR U19924 ( .A(n18462), .B(n18463), .Z(n18456) );
  AND U19925 ( .A(n18464), .B(n18465), .Z(n18462) );
  XOR U19926 ( .A(n18463), .B(n11161), .Z(n18465) );
  XNOR U19927 ( .A(n18466), .B(n18467), .Z(n11161) );
  XNOR U19928 ( .A(n[436]), .B(n18468), .Z(n18464) );
  IV U19929 ( .A(n18463), .Z(n18468) );
  XOR U19930 ( .A(n18469), .B(n18470), .Z(n18463) );
  AND U19931 ( .A(n18471), .B(n18472), .Z(n18469) );
  XOR U19932 ( .A(n18470), .B(n11166), .Z(n18472) );
  XNOR U19933 ( .A(n18473), .B(n18474), .Z(n11166) );
  XNOR U19934 ( .A(n[435]), .B(n18475), .Z(n18471) );
  IV U19935 ( .A(n18470), .Z(n18475) );
  XOR U19936 ( .A(n18476), .B(n18477), .Z(n18470) );
  AND U19937 ( .A(n18478), .B(n18479), .Z(n18476) );
  XOR U19938 ( .A(n18477), .B(n11171), .Z(n18479) );
  XNOR U19939 ( .A(n18480), .B(n18481), .Z(n11171) );
  XNOR U19940 ( .A(n[434]), .B(n18482), .Z(n18478) );
  IV U19941 ( .A(n18477), .Z(n18482) );
  XOR U19942 ( .A(n18483), .B(n18484), .Z(n18477) );
  AND U19943 ( .A(n18485), .B(n18486), .Z(n18483) );
  XOR U19944 ( .A(n18484), .B(n11176), .Z(n18486) );
  XNOR U19945 ( .A(n18487), .B(n18488), .Z(n11176) );
  XNOR U19946 ( .A(n[433]), .B(n18489), .Z(n18485) );
  IV U19947 ( .A(n18484), .Z(n18489) );
  XOR U19948 ( .A(n18490), .B(n18491), .Z(n18484) );
  AND U19949 ( .A(n18492), .B(n18493), .Z(n18490) );
  XOR U19950 ( .A(n18491), .B(n11181), .Z(n18493) );
  XNOR U19951 ( .A(n18494), .B(n18495), .Z(n11181) );
  XNOR U19952 ( .A(n[432]), .B(n18496), .Z(n18492) );
  IV U19953 ( .A(n18491), .Z(n18496) );
  XOR U19954 ( .A(n18497), .B(n18498), .Z(n18491) );
  AND U19955 ( .A(n18499), .B(n18500), .Z(n18497) );
  XOR U19956 ( .A(n18498), .B(n11186), .Z(n18500) );
  XNOR U19957 ( .A(n18501), .B(n18502), .Z(n11186) );
  XNOR U19958 ( .A(n[431]), .B(n18503), .Z(n18499) );
  IV U19959 ( .A(n18498), .Z(n18503) );
  XOR U19960 ( .A(n18504), .B(n18505), .Z(n18498) );
  AND U19961 ( .A(n18506), .B(n18507), .Z(n18504) );
  XOR U19962 ( .A(n18505), .B(n11191), .Z(n18507) );
  XNOR U19963 ( .A(n18508), .B(n18509), .Z(n11191) );
  XNOR U19964 ( .A(n[430]), .B(n18510), .Z(n18506) );
  IV U19965 ( .A(n18505), .Z(n18510) );
  XOR U19966 ( .A(n18511), .B(n18512), .Z(n18505) );
  AND U19967 ( .A(n18513), .B(n18514), .Z(n18511) );
  XOR U19968 ( .A(n18512), .B(n11196), .Z(n18514) );
  XNOR U19969 ( .A(n18515), .B(n18516), .Z(n11196) );
  XNOR U19970 ( .A(n[429]), .B(n18517), .Z(n18513) );
  IV U19971 ( .A(n18512), .Z(n18517) );
  XOR U19972 ( .A(n18518), .B(n18519), .Z(n18512) );
  AND U19973 ( .A(n18520), .B(n18521), .Z(n18518) );
  XOR U19974 ( .A(n18519), .B(n11201), .Z(n18521) );
  XNOR U19975 ( .A(n18522), .B(n18523), .Z(n11201) );
  XNOR U19976 ( .A(n[428]), .B(n18524), .Z(n18520) );
  IV U19977 ( .A(n18519), .Z(n18524) );
  XOR U19978 ( .A(n18525), .B(n18526), .Z(n18519) );
  AND U19979 ( .A(n18527), .B(n18528), .Z(n18525) );
  XOR U19980 ( .A(n18526), .B(n11206), .Z(n18528) );
  XNOR U19981 ( .A(n18529), .B(n18530), .Z(n11206) );
  XNOR U19982 ( .A(n[427]), .B(n18531), .Z(n18527) );
  IV U19983 ( .A(n18526), .Z(n18531) );
  XOR U19984 ( .A(n18532), .B(n18533), .Z(n18526) );
  AND U19985 ( .A(n18534), .B(n18535), .Z(n18532) );
  XOR U19986 ( .A(n18533), .B(n11211), .Z(n18535) );
  XNOR U19987 ( .A(n18536), .B(n18537), .Z(n11211) );
  XNOR U19988 ( .A(n[426]), .B(n18538), .Z(n18534) );
  IV U19989 ( .A(n18533), .Z(n18538) );
  XOR U19990 ( .A(n18539), .B(n18540), .Z(n18533) );
  AND U19991 ( .A(n18541), .B(n18542), .Z(n18539) );
  XOR U19992 ( .A(n18540), .B(n11216), .Z(n18542) );
  XNOR U19993 ( .A(n18543), .B(n18544), .Z(n11216) );
  XNOR U19994 ( .A(n[425]), .B(n18545), .Z(n18541) );
  IV U19995 ( .A(n18540), .Z(n18545) );
  XOR U19996 ( .A(n18546), .B(n18547), .Z(n18540) );
  AND U19997 ( .A(n18548), .B(n18549), .Z(n18546) );
  XOR U19998 ( .A(n18547), .B(n11221), .Z(n18549) );
  XNOR U19999 ( .A(n18550), .B(n18551), .Z(n11221) );
  XNOR U20000 ( .A(n[424]), .B(n18552), .Z(n18548) );
  IV U20001 ( .A(n18547), .Z(n18552) );
  XOR U20002 ( .A(n18553), .B(n18554), .Z(n18547) );
  AND U20003 ( .A(n18555), .B(n18556), .Z(n18553) );
  XOR U20004 ( .A(n18554), .B(n11226), .Z(n18556) );
  XNOR U20005 ( .A(n18557), .B(n18558), .Z(n11226) );
  XNOR U20006 ( .A(n[423]), .B(n18559), .Z(n18555) );
  IV U20007 ( .A(n18554), .Z(n18559) );
  XOR U20008 ( .A(n18560), .B(n18561), .Z(n18554) );
  AND U20009 ( .A(n18562), .B(n18563), .Z(n18560) );
  XOR U20010 ( .A(n18561), .B(n11231), .Z(n18563) );
  XNOR U20011 ( .A(n18564), .B(n18565), .Z(n11231) );
  XNOR U20012 ( .A(n[422]), .B(n18566), .Z(n18562) );
  IV U20013 ( .A(n18561), .Z(n18566) );
  XOR U20014 ( .A(n18567), .B(n18568), .Z(n18561) );
  AND U20015 ( .A(n18569), .B(n18570), .Z(n18567) );
  XOR U20016 ( .A(n18568), .B(n11236), .Z(n18570) );
  XNOR U20017 ( .A(n18571), .B(n18572), .Z(n11236) );
  XNOR U20018 ( .A(n[421]), .B(n18573), .Z(n18569) );
  IV U20019 ( .A(n18568), .Z(n18573) );
  XOR U20020 ( .A(n18574), .B(n18575), .Z(n18568) );
  AND U20021 ( .A(n18576), .B(n18577), .Z(n18574) );
  XOR U20022 ( .A(n18575), .B(n11241), .Z(n18577) );
  XNOR U20023 ( .A(n18578), .B(n18579), .Z(n11241) );
  XNOR U20024 ( .A(n[420]), .B(n18580), .Z(n18576) );
  IV U20025 ( .A(n18575), .Z(n18580) );
  XOR U20026 ( .A(n18581), .B(n18582), .Z(n18575) );
  AND U20027 ( .A(n18583), .B(n18584), .Z(n18581) );
  XOR U20028 ( .A(n18582), .B(n11246), .Z(n18584) );
  XNOR U20029 ( .A(n18585), .B(n18586), .Z(n11246) );
  XNOR U20030 ( .A(n[419]), .B(n18587), .Z(n18583) );
  IV U20031 ( .A(n18582), .Z(n18587) );
  XOR U20032 ( .A(n18588), .B(n18589), .Z(n18582) );
  AND U20033 ( .A(n18590), .B(n18591), .Z(n18588) );
  XOR U20034 ( .A(n18589), .B(n11251), .Z(n18591) );
  XNOR U20035 ( .A(n18592), .B(n18593), .Z(n11251) );
  XNOR U20036 ( .A(n[418]), .B(n18594), .Z(n18590) );
  IV U20037 ( .A(n18589), .Z(n18594) );
  XOR U20038 ( .A(n18595), .B(n18596), .Z(n18589) );
  AND U20039 ( .A(n18597), .B(n18598), .Z(n18595) );
  XOR U20040 ( .A(n18596), .B(n11256), .Z(n18598) );
  XNOR U20041 ( .A(n18599), .B(n18600), .Z(n11256) );
  XNOR U20042 ( .A(n[417]), .B(n18601), .Z(n18597) );
  IV U20043 ( .A(n18596), .Z(n18601) );
  XOR U20044 ( .A(n18602), .B(n18603), .Z(n18596) );
  AND U20045 ( .A(n18604), .B(n18605), .Z(n18602) );
  XOR U20046 ( .A(n18603), .B(n11261), .Z(n18605) );
  XNOR U20047 ( .A(n18606), .B(n18607), .Z(n11261) );
  XNOR U20048 ( .A(n[416]), .B(n18608), .Z(n18604) );
  IV U20049 ( .A(n18603), .Z(n18608) );
  XOR U20050 ( .A(n18609), .B(n18610), .Z(n18603) );
  AND U20051 ( .A(n18611), .B(n18612), .Z(n18609) );
  XOR U20052 ( .A(n18610), .B(n11266), .Z(n18612) );
  XNOR U20053 ( .A(n18613), .B(n18614), .Z(n11266) );
  XNOR U20054 ( .A(n[415]), .B(n18615), .Z(n18611) );
  IV U20055 ( .A(n18610), .Z(n18615) );
  XOR U20056 ( .A(n18616), .B(n18617), .Z(n18610) );
  AND U20057 ( .A(n18618), .B(n18619), .Z(n18616) );
  XOR U20058 ( .A(n18617), .B(n11271), .Z(n18619) );
  XNOR U20059 ( .A(n18620), .B(n18621), .Z(n11271) );
  XNOR U20060 ( .A(n[414]), .B(n18622), .Z(n18618) );
  IV U20061 ( .A(n18617), .Z(n18622) );
  XOR U20062 ( .A(n18623), .B(n18624), .Z(n18617) );
  AND U20063 ( .A(n18625), .B(n18626), .Z(n18623) );
  XOR U20064 ( .A(n18624), .B(n11276), .Z(n18626) );
  XNOR U20065 ( .A(n18627), .B(n18628), .Z(n11276) );
  XNOR U20066 ( .A(n[413]), .B(n18629), .Z(n18625) );
  IV U20067 ( .A(n18624), .Z(n18629) );
  XOR U20068 ( .A(n18630), .B(n18631), .Z(n18624) );
  AND U20069 ( .A(n18632), .B(n18633), .Z(n18630) );
  XOR U20070 ( .A(n18631), .B(n11281), .Z(n18633) );
  XNOR U20071 ( .A(n18634), .B(n18635), .Z(n11281) );
  XNOR U20072 ( .A(n[412]), .B(n18636), .Z(n18632) );
  IV U20073 ( .A(n18631), .Z(n18636) );
  XOR U20074 ( .A(n18637), .B(n18638), .Z(n18631) );
  AND U20075 ( .A(n18639), .B(n18640), .Z(n18637) );
  XOR U20076 ( .A(n18638), .B(n11286), .Z(n18640) );
  XNOR U20077 ( .A(n18641), .B(n18642), .Z(n11286) );
  XNOR U20078 ( .A(n[411]), .B(n18643), .Z(n18639) );
  IV U20079 ( .A(n18638), .Z(n18643) );
  XOR U20080 ( .A(n18644), .B(n18645), .Z(n18638) );
  AND U20081 ( .A(n18646), .B(n18647), .Z(n18644) );
  XOR U20082 ( .A(n18645), .B(n11291), .Z(n18647) );
  XNOR U20083 ( .A(n18648), .B(n18649), .Z(n11291) );
  XNOR U20084 ( .A(n[410]), .B(n18650), .Z(n18646) );
  IV U20085 ( .A(n18645), .Z(n18650) );
  XOR U20086 ( .A(n18651), .B(n18652), .Z(n18645) );
  AND U20087 ( .A(n18653), .B(n18654), .Z(n18651) );
  XOR U20088 ( .A(n18652), .B(n11296), .Z(n18654) );
  XNOR U20089 ( .A(n18655), .B(n18656), .Z(n11296) );
  XNOR U20090 ( .A(n[409]), .B(n18657), .Z(n18653) );
  IV U20091 ( .A(n18652), .Z(n18657) );
  XOR U20092 ( .A(n18658), .B(n18659), .Z(n18652) );
  AND U20093 ( .A(n18660), .B(n18661), .Z(n18658) );
  XOR U20094 ( .A(n18659), .B(n11301), .Z(n18661) );
  XNOR U20095 ( .A(n18662), .B(n18663), .Z(n11301) );
  XNOR U20096 ( .A(n[408]), .B(n18664), .Z(n18660) );
  IV U20097 ( .A(n18659), .Z(n18664) );
  XOR U20098 ( .A(n18665), .B(n18666), .Z(n18659) );
  AND U20099 ( .A(n18667), .B(n18668), .Z(n18665) );
  XOR U20100 ( .A(n18666), .B(n11306), .Z(n18668) );
  XNOR U20101 ( .A(n18669), .B(n18670), .Z(n11306) );
  XNOR U20102 ( .A(n[407]), .B(n18671), .Z(n18667) );
  IV U20103 ( .A(n18666), .Z(n18671) );
  XOR U20104 ( .A(n18672), .B(n18673), .Z(n18666) );
  AND U20105 ( .A(n18674), .B(n18675), .Z(n18672) );
  XOR U20106 ( .A(n18673), .B(n11311), .Z(n18675) );
  XNOR U20107 ( .A(n18676), .B(n18677), .Z(n11311) );
  XNOR U20108 ( .A(n[406]), .B(n18678), .Z(n18674) );
  IV U20109 ( .A(n18673), .Z(n18678) );
  XOR U20110 ( .A(n18679), .B(n18680), .Z(n18673) );
  AND U20111 ( .A(n18681), .B(n18682), .Z(n18679) );
  XOR U20112 ( .A(n18680), .B(n11316), .Z(n18682) );
  XNOR U20113 ( .A(n18683), .B(n18684), .Z(n11316) );
  XNOR U20114 ( .A(n[405]), .B(n18685), .Z(n18681) );
  IV U20115 ( .A(n18680), .Z(n18685) );
  XOR U20116 ( .A(n18686), .B(n18687), .Z(n18680) );
  AND U20117 ( .A(n18688), .B(n18689), .Z(n18686) );
  XOR U20118 ( .A(n18687), .B(n11321), .Z(n18689) );
  XNOR U20119 ( .A(n18690), .B(n18691), .Z(n11321) );
  XNOR U20120 ( .A(n[404]), .B(n18692), .Z(n18688) );
  IV U20121 ( .A(n18687), .Z(n18692) );
  XOR U20122 ( .A(n18693), .B(n18694), .Z(n18687) );
  AND U20123 ( .A(n18695), .B(n18696), .Z(n18693) );
  XOR U20124 ( .A(n18694), .B(n11326), .Z(n18696) );
  XNOR U20125 ( .A(n18697), .B(n18698), .Z(n11326) );
  XNOR U20126 ( .A(n[403]), .B(n18699), .Z(n18695) );
  IV U20127 ( .A(n18694), .Z(n18699) );
  XOR U20128 ( .A(n18700), .B(n18701), .Z(n18694) );
  AND U20129 ( .A(n18702), .B(n18703), .Z(n18700) );
  XOR U20130 ( .A(n18701), .B(n11331), .Z(n18703) );
  XNOR U20131 ( .A(n18704), .B(n18705), .Z(n11331) );
  XNOR U20132 ( .A(n[402]), .B(n18706), .Z(n18702) );
  IV U20133 ( .A(n18701), .Z(n18706) );
  XOR U20134 ( .A(n18707), .B(n18708), .Z(n18701) );
  AND U20135 ( .A(n18709), .B(n18710), .Z(n18707) );
  XOR U20136 ( .A(n18708), .B(n11336), .Z(n18710) );
  XNOR U20137 ( .A(n18711), .B(n18712), .Z(n11336) );
  XNOR U20138 ( .A(n[401]), .B(n18713), .Z(n18709) );
  IV U20139 ( .A(n18708), .Z(n18713) );
  XOR U20140 ( .A(n18714), .B(n18715), .Z(n18708) );
  AND U20141 ( .A(n18716), .B(n18717), .Z(n18714) );
  XOR U20142 ( .A(n18715), .B(n11341), .Z(n18717) );
  XNOR U20143 ( .A(n18718), .B(n18719), .Z(n11341) );
  XNOR U20144 ( .A(n[400]), .B(n18720), .Z(n18716) );
  IV U20145 ( .A(n18715), .Z(n18720) );
  XOR U20146 ( .A(n18721), .B(n18722), .Z(n18715) );
  AND U20147 ( .A(n18723), .B(n18724), .Z(n18721) );
  XOR U20148 ( .A(n18722), .B(n11346), .Z(n18724) );
  XNOR U20149 ( .A(n18725), .B(n18726), .Z(n11346) );
  XNOR U20150 ( .A(n[399]), .B(n18727), .Z(n18723) );
  IV U20151 ( .A(n18722), .Z(n18727) );
  XOR U20152 ( .A(n18728), .B(n18729), .Z(n18722) );
  AND U20153 ( .A(n18730), .B(n18731), .Z(n18728) );
  XOR U20154 ( .A(n18729), .B(n11351), .Z(n18731) );
  XNOR U20155 ( .A(n18732), .B(n18733), .Z(n11351) );
  XNOR U20156 ( .A(n[398]), .B(n18734), .Z(n18730) );
  IV U20157 ( .A(n18729), .Z(n18734) );
  XOR U20158 ( .A(n18735), .B(n18736), .Z(n18729) );
  AND U20159 ( .A(n18737), .B(n18738), .Z(n18735) );
  XOR U20160 ( .A(n18736), .B(n11356), .Z(n18738) );
  XNOR U20161 ( .A(n18739), .B(n18740), .Z(n11356) );
  XNOR U20162 ( .A(n[397]), .B(n18741), .Z(n18737) );
  IV U20163 ( .A(n18736), .Z(n18741) );
  XOR U20164 ( .A(n18742), .B(n18743), .Z(n18736) );
  AND U20165 ( .A(n18744), .B(n18745), .Z(n18742) );
  XOR U20166 ( .A(n18743), .B(n11361), .Z(n18745) );
  XNOR U20167 ( .A(n18746), .B(n18747), .Z(n11361) );
  XNOR U20168 ( .A(n[396]), .B(n18748), .Z(n18744) );
  IV U20169 ( .A(n18743), .Z(n18748) );
  XOR U20170 ( .A(n18749), .B(n18750), .Z(n18743) );
  AND U20171 ( .A(n18751), .B(n18752), .Z(n18749) );
  XOR U20172 ( .A(n18750), .B(n11366), .Z(n18752) );
  XNOR U20173 ( .A(n18753), .B(n18754), .Z(n11366) );
  XNOR U20174 ( .A(n[395]), .B(n18755), .Z(n18751) );
  IV U20175 ( .A(n18750), .Z(n18755) );
  XOR U20176 ( .A(n18756), .B(n18757), .Z(n18750) );
  AND U20177 ( .A(n18758), .B(n18759), .Z(n18756) );
  XOR U20178 ( .A(n18757), .B(n11371), .Z(n18759) );
  XNOR U20179 ( .A(n18760), .B(n18761), .Z(n11371) );
  XNOR U20180 ( .A(n[394]), .B(n18762), .Z(n18758) );
  IV U20181 ( .A(n18757), .Z(n18762) );
  XOR U20182 ( .A(n18763), .B(n18764), .Z(n18757) );
  AND U20183 ( .A(n18765), .B(n18766), .Z(n18763) );
  XOR U20184 ( .A(n18764), .B(n11376), .Z(n18766) );
  XNOR U20185 ( .A(n18767), .B(n18768), .Z(n11376) );
  XNOR U20186 ( .A(n[393]), .B(n18769), .Z(n18765) );
  IV U20187 ( .A(n18764), .Z(n18769) );
  XOR U20188 ( .A(n18770), .B(n18771), .Z(n18764) );
  AND U20189 ( .A(n18772), .B(n18773), .Z(n18770) );
  XOR U20190 ( .A(n18771), .B(n11381), .Z(n18773) );
  XNOR U20191 ( .A(n18774), .B(n18775), .Z(n11381) );
  XNOR U20192 ( .A(n[392]), .B(n18776), .Z(n18772) );
  IV U20193 ( .A(n18771), .Z(n18776) );
  XOR U20194 ( .A(n18777), .B(n18778), .Z(n18771) );
  AND U20195 ( .A(n18779), .B(n18780), .Z(n18777) );
  XOR U20196 ( .A(n18778), .B(n11386), .Z(n18780) );
  XNOR U20197 ( .A(n18781), .B(n18782), .Z(n11386) );
  XNOR U20198 ( .A(n[391]), .B(n18783), .Z(n18779) );
  IV U20199 ( .A(n18778), .Z(n18783) );
  XOR U20200 ( .A(n18784), .B(n18785), .Z(n18778) );
  AND U20201 ( .A(n18786), .B(n18787), .Z(n18784) );
  XOR U20202 ( .A(n18785), .B(n11391), .Z(n18787) );
  XNOR U20203 ( .A(n18788), .B(n18789), .Z(n11391) );
  XNOR U20204 ( .A(n[390]), .B(n18790), .Z(n18786) );
  IV U20205 ( .A(n18785), .Z(n18790) );
  XOR U20206 ( .A(n18791), .B(n18792), .Z(n18785) );
  AND U20207 ( .A(n18793), .B(n18794), .Z(n18791) );
  XOR U20208 ( .A(n18792), .B(n11396), .Z(n18794) );
  XNOR U20209 ( .A(n18795), .B(n18796), .Z(n11396) );
  XNOR U20210 ( .A(n[389]), .B(n18797), .Z(n18793) );
  IV U20211 ( .A(n18792), .Z(n18797) );
  XOR U20212 ( .A(n18798), .B(n18799), .Z(n18792) );
  AND U20213 ( .A(n18800), .B(n18801), .Z(n18798) );
  XOR U20214 ( .A(n18799), .B(n11401), .Z(n18801) );
  XNOR U20215 ( .A(n18802), .B(n18803), .Z(n11401) );
  XNOR U20216 ( .A(n[388]), .B(n18804), .Z(n18800) );
  IV U20217 ( .A(n18799), .Z(n18804) );
  XOR U20218 ( .A(n18805), .B(n18806), .Z(n18799) );
  AND U20219 ( .A(n18807), .B(n18808), .Z(n18805) );
  XOR U20220 ( .A(n18806), .B(n11406), .Z(n18808) );
  XNOR U20221 ( .A(n18809), .B(n18810), .Z(n11406) );
  XNOR U20222 ( .A(n[387]), .B(n18811), .Z(n18807) );
  IV U20223 ( .A(n18806), .Z(n18811) );
  XOR U20224 ( .A(n18812), .B(n18813), .Z(n18806) );
  AND U20225 ( .A(n18814), .B(n18815), .Z(n18812) );
  XOR U20226 ( .A(n18813), .B(n11411), .Z(n18815) );
  XNOR U20227 ( .A(n18816), .B(n18817), .Z(n11411) );
  XNOR U20228 ( .A(n[386]), .B(n18818), .Z(n18814) );
  IV U20229 ( .A(n18813), .Z(n18818) );
  XOR U20230 ( .A(n18819), .B(n18820), .Z(n18813) );
  AND U20231 ( .A(n18821), .B(n18822), .Z(n18819) );
  XOR U20232 ( .A(n18820), .B(n11416), .Z(n18822) );
  XNOR U20233 ( .A(n18823), .B(n18824), .Z(n11416) );
  XNOR U20234 ( .A(n[385]), .B(n18825), .Z(n18821) );
  IV U20235 ( .A(n18820), .Z(n18825) );
  XOR U20236 ( .A(n18826), .B(n18827), .Z(n18820) );
  AND U20237 ( .A(n18828), .B(n18829), .Z(n18826) );
  XOR U20238 ( .A(n18827), .B(n11421), .Z(n18829) );
  XNOR U20239 ( .A(n18830), .B(n18831), .Z(n11421) );
  XNOR U20240 ( .A(n[384]), .B(n18832), .Z(n18828) );
  IV U20241 ( .A(n18827), .Z(n18832) );
  XOR U20242 ( .A(n18833), .B(n18834), .Z(n18827) );
  AND U20243 ( .A(n18835), .B(n18836), .Z(n18833) );
  XOR U20244 ( .A(n18834), .B(n11426), .Z(n18836) );
  XNOR U20245 ( .A(n18837), .B(n18838), .Z(n11426) );
  XNOR U20246 ( .A(n[383]), .B(n18839), .Z(n18835) );
  IV U20247 ( .A(n18834), .Z(n18839) );
  XOR U20248 ( .A(n18840), .B(n18841), .Z(n18834) );
  AND U20249 ( .A(n18842), .B(n18843), .Z(n18840) );
  XOR U20250 ( .A(n18841), .B(n11431), .Z(n18843) );
  XNOR U20251 ( .A(n18844), .B(n18845), .Z(n11431) );
  XNOR U20252 ( .A(n[382]), .B(n18846), .Z(n18842) );
  IV U20253 ( .A(n18841), .Z(n18846) );
  XOR U20254 ( .A(n18847), .B(n18848), .Z(n18841) );
  AND U20255 ( .A(n18849), .B(n18850), .Z(n18847) );
  XOR U20256 ( .A(n18848), .B(n11436), .Z(n18850) );
  XNOR U20257 ( .A(n18851), .B(n18852), .Z(n11436) );
  XNOR U20258 ( .A(n[381]), .B(n18853), .Z(n18849) );
  IV U20259 ( .A(n18848), .Z(n18853) );
  XOR U20260 ( .A(n18854), .B(n18855), .Z(n18848) );
  AND U20261 ( .A(n18856), .B(n18857), .Z(n18854) );
  XOR U20262 ( .A(n18855), .B(n11441), .Z(n18857) );
  XNOR U20263 ( .A(n18858), .B(n18859), .Z(n11441) );
  XNOR U20264 ( .A(n[380]), .B(n18860), .Z(n18856) );
  IV U20265 ( .A(n18855), .Z(n18860) );
  XOR U20266 ( .A(n18861), .B(n18862), .Z(n18855) );
  AND U20267 ( .A(n18863), .B(n18864), .Z(n18861) );
  XOR U20268 ( .A(n18862), .B(n11446), .Z(n18864) );
  XNOR U20269 ( .A(n18865), .B(n18866), .Z(n11446) );
  XNOR U20270 ( .A(n[379]), .B(n18867), .Z(n18863) );
  IV U20271 ( .A(n18862), .Z(n18867) );
  XOR U20272 ( .A(n18868), .B(n18869), .Z(n18862) );
  AND U20273 ( .A(n18870), .B(n18871), .Z(n18868) );
  XOR U20274 ( .A(n18869), .B(n11451), .Z(n18871) );
  XNOR U20275 ( .A(n18872), .B(n18873), .Z(n11451) );
  XNOR U20276 ( .A(n[378]), .B(n18874), .Z(n18870) );
  IV U20277 ( .A(n18869), .Z(n18874) );
  XOR U20278 ( .A(n18875), .B(n18876), .Z(n18869) );
  AND U20279 ( .A(n18877), .B(n18878), .Z(n18875) );
  XOR U20280 ( .A(n18876), .B(n11456), .Z(n18878) );
  XNOR U20281 ( .A(n18879), .B(n18880), .Z(n11456) );
  XNOR U20282 ( .A(n[377]), .B(n18881), .Z(n18877) );
  IV U20283 ( .A(n18876), .Z(n18881) );
  XOR U20284 ( .A(n18882), .B(n18883), .Z(n18876) );
  AND U20285 ( .A(n18884), .B(n18885), .Z(n18882) );
  XOR U20286 ( .A(n18883), .B(n11461), .Z(n18885) );
  XNOR U20287 ( .A(n18886), .B(n18887), .Z(n11461) );
  XNOR U20288 ( .A(n[376]), .B(n18888), .Z(n18884) );
  IV U20289 ( .A(n18883), .Z(n18888) );
  XOR U20290 ( .A(n18889), .B(n18890), .Z(n18883) );
  AND U20291 ( .A(n18891), .B(n18892), .Z(n18889) );
  XOR U20292 ( .A(n18890), .B(n11466), .Z(n18892) );
  XNOR U20293 ( .A(n18893), .B(n18894), .Z(n11466) );
  XNOR U20294 ( .A(n[375]), .B(n18895), .Z(n18891) );
  IV U20295 ( .A(n18890), .Z(n18895) );
  XOR U20296 ( .A(n18896), .B(n18897), .Z(n18890) );
  AND U20297 ( .A(n18898), .B(n18899), .Z(n18896) );
  XOR U20298 ( .A(n18897), .B(n11471), .Z(n18899) );
  XNOR U20299 ( .A(n18900), .B(n18901), .Z(n11471) );
  XNOR U20300 ( .A(n[374]), .B(n18902), .Z(n18898) );
  IV U20301 ( .A(n18897), .Z(n18902) );
  XOR U20302 ( .A(n18903), .B(n18904), .Z(n18897) );
  AND U20303 ( .A(n18905), .B(n18906), .Z(n18903) );
  XOR U20304 ( .A(n18904), .B(n11476), .Z(n18906) );
  XNOR U20305 ( .A(n18907), .B(n18908), .Z(n11476) );
  XNOR U20306 ( .A(n[373]), .B(n18909), .Z(n18905) );
  IV U20307 ( .A(n18904), .Z(n18909) );
  XOR U20308 ( .A(n18910), .B(n18911), .Z(n18904) );
  AND U20309 ( .A(n18912), .B(n18913), .Z(n18910) );
  XOR U20310 ( .A(n18911), .B(n11481), .Z(n18913) );
  XNOR U20311 ( .A(n18914), .B(n18915), .Z(n11481) );
  XNOR U20312 ( .A(n[372]), .B(n18916), .Z(n18912) );
  IV U20313 ( .A(n18911), .Z(n18916) );
  XOR U20314 ( .A(n18917), .B(n18918), .Z(n18911) );
  AND U20315 ( .A(n18919), .B(n18920), .Z(n18917) );
  XOR U20316 ( .A(n18918), .B(n11486), .Z(n18920) );
  XNOR U20317 ( .A(n18921), .B(n18922), .Z(n11486) );
  XNOR U20318 ( .A(n[371]), .B(n18923), .Z(n18919) );
  IV U20319 ( .A(n18918), .Z(n18923) );
  XOR U20320 ( .A(n18924), .B(n18925), .Z(n18918) );
  AND U20321 ( .A(n18926), .B(n18927), .Z(n18924) );
  XOR U20322 ( .A(n18925), .B(n11491), .Z(n18927) );
  XNOR U20323 ( .A(n18928), .B(n18929), .Z(n11491) );
  XNOR U20324 ( .A(n[370]), .B(n18930), .Z(n18926) );
  IV U20325 ( .A(n18925), .Z(n18930) );
  XOR U20326 ( .A(n18931), .B(n18932), .Z(n18925) );
  AND U20327 ( .A(n18933), .B(n18934), .Z(n18931) );
  XOR U20328 ( .A(n18932), .B(n11496), .Z(n18934) );
  XNOR U20329 ( .A(n18935), .B(n18936), .Z(n11496) );
  XNOR U20330 ( .A(n[369]), .B(n18937), .Z(n18933) );
  IV U20331 ( .A(n18932), .Z(n18937) );
  XOR U20332 ( .A(n18938), .B(n18939), .Z(n18932) );
  AND U20333 ( .A(n18940), .B(n18941), .Z(n18938) );
  XOR U20334 ( .A(n18939), .B(n11501), .Z(n18941) );
  XNOR U20335 ( .A(n18942), .B(n18943), .Z(n11501) );
  XNOR U20336 ( .A(n[368]), .B(n18944), .Z(n18940) );
  IV U20337 ( .A(n18939), .Z(n18944) );
  XOR U20338 ( .A(n18945), .B(n18946), .Z(n18939) );
  AND U20339 ( .A(n18947), .B(n18948), .Z(n18945) );
  XOR U20340 ( .A(n18946), .B(n11506), .Z(n18948) );
  XNOR U20341 ( .A(n18949), .B(n18950), .Z(n11506) );
  XNOR U20342 ( .A(n[367]), .B(n18951), .Z(n18947) );
  IV U20343 ( .A(n18946), .Z(n18951) );
  XOR U20344 ( .A(n18952), .B(n18953), .Z(n18946) );
  AND U20345 ( .A(n18954), .B(n18955), .Z(n18952) );
  XOR U20346 ( .A(n18953), .B(n11511), .Z(n18955) );
  XNOR U20347 ( .A(n18956), .B(n18957), .Z(n11511) );
  XNOR U20348 ( .A(n[366]), .B(n18958), .Z(n18954) );
  IV U20349 ( .A(n18953), .Z(n18958) );
  XOR U20350 ( .A(n18959), .B(n18960), .Z(n18953) );
  AND U20351 ( .A(n18961), .B(n18962), .Z(n18959) );
  XOR U20352 ( .A(n18960), .B(n11516), .Z(n18962) );
  XNOR U20353 ( .A(n18963), .B(n18964), .Z(n11516) );
  XNOR U20354 ( .A(n[365]), .B(n18965), .Z(n18961) );
  IV U20355 ( .A(n18960), .Z(n18965) );
  XOR U20356 ( .A(n18966), .B(n18967), .Z(n18960) );
  AND U20357 ( .A(n18968), .B(n18969), .Z(n18966) );
  XOR U20358 ( .A(n18967), .B(n11521), .Z(n18969) );
  XNOR U20359 ( .A(n18970), .B(n18971), .Z(n11521) );
  XNOR U20360 ( .A(n[364]), .B(n18972), .Z(n18968) );
  IV U20361 ( .A(n18967), .Z(n18972) );
  XOR U20362 ( .A(n18973), .B(n18974), .Z(n18967) );
  AND U20363 ( .A(n18975), .B(n18976), .Z(n18973) );
  XOR U20364 ( .A(n18974), .B(n11526), .Z(n18976) );
  XNOR U20365 ( .A(n18977), .B(n18978), .Z(n11526) );
  XNOR U20366 ( .A(n[363]), .B(n18979), .Z(n18975) );
  IV U20367 ( .A(n18974), .Z(n18979) );
  XOR U20368 ( .A(n18980), .B(n18981), .Z(n18974) );
  AND U20369 ( .A(n18982), .B(n18983), .Z(n18980) );
  XOR U20370 ( .A(n18981), .B(n11531), .Z(n18983) );
  XNOR U20371 ( .A(n18984), .B(n18985), .Z(n11531) );
  XNOR U20372 ( .A(n[362]), .B(n18986), .Z(n18982) );
  IV U20373 ( .A(n18981), .Z(n18986) );
  XOR U20374 ( .A(n18987), .B(n18988), .Z(n18981) );
  AND U20375 ( .A(n18989), .B(n18990), .Z(n18987) );
  XOR U20376 ( .A(n18988), .B(n11536), .Z(n18990) );
  XNOR U20377 ( .A(n18991), .B(n18992), .Z(n11536) );
  XNOR U20378 ( .A(n[361]), .B(n18993), .Z(n18989) );
  IV U20379 ( .A(n18988), .Z(n18993) );
  XOR U20380 ( .A(n18994), .B(n18995), .Z(n18988) );
  AND U20381 ( .A(n18996), .B(n18997), .Z(n18994) );
  XOR U20382 ( .A(n18995), .B(n11541), .Z(n18997) );
  XNOR U20383 ( .A(n18998), .B(n18999), .Z(n11541) );
  XNOR U20384 ( .A(n[360]), .B(n19000), .Z(n18996) );
  IV U20385 ( .A(n18995), .Z(n19000) );
  XOR U20386 ( .A(n19001), .B(n19002), .Z(n18995) );
  AND U20387 ( .A(n19003), .B(n19004), .Z(n19001) );
  XOR U20388 ( .A(n19002), .B(n11546), .Z(n19004) );
  XNOR U20389 ( .A(n19005), .B(n19006), .Z(n11546) );
  XNOR U20390 ( .A(n[359]), .B(n19007), .Z(n19003) );
  IV U20391 ( .A(n19002), .Z(n19007) );
  XOR U20392 ( .A(n19008), .B(n19009), .Z(n19002) );
  AND U20393 ( .A(n19010), .B(n19011), .Z(n19008) );
  XOR U20394 ( .A(n19009), .B(n11551), .Z(n19011) );
  XNOR U20395 ( .A(n19012), .B(n19013), .Z(n11551) );
  XNOR U20396 ( .A(n[358]), .B(n19014), .Z(n19010) );
  IV U20397 ( .A(n19009), .Z(n19014) );
  XOR U20398 ( .A(n19015), .B(n19016), .Z(n19009) );
  AND U20399 ( .A(n19017), .B(n19018), .Z(n19015) );
  XOR U20400 ( .A(n19016), .B(n11556), .Z(n19018) );
  XNOR U20401 ( .A(n19019), .B(n19020), .Z(n11556) );
  XNOR U20402 ( .A(n[357]), .B(n19021), .Z(n19017) );
  IV U20403 ( .A(n19016), .Z(n19021) );
  XOR U20404 ( .A(n19022), .B(n19023), .Z(n19016) );
  AND U20405 ( .A(n19024), .B(n19025), .Z(n19022) );
  XOR U20406 ( .A(n19023), .B(n11561), .Z(n19025) );
  XNOR U20407 ( .A(n19026), .B(n19027), .Z(n11561) );
  XNOR U20408 ( .A(n[356]), .B(n19028), .Z(n19024) );
  IV U20409 ( .A(n19023), .Z(n19028) );
  XOR U20410 ( .A(n19029), .B(n19030), .Z(n19023) );
  AND U20411 ( .A(n19031), .B(n19032), .Z(n19029) );
  XOR U20412 ( .A(n19030), .B(n11566), .Z(n19032) );
  XNOR U20413 ( .A(n19033), .B(n19034), .Z(n11566) );
  XNOR U20414 ( .A(n[355]), .B(n19035), .Z(n19031) );
  IV U20415 ( .A(n19030), .Z(n19035) );
  XOR U20416 ( .A(n19036), .B(n19037), .Z(n19030) );
  AND U20417 ( .A(n19038), .B(n19039), .Z(n19036) );
  XOR U20418 ( .A(n19037), .B(n11571), .Z(n19039) );
  XNOR U20419 ( .A(n19040), .B(n19041), .Z(n11571) );
  XNOR U20420 ( .A(n[354]), .B(n19042), .Z(n19038) );
  IV U20421 ( .A(n19037), .Z(n19042) );
  XOR U20422 ( .A(n19043), .B(n19044), .Z(n19037) );
  AND U20423 ( .A(n19045), .B(n19046), .Z(n19043) );
  XOR U20424 ( .A(n19044), .B(n11576), .Z(n19046) );
  XNOR U20425 ( .A(n19047), .B(n19048), .Z(n11576) );
  XNOR U20426 ( .A(n[353]), .B(n19049), .Z(n19045) );
  IV U20427 ( .A(n19044), .Z(n19049) );
  XOR U20428 ( .A(n19050), .B(n19051), .Z(n19044) );
  AND U20429 ( .A(n19052), .B(n19053), .Z(n19050) );
  XOR U20430 ( .A(n19051), .B(n11581), .Z(n19053) );
  XNOR U20431 ( .A(n19054), .B(n19055), .Z(n11581) );
  XNOR U20432 ( .A(n[352]), .B(n19056), .Z(n19052) );
  IV U20433 ( .A(n19051), .Z(n19056) );
  XOR U20434 ( .A(n19057), .B(n19058), .Z(n19051) );
  AND U20435 ( .A(n19059), .B(n19060), .Z(n19057) );
  XOR U20436 ( .A(n19058), .B(n11586), .Z(n19060) );
  XNOR U20437 ( .A(n19061), .B(n19062), .Z(n11586) );
  XNOR U20438 ( .A(n[351]), .B(n19063), .Z(n19059) );
  IV U20439 ( .A(n19058), .Z(n19063) );
  XOR U20440 ( .A(n19064), .B(n19065), .Z(n19058) );
  AND U20441 ( .A(n19066), .B(n19067), .Z(n19064) );
  XOR U20442 ( .A(n19065), .B(n11591), .Z(n19067) );
  XNOR U20443 ( .A(n19068), .B(n19069), .Z(n11591) );
  XNOR U20444 ( .A(n[350]), .B(n19070), .Z(n19066) );
  IV U20445 ( .A(n19065), .Z(n19070) );
  XOR U20446 ( .A(n19071), .B(n19072), .Z(n19065) );
  AND U20447 ( .A(n19073), .B(n19074), .Z(n19071) );
  XOR U20448 ( .A(n19072), .B(n11596), .Z(n19074) );
  XNOR U20449 ( .A(n19075), .B(n19076), .Z(n11596) );
  XNOR U20450 ( .A(n[349]), .B(n19077), .Z(n19073) );
  IV U20451 ( .A(n19072), .Z(n19077) );
  XOR U20452 ( .A(n19078), .B(n19079), .Z(n19072) );
  AND U20453 ( .A(n19080), .B(n19081), .Z(n19078) );
  XOR U20454 ( .A(n19079), .B(n11601), .Z(n19081) );
  XNOR U20455 ( .A(n19082), .B(n19083), .Z(n11601) );
  XNOR U20456 ( .A(n[348]), .B(n19084), .Z(n19080) );
  IV U20457 ( .A(n19079), .Z(n19084) );
  XOR U20458 ( .A(n19085), .B(n19086), .Z(n19079) );
  AND U20459 ( .A(n19087), .B(n19088), .Z(n19085) );
  XOR U20460 ( .A(n19086), .B(n11606), .Z(n19088) );
  XNOR U20461 ( .A(n19089), .B(n19090), .Z(n11606) );
  XNOR U20462 ( .A(n[347]), .B(n19091), .Z(n19087) );
  IV U20463 ( .A(n19086), .Z(n19091) );
  XOR U20464 ( .A(n19092), .B(n19093), .Z(n19086) );
  AND U20465 ( .A(n19094), .B(n19095), .Z(n19092) );
  XOR U20466 ( .A(n19093), .B(n11611), .Z(n19095) );
  XNOR U20467 ( .A(n19096), .B(n19097), .Z(n11611) );
  XNOR U20468 ( .A(n[346]), .B(n19098), .Z(n19094) );
  IV U20469 ( .A(n19093), .Z(n19098) );
  XOR U20470 ( .A(n19099), .B(n19100), .Z(n19093) );
  AND U20471 ( .A(n19101), .B(n19102), .Z(n19099) );
  XOR U20472 ( .A(n19100), .B(n11616), .Z(n19102) );
  XNOR U20473 ( .A(n19103), .B(n19104), .Z(n11616) );
  XNOR U20474 ( .A(n[345]), .B(n19105), .Z(n19101) );
  IV U20475 ( .A(n19100), .Z(n19105) );
  XOR U20476 ( .A(n19106), .B(n19107), .Z(n19100) );
  AND U20477 ( .A(n19108), .B(n19109), .Z(n19106) );
  XOR U20478 ( .A(n19107), .B(n11621), .Z(n19109) );
  XNOR U20479 ( .A(n19110), .B(n19111), .Z(n11621) );
  XNOR U20480 ( .A(n[344]), .B(n19112), .Z(n19108) );
  IV U20481 ( .A(n19107), .Z(n19112) );
  XOR U20482 ( .A(n19113), .B(n19114), .Z(n19107) );
  AND U20483 ( .A(n19115), .B(n19116), .Z(n19113) );
  XOR U20484 ( .A(n19114), .B(n11626), .Z(n19116) );
  XNOR U20485 ( .A(n19117), .B(n19118), .Z(n11626) );
  XNOR U20486 ( .A(n[343]), .B(n19119), .Z(n19115) );
  IV U20487 ( .A(n19114), .Z(n19119) );
  XOR U20488 ( .A(n19120), .B(n19121), .Z(n19114) );
  AND U20489 ( .A(n19122), .B(n19123), .Z(n19120) );
  XOR U20490 ( .A(n19121), .B(n11631), .Z(n19123) );
  XNOR U20491 ( .A(n19124), .B(n19125), .Z(n11631) );
  XNOR U20492 ( .A(n[342]), .B(n19126), .Z(n19122) );
  IV U20493 ( .A(n19121), .Z(n19126) );
  XOR U20494 ( .A(n19127), .B(n19128), .Z(n19121) );
  AND U20495 ( .A(n19129), .B(n19130), .Z(n19127) );
  XOR U20496 ( .A(n19128), .B(n11636), .Z(n19130) );
  XNOR U20497 ( .A(n19131), .B(n19132), .Z(n11636) );
  XNOR U20498 ( .A(n[341]), .B(n19133), .Z(n19129) );
  IV U20499 ( .A(n19128), .Z(n19133) );
  XOR U20500 ( .A(n19134), .B(n19135), .Z(n19128) );
  AND U20501 ( .A(n19136), .B(n19137), .Z(n19134) );
  XOR U20502 ( .A(n19135), .B(n11641), .Z(n19137) );
  XNOR U20503 ( .A(n19138), .B(n19139), .Z(n11641) );
  XNOR U20504 ( .A(n[340]), .B(n19140), .Z(n19136) );
  IV U20505 ( .A(n19135), .Z(n19140) );
  XOR U20506 ( .A(n19141), .B(n19142), .Z(n19135) );
  AND U20507 ( .A(n19143), .B(n19144), .Z(n19141) );
  XOR U20508 ( .A(n19142), .B(n11646), .Z(n19144) );
  XNOR U20509 ( .A(n19145), .B(n19146), .Z(n11646) );
  XNOR U20510 ( .A(n[339]), .B(n19147), .Z(n19143) );
  IV U20511 ( .A(n19142), .Z(n19147) );
  XOR U20512 ( .A(n19148), .B(n19149), .Z(n19142) );
  AND U20513 ( .A(n19150), .B(n19151), .Z(n19148) );
  XOR U20514 ( .A(n19149), .B(n11651), .Z(n19151) );
  XNOR U20515 ( .A(n19152), .B(n19153), .Z(n11651) );
  XNOR U20516 ( .A(n[338]), .B(n19154), .Z(n19150) );
  IV U20517 ( .A(n19149), .Z(n19154) );
  XOR U20518 ( .A(n19155), .B(n19156), .Z(n19149) );
  AND U20519 ( .A(n19157), .B(n19158), .Z(n19155) );
  XOR U20520 ( .A(n19156), .B(n11656), .Z(n19158) );
  XNOR U20521 ( .A(n19159), .B(n19160), .Z(n11656) );
  XNOR U20522 ( .A(n[337]), .B(n19161), .Z(n19157) );
  IV U20523 ( .A(n19156), .Z(n19161) );
  XOR U20524 ( .A(n19162), .B(n19163), .Z(n19156) );
  AND U20525 ( .A(n19164), .B(n19165), .Z(n19162) );
  XOR U20526 ( .A(n19163), .B(n11661), .Z(n19165) );
  XNOR U20527 ( .A(n19166), .B(n19167), .Z(n11661) );
  XNOR U20528 ( .A(n[336]), .B(n19168), .Z(n19164) );
  IV U20529 ( .A(n19163), .Z(n19168) );
  XOR U20530 ( .A(n19169), .B(n19170), .Z(n19163) );
  AND U20531 ( .A(n19171), .B(n19172), .Z(n19169) );
  XOR U20532 ( .A(n19170), .B(n11666), .Z(n19172) );
  XNOR U20533 ( .A(n19173), .B(n19174), .Z(n11666) );
  XNOR U20534 ( .A(n[335]), .B(n19175), .Z(n19171) );
  IV U20535 ( .A(n19170), .Z(n19175) );
  XOR U20536 ( .A(n19176), .B(n19177), .Z(n19170) );
  AND U20537 ( .A(n19178), .B(n19179), .Z(n19176) );
  XOR U20538 ( .A(n19177), .B(n11671), .Z(n19179) );
  XNOR U20539 ( .A(n19180), .B(n19181), .Z(n11671) );
  XNOR U20540 ( .A(n[334]), .B(n19182), .Z(n19178) );
  IV U20541 ( .A(n19177), .Z(n19182) );
  XOR U20542 ( .A(n19183), .B(n19184), .Z(n19177) );
  AND U20543 ( .A(n19185), .B(n19186), .Z(n19183) );
  XOR U20544 ( .A(n19184), .B(n11676), .Z(n19186) );
  XNOR U20545 ( .A(n19187), .B(n19188), .Z(n11676) );
  XNOR U20546 ( .A(n[333]), .B(n19189), .Z(n19185) );
  IV U20547 ( .A(n19184), .Z(n19189) );
  XOR U20548 ( .A(n19190), .B(n19191), .Z(n19184) );
  AND U20549 ( .A(n19192), .B(n19193), .Z(n19190) );
  XOR U20550 ( .A(n19191), .B(n11681), .Z(n19193) );
  XNOR U20551 ( .A(n19194), .B(n19195), .Z(n11681) );
  XNOR U20552 ( .A(n[332]), .B(n19196), .Z(n19192) );
  IV U20553 ( .A(n19191), .Z(n19196) );
  XOR U20554 ( .A(n19197), .B(n19198), .Z(n19191) );
  AND U20555 ( .A(n19199), .B(n19200), .Z(n19197) );
  XOR U20556 ( .A(n19198), .B(n11686), .Z(n19200) );
  XNOR U20557 ( .A(n19201), .B(n19202), .Z(n11686) );
  XNOR U20558 ( .A(n[331]), .B(n19203), .Z(n19199) );
  IV U20559 ( .A(n19198), .Z(n19203) );
  XOR U20560 ( .A(n19204), .B(n19205), .Z(n19198) );
  AND U20561 ( .A(n19206), .B(n19207), .Z(n19204) );
  XOR U20562 ( .A(n19205), .B(n11691), .Z(n19207) );
  XNOR U20563 ( .A(n19208), .B(n19209), .Z(n11691) );
  XNOR U20564 ( .A(n[330]), .B(n19210), .Z(n19206) );
  IV U20565 ( .A(n19205), .Z(n19210) );
  XOR U20566 ( .A(n19211), .B(n19212), .Z(n19205) );
  AND U20567 ( .A(n19213), .B(n19214), .Z(n19211) );
  XOR U20568 ( .A(n19212), .B(n11696), .Z(n19214) );
  XNOR U20569 ( .A(n19215), .B(n19216), .Z(n11696) );
  XNOR U20570 ( .A(n[329]), .B(n19217), .Z(n19213) );
  IV U20571 ( .A(n19212), .Z(n19217) );
  XOR U20572 ( .A(n19218), .B(n19219), .Z(n19212) );
  AND U20573 ( .A(n19220), .B(n19221), .Z(n19218) );
  XOR U20574 ( .A(n19219), .B(n11701), .Z(n19221) );
  XNOR U20575 ( .A(n19222), .B(n19223), .Z(n11701) );
  XNOR U20576 ( .A(n[328]), .B(n19224), .Z(n19220) );
  IV U20577 ( .A(n19219), .Z(n19224) );
  XOR U20578 ( .A(n19225), .B(n19226), .Z(n19219) );
  AND U20579 ( .A(n19227), .B(n19228), .Z(n19225) );
  XOR U20580 ( .A(n19226), .B(n11706), .Z(n19228) );
  XNOR U20581 ( .A(n19229), .B(n19230), .Z(n11706) );
  XNOR U20582 ( .A(n[327]), .B(n19231), .Z(n19227) );
  IV U20583 ( .A(n19226), .Z(n19231) );
  XOR U20584 ( .A(n19232), .B(n19233), .Z(n19226) );
  AND U20585 ( .A(n19234), .B(n19235), .Z(n19232) );
  XOR U20586 ( .A(n19233), .B(n11711), .Z(n19235) );
  XNOR U20587 ( .A(n19236), .B(n19237), .Z(n11711) );
  XNOR U20588 ( .A(n[326]), .B(n19238), .Z(n19234) );
  IV U20589 ( .A(n19233), .Z(n19238) );
  XOR U20590 ( .A(n19239), .B(n19240), .Z(n19233) );
  AND U20591 ( .A(n19241), .B(n19242), .Z(n19239) );
  XOR U20592 ( .A(n19240), .B(n11716), .Z(n19242) );
  XNOR U20593 ( .A(n19243), .B(n19244), .Z(n11716) );
  XNOR U20594 ( .A(n[325]), .B(n19245), .Z(n19241) );
  IV U20595 ( .A(n19240), .Z(n19245) );
  XOR U20596 ( .A(n19246), .B(n19247), .Z(n19240) );
  AND U20597 ( .A(n19248), .B(n19249), .Z(n19246) );
  XOR U20598 ( .A(n19247), .B(n11721), .Z(n19249) );
  XNOR U20599 ( .A(n19250), .B(n19251), .Z(n11721) );
  XNOR U20600 ( .A(n[324]), .B(n19252), .Z(n19248) );
  IV U20601 ( .A(n19247), .Z(n19252) );
  XOR U20602 ( .A(n19253), .B(n19254), .Z(n19247) );
  AND U20603 ( .A(n19255), .B(n19256), .Z(n19253) );
  XOR U20604 ( .A(n19254), .B(n11726), .Z(n19256) );
  XNOR U20605 ( .A(n19257), .B(n19258), .Z(n11726) );
  XNOR U20606 ( .A(n[323]), .B(n19259), .Z(n19255) );
  IV U20607 ( .A(n19254), .Z(n19259) );
  XOR U20608 ( .A(n19260), .B(n19261), .Z(n19254) );
  AND U20609 ( .A(n19262), .B(n19263), .Z(n19260) );
  XOR U20610 ( .A(n19261), .B(n11731), .Z(n19263) );
  XNOR U20611 ( .A(n19264), .B(n19265), .Z(n11731) );
  XNOR U20612 ( .A(n[322]), .B(n19266), .Z(n19262) );
  IV U20613 ( .A(n19261), .Z(n19266) );
  XOR U20614 ( .A(n19267), .B(n19268), .Z(n19261) );
  AND U20615 ( .A(n19269), .B(n19270), .Z(n19267) );
  XOR U20616 ( .A(n19268), .B(n11736), .Z(n19270) );
  XNOR U20617 ( .A(n19271), .B(n19272), .Z(n11736) );
  XNOR U20618 ( .A(n[321]), .B(n19273), .Z(n19269) );
  IV U20619 ( .A(n19268), .Z(n19273) );
  XOR U20620 ( .A(n19274), .B(n19275), .Z(n19268) );
  AND U20621 ( .A(n19276), .B(n19277), .Z(n19274) );
  XOR U20622 ( .A(n19275), .B(n11741), .Z(n19277) );
  XNOR U20623 ( .A(n19278), .B(n19279), .Z(n11741) );
  XNOR U20624 ( .A(n[320]), .B(n19280), .Z(n19276) );
  IV U20625 ( .A(n19275), .Z(n19280) );
  XOR U20626 ( .A(n19281), .B(n19282), .Z(n19275) );
  AND U20627 ( .A(n19283), .B(n19284), .Z(n19281) );
  XOR U20628 ( .A(n19282), .B(n11746), .Z(n19284) );
  XNOR U20629 ( .A(n19285), .B(n19286), .Z(n11746) );
  XNOR U20630 ( .A(n[319]), .B(n19287), .Z(n19283) );
  IV U20631 ( .A(n19282), .Z(n19287) );
  XOR U20632 ( .A(n19288), .B(n19289), .Z(n19282) );
  AND U20633 ( .A(n19290), .B(n19291), .Z(n19288) );
  XOR U20634 ( .A(n19289), .B(n11751), .Z(n19291) );
  XNOR U20635 ( .A(n19292), .B(n19293), .Z(n11751) );
  XNOR U20636 ( .A(n[318]), .B(n19294), .Z(n19290) );
  IV U20637 ( .A(n19289), .Z(n19294) );
  XOR U20638 ( .A(n19295), .B(n19296), .Z(n19289) );
  AND U20639 ( .A(n19297), .B(n19298), .Z(n19295) );
  XOR U20640 ( .A(n19296), .B(n11756), .Z(n19298) );
  XNOR U20641 ( .A(n19299), .B(n19300), .Z(n11756) );
  XNOR U20642 ( .A(n[317]), .B(n19301), .Z(n19297) );
  IV U20643 ( .A(n19296), .Z(n19301) );
  XOR U20644 ( .A(n19302), .B(n19303), .Z(n19296) );
  AND U20645 ( .A(n19304), .B(n19305), .Z(n19302) );
  XOR U20646 ( .A(n19303), .B(n11761), .Z(n19305) );
  XNOR U20647 ( .A(n19306), .B(n19307), .Z(n11761) );
  XNOR U20648 ( .A(n[316]), .B(n19308), .Z(n19304) );
  IV U20649 ( .A(n19303), .Z(n19308) );
  XOR U20650 ( .A(n19309), .B(n19310), .Z(n19303) );
  AND U20651 ( .A(n19311), .B(n19312), .Z(n19309) );
  XOR U20652 ( .A(n19310), .B(n11766), .Z(n19312) );
  XNOR U20653 ( .A(n19313), .B(n19314), .Z(n11766) );
  XNOR U20654 ( .A(n[315]), .B(n19315), .Z(n19311) );
  IV U20655 ( .A(n19310), .Z(n19315) );
  XOR U20656 ( .A(n19316), .B(n19317), .Z(n19310) );
  AND U20657 ( .A(n19318), .B(n19319), .Z(n19316) );
  XOR U20658 ( .A(n19317), .B(n11771), .Z(n19319) );
  XNOR U20659 ( .A(n19320), .B(n19321), .Z(n11771) );
  XNOR U20660 ( .A(n[314]), .B(n19322), .Z(n19318) );
  IV U20661 ( .A(n19317), .Z(n19322) );
  XOR U20662 ( .A(n19323), .B(n19324), .Z(n19317) );
  AND U20663 ( .A(n19325), .B(n19326), .Z(n19323) );
  XOR U20664 ( .A(n19324), .B(n11776), .Z(n19326) );
  XNOR U20665 ( .A(n19327), .B(n19328), .Z(n11776) );
  XNOR U20666 ( .A(n[313]), .B(n19329), .Z(n19325) );
  IV U20667 ( .A(n19324), .Z(n19329) );
  XOR U20668 ( .A(n19330), .B(n19331), .Z(n19324) );
  AND U20669 ( .A(n19332), .B(n19333), .Z(n19330) );
  XOR U20670 ( .A(n19331), .B(n11781), .Z(n19333) );
  XNOR U20671 ( .A(n19334), .B(n19335), .Z(n11781) );
  XNOR U20672 ( .A(n[312]), .B(n19336), .Z(n19332) );
  IV U20673 ( .A(n19331), .Z(n19336) );
  XOR U20674 ( .A(n19337), .B(n19338), .Z(n19331) );
  AND U20675 ( .A(n19339), .B(n19340), .Z(n19337) );
  XOR U20676 ( .A(n19338), .B(n11786), .Z(n19340) );
  XNOR U20677 ( .A(n19341), .B(n19342), .Z(n11786) );
  XNOR U20678 ( .A(n[311]), .B(n19343), .Z(n19339) );
  IV U20679 ( .A(n19338), .Z(n19343) );
  XOR U20680 ( .A(n19344), .B(n19345), .Z(n19338) );
  AND U20681 ( .A(n19346), .B(n19347), .Z(n19344) );
  XOR U20682 ( .A(n19345), .B(n11791), .Z(n19347) );
  XNOR U20683 ( .A(n19348), .B(n19349), .Z(n11791) );
  XNOR U20684 ( .A(n[310]), .B(n19350), .Z(n19346) );
  IV U20685 ( .A(n19345), .Z(n19350) );
  XOR U20686 ( .A(n19351), .B(n19352), .Z(n19345) );
  AND U20687 ( .A(n19353), .B(n19354), .Z(n19351) );
  XOR U20688 ( .A(n19352), .B(n11796), .Z(n19354) );
  XNOR U20689 ( .A(n19355), .B(n19356), .Z(n11796) );
  XNOR U20690 ( .A(n[309]), .B(n19357), .Z(n19353) );
  IV U20691 ( .A(n19352), .Z(n19357) );
  XOR U20692 ( .A(n19358), .B(n19359), .Z(n19352) );
  AND U20693 ( .A(n19360), .B(n19361), .Z(n19358) );
  XOR U20694 ( .A(n19359), .B(n11801), .Z(n19361) );
  XNOR U20695 ( .A(n19362), .B(n19363), .Z(n11801) );
  XNOR U20696 ( .A(n[308]), .B(n19364), .Z(n19360) );
  IV U20697 ( .A(n19359), .Z(n19364) );
  XOR U20698 ( .A(n19365), .B(n19366), .Z(n19359) );
  AND U20699 ( .A(n19367), .B(n19368), .Z(n19365) );
  XOR U20700 ( .A(n19366), .B(n11806), .Z(n19368) );
  XNOR U20701 ( .A(n19369), .B(n19370), .Z(n11806) );
  XNOR U20702 ( .A(n[307]), .B(n19371), .Z(n19367) );
  IV U20703 ( .A(n19366), .Z(n19371) );
  XOR U20704 ( .A(n19372), .B(n19373), .Z(n19366) );
  AND U20705 ( .A(n19374), .B(n19375), .Z(n19372) );
  XOR U20706 ( .A(n19373), .B(n11811), .Z(n19375) );
  XNOR U20707 ( .A(n19376), .B(n19377), .Z(n11811) );
  XNOR U20708 ( .A(n[306]), .B(n19378), .Z(n19374) );
  IV U20709 ( .A(n19373), .Z(n19378) );
  XOR U20710 ( .A(n19379), .B(n19380), .Z(n19373) );
  AND U20711 ( .A(n19381), .B(n19382), .Z(n19379) );
  XOR U20712 ( .A(n19380), .B(n11816), .Z(n19382) );
  XNOR U20713 ( .A(n19383), .B(n19384), .Z(n11816) );
  XNOR U20714 ( .A(n[305]), .B(n19385), .Z(n19381) );
  IV U20715 ( .A(n19380), .Z(n19385) );
  XOR U20716 ( .A(n19386), .B(n19387), .Z(n19380) );
  AND U20717 ( .A(n19388), .B(n19389), .Z(n19386) );
  XOR U20718 ( .A(n19387), .B(n11821), .Z(n19389) );
  XNOR U20719 ( .A(n19390), .B(n19391), .Z(n11821) );
  XNOR U20720 ( .A(n[304]), .B(n19392), .Z(n19388) );
  IV U20721 ( .A(n19387), .Z(n19392) );
  XOR U20722 ( .A(n19393), .B(n19394), .Z(n19387) );
  AND U20723 ( .A(n19395), .B(n19396), .Z(n19393) );
  XOR U20724 ( .A(n19394), .B(n11826), .Z(n19396) );
  XNOR U20725 ( .A(n19397), .B(n19398), .Z(n11826) );
  XNOR U20726 ( .A(n[303]), .B(n19399), .Z(n19395) );
  IV U20727 ( .A(n19394), .Z(n19399) );
  XOR U20728 ( .A(n19400), .B(n19401), .Z(n19394) );
  AND U20729 ( .A(n19402), .B(n19403), .Z(n19400) );
  XOR U20730 ( .A(n19401), .B(n11831), .Z(n19403) );
  XNOR U20731 ( .A(n19404), .B(n19405), .Z(n11831) );
  XNOR U20732 ( .A(n[302]), .B(n19406), .Z(n19402) );
  IV U20733 ( .A(n19401), .Z(n19406) );
  XOR U20734 ( .A(n19407), .B(n19408), .Z(n19401) );
  AND U20735 ( .A(n19409), .B(n19410), .Z(n19407) );
  XOR U20736 ( .A(n19408), .B(n11836), .Z(n19410) );
  XNOR U20737 ( .A(n19411), .B(n19412), .Z(n11836) );
  XNOR U20738 ( .A(n[301]), .B(n19413), .Z(n19409) );
  IV U20739 ( .A(n19408), .Z(n19413) );
  XOR U20740 ( .A(n19414), .B(n19415), .Z(n19408) );
  AND U20741 ( .A(n19416), .B(n19417), .Z(n19414) );
  XOR U20742 ( .A(n19415), .B(n11841), .Z(n19417) );
  XNOR U20743 ( .A(n19418), .B(n19419), .Z(n11841) );
  XNOR U20744 ( .A(n[300]), .B(n19420), .Z(n19416) );
  IV U20745 ( .A(n19415), .Z(n19420) );
  XOR U20746 ( .A(n19421), .B(n19422), .Z(n19415) );
  AND U20747 ( .A(n19423), .B(n19424), .Z(n19421) );
  XOR U20748 ( .A(n19422), .B(n11846), .Z(n19424) );
  XNOR U20749 ( .A(n19425), .B(n19426), .Z(n11846) );
  XNOR U20750 ( .A(n[299]), .B(n19427), .Z(n19423) );
  IV U20751 ( .A(n19422), .Z(n19427) );
  XOR U20752 ( .A(n19428), .B(n19429), .Z(n19422) );
  AND U20753 ( .A(n19430), .B(n19431), .Z(n19428) );
  XOR U20754 ( .A(n19429), .B(n11851), .Z(n19431) );
  XNOR U20755 ( .A(n19432), .B(n19433), .Z(n11851) );
  XNOR U20756 ( .A(n[298]), .B(n19434), .Z(n19430) );
  IV U20757 ( .A(n19429), .Z(n19434) );
  XOR U20758 ( .A(n19435), .B(n19436), .Z(n19429) );
  AND U20759 ( .A(n19437), .B(n19438), .Z(n19435) );
  XOR U20760 ( .A(n19436), .B(n11856), .Z(n19438) );
  XNOR U20761 ( .A(n19439), .B(n19440), .Z(n11856) );
  XNOR U20762 ( .A(n[297]), .B(n19441), .Z(n19437) );
  IV U20763 ( .A(n19436), .Z(n19441) );
  XOR U20764 ( .A(n19442), .B(n19443), .Z(n19436) );
  AND U20765 ( .A(n19444), .B(n19445), .Z(n19442) );
  XOR U20766 ( .A(n19443), .B(n11861), .Z(n19445) );
  XNOR U20767 ( .A(n19446), .B(n19447), .Z(n11861) );
  XNOR U20768 ( .A(n[296]), .B(n19448), .Z(n19444) );
  IV U20769 ( .A(n19443), .Z(n19448) );
  XOR U20770 ( .A(n19449), .B(n19450), .Z(n19443) );
  AND U20771 ( .A(n19451), .B(n19452), .Z(n19449) );
  XOR U20772 ( .A(n19450), .B(n11866), .Z(n19452) );
  XNOR U20773 ( .A(n19453), .B(n19454), .Z(n11866) );
  XNOR U20774 ( .A(n[295]), .B(n19455), .Z(n19451) );
  IV U20775 ( .A(n19450), .Z(n19455) );
  XOR U20776 ( .A(n19456), .B(n19457), .Z(n19450) );
  AND U20777 ( .A(n19458), .B(n19459), .Z(n19456) );
  XOR U20778 ( .A(n19457), .B(n11871), .Z(n19459) );
  XNOR U20779 ( .A(n19460), .B(n19461), .Z(n11871) );
  XNOR U20780 ( .A(n[294]), .B(n19462), .Z(n19458) );
  IV U20781 ( .A(n19457), .Z(n19462) );
  XOR U20782 ( .A(n19463), .B(n19464), .Z(n19457) );
  AND U20783 ( .A(n19465), .B(n19466), .Z(n19463) );
  XOR U20784 ( .A(n19464), .B(n11876), .Z(n19466) );
  XNOR U20785 ( .A(n19467), .B(n19468), .Z(n11876) );
  XNOR U20786 ( .A(n[293]), .B(n19469), .Z(n19465) );
  IV U20787 ( .A(n19464), .Z(n19469) );
  XOR U20788 ( .A(n19470), .B(n19471), .Z(n19464) );
  AND U20789 ( .A(n19472), .B(n19473), .Z(n19470) );
  XOR U20790 ( .A(n19471), .B(n11881), .Z(n19473) );
  XNOR U20791 ( .A(n19474), .B(n19475), .Z(n11881) );
  XNOR U20792 ( .A(n[292]), .B(n19476), .Z(n19472) );
  IV U20793 ( .A(n19471), .Z(n19476) );
  XOR U20794 ( .A(n19477), .B(n19478), .Z(n19471) );
  AND U20795 ( .A(n19479), .B(n19480), .Z(n19477) );
  XOR U20796 ( .A(n19478), .B(n11886), .Z(n19480) );
  XNOR U20797 ( .A(n19481), .B(n19482), .Z(n11886) );
  XNOR U20798 ( .A(n[291]), .B(n19483), .Z(n19479) );
  IV U20799 ( .A(n19478), .Z(n19483) );
  XOR U20800 ( .A(n19484), .B(n19485), .Z(n19478) );
  AND U20801 ( .A(n19486), .B(n19487), .Z(n19484) );
  XOR U20802 ( .A(n19485), .B(n11891), .Z(n19487) );
  XNOR U20803 ( .A(n19488), .B(n19489), .Z(n11891) );
  XNOR U20804 ( .A(n[290]), .B(n19490), .Z(n19486) );
  IV U20805 ( .A(n19485), .Z(n19490) );
  XOR U20806 ( .A(n19491), .B(n19492), .Z(n19485) );
  AND U20807 ( .A(n19493), .B(n19494), .Z(n19491) );
  XOR U20808 ( .A(n19492), .B(n11896), .Z(n19494) );
  XNOR U20809 ( .A(n19495), .B(n19496), .Z(n11896) );
  XNOR U20810 ( .A(n[289]), .B(n19497), .Z(n19493) );
  IV U20811 ( .A(n19492), .Z(n19497) );
  XOR U20812 ( .A(n19498), .B(n19499), .Z(n19492) );
  AND U20813 ( .A(n19500), .B(n19501), .Z(n19498) );
  XOR U20814 ( .A(n19499), .B(n11901), .Z(n19501) );
  XNOR U20815 ( .A(n19502), .B(n19503), .Z(n11901) );
  XNOR U20816 ( .A(n[288]), .B(n19504), .Z(n19500) );
  IV U20817 ( .A(n19499), .Z(n19504) );
  XOR U20818 ( .A(n19505), .B(n19506), .Z(n19499) );
  AND U20819 ( .A(n19507), .B(n19508), .Z(n19505) );
  XOR U20820 ( .A(n19506), .B(n11906), .Z(n19508) );
  XNOR U20821 ( .A(n19509), .B(n19510), .Z(n11906) );
  XNOR U20822 ( .A(n[287]), .B(n19511), .Z(n19507) );
  IV U20823 ( .A(n19506), .Z(n19511) );
  XOR U20824 ( .A(n19512), .B(n19513), .Z(n19506) );
  AND U20825 ( .A(n19514), .B(n19515), .Z(n19512) );
  XOR U20826 ( .A(n19513), .B(n11911), .Z(n19515) );
  XNOR U20827 ( .A(n19516), .B(n19517), .Z(n11911) );
  XNOR U20828 ( .A(n[286]), .B(n19518), .Z(n19514) );
  IV U20829 ( .A(n19513), .Z(n19518) );
  XOR U20830 ( .A(n19519), .B(n19520), .Z(n19513) );
  AND U20831 ( .A(n19521), .B(n19522), .Z(n19519) );
  XOR U20832 ( .A(n19520), .B(n11916), .Z(n19522) );
  XNOR U20833 ( .A(n19523), .B(n19524), .Z(n11916) );
  XNOR U20834 ( .A(n[285]), .B(n19525), .Z(n19521) );
  IV U20835 ( .A(n19520), .Z(n19525) );
  XOR U20836 ( .A(n19526), .B(n19527), .Z(n19520) );
  AND U20837 ( .A(n19528), .B(n19529), .Z(n19526) );
  XOR U20838 ( .A(n19527), .B(n11921), .Z(n19529) );
  XNOR U20839 ( .A(n19530), .B(n19531), .Z(n11921) );
  XNOR U20840 ( .A(n[284]), .B(n19532), .Z(n19528) );
  IV U20841 ( .A(n19527), .Z(n19532) );
  XOR U20842 ( .A(n19533), .B(n19534), .Z(n19527) );
  AND U20843 ( .A(n19535), .B(n19536), .Z(n19533) );
  XOR U20844 ( .A(n19534), .B(n11926), .Z(n19536) );
  XNOR U20845 ( .A(n19537), .B(n19538), .Z(n11926) );
  XNOR U20846 ( .A(n[283]), .B(n19539), .Z(n19535) );
  IV U20847 ( .A(n19534), .Z(n19539) );
  XOR U20848 ( .A(n19540), .B(n19541), .Z(n19534) );
  AND U20849 ( .A(n19542), .B(n19543), .Z(n19540) );
  XOR U20850 ( .A(n19541), .B(n11931), .Z(n19543) );
  XNOR U20851 ( .A(n19544), .B(n19545), .Z(n11931) );
  XNOR U20852 ( .A(n[282]), .B(n19546), .Z(n19542) );
  IV U20853 ( .A(n19541), .Z(n19546) );
  XOR U20854 ( .A(n19547), .B(n19548), .Z(n19541) );
  AND U20855 ( .A(n19549), .B(n19550), .Z(n19547) );
  XOR U20856 ( .A(n19548), .B(n11936), .Z(n19550) );
  XNOR U20857 ( .A(n19551), .B(n19552), .Z(n11936) );
  XNOR U20858 ( .A(n[281]), .B(n19553), .Z(n19549) );
  IV U20859 ( .A(n19548), .Z(n19553) );
  XOR U20860 ( .A(n19554), .B(n19555), .Z(n19548) );
  AND U20861 ( .A(n19556), .B(n19557), .Z(n19554) );
  XOR U20862 ( .A(n19555), .B(n11941), .Z(n19557) );
  XNOR U20863 ( .A(n19558), .B(n19559), .Z(n11941) );
  XNOR U20864 ( .A(n[280]), .B(n19560), .Z(n19556) );
  IV U20865 ( .A(n19555), .Z(n19560) );
  XOR U20866 ( .A(n19561), .B(n19562), .Z(n19555) );
  AND U20867 ( .A(n19563), .B(n19564), .Z(n19561) );
  XOR U20868 ( .A(n19562), .B(n11946), .Z(n19564) );
  XNOR U20869 ( .A(n19565), .B(n19566), .Z(n11946) );
  XNOR U20870 ( .A(n[279]), .B(n19567), .Z(n19563) );
  IV U20871 ( .A(n19562), .Z(n19567) );
  XOR U20872 ( .A(n19568), .B(n19569), .Z(n19562) );
  AND U20873 ( .A(n19570), .B(n19571), .Z(n19568) );
  XOR U20874 ( .A(n19569), .B(n11951), .Z(n19571) );
  XNOR U20875 ( .A(n19572), .B(n19573), .Z(n11951) );
  XNOR U20876 ( .A(n[278]), .B(n19574), .Z(n19570) );
  IV U20877 ( .A(n19569), .Z(n19574) );
  XOR U20878 ( .A(n19575), .B(n19576), .Z(n19569) );
  AND U20879 ( .A(n19577), .B(n19578), .Z(n19575) );
  XOR U20880 ( .A(n19576), .B(n11956), .Z(n19578) );
  XNOR U20881 ( .A(n19579), .B(n19580), .Z(n11956) );
  XNOR U20882 ( .A(n[277]), .B(n19581), .Z(n19577) );
  IV U20883 ( .A(n19576), .Z(n19581) );
  XOR U20884 ( .A(n19582), .B(n19583), .Z(n19576) );
  AND U20885 ( .A(n19584), .B(n19585), .Z(n19582) );
  XOR U20886 ( .A(n19583), .B(n11961), .Z(n19585) );
  XNOR U20887 ( .A(n19586), .B(n19587), .Z(n11961) );
  XNOR U20888 ( .A(n[276]), .B(n19588), .Z(n19584) );
  IV U20889 ( .A(n19583), .Z(n19588) );
  XOR U20890 ( .A(n19589), .B(n19590), .Z(n19583) );
  AND U20891 ( .A(n19591), .B(n19592), .Z(n19589) );
  XOR U20892 ( .A(n19590), .B(n11966), .Z(n19592) );
  XNOR U20893 ( .A(n19593), .B(n19594), .Z(n11966) );
  XNOR U20894 ( .A(n[275]), .B(n19595), .Z(n19591) );
  IV U20895 ( .A(n19590), .Z(n19595) );
  XOR U20896 ( .A(n19596), .B(n19597), .Z(n19590) );
  AND U20897 ( .A(n19598), .B(n19599), .Z(n19596) );
  XOR U20898 ( .A(n19597), .B(n11971), .Z(n19599) );
  XNOR U20899 ( .A(n19600), .B(n19601), .Z(n11971) );
  XNOR U20900 ( .A(n[274]), .B(n19602), .Z(n19598) );
  IV U20901 ( .A(n19597), .Z(n19602) );
  XOR U20902 ( .A(n19603), .B(n19604), .Z(n19597) );
  AND U20903 ( .A(n19605), .B(n19606), .Z(n19603) );
  XOR U20904 ( .A(n19604), .B(n11976), .Z(n19606) );
  XNOR U20905 ( .A(n19607), .B(n19608), .Z(n11976) );
  XNOR U20906 ( .A(n[273]), .B(n19609), .Z(n19605) );
  IV U20907 ( .A(n19604), .Z(n19609) );
  XOR U20908 ( .A(n19610), .B(n19611), .Z(n19604) );
  AND U20909 ( .A(n19612), .B(n19613), .Z(n19610) );
  XOR U20910 ( .A(n19611), .B(n11981), .Z(n19613) );
  XNOR U20911 ( .A(n19614), .B(n19615), .Z(n11981) );
  XNOR U20912 ( .A(n[272]), .B(n19616), .Z(n19612) );
  IV U20913 ( .A(n19611), .Z(n19616) );
  XOR U20914 ( .A(n19617), .B(n19618), .Z(n19611) );
  AND U20915 ( .A(n19619), .B(n19620), .Z(n19617) );
  XOR U20916 ( .A(n19618), .B(n11986), .Z(n19620) );
  XNOR U20917 ( .A(n19621), .B(n19622), .Z(n11986) );
  XNOR U20918 ( .A(n[271]), .B(n19623), .Z(n19619) );
  IV U20919 ( .A(n19618), .Z(n19623) );
  XOR U20920 ( .A(n19624), .B(n19625), .Z(n19618) );
  AND U20921 ( .A(n19626), .B(n19627), .Z(n19624) );
  XOR U20922 ( .A(n19625), .B(n11991), .Z(n19627) );
  XNOR U20923 ( .A(n19628), .B(n19629), .Z(n11991) );
  XNOR U20924 ( .A(n[270]), .B(n19630), .Z(n19626) );
  IV U20925 ( .A(n19625), .Z(n19630) );
  XOR U20926 ( .A(n19631), .B(n19632), .Z(n19625) );
  AND U20927 ( .A(n19633), .B(n19634), .Z(n19631) );
  XOR U20928 ( .A(n19632), .B(n11996), .Z(n19634) );
  XNOR U20929 ( .A(n19635), .B(n19636), .Z(n11996) );
  XNOR U20930 ( .A(n[269]), .B(n19637), .Z(n19633) );
  IV U20931 ( .A(n19632), .Z(n19637) );
  XOR U20932 ( .A(n19638), .B(n19639), .Z(n19632) );
  AND U20933 ( .A(n19640), .B(n19641), .Z(n19638) );
  XOR U20934 ( .A(n19639), .B(n12001), .Z(n19641) );
  XNOR U20935 ( .A(n19642), .B(n19643), .Z(n12001) );
  XNOR U20936 ( .A(n[268]), .B(n19644), .Z(n19640) );
  IV U20937 ( .A(n19639), .Z(n19644) );
  XOR U20938 ( .A(n19645), .B(n19646), .Z(n19639) );
  AND U20939 ( .A(n19647), .B(n19648), .Z(n19645) );
  XOR U20940 ( .A(n19646), .B(n12006), .Z(n19648) );
  XNOR U20941 ( .A(n19649), .B(n19650), .Z(n12006) );
  XNOR U20942 ( .A(n[267]), .B(n19651), .Z(n19647) );
  IV U20943 ( .A(n19646), .Z(n19651) );
  XOR U20944 ( .A(n19652), .B(n19653), .Z(n19646) );
  AND U20945 ( .A(n19654), .B(n19655), .Z(n19652) );
  XOR U20946 ( .A(n19653), .B(n12011), .Z(n19655) );
  XNOR U20947 ( .A(n19656), .B(n19657), .Z(n12011) );
  XNOR U20948 ( .A(n[266]), .B(n19658), .Z(n19654) );
  IV U20949 ( .A(n19653), .Z(n19658) );
  XOR U20950 ( .A(n19659), .B(n19660), .Z(n19653) );
  AND U20951 ( .A(n19661), .B(n19662), .Z(n19659) );
  XOR U20952 ( .A(n19660), .B(n12016), .Z(n19662) );
  XNOR U20953 ( .A(n19663), .B(n19664), .Z(n12016) );
  XNOR U20954 ( .A(n[265]), .B(n19665), .Z(n19661) );
  IV U20955 ( .A(n19660), .Z(n19665) );
  XOR U20956 ( .A(n19666), .B(n19667), .Z(n19660) );
  AND U20957 ( .A(n19668), .B(n19669), .Z(n19666) );
  XOR U20958 ( .A(n19667), .B(n12021), .Z(n19669) );
  XNOR U20959 ( .A(n19670), .B(n19671), .Z(n12021) );
  XNOR U20960 ( .A(n[264]), .B(n19672), .Z(n19668) );
  IV U20961 ( .A(n19667), .Z(n19672) );
  XOR U20962 ( .A(n19673), .B(n19674), .Z(n19667) );
  AND U20963 ( .A(n19675), .B(n19676), .Z(n19673) );
  XOR U20964 ( .A(n19674), .B(n12026), .Z(n19676) );
  XNOR U20965 ( .A(n19677), .B(n19678), .Z(n12026) );
  XNOR U20966 ( .A(n[263]), .B(n19679), .Z(n19675) );
  IV U20967 ( .A(n19674), .Z(n19679) );
  XOR U20968 ( .A(n19680), .B(n19681), .Z(n19674) );
  AND U20969 ( .A(n19682), .B(n19683), .Z(n19680) );
  XOR U20970 ( .A(n19681), .B(n12031), .Z(n19683) );
  XNOR U20971 ( .A(n19684), .B(n19685), .Z(n12031) );
  XNOR U20972 ( .A(n[262]), .B(n19686), .Z(n19682) );
  IV U20973 ( .A(n19681), .Z(n19686) );
  XOR U20974 ( .A(n19687), .B(n19688), .Z(n19681) );
  AND U20975 ( .A(n19689), .B(n19690), .Z(n19687) );
  XOR U20976 ( .A(n19688), .B(n12036), .Z(n19690) );
  XNOR U20977 ( .A(n19691), .B(n19692), .Z(n12036) );
  XNOR U20978 ( .A(n[261]), .B(n19693), .Z(n19689) );
  IV U20979 ( .A(n19688), .Z(n19693) );
  XOR U20980 ( .A(n19694), .B(n19695), .Z(n19688) );
  AND U20981 ( .A(n19696), .B(n19697), .Z(n19694) );
  XOR U20982 ( .A(n19695), .B(n12041), .Z(n19697) );
  XNOR U20983 ( .A(n19698), .B(n19699), .Z(n12041) );
  XNOR U20984 ( .A(n[260]), .B(n19700), .Z(n19696) );
  IV U20985 ( .A(n19695), .Z(n19700) );
  XOR U20986 ( .A(n19701), .B(n19702), .Z(n19695) );
  AND U20987 ( .A(n19703), .B(n19704), .Z(n19701) );
  XOR U20988 ( .A(n19702), .B(n12046), .Z(n19704) );
  XNOR U20989 ( .A(n19705), .B(n19706), .Z(n12046) );
  XNOR U20990 ( .A(n[259]), .B(n19707), .Z(n19703) );
  IV U20991 ( .A(n19702), .Z(n19707) );
  XOR U20992 ( .A(n19708), .B(n19709), .Z(n19702) );
  AND U20993 ( .A(n19710), .B(n19711), .Z(n19708) );
  XOR U20994 ( .A(n19709), .B(n12051), .Z(n19711) );
  XNOR U20995 ( .A(n19712), .B(n19713), .Z(n12051) );
  XNOR U20996 ( .A(n[258]), .B(n19714), .Z(n19710) );
  IV U20997 ( .A(n19709), .Z(n19714) );
  XOR U20998 ( .A(n19715), .B(n19716), .Z(n19709) );
  AND U20999 ( .A(n19717), .B(n19718), .Z(n19715) );
  XOR U21000 ( .A(n19716), .B(n12056), .Z(n19718) );
  XNOR U21001 ( .A(n19719), .B(n19720), .Z(n12056) );
  XNOR U21002 ( .A(n[257]), .B(n19721), .Z(n19717) );
  IV U21003 ( .A(n19716), .Z(n19721) );
  XOR U21004 ( .A(n19722), .B(n19723), .Z(n19716) );
  AND U21005 ( .A(n19724), .B(n19725), .Z(n19722) );
  XOR U21006 ( .A(n19723), .B(n12061), .Z(n19725) );
  XNOR U21007 ( .A(n19726), .B(n19727), .Z(n12061) );
  XNOR U21008 ( .A(n[256]), .B(n19728), .Z(n19724) );
  IV U21009 ( .A(n19723), .Z(n19728) );
  XOR U21010 ( .A(n19729), .B(n19730), .Z(n19723) );
  AND U21011 ( .A(n19731), .B(n19732), .Z(n19729) );
  XOR U21012 ( .A(n19730), .B(n12066), .Z(n19732) );
  XNOR U21013 ( .A(n19733), .B(n19734), .Z(n12066) );
  XNOR U21014 ( .A(n[255]), .B(n19735), .Z(n19731) );
  IV U21015 ( .A(n19730), .Z(n19735) );
  XOR U21016 ( .A(n19736), .B(n19737), .Z(n19730) );
  AND U21017 ( .A(n19738), .B(n19739), .Z(n19736) );
  XOR U21018 ( .A(n19737), .B(n12071), .Z(n19739) );
  XNOR U21019 ( .A(n19740), .B(n19741), .Z(n12071) );
  XNOR U21020 ( .A(n[254]), .B(n19742), .Z(n19738) );
  IV U21021 ( .A(n19737), .Z(n19742) );
  XOR U21022 ( .A(n19743), .B(n19744), .Z(n19737) );
  AND U21023 ( .A(n19745), .B(n19746), .Z(n19743) );
  XOR U21024 ( .A(n19744), .B(n12076), .Z(n19746) );
  XNOR U21025 ( .A(n19747), .B(n19748), .Z(n12076) );
  XNOR U21026 ( .A(n[253]), .B(n19749), .Z(n19745) );
  IV U21027 ( .A(n19744), .Z(n19749) );
  XOR U21028 ( .A(n19750), .B(n19751), .Z(n19744) );
  AND U21029 ( .A(n19752), .B(n19753), .Z(n19750) );
  XOR U21030 ( .A(n19751), .B(n12081), .Z(n19753) );
  XNOR U21031 ( .A(n19754), .B(n19755), .Z(n12081) );
  XNOR U21032 ( .A(n[252]), .B(n19756), .Z(n19752) );
  IV U21033 ( .A(n19751), .Z(n19756) );
  XOR U21034 ( .A(n19757), .B(n19758), .Z(n19751) );
  AND U21035 ( .A(n19759), .B(n19760), .Z(n19757) );
  XOR U21036 ( .A(n19758), .B(n12086), .Z(n19760) );
  XNOR U21037 ( .A(n19761), .B(n19762), .Z(n12086) );
  XNOR U21038 ( .A(n[251]), .B(n19763), .Z(n19759) );
  IV U21039 ( .A(n19758), .Z(n19763) );
  XOR U21040 ( .A(n19764), .B(n19765), .Z(n19758) );
  AND U21041 ( .A(n19766), .B(n19767), .Z(n19764) );
  XOR U21042 ( .A(n19765), .B(n12091), .Z(n19767) );
  XNOR U21043 ( .A(n19768), .B(n19769), .Z(n12091) );
  XNOR U21044 ( .A(n[250]), .B(n19770), .Z(n19766) );
  IV U21045 ( .A(n19765), .Z(n19770) );
  XOR U21046 ( .A(n19771), .B(n19772), .Z(n19765) );
  AND U21047 ( .A(n19773), .B(n19774), .Z(n19771) );
  XOR U21048 ( .A(n19772), .B(n12096), .Z(n19774) );
  XNOR U21049 ( .A(n19775), .B(n19776), .Z(n12096) );
  XNOR U21050 ( .A(n[249]), .B(n19777), .Z(n19773) );
  IV U21051 ( .A(n19772), .Z(n19777) );
  XOR U21052 ( .A(n19778), .B(n19779), .Z(n19772) );
  AND U21053 ( .A(n19780), .B(n19781), .Z(n19778) );
  XOR U21054 ( .A(n19779), .B(n12101), .Z(n19781) );
  XNOR U21055 ( .A(n19782), .B(n19783), .Z(n12101) );
  XNOR U21056 ( .A(n[248]), .B(n19784), .Z(n19780) );
  IV U21057 ( .A(n19779), .Z(n19784) );
  XOR U21058 ( .A(n19785), .B(n19786), .Z(n19779) );
  AND U21059 ( .A(n19787), .B(n19788), .Z(n19785) );
  XOR U21060 ( .A(n19786), .B(n12106), .Z(n19788) );
  XNOR U21061 ( .A(n19789), .B(n19790), .Z(n12106) );
  XNOR U21062 ( .A(n[247]), .B(n19791), .Z(n19787) );
  IV U21063 ( .A(n19786), .Z(n19791) );
  XOR U21064 ( .A(n19792), .B(n19793), .Z(n19786) );
  AND U21065 ( .A(n19794), .B(n19795), .Z(n19792) );
  XOR U21066 ( .A(n19793), .B(n12111), .Z(n19795) );
  XNOR U21067 ( .A(n19796), .B(n19797), .Z(n12111) );
  XNOR U21068 ( .A(n[246]), .B(n19798), .Z(n19794) );
  IV U21069 ( .A(n19793), .Z(n19798) );
  XOR U21070 ( .A(n19799), .B(n19800), .Z(n19793) );
  AND U21071 ( .A(n19801), .B(n19802), .Z(n19799) );
  XOR U21072 ( .A(n19800), .B(n12116), .Z(n19802) );
  XNOR U21073 ( .A(n19803), .B(n19804), .Z(n12116) );
  XNOR U21074 ( .A(n[245]), .B(n19805), .Z(n19801) );
  IV U21075 ( .A(n19800), .Z(n19805) );
  XOR U21076 ( .A(n19806), .B(n19807), .Z(n19800) );
  AND U21077 ( .A(n19808), .B(n19809), .Z(n19806) );
  XOR U21078 ( .A(n19807), .B(n12121), .Z(n19809) );
  XNOR U21079 ( .A(n19810), .B(n19811), .Z(n12121) );
  XNOR U21080 ( .A(n[244]), .B(n19812), .Z(n19808) );
  IV U21081 ( .A(n19807), .Z(n19812) );
  XOR U21082 ( .A(n19813), .B(n19814), .Z(n19807) );
  AND U21083 ( .A(n19815), .B(n19816), .Z(n19813) );
  XOR U21084 ( .A(n19814), .B(n12126), .Z(n19816) );
  XNOR U21085 ( .A(n19817), .B(n19818), .Z(n12126) );
  XNOR U21086 ( .A(n[243]), .B(n19819), .Z(n19815) );
  IV U21087 ( .A(n19814), .Z(n19819) );
  XOR U21088 ( .A(n19820), .B(n19821), .Z(n19814) );
  AND U21089 ( .A(n19822), .B(n19823), .Z(n19820) );
  XOR U21090 ( .A(n19821), .B(n12131), .Z(n19823) );
  XNOR U21091 ( .A(n19824), .B(n19825), .Z(n12131) );
  XNOR U21092 ( .A(n[242]), .B(n19826), .Z(n19822) );
  IV U21093 ( .A(n19821), .Z(n19826) );
  XOR U21094 ( .A(n19827), .B(n19828), .Z(n19821) );
  AND U21095 ( .A(n19829), .B(n19830), .Z(n19827) );
  XOR U21096 ( .A(n19828), .B(n12136), .Z(n19830) );
  XNOR U21097 ( .A(n19831), .B(n19832), .Z(n12136) );
  XNOR U21098 ( .A(n[241]), .B(n19833), .Z(n19829) );
  IV U21099 ( .A(n19828), .Z(n19833) );
  XOR U21100 ( .A(n19834), .B(n19835), .Z(n19828) );
  AND U21101 ( .A(n19836), .B(n19837), .Z(n19834) );
  XOR U21102 ( .A(n19835), .B(n12141), .Z(n19837) );
  XNOR U21103 ( .A(n19838), .B(n19839), .Z(n12141) );
  XNOR U21104 ( .A(n[240]), .B(n19840), .Z(n19836) );
  IV U21105 ( .A(n19835), .Z(n19840) );
  XOR U21106 ( .A(n19841), .B(n19842), .Z(n19835) );
  AND U21107 ( .A(n19843), .B(n19844), .Z(n19841) );
  XOR U21108 ( .A(n19842), .B(n12146), .Z(n19844) );
  XNOR U21109 ( .A(n19845), .B(n19846), .Z(n12146) );
  XNOR U21110 ( .A(n[239]), .B(n19847), .Z(n19843) );
  IV U21111 ( .A(n19842), .Z(n19847) );
  XOR U21112 ( .A(n19848), .B(n19849), .Z(n19842) );
  AND U21113 ( .A(n19850), .B(n19851), .Z(n19848) );
  XOR U21114 ( .A(n19849), .B(n12151), .Z(n19851) );
  XNOR U21115 ( .A(n19852), .B(n19853), .Z(n12151) );
  XNOR U21116 ( .A(n[238]), .B(n19854), .Z(n19850) );
  IV U21117 ( .A(n19849), .Z(n19854) );
  XOR U21118 ( .A(n19855), .B(n19856), .Z(n19849) );
  AND U21119 ( .A(n19857), .B(n19858), .Z(n19855) );
  XOR U21120 ( .A(n19856), .B(n12156), .Z(n19858) );
  XNOR U21121 ( .A(n19859), .B(n19860), .Z(n12156) );
  XNOR U21122 ( .A(n[237]), .B(n19861), .Z(n19857) );
  IV U21123 ( .A(n19856), .Z(n19861) );
  XOR U21124 ( .A(n19862), .B(n19863), .Z(n19856) );
  AND U21125 ( .A(n19864), .B(n19865), .Z(n19862) );
  XOR U21126 ( .A(n19863), .B(n12161), .Z(n19865) );
  XNOR U21127 ( .A(n19866), .B(n19867), .Z(n12161) );
  XNOR U21128 ( .A(n[236]), .B(n19868), .Z(n19864) );
  IV U21129 ( .A(n19863), .Z(n19868) );
  XOR U21130 ( .A(n19869), .B(n19870), .Z(n19863) );
  AND U21131 ( .A(n19871), .B(n19872), .Z(n19869) );
  XOR U21132 ( .A(n19870), .B(n12166), .Z(n19872) );
  XNOR U21133 ( .A(n19873), .B(n19874), .Z(n12166) );
  XNOR U21134 ( .A(n[235]), .B(n19875), .Z(n19871) );
  IV U21135 ( .A(n19870), .Z(n19875) );
  XOR U21136 ( .A(n19876), .B(n19877), .Z(n19870) );
  AND U21137 ( .A(n19878), .B(n19879), .Z(n19876) );
  XOR U21138 ( .A(n19877), .B(n12171), .Z(n19879) );
  XNOR U21139 ( .A(n19880), .B(n19881), .Z(n12171) );
  XNOR U21140 ( .A(n[234]), .B(n19882), .Z(n19878) );
  IV U21141 ( .A(n19877), .Z(n19882) );
  XOR U21142 ( .A(n19883), .B(n19884), .Z(n19877) );
  AND U21143 ( .A(n19885), .B(n19886), .Z(n19883) );
  XOR U21144 ( .A(n19884), .B(n12176), .Z(n19886) );
  XNOR U21145 ( .A(n19887), .B(n19888), .Z(n12176) );
  XNOR U21146 ( .A(n[233]), .B(n19889), .Z(n19885) );
  IV U21147 ( .A(n19884), .Z(n19889) );
  XOR U21148 ( .A(n19890), .B(n19891), .Z(n19884) );
  AND U21149 ( .A(n19892), .B(n19893), .Z(n19890) );
  XOR U21150 ( .A(n19891), .B(n12181), .Z(n19893) );
  XNOR U21151 ( .A(n19894), .B(n19895), .Z(n12181) );
  XNOR U21152 ( .A(n[232]), .B(n19896), .Z(n19892) );
  IV U21153 ( .A(n19891), .Z(n19896) );
  XOR U21154 ( .A(n19897), .B(n19898), .Z(n19891) );
  AND U21155 ( .A(n19899), .B(n19900), .Z(n19897) );
  XOR U21156 ( .A(n19898), .B(n12186), .Z(n19900) );
  XNOR U21157 ( .A(n19901), .B(n19902), .Z(n12186) );
  XNOR U21158 ( .A(n[231]), .B(n19903), .Z(n19899) );
  IV U21159 ( .A(n19898), .Z(n19903) );
  XOR U21160 ( .A(n19904), .B(n19905), .Z(n19898) );
  AND U21161 ( .A(n19906), .B(n19907), .Z(n19904) );
  XOR U21162 ( .A(n19905), .B(n12191), .Z(n19907) );
  XNOR U21163 ( .A(n19908), .B(n19909), .Z(n12191) );
  XNOR U21164 ( .A(n[230]), .B(n19910), .Z(n19906) );
  IV U21165 ( .A(n19905), .Z(n19910) );
  XOR U21166 ( .A(n19911), .B(n19912), .Z(n19905) );
  AND U21167 ( .A(n19913), .B(n19914), .Z(n19911) );
  XOR U21168 ( .A(n19912), .B(n12196), .Z(n19914) );
  XNOR U21169 ( .A(n19915), .B(n19916), .Z(n12196) );
  XNOR U21170 ( .A(n[229]), .B(n19917), .Z(n19913) );
  IV U21171 ( .A(n19912), .Z(n19917) );
  XOR U21172 ( .A(n19918), .B(n19919), .Z(n19912) );
  AND U21173 ( .A(n19920), .B(n19921), .Z(n19918) );
  XOR U21174 ( .A(n19919), .B(n12201), .Z(n19921) );
  XNOR U21175 ( .A(n19922), .B(n19923), .Z(n12201) );
  XNOR U21176 ( .A(n[228]), .B(n19924), .Z(n19920) );
  IV U21177 ( .A(n19919), .Z(n19924) );
  XOR U21178 ( .A(n19925), .B(n19926), .Z(n19919) );
  AND U21179 ( .A(n19927), .B(n19928), .Z(n19925) );
  XOR U21180 ( .A(n19926), .B(n12206), .Z(n19928) );
  XNOR U21181 ( .A(n19929), .B(n19930), .Z(n12206) );
  XNOR U21182 ( .A(n[227]), .B(n19931), .Z(n19927) );
  IV U21183 ( .A(n19926), .Z(n19931) );
  XOR U21184 ( .A(n19932), .B(n19933), .Z(n19926) );
  AND U21185 ( .A(n19934), .B(n19935), .Z(n19932) );
  XOR U21186 ( .A(n19933), .B(n12211), .Z(n19935) );
  XNOR U21187 ( .A(n19936), .B(n19937), .Z(n12211) );
  XNOR U21188 ( .A(n[226]), .B(n19938), .Z(n19934) );
  IV U21189 ( .A(n19933), .Z(n19938) );
  XOR U21190 ( .A(n19939), .B(n19940), .Z(n19933) );
  AND U21191 ( .A(n19941), .B(n19942), .Z(n19939) );
  XOR U21192 ( .A(n19940), .B(n12216), .Z(n19942) );
  XNOR U21193 ( .A(n19943), .B(n19944), .Z(n12216) );
  XNOR U21194 ( .A(n[225]), .B(n19945), .Z(n19941) );
  IV U21195 ( .A(n19940), .Z(n19945) );
  XOR U21196 ( .A(n19946), .B(n19947), .Z(n19940) );
  AND U21197 ( .A(n19948), .B(n19949), .Z(n19946) );
  XOR U21198 ( .A(n19947), .B(n12221), .Z(n19949) );
  XNOR U21199 ( .A(n19950), .B(n19951), .Z(n12221) );
  XNOR U21200 ( .A(n[224]), .B(n19952), .Z(n19948) );
  IV U21201 ( .A(n19947), .Z(n19952) );
  XOR U21202 ( .A(n19953), .B(n19954), .Z(n19947) );
  AND U21203 ( .A(n19955), .B(n19956), .Z(n19953) );
  XOR U21204 ( .A(n19954), .B(n12226), .Z(n19956) );
  XNOR U21205 ( .A(n19957), .B(n19958), .Z(n12226) );
  XNOR U21206 ( .A(n[223]), .B(n19959), .Z(n19955) );
  IV U21207 ( .A(n19954), .Z(n19959) );
  XOR U21208 ( .A(n19960), .B(n19961), .Z(n19954) );
  AND U21209 ( .A(n19962), .B(n19963), .Z(n19960) );
  XOR U21210 ( .A(n19961), .B(n12231), .Z(n19963) );
  XNOR U21211 ( .A(n19964), .B(n19965), .Z(n12231) );
  XNOR U21212 ( .A(n[222]), .B(n19966), .Z(n19962) );
  IV U21213 ( .A(n19961), .Z(n19966) );
  XOR U21214 ( .A(n19967), .B(n19968), .Z(n19961) );
  AND U21215 ( .A(n19969), .B(n19970), .Z(n19967) );
  XOR U21216 ( .A(n19968), .B(n12236), .Z(n19970) );
  XNOR U21217 ( .A(n19971), .B(n19972), .Z(n12236) );
  XNOR U21218 ( .A(n[221]), .B(n19973), .Z(n19969) );
  IV U21219 ( .A(n19968), .Z(n19973) );
  XOR U21220 ( .A(n19974), .B(n19975), .Z(n19968) );
  AND U21221 ( .A(n19976), .B(n19977), .Z(n19974) );
  XOR U21222 ( .A(n19975), .B(n12241), .Z(n19977) );
  XNOR U21223 ( .A(n19978), .B(n19979), .Z(n12241) );
  XNOR U21224 ( .A(n[220]), .B(n19980), .Z(n19976) );
  IV U21225 ( .A(n19975), .Z(n19980) );
  XOR U21226 ( .A(n19981), .B(n19982), .Z(n19975) );
  AND U21227 ( .A(n19983), .B(n19984), .Z(n19981) );
  XOR U21228 ( .A(n19982), .B(n12246), .Z(n19984) );
  XNOR U21229 ( .A(n19985), .B(n19986), .Z(n12246) );
  XNOR U21230 ( .A(n[219]), .B(n19987), .Z(n19983) );
  IV U21231 ( .A(n19982), .Z(n19987) );
  XOR U21232 ( .A(n19988), .B(n19989), .Z(n19982) );
  AND U21233 ( .A(n19990), .B(n19991), .Z(n19988) );
  XOR U21234 ( .A(n19989), .B(n12251), .Z(n19991) );
  XNOR U21235 ( .A(n19992), .B(n19993), .Z(n12251) );
  XNOR U21236 ( .A(n[218]), .B(n19994), .Z(n19990) );
  IV U21237 ( .A(n19989), .Z(n19994) );
  XOR U21238 ( .A(n19995), .B(n19996), .Z(n19989) );
  AND U21239 ( .A(n19997), .B(n19998), .Z(n19995) );
  XOR U21240 ( .A(n19996), .B(n12256), .Z(n19998) );
  XNOR U21241 ( .A(n19999), .B(n20000), .Z(n12256) );
  XNOR U21242 ( .A(n[217]), .B(n20001), .Z(n19997) );
  IV U21243 ( .A(n19996), .Z(n20001) );
  XOR U21244 ( .A(n20002), .B(n20003), .Z(n19996) );
  AND U21245 ( .A(n20004), .B(n20005), .Z(n20002) );
  XOR U21246 ( .A(n20003), .B(n12261), .Z(n20005) );
  XNOR U21247 ( .A(n20006), .B(n20007), .Z(n12261) );
  XNOR U21248 ( .A(n[216]), .B(n20008), .Z(n20004) );
  IV U21249 ( .A(n20003), .Z(n20008) );
  XOR U21250 ( .A(n20009), .B(n20010), .Z(n20003) );
  AND U21251 ( .A(n20011), .B(n20012), .Z(n20009) );
  XOR U21252 ( .A(n20010), .B(n12266), .Z(n20012) );
  XNOR U21253 ( .A(n20013), .B(n20014), .Z(n12266) );
  XNOR U21254 ( .A(n[215]), .B(n20015), .Z(n20011) );
  IV U21255 ( .A(n20010), .Z(n20015) );
  XOR U21256 ( .A(n20016), .B(n20017), .Z(n20010) );
  AND U21257 ( .A(n20018), .B(n20019), .Z(n20016) );
  XOR U21258 ( .A(n20017), .B(n12271), .Z(n20019) );
  XNOR U21259 ( .A(n20020), .B(n20021), .Z(n12271) );
  XNOR U21260 ( .A(n[214]), .B(n20022), .Z(n20018) );
  IV U21261 ( .A(n20017), .Z(n20022) );
  XOR U21262 ( .A(n20023), .B(n20024), .Z(n20017) );
  AND U21263 ( .A(n20025), .B(n20026), .Z(n20023) );
  XOR U21264 ( .A(n20024), .B(n12276), .Z(n20026) );
  XNOR U21265 ( .A(n20027), .B(n20028), .Z(n12276) );
  XNOR U21266 ( .A(n[213]), .B(n20029), .Z(n20025) );
  IV U21267 ( .A(n20024), .Z(n20029) );
  XOR U21268 ( .A(n20030), .B(n20031), .Z(n20024) );
  AND U21269 ( .A(n20032), .B(n20033), .Z(n20030) );
  XOR U21270 ( .A(n20031), .B(n12281), .Z(n20033) );
  XNOR U21271 ( .A(n20034), .B(n20035), .Z(n12281) );
  XNOR U21272 ( .A(n[212]), .B(n20036), .Z(n20032) );
  IV U21273 ( .A(n20031), .Z(n20036) );
  XOR U21274 ( .A(n20037), .B(n20038), .Z(n20031) );
  AND U21275 ( .A(n20039), .B(n20040), .Z(n20037) );
  XOR U21276 ( .A(n20038), .B(n12286), .Z(n20040) );
  XNOR U21277 ( .A(n20041), .B(n20042), .Z(n12286) );
  XNOR U21278 ( .A(n[211]), .B(n20043), .Z(n20039) );
  IV U21279 ( .A(n20038), .Z(n20043) );
  XOR U21280 ( .A(n20044), .B(n20045), .Z(n20038) );
  AND U21281 ( .A(n20046), .B(n20047), .Z(n20044) );
  XOR U21282 ( .A(n20045), .B(n12291), .Z(n20047) );
  XNOR U21283 ( .A(n20048), .B(n20049), .Z(n12291) );
  XNOR U21284 ( .A(n[210]), .B(n20050), .Z(n20046) );
  IV U21285 ( .A(n20045), .Z(n20050) );
  XOR U21286 ( .A(n20051), .B(n20052), .Z(n20045) );
  AND U21287 ( .A(n20053), .B(n20054), .Z(n20051) );
  XOR U21288 ( .A(n20052), .B(n12296), .Z(n20054) );
  XNOR U21289 ( .A(n20055), .B(n20056), .Z(n12296) );
  XNOR U21290 ( .A(n[209]), .B(n20057), .Z(n20053) );
  IV U21291 ( .A(n20052), .Z(n20057) );
  XOR U21292 ( .A(n20058), .B(n20059), .Z(n20052) );
  AND U21293 ( .A(n20060), .B(n20061), .Z(n20058) );
  XOR U21294 ( .A(n20059), .B(n12301), .Z(n20061) );
  XNOR U21295 ( .A(n20062), .B(n20063), .Z(n12301) );
  XNOR U21296 ( .A(n[208]), .B(n20064), .Z(n20060) );
  IV U21297 ( .A(n20059), .Z(n20064) );
  XOR U21298 ( .A(n20065), .B(n20066), .Z(n20059) );
  AND U21299 ( .A(n20067), .B(n20068), .Z(n20065) );
  XOR U21300 ( .A(n20066), .B(n12306), .Z(n20068) );
  XNOR U21301 ( .A(n20069), .B(n20070), .Z(n12306) );
  XNOR U21302 ( .A(n[207]), .B(n20071), .Z(n20067) );
  IV U21303 ( .A(n20066), .Z(n20071) );
  XOR U21304 ( .A(n20072), .B(n20073), .Z(n20066) );
  AND U21305 ( .A(n20074), .B(n20075), .Z(n20072) );
  XOR U21306 ( .A(n20073), .B(n12311), .Z(n20075) );
  XNOR U21307 ( .A(n20076), .B(n20077), .Z(n12311) );
  XNOR U21308 ( .A(n[206]), .B(n20078), .Z(n20074) );
  IV U21309 ( .A(n20073), .Z(n20078) );
  XOR U21310 ( .A(n20079), .B(n20080), .Z(n20073) );
  AND U21311 ( .A(n20081), .B(n20082), .Z(n20079) );
  XOR U21312 ( .A(n20080), .B(n12316), .Z(n20082) );
  XNOR U21313 ( .A(n20083), .B(n20084), .Z(n12316) );
  XNOR U21314 ( .A(n[205]), .B(n20085), .Z(n20081) );
  IV U21315 ( .A(n20080), .Z(n20085) );
  XOR U21316 ( .A(n20086), .B(n20087), .Z(n20080) );
  AND U21317 ( .A(n20088), .B(n20089), .Z(n20086) );
  XOR U21318 ( .A(n20087), .B(n12321), .Z(n20089) );
  XNOR U21319 ( .A(n20090), .B(n20091), .Z(n12321) );
  XNOR U21320 ( .A(n[204]), .B(n20092), .Z(n20088) );
  IV U21321 ( .A(n20087), .Z(n20092) );
  XOR U21322 ( .A(n20093), .B(n20094), .Z(n20087) );
  AND U21323 ( .A(n20095), .B(n20096), .Z(n20093) );
  XOR U21324 ( .A(n20094), .B(n12326), .Z(n20096) );
  XNOR U21325 ( .A(n20097), .B(n20098), .Z(n12326) );
  XNOR U21326 ( .A(n[203]), .B(n20099), .Z(n20095) );
  IV U21327 ( .A(n20094), .Z(n20099) );
  XOR U21328 ( .A(n20100), .B(n20101), .Z(n20094) );
  AND U21329 ( .A(n20102), .B(n20103), .Z(n20100) );
  XOR U21330 ( .A(n20101), .B(n12331), .Z(n20103) );
  XNOR U21331 ( .A(n20104), .B(n20105), .Z(n12331) );
  XNOR U21332 ( .A(n[202]), .B(n20106), .Z(n20102) );
  IV U21333 ( .A(n20101), .Z(n20106) );
  XOR U21334 ( .A(n20107), .B(n20108), .Z(n20101) );
  AND U21335 ( .A(n20109), .B(n20110), .Z(n20107) );
  XOR U21336 ( .A(n20108), .B(n12336), .Z(n20110) );
  XNOR U21337 ( .A(n20111), .B(n20112), .Z(n12336) );
  XNOR U21338 ( .A(n[201]), .B(n20113), .Z(n20109) );
  IV U21339 ( .A(n20108), .Z(n20113) );
  XOR U21340 ( .A(n20114), .B(n20115), .Z(n20108) );
  AND U21341 ( .A(n20116), .B(n20117), .Z(n20114) );
  XOR U21342 ( .A(n20115), .B(n12341), .Z(n20117) );
  XNOR U21343 ( .A(n20118), .B(n20119), .Z(n12341) );
  XNOR U21344 ( .A(n[200]), .B(n20120), .Z(n20116) );
  IV U21345 ( .A(n20115), .Z(n20120) );
  XOR U21346 ( .A(n20121), .B(n20122), .Z(n20115) );
  AND U21347 ( .A(n20123), .B(n20124), .Z(n20121) );
  XOR U21348 ( .A(n20122), .B(n12346), .Z(n20124) );
  XNOR U21349 ( .A(n20125), .B(n20126), .Z(n12346) );
  XNOR U21350 ( .A(n[199]), .B(n20127), .Z(n20123) );
  IV U21351 ( .A(n20122), .Z(n20127) );
  XOR U21352 ( .A(n20128), .B(n20129), .Z(n20122) );
  AND U21353 ( .A(n20130), .B(n20131), .Z(n20128) );
  XOR U21354 ( .A(n20129), .B(n12351), .Z(n20131) );
  XNOR U21355 ( .A(n20132), .B(n20133), .Z(n12351) );
  XNOR U21356 ( .A(n[198]), .B(n20134), .Z(n20130) );
  IV U21357 ( .A(n20129), .Z(n20134) );
  XOR U21358 ( .A(n20135), .B(n20136), .Z(n20129) );
  AND U21359 ( .A(n20137), .B(n20138), .Z(n20135) );
  XOR U21360 ( .A(n20136), .B(n12356), .Z(n20138) );
  XNOR U21361 ( .A(n20139), .B(n20140), .Z(n12356) );
  XNOR U21362 ( .A(n[197]), .B(n20141), .Z(n20137) );
  IV U21363 ( .A(n20136), .Z(n20141) );
  XOR U21364 ( .A(n20142), .B(n20143), .Z(n20136) );
  AND U21365 ( .A(n20144), .B(n20145), .Z(n20142) );
  XOR U21366 ( .A(n20143), .B(n12361), .Z(n20145) );
  XNOR U21367 ( .A(n20146), .B(n20147), .Z(n12361) );
  XNOR U21368 ( .A(n[196]), .B(n20148), .Z(n20144) );
  IV U21369 ( .A(n20143), .Z(n20148) );
  XOR U21370 ( .A(n20149), .B(n20150), .Z(n20143) );
  AND U21371 ( .A(n20151), .B(n20152), .Z(n20149) );
  XOR U21372 ( .A(n20150), .B(n12366), .Z(n20152) );
  XNOR U21373 ( .A(n20153), .B(n20154), .Z(n12366) );
  XNOR U21374 ( .A(n[195]), .B(n20155), .Z(n20151) );
  IV U21375 ( .A(n20150), .Z(n20155) );
  XOR U21376 ( .A(n20156), .B(n20157), .Z(n20150) );
  AND U21377 ( .A(n20158), .B(n20159), .Z(n20156) );
  XOR U21378 ( .A(n20157), .B(n12371), .Z(n20159) );
  XNOR U21379 ( .A(n20160), .B(n20161), .Z(n12371) );
  XNOR U21380 ( .A(n[194]), .B(n20162), .Z(n20158) );
  IV U21381 ( .A(n20157), .Z(n20162) );
  XOR U21382 ( .A(n20163), .B(n20164), .Z(n20157) );
  AND U21383 ( .A(n20165), .B(n20166), .Z(n20163) );
  XOR U21384 ( .A(n20164), .B(n12376), .Z(n20166) );
  XNOR U21385 ( .A(n20167), .B(n20168), .Z(n12376) );
  XNOR U21386 ( .A(n[193]), .B(n20169), .Z(n20165) );
  IV U21387 ( .A(n20164), .Z(n20169) );
  XOR U21388 ( .A(n20170), .B(n20171), .Z(n20164) );
  AND U21389 ( .A(n20172), .B(n20173), .Z(n20170) );
  XOR U21390 ( .A(n20171), .B(n12381), .Z(n20173) );
  XNOR U21391 ( .A(n20174), .B(n20175), .Z(n12381) );
  XNOR U21392 ( .A(n[192]), .B(n20176), .Z(n20172) );
  IV U21393 ( .A(n20171), .Z(n20176) );
  XOR U21394 ( .A(n20177), .B(n20178), .Z(n20171) );
  AND U21395 ( .A(n20179), .B(n20180), .Z(n20177) );
  XOR U21396 ( .A(n20178), .B(n12386), .Z(n20180) );
  XNOR U21397 ( .A(n20181), .B(n20182), .Z(n12386) );
  XNOR U21398 ( .A(n[191]), .B(n20183), .Z(n20179) );
  IV U21399 ( .A(n20178), .Z(n20183) );
  XOR U21400 ( .A(n20184), .B(n20185), .Z(n20178) );
  AND U21401 ( .A(n20186), .B(n20187), .Z(n20184) );
  XOR U21402 ( .A(n20185), .B(n12391), .Z(n20187) );
  XNOR U21403 ( .A(n20188), .B(n20189), .Z(n12391) );
  XNOR U21404 ( .A(n[190]), .B(n20190), .Z(n20186) );
  IV U21405 ( .A(n20185), .Z(n20190) );
  XOR U21406 ( .A(n20191), .B(n20192), .Z(n20185) );
  AND U21407 ( .A(n20193), .B(n20194), .Z(n20191) );
  XOR U21408 ( .A(n20192), .B(n12396), .Z(n20194) );
  XNOR U21409 ( .A(n20195), .B(n20196), .Z(n12396) );
  XNOR U21410 ( .A(n[189]), .B(n20197), .Z(n20193) );
  IV U21411 ( .A(n20192), .Z(n20197) );
  XOR U21412 ( .A(n20198), .B(n20199), .Z(n20192) );
  AND U21413 ( .A(n20200), .B(n20201), .Z(n20198) );
  XOR U21414 ( .A(n20199), .B(n12401), .Z(n20201) );
  XNOR U21415 ( .A(n20202), .B(n20203), .Z(n12401) );
  XNOR U21416 ( .A(n[188]), .B(n20204), .Z(n20200) );
  IV U21417 ( .A(n20199), .Z(n20204) );
  XOR U21418 ( .A(n20205), .B(n20206), .Z(n20199) );
  AND U21419 ( .A(n20207), .B(n20208), .Z(n20205) );
  XOR U21420 ( .A(n20206), .B(n12406), .Z(n20208) );
  XNOR U21421 ( .A(n20209), .B(n20210), .Z(n12406) );
  XNOR U21422 ( .A(n[187]), .B(n20211), .Z(n20207) );
  IV U21423 ( .A(n20206), .Z(n20211) );
  XOR U21424 ( .A(n20212), .B(n20213), .Z(n20206) );
  AND U21425 ( .A(n20214), .B(n20215), .Z(n20212) );
  XOR U21426 ( .A(n20213), .B(n12411), .Z(n20215) );
  XNOR U21427 ( .A(n20216), .B(n20217), .Z(n12411) );
  XNOR U21428 ( .A(n[186]), .B(n20218), .Z(n20214) );
  IV U21429 ( .A(n20213), .Z(n20218) );
  XOR U21430 ( .A(n20219), .B(n20220), .Z(n20213) );
  AND U21431 ( .A(n20221), .B(n20222), .Z(n20219) );
  XOR U21432 ( .A(n20220), .B(n12416), .Z(n20222) );
  XNOR U21433 ( .A(n20223), .B(n20224), .Z(n12416) );
  XNOR U21434 ( .A(n[185]), .B(n20225), .Z(n20221) );
  IV U21435 ( .A(n20220), .Z(n20225) );
  XOR U21436 ( .A(n20226), .B(n20227), .Z(n20220) );
  AND U21437 ( .A(n20228), .B(n20229), .Z(n20226) );
  XOR U21438 ( .A(n20227), .B(n12421), .Z(n20229) );
  XNOR U21439 ( .A(n20230), .B(n20231), .Z(n12421) );
  XNOR U21440 ( .A(n[184]), .B(n20232), .Z(n20228) );
  IV U21441 ( .A(n20227), .Z(n20232) );
  XOR U21442 ( .A(n20233), .B(n20234), .Z(n20227) );
  AND U21443 ( .A(n20235), .B(n20236), .Z(n20233) );
  XOR U21444 ( .A(n20234), .B(n12426), .Z(n20236) );
  XNOR U21445 ( .A(n20237), .B(n20238), .Z(n12426) );
  XNOR U21446 ( .A(n[183]), .B(n20239), .Z(n20235) );
  IV U21447 ( .A(n20234), .Z(n20239) );
  XOR U21448 ( .A(n20240), .B(n20241), .Z(n20234) );
  AND U21449 ( .A(n20242), .B(n20243), .Z(n20240) );
  XOR U21450 ( .A(n20241), .B(n12431), .Z(n20243) );
  XNOR U21451 ( .A(n20244), .B(n20245), .Z(n12431) );
  XNOR U21452 ( .A(n[182]), .B(n20246), .Z(n20242) );
  IV U21453 ( .A(n20241), .Z(n20246) );
  XOR U21454 ( .A(n20247), .B(n20248), .Z(n20241) );
  AND U21455 ( .A(n20249), .B(n20250), .Z(n20247) );
  XOR U21456 ( .A(n20248), .B(n12436), .Z(n20250) );
  XNOR U21457 ( .A(n20251), .B(n20252), .Z(n12436) );
  XNOR U21458 ( .A(n[181]), .B(n20253), .Z(n20249) );
  IV U21459 ( .A(n20248), .Z(n20253) );
  XOR U21460 ( .A(n20254), .B(n20255), .Z(n20248) );
  AND U21461 ( .A(n20256), .B(n20257), .Z(n20254) );
  XOR U21462 ( .A(n20255), .B(n12441), .Z(n20257) );
  XNOR U21463 ( .A(n20258), .B(n20259), .Z(n12441) );
  XNOR U21464 ( .A(n[180]), .B(n20260), .Z(n20256) );
  IV U21465 ( .A(n20255), .Z(n20260) );
  XOR U21466 ( .A(n20261), .B(n20262), .Z(n20255) );
  AND U21467 ( .A(n20263), .B(n20264), .Z(n20261) );
  XOR U21468 ( .A(n20262), .B(n12446), .Z(n20264) );
  XNOR U21469 ( .A(n20265), .B(n20266), .Z(n12446) );
  XNOR U21470 ( .A(n[179]), .B(n20267), .Z(n20263) );
  IV U21471 ( .A(n20262), .Z(n20267) );
  XOR U21472 ( .A(n20268), .B(n20269), .Z(n20262) );
  AND U21473 ( .A(n20270), .B(n20271), .Z(n20268) );
  XOR U21474 ( .A(n20269), .B(n12451), .Z(n20271) );
  XNOR U21475 ( .A(n20272), .B(n20273), .Z(n12451) );
  XNOR U21476 ( .A(n[178]), .B(n20274), .Z(n20270) );
  IV U21477 ( .A(n20269), .Z(n20274) );
  XOR U21478 ( .A(n20275), .B(n20276), .Z(n20269) );
  AND U21479 ( .A(n20277), .B(n20278), .Z(n20275) );
  XOR U21480 ( .A(n20276), .B(n12456), .Z(n20278) );
  XNOR U21481 ( .A(n20279), .B(n20280), .Z(n12456) );
  XNOR U21482 ( .A(n[177]), .B(n20281), .Z(n20277) );
  IV U21483 ( .A(n20276), .Z(n20281) );
  XOR U21484 ( .A(n20282), .B(n20283), .Z(n20276) );
  AND U21485 ( .A(n20284), .B(n20285), .Z(n20282) );
  XOR U21486 ( .A(n20283), .B(n12461), .Z(n20285) );
  XNOR U21487 ( .A(n20286), .B(n20287), .Z(n12461) );
  XNOR U21488 ( .A(n[176]), .B(n20288), .Z(n20284) );
  IV U21489 ( .A(n20283), .Z(n20288) );
  XOR U21490 ( .A(n20289), .B(n20290), .Z(n20283) );
  AND U21491 ( .A(n20291), .B(n20292), .Z(n20289) );
  XOR U21492 ( .A(n20290), .B(n12466), .Z(n20292) );
  XNOR U21493 ( .A(n20293), .B(n20294), .Z(n12466) );
  XNOR U21494 ( .A(n[175]), .B(n20295), .Z(n20291) );
  IV U21495 ( .A(n20290), .Z(n20295) );
  XOR U21496 ( .A(n20296), .B(n20297), .Z(n20290) );
  AND U21497 ( .A(n20298), .B(n20299), .Z(n20296) );
  XOR U21498 ( .A(n20297), .B(n12471), .Z(n20299) );
  XNOR U21499 ( .A(n20300), .B(n20301), .Z(n12471) );
  XNOR U21500 ( .A(n[174]), .B(n20302), .Z(n20298) );
  IV U21501 ( .A(n20297), .Z(n20302) );
  XOR U21502 ( .A(n20303), .B(n20304), .Z(n20297) );
  AND U21503 ( .A(n20305), .B(n20306), .Z(n20303) );
  XOR U21504 ( .A(n20304), .B(n12476), .Z(n20306) );
  XNOR U21505 ( .A(n20307), .B(n20308), .Z(n12476) );
  XNOR U21506 ( .A(n[173]), .B(n20309), .Z(n20305) );
  IV U21507 ( .A(n20304), .Z(n20309) );
  XOR U21508 ( .A(n20310), .B(n20311), .Z(n20304) );
  AND U21509 ( .A(n20312), .B(n20313), .Z(n20310) );
  XOR U21510 ( .A(n20311), .B(n12481), .Z(n20313) );
  XNOR U21511 ( .A(n20314), .B(n20315), .Z(n12481) );
  XNOR U21512 ( .A(n[172]), .B(n20316), .Z(n20312) );
  IV U21513 ( .A(n20311), .Z(n20316) );
  XOR U21514 ( .A(n20317), .B(n20318), .Z(n20311) );
  AND U21515 ( .A(n20319), .B(n20320), .Z(n20317) );
  XOR U21516 ( .A(n20318), .B(n12486), .Z(n20320) );
  XNOR U21517 ( .A(n20321), .B(n20322), .Z(n12486) );
  XNOR U21518 ( .A(n[171]), .B(n20323), .Z(n20319) );
  IV U21519 ( .A(n20318), .Z(n20323) );
  XOR U21520 ( .A(n20324), .B(n20325), .Z(n20318) );
  AND U21521 ( .A(n20326), .B(n20327), .Z(n20324) );
  XOR U21522 ( .A(n20325), .B(n12491), .Z(n20327) );
  XNOR U21523 ( .A(n20328), .B(n20329), .Z(n12491) );
  XNOR U21524 ( .A(n[170]), .B(n20330), .Z(n20326) );
  IV U21525 ( .A(n20325), .Z(n20330) );
  XOR U21526 ( .A(n20331), .B(n20332), .Z(n20325) );
  AND U21527 ( .A(n20333), .B(n20334), .Z(n20331) );
  XOR U21528 ( .A(n20332), .B(n12496), .Z(n20334) );
  XNOR U21529 ( .A(n20335), .B(n20336), .Z(n12496) );
  XNOR U21530 ( .A(n[169]), .B(n20337), .Z(n20333) );
  IV U21531 ( .A(n20332), .Z(n20337) );
  XOR U21532 ( .A(n20338), .B(n20339), .Z(n20332) );
  AND U21533 ( .A(n20340), .B(n20341), .Z(n20338) );
  XOR U21534 ( .A(n20339), .B(n12501), .Z(n20341) );
  XNOR U21535 ( .A(n20342), .B(n20343), .Z(n12501) );
  XNOR U21536 ( .A(n[168]), .B(n20344), .Z(n20340) );
  IV U21537 ( .A(n20339), .Z(n20344) );
  XOR U21538 ( .A(n20345), .B(n20346), .Z(n20339) );
  AND U21539 ( .A(n20347), .B(n20348), .Z(n20345) );
  XOR U21540 ( .A(n20346), .B(n12506), .Z(n20348) );
  XNOR U21541 ( .A(n20349), .B(n20350), .Z(n12506) );
  XNOR U21542 ( .A(n[167]), .B(n20351), .Z(n20347) );
  IV U21543 ( .A(n20346), .Z(n20351) );
  XOR U21544 ( .A(n20352), .B(n20353), .Z(n20346) );
  AND U21545 ( .A(n20354), .B(n20355), .Z(n20352) );
  XOR U21546 ( .A(n20353), .B(n12511), .Z(n20355) );
  XNOR U21547 ( .A(n20356), .B(n20357), .Z(n12511) );
  XNOR U21548 ( .A(n[166]), .B(n20358), .Z(n20354) );
  IV U21549 ( .A(n20353), .Z(n20358) );
  XOR U21550 ( .A(n20359), .B(n20360), .Z(n20353) );
  AND U21551 ( .A(n20361), .B(n20362), .Z(n20359) );
  XOR U21552 ( .A(n20360), .B(n12516), .Z(n20362) );
  XNOR U21553 ( .A(n20363), .B(n20364), .Z(n12516) );
  XNOR U21554 ( .A(n[165]), .B(n20365), .Z(n20361) );
  IV U21555 ( .A(n20360), .Z(n20365) );
  XOR U21556 ( .A(n20366), .B(n20367), .Z(n20360) );
  AND U21557 ( .A(n20368), .B(n20369), .Z(n20366) );
  XOR U21558 ( .A(n20367), .B(n12521), .Z(n20369) );
  XNOR U21559 ( .A(n20370), .B(n20371), .Z(n12521) );
  XNOR U21560 ( .A(n[164]), .B(n20372), .Z(n20368) );
  IV U21561 ( .A(n20367), .Z(n20372) );
  XOR U21562 ( .A(n20373), .B(n20374), .Z(n20367) );
  AND U21563 ( .A(n20375), .B(n20376), .Z(n20373) );
  XOR U21564 ( .A(n20374), .B(n12526), .Z(n20376) );
  XNOR U21565 ( .A(n20377), .B(n20378), .Z(n12526) );
  XNOR U21566 ( .A(n[163]), .B(n20379), .Z(n20375) );
  IV U21567 ( .A(n20374), .Z(n20379) );
  XOR U21568 ( .A(n20380), .B(n20381), .Z(n20374) );
  AND U21569 ( .A(n20382), .B(n20383), .Z(n20380) );
  XOR U21570 ( .A(n20381), .B(n12531), .Z(n20383) );
  XNOR U21571 ( .A(n20384), .B(n20385), .Z(n12531) );
  XNOR U21572 ( .A(n[162]), .B(n20386), .Z(n20382) );
  IV U21573 ( .A(n20381), .Z(n20386) );
  XOR U21574 ( .A(n20387), .B(n20388), .Z(n20381) );
  AND U21575 ( .A(n20389), .B(n20390), .Z(n20387) );
  XOR U21576 ( .A(n20388), .B(n12536), .Z(n20390) );
  XNOR U21577 ( .A(n20391), .B(n20392), .Z(n12536) );
  XNOR U21578 ( .A(n[161]), .B(n20393), .Z(n20389) );
  IV U21579 ( .A(n20388), .Z(n20393) );
  XOR U21580 ( .A(n20394), .B(n20395), .Z(n20388) );
  AND U21581 ( .A(n20396), .B(n20397), .Z(n20394) );
  XOR U21582 ( .A(n20395), .B(n12541), .Z(n20397) );
  XNOR U21583 ( .A(n20398), .B(n20399), .Z(n12541) );
  XNOR U21584 ( .A(n[160]), .B(n20400), .Z(n20396) );
  IV U21585 ( .A(n20395), .Z(n20400) );
  XOR U21586 ( .A(n20401), .B(n20402), .Z(n20395) );
  AND U21587 ( .A(n20403), .B(n20404), .Z(n20401) );
  XOR U21588 ( .A(n20402), .B(n12546), .Z(n20404) );
  XNOR U21589 ( .A(n20405), .B(n20406), .Z(n12546) );
  XNOR U21590 ( .A(n[159]), .B(n20407), .Z(n20403) );
  IV U21591 ( .A(n20402), .Z(n20407) );
  XOR U21592 ( .A(n20408), .B(n20409), .Z(n20402) );
  AND U21593 ( .A(n20410), .B(n20411), .Z(n20408) );
  XOR U21594 ( .A(n20409), .B(n12551), .Z(n20411) );
  XNOR U21595 ( .A(n20412), .B(n20413), .Z(n12551) );
  XNOR U21596 ( .A(n[158]), .B(n20414), .Z(n20410) );
  IV U21597 ( .A(n20409), .Z(n20414) );
  XOR U21598 ( .A(n20415), .B(n20416), .Z(n20409) );
  AND U21599 ( .A(n20417), .B(n20418), .Z(n20415) );
  XOR U21600 ( .A(n20416), .B(n12556), .Z(n20418) );
  XNOR U21601 ( .A(n20419), .B(n20420), .Z(n12556) );
  XNOR U21602 ( .A(n[157]), .B(n20421), .Z(n20417) );
  IV U21603 ( .A(n20416), .Z(n20421) );
  XOR U21604 ( .A(n20422), .B(n20423), .Z(n20416) );
  AND U21605 ( .A(n20424), .B(n20425), .Z(n20422) );
  XOR U21606 ( .A(n20423), .B(n12561), .Z(n20425) );
  XNOR U21607 ( .A(n20426), .B(n20427), .Z(n12561) );
  XNOR U21608 ( .A(n[156]), .B(n20428), .Z(n20424) );
  IV U21609 ( .A(n20423), .Z(n20428) );
  XOR U21610 ( .A(n20429), .B(n20430), .Z(n20423) );
  AND U21611 ( .A(n20431), .B(n20432), .Z(n20429) );
  XOR U21612 ( .A(n20430), .B(n12566), .Z(n20432) );
  XNOR U21613 ( .A(n20433), .B(n20434), .Z(n12566) );
  XNOR U21614 ( .A(n[155]), .B(n20435), .Z(n20431) );
  IV U21615 ( .A(n20430), .Z(n20435) );
  XOR U21616 ( .A(n20436), .B(n20437), .Z(n20430) );
  AND U21617 ( .A(n20438), .B(n20439), .Z(n20436) );
  XOR U21618 ( .A(n20437), .B(n12571), .Z(n20439) );
  XNOR U21619 ( .A(n20440), .B(n20441), .Z(n12571) );
  XNOR U21620 ( .A(n[154]), .B(n20442), .Z(n20438) );
  IV U21621 ( .A(n20437), .Z(n20442) );
  XOR U21622 ( .A(n20443), .B(n20444), .Z(n20437) );
  AND U21623 ( .A(n20445), .B(n20446), .Z(n20443) );
  XOR U21624 ( .A(n20444), .B(n12576), .Z(n20446) );
  XNOR U21625 ( .A(n20447), .B(n20448), .Z(n12576) );
  XNOR U21626 ( .A(n[153]), .B(n20449), .Z(n20445) );
  IV U21627 ( .A(n20444), .Z(n20449) );
  XOR U21628 ( .A(n20450), .B(n20451), .Z(n20444) );
  AND U21629 ( .A(n20452), .B(n20453), .Z(n20450) );
  XOR U21630 ( .A(n20451), .B(n12581), .Z(n20453) );
  XNOR U21631 ( .A(n20454), .B(n20455), .Z(n12581) );
  XNOR U21632 ( .A(n[152]), .B(n20456), .Z(n20452) );
  IV U21633 ( .A(n20451), .Z(n20456) );
  XOR U21634 ( .A(n20457), .B(n20458), .Z(n20451) );
  AND U21635 ( .A(n20459), .B(n20460), .Z(n20457) );
  XOR U21636 ( .A(n20458), .B(n12586), .Z(n20460) );
  XNOR U21637 ( .A(n20461), .B(n20462), .Z(n12586) );
  XNOR U21638 ( .A(n[151]), .B(n20463), .Z(n20459) );
  IV U21639 ( .A(n20458), .Z(n20463) );
  XOR U21640 ( .A(n20464), .B(n20465), .Z(n20458) );
  AND U21641 ( .A(n20466), .B(n20467), .Z(n20464) );
  XOR U21642 ( .A(n20465), .B(n12591), .Z(n20467) );
  XNOR U21643 ( .A(n20468), .B(n20469), .Z(n12591) );
  XNOR U21644 ( .A(n[150]), .B(n20470), .Z(n20466) );
  IV U21645 ( .A(n20465), .Z(n20470) );
  XOR U21646 ( .A(n20471), .B(n20472), .Z(n20465) );
  AND U21647 ( .A(n20473), .B(n20474), .Z(n20471) );
  XOR U21648 ( .A(n20472), .B(n12596), .Z(n20474) );
  XNOR U21649 ( .A(n20475), .B(n20476), .Z(n12596) );
  XNOR U21650 ( .A(n[149]), .B(n20477), .Z(n20473) );
  IV U21651 ( .A(n20472), .Z(n20477) );
  XOR U21652 ( .A(n20478), .B(n20479), .Z(n20472) );
  AND U21653 ( .A(n20480), .B(n20481), .Z(n20478) );
  XOR U21654 ( .A(n20479), .B(n12601), .Z(n20481) );
  XNOR U21655 ( .A(n20482), .B(n20483), .Z(n12601) );
  XNOR U21656 ( .A(n[148]), .B(n20484), .Z(n20480) );
  IV U21657 ( .A(n20479), .Z(n20484) );
  XOR U21658 ( .A(n20485), .B(n20486), .Z(n20479) );
  AND U21659 ( .A(n20487), .B(n20488), .Z(n20485) );
  XOR U21660 ( .A(n20486), .B(n12606), .Z(n20488) );
  XNOR U21661 ( .A(n20489), .B(n20490), .Z(n12606) );
  XNOR U21662 ( .A(n[147]), .B(n20491), .Z(n20487) );
  IV U21663 ( .A(n20486), .Z(n20491) );
  XOR U21664 ( .A(n20492), .B(n20493), .Z(n20486) );
  AND U21665 ( .A(n20494), .B(n20495), .Z(n20492) );
  XOR U21666 ( .A(n20493), .B(n12611), .Z(n20495) );
  XNOR U21667 ( .A(n20496), .B(n20497), .Z(n12611) );
  XNOR U21668 ( .A(n[146]), .B(n20498), .Z(n20494) );
  IV U21669 ( .A(n20493), .Z(n20498) );
  XOR U21670 ( .A(n20499), .B(n20500), .Z(n20493) );
  AND U21671 ( .A(n20501), .B(n20502), .Z(n20499) );
  XOR U21672 ( .A(n20500), .B(n12616), .Z(n20502) );
  XNOR U21673 ( .A(n20503), .B(n20504), .Z(n12616) );
  XNOR U21674 ( .A(n[145]), .B(n20505), .Z(n20501) );
  IV U21675 ( .A(n20500), .Z(n20505) );
  XOR U21676 ( .A(n20506), .B(n20507), .Z(n20500) );
  AND U21677 ( .A(n20508), .B(n20509), .Z(n20506) );
  XOR U21678 ( .A(n20507), .B(n12621), .Z(n20509) );
  XNOR U21679 ( .A(n20510), .B(n20511), .Z(n12621) );
  XNOR U21680 ( .A(n[144]), .B(n20512), .Z(n20508) );
  IV U21681 ( .A(n20507), .Z(n20512) );
  XOR U21682 ( .A(n20513), .B(n20514), .Z(n20507) );
  AND U21683 ( .A(n20515), .B(n20516), .Z(n20513) );
  XOR U21684 ( .A(n20514), .B(n12626), .Z(n20516) );
  XNOR U21685 ( .A(n20517), .B(n20518), .Z(n12626) );
  XNOR U21686 ( .A(n[143]), .B(n20519), .Z(n20515) );
  IV U21687 ( .A(n20514), .Z(n20519) );
  XOR U21688 ( .A(n20520), .B(n20521), .Z(n20514) );
  AND U21689 ( .A(n20522), .B(n20523), .Z(n20520) );
  XOR U21690 ( .A(n20521), .B(n12631), .Z(n20523) );
  XNOR U21691 ( .A(n20524), .B(n20525), .Z(n12631) );
  XNOR U21692 ( .A(n[142]), .B(n20526), .Z(n20522) );
  IV U21693 ( .A(n20521), .Z(n20526) );
  XOR U21694 ( .A(n20527), .B(n20528), .Z(n20521) );
  AND U21695 ( .A(n20529), .B(n20530), .Z(n20527) );
  XOR U21696 ( .A(n20528), .B(n12636), .Z(n20530) );
  XNOR U21697 ( .A(n20531), .B(n20532), .Z(n12636) );
  XNOR U21698 ( .A(n[141]), .B(n20533), .Z(n20529) );
  IV U21699 ( .A(n20528), .Z(n20533) );
  XOR U21700 ( .A(n20534), .B(n20535), .Z(n20528) );
  AND U21701 ( .A(n20536), .B(n20537), .Z(n20534) );
  XOR U21702 ( .A(n20535), .B(n12641), .Z(n20537) );
  XNOR U21703 ( .A(n20538), .B(n20539), .Z(n12641) );
  XNOR U21704 ( .A(n[140]), .B(n20540), .Z(n20536) );
  IV U21705 ( .A(n20535), .Z(n20540) );
  XOR U21706 ( .A(n20541), .B(n20542), .Z(n20535) );
  AND U21707 ( .A(n20543), .B(n20544), .Z(n20541) );
  XOR U21708 ( .A(n20542), .B(n12646), .Z(n20544) );
  XNOR U21709 ( .A(n20545), .B(n20546), .Z(n12646) );
  XNOR U21710 ( .A(n[139]), .B(n20547), .Z(n20543) );
  IV U21711 ( .A(n20542), .Z(n20547) );
  XOR U21712 ( .A(n20548), .B(n20549), .Z(n20542) );
  AND U21713 ( .A(n20550), .B(n20551), .Z(n20548) );
  XOR U21714 ( .A(n20549), .B(n12651), .Z(n20551) );
  XNOR U21715 ( .A(n20552), .B(n20553), .Z(n12651) );
  XNOR U21716 ( .A(n[138]), .B(n20554), .Z(n20550) );
  IV U21717 ( .A(n20549), .Z(n20554) );
  XOR U21718 ( .A(n20555), .B(n20556), .Z(n20549) );
  AND U21719 ( .A(n20557), .B(n20558), .Z(n20555) );
  XOR U21720 ( .A(n20556), .B(n12656), .Z(n20558) );
  XNOR U21721 ( .A(n20559), .B(n20560), .Z(n12656) );
  XNOR U21722 ( .A(n[137]), .B(n20561), .Z(n20557) );
  IV U21723 ( .A(n20556), .Z(n20561) );
  XOR U21724 ( .A(n20562), .B(n20563), .Z(n20556) );
  AND U21725 ( .A(n20564), .B(n20565), .Z(n20562) );
  XOR U21726 ( .A(n20563), .B(n12661), .Z(n20565) );
  XNOR U21727 ( .A(n20566), .B(n20567), .Z(n12661) );
  XNOR U21728 ( .A(n[136]), .B(n20568), .Z(n20564) );
  IV U21729 ( .A(n20563), .Z(n20568) );
  XOR U21730 ( .A(n20569), .B(n20570), .Z(n20563) );
  AND U21731 ( .A(n20571), .B(n20572), .Z(n20569) );
  XOR U21732 ( .A(n20570), .B(n12666), .Z(n20572) );
  XNOR U21733 ( .A(n20573), .B(n20574), .Z(n12666) );
  XNOR U21734 ( .A(n[135]), .B(n20575), .Z(n20571) );
  IV U21735 ( .A(n20570), .Z(n20575) );
  XOR U21736 ( .A(n20576), .B(n20577), .Z(n20570) );
  AND U21737 ( .A(n20578), .B(n20579), .Z(n20576) );
  XOR U21738 ( .A(n20577), .B(n12671), .Z(n20579) );
  XNOR U21739 ( .A(n20580), .B(n20581), .Z(n12671) );
  XNOR U21740 ( .A(n[134]), .B(n20582), .Z(n20578) );
  IV U21741 ( .A(n20577), .Z(n20582) );
  XOR U21742 ( .A(n20583), .B(n20584), .Z(n20577) );
  AND U21743 ( .A(n20585), .B(n20586), .Z(n20583) );
  XOR U21744 ( .A(n20584), .B(n12676), .Z(n20586) );
  XNOR U21745 ( .A(n20587), .B(n20588), .Z(n12676) );
  XNOR U21746 ( .A(n[133]), .B(n20589), .Z(n20585) );
  IV U21747 ( .A(n20584), .Z(n20589) );
  XOR U21748 ( .A(n20590), .B(n20591), .Z(n20584) );
  AND U21749 ( .A(n20592), .B(n20593), .Z(n20590) );
  XOR U21750 ( .A(n20591), .B(n12681), .Z(n20593) );
  XNOR U21751 ( .A(n20594), .B(n20595), .Z(n12681) );
  XNOR U21752 ( .A(n[132]), .B(n20596), .Z(n20592) );
  IV U21753 ( .A(n20591), .Z(n20596) );
  XOR U21754 ( .A(n20597), .B(n20598), .Z(n20591) );
  AND U21755 ( .A(n20599), .B(n20600), .Z(n20597) );
  XOR U21756 ( .A(n20598), .B(n12686), .Z(n20600) );
  XNOR U21757 ( .A(n20601), .B(n20602), .Z(n12686) );
  XNOR U21758 ( .A(n[131]), .B(n20603), .Z(n20599) );
  IV U21759 ( .A(n20598), .Z(n20603) );
  XOR U21760 ( .A(n20604), .B(n20605), .Z(n20598) );
  AND U21761 ( .A(n20606), .B(n20607), .Z(n20604) );
  XOR U21762 ( .A(n20605), .B(n12691), .Z(n20607) );
  XNOR U21763 ( .A(n20608), .B(n20609), .Z(n12691) );
  XNOR U21764 ( .A(n[130]), .B(n20610), .Z(n20606) );
  IV U21765 ( .A(n20605), .Z(n20610) );
  XOR U21766 ( .A(n20611), .B(n20612), .Z(n20605) );
  AND U21767 ( .A(n20613), .B(n20614), .Z(n20611) );
  XOR U21768 ( .A(n20612), .B(n12696), .Z(n20614) );
  XNOR U21769 ( .A(n20615), .B(n20616), .Z(n12696) );
  XNOR U21770 ( .A(n[129]), .B(n20617), .Z(n20613) );
  IV U21771 ( .A(n20612), .Z(n20617) );
  XOR U21772 ( .A(n20618), .B(n20619), .Z(n20612) );
  AND U21773 ( .A(n20620), .B(n20621), .Z(n20618) );
  XOR U21774 ( .A(n20619), .B(n12701), .Z(n20621) );
  XNOR U21775 ( .A(n20622), .B(n20623), .Z(n12701) );
  XNOR U21776 ( .A(n[128]), .B(n20624), .Z(n20620) );
  IV U21777 ( .A(n20619), .Z(n20624) );
  XOR U21778 ( .A(n20625), .B(n20626), .Z(n20619) );
  AND U21779 ( .A(n20627), .B(n20628), .Z(n20625) );
  XOR U21780 ( .A(n20626), .B(n12706), .Z(n20628) );
  XNOR U21781 ( .A(n20629), .B(n20630), .Z(n12706) );
  XNOR U21782 ( .A(n[127]), .B(n20631), .Z(n20627) );
  IV U21783 ( .A(n20626), .Z(n20631) );
  XOR U21784 ( .A(n20632), .B(n20633), .Z(n20626) );
  AND U21785 ( .A(n20634), .B(n20635), .Z(n20632) );
  XOR U21786 ( .A(n20633), .B(n12711), .Z(n20635) );
  XNOR U21787 ( .A(n20636), .B(n20637), .Z(n12711) );
  XNOR U21788 ( .A(n[126]), .B(n20638), .Z(n20634) );
  IV U21789 ( .A(n20633), .Z(n20638) );
  XOR U21790 ( .A(n20639), .B(n20640), .Z(n20633) );
  AND U21791 ( .A(n20641), .B(n20642), .Z(n20639) );
  XOR U21792 ( .A(n20640), .B(n12716), .Z(n20642) );
  XNOR U21793 ( .A(n20643), .B(n20644), .Z(n12716) );
  XNOR U21794 ( .A(n[125]), .B(n20645), .Z(n20641) );
  IV U21795 ( .A(n20640), .Z(n20645) );
  XOR U21796 ( .A(n20646), .B(n20647), .Z(n20640) );
  AND U21797 ( .A(n20648), .B(n20649), .Z(n20646) );
  XOR U21798 ( .A(n20647), .B(n12721), .Z(n20649) );
  XNOR U21799 ( .A(n20650), .B(n20651), .Z(n12721) );
  XNOR U21800 ( .A(n[124]), .B(n20652), .Z(n20648) );
  IV U21801 ( .A(n20647), .Z(n20652) );
  XOR U21802 ( .A(n20653), .B(n20654), .Z(n20647) );
  AND U21803 ( .A(n20655), .B(n20656), .Z(n20653) );
  XOR U21804 ( .A(n20654), .B(n12726), .Z(n20656) );
  XNOR U21805 ( .A(n20657), .B(n20658), .Z(n12726) );
  XNOR U21806 ( .A(n[123]), .B(n20659), .Z(n20655) );
  IV U21807 ( .A(n20654), .Z(n20659) );
  XOR U21808 ( .A(n20660), .B(n20661), .Z(n20654) );
  AND U21809 ( .A(n20662), .B(n20663), .Z(n20660) );
  XOR U21810 ( .A(n20661), .B(n12731), .Z(n20663) );
  XNOR U21811 ( .A(n20664), .B(n20665), .Z(n12731) );
  XNOR U21812 ( .A(n[122]), .B(n20666), .Z(n20662) );
  IV U21813 ( .A(n20661), .Z(n20666) );
  XOR U21814 ( .A(n20667), .B(n20668), .Z(n20661) );
  AND U21815 ( .A(n20669), .B(n20670), .Z(n20667) );
  XOR U21816 ( .A(n20668), .B(n12736), .Z(n20670) );
  XNOR U21817 ( .A(n20671), .B(n20672), .Z(n12736) );
  XNOR U21818 ( .A(n[121]), .B(n20673), .Z(n20669) );
  IV U21819 ( .A(n20668), .Z(n20673) );
  XOR U21820 ( .A(n20674), .B(n20675), .Z(n20668) );
  AND U21821 ( .A(n20676), .B(n20677), .Z(n20674) );
  XOR U21822 ( .A(n20675), .B(n12741), .Z(n20677) );
  XNOR U21823 ( .A(n20678), .B(n20679), .Z(n12741) );
  XNOR U21824 ( .A(n[120]), .B(n20680), .Z(n20676) );
  IV U21825 ( .A(n20675), .Z(n20680) );
  XOR U21826 ( .A(n20681), .B(n20682), .Z(n20675) );
  AND U21827 ( .A(n20683), .B(n20684), .Z(n20681) );
  XOR U21828 ( .A(n20682), .B(n12746), .Z(n20684) );
  XNOR U21829 ( .A(n20685), .B(n20686), .Z(n12746) );
  XNOR U21830 ( .A(n[119]), .B(n20687), .Z(n20683) );
  IV U21831 ( .A(n20682), .Z(n20687) );
  XOR U21832 ( .A(n20688), .B(n20689), .Z(n20682) );
  AND U21833 ( .A(n20690), .B(n20691), .Z(n20688) );
  XOR U21834 ( .A(n20689), .B(n12751), .Z(n20691) );
  XNOR U21835 ( .A(n20692), .B(n20693), .Z(n12751) );
  XNOR U21836 ( .A(n[118]), .B(n20694), .Z(n20690) );
  IV U21837 ( .A(n20689), .Z(n20694) );
  XOR U21838 ( .A(n20695), .B(n20696), .Z(n20689) );
  AND U21839 ( .A(n20697), .B(n20698), .Z(n20695) );
  XOR U21840 ( .A(n20696), .B(n12756), .Z(n20698) );
  XNOR U21841 ( .A(n20699), .B(n20700), .Z(n12756) );
  XNOR U21842 ( .A(n[117]), .B(n20701), .Z(n20697) );
  IV U21843 ( .A(n20696), .Z(n20701) );
  XOR U21844 ( .A(n20702), .B(n20703), .Z(n20696) );
  AND U21845 ( .A(n20704), .B(n20705), .Z(n20702) );
  XOR U21846 ( .A(n20703), .B(n12761), .Z(n20705) );
  XNOR U21847 ( .A(n20706), .B(n20707), .Z(n12761) );
  XNOR U21848 ( .A(n[116]), .B(n20708), .Z(n20704) );
  IV U21849 ( .A(n20703), .Z(n20708) );
  XOR U21850 ( .A(n20709), .B(n20710), .Z(n20703) );
  AND U21851 ( .A(n20711), .B(n20712), .Z(n20709) );
  XOR U21852 ( .A(n20710), .B(n12766), .Z(n20712) );
  XNOR U21853 ( .A(n20713), .B(n20714), .Z(n12766) );
  XNOR U21854 ( .A(n[115]), .B(n20715), .Z(n20711) );
  IV U21855 ( .A(n20710), .Z(n20715) );
  XOR U21856 ( .A(n20716), .B(n20717), .Z(n20710) );
  AND U21857 ( .A(n20718), .B(n20719), .Z(n20716) );
  XOR U21858 ( .A(n20717), .B(n12771), .Z(n20719) );
  XNOR U21859 ( .A(n20720), .B(n20721), .Z(n12771) );
  XNOR U21860 ( .A(n[114]), .B(n20722), .Z(n20718) );
  IV U21861 ( .A(n20717), .Z(n20722) );
  XOR U21862 ( .A(n20723), .B(n20724), .Z(n20717) );
  AND U21863 ( .A(n20725), .B(n20726), .Z(n20723) );
  XOR U21864 ( .A(n20724), .B(n12776), .Z(n20726) );
  XNOR U21865 ( .A(n20727), .B(n20728), .Z(n12776) );
  XNOR U21866 ( .A(n[113]), .B(n20729), .Z(n20725) );
  IV U21867 ( .A(n20724), .Z(n20729) );
  XOR U21868 ( .A(n20730), .B(n20731), .Z(n20724) );
  AND U21869 ( .A(n20732), .B(n20733), .Z(n20730) );
  XOR U21870 ( .A(n20731), .B(n12781), .Z(n20733) );
  XNOR U21871 ( .A(n20734), .B(n20735), .Z(n12781) );
  XNOR U21872 ( .A(n[112]), .B(n20736), .Z(n20732) );
  IV U21873 ( .A(n20731), .Z(n20736) );
  XOR U21874 ( .A(n20737), .B(n20738), .Z(n20731) );
  AND U21875 ( .A(n20739), .B(n20740), .Z(n20737) );
  XOR U21876 ( .A(n20738), .B(n12786), .Z(n20740) );
  XNOR U21877 ( .A(n20741), .B(n20742), .Z(n12786) );
  XNOR U21878 ( .A(n[111]), .B(n20743), .Z(n20739) );
  IV U21879 ( .A(n20738), .Z(n20743) );
  XOR U21880 ( .A(n20744), .B(n20745), .Z(n20738) );
  AND U21881 ( .A(n20746), .B(n20747), .Z(n20744) );
  XOR U21882 ( .A(n20745), .B(n12791), .Z(n20747) );
  XNOR U21883 ( .A(n20748), .B(n20749), .Z(n12791) );
  XNOR U21884 ( .A(n[110]), .B(n20750), .Z(n20746) );
  IV U21885 ( .A(n20745), .Z(n20750) );
  XOR U21886 ( .A(n20751), .B(n20752), .Z(n20745) );
  AND U21887 ( .A(n20753), .B(n20754), .Z(n20751) );
  XOR U21888 ( .A(n20752), .B(n12796), .Z(n20754) );
  XNOR U21889 ( .A(n20755), .B(n20756), .Z(n12796) );
  XNOR U21890 ( .A(n[109]), .B(n20757), .Z(n20753) );
  IV U21891 ( .A(n20752), .Z(n20757) );
  XOR U21892 ( .A(n20758), .B(n20759), .Z(n20752) );
  AND U21893 ( .A(n20760), .B(n20761), .Z(n20758) );
  XOR U21894 ( .A(n20759), .B(n12801), .Z(n20761) );
  XNOR U21895 ( .A(n20762), .B(n20763), .Z(n12801) );
  XNOR U21896 ( .A(n[108]), .B(n20764), .Z(n20760) );
  IV U21897 ( .A(n20759), .Z(n20764) );
  XOR U21898 ( .A(n20765), .B(n20766), .Z(n20759) );
  AND U21899 ( .A(n20767), .B(n20768), .Z(n20765) );
  XOR U21900 ( .A(n20766), .B(n12806), .Z(n20768) );
  XNOR U21901 ( .A(n20769), .B(n20770), .Z(n12806) );
  XNOR U21902 ( .A(n[107]), .B(n20771), .Z(n20767) );
  IV U21903 ( .A(n20766), .Z(n20771) );
  XOR U21904 ( .A(n20772), .B(n20773), .Z(n20766) );
  AND U21905 ( .A(n20774), .B(n20775), .Z(n20772) );
  XOR U21906 ( .A(n20773), .B(n12811), .Z(n20775) );
  XNOR U21907 ( .A(n20776), .B(n20777), .Z(n12811) );
  XNOR U21908 ( .A(n[106]), .B(n20778), .Z(n20774) );
  IV U21909 ( .A(n20773), .Z(n20778) );
  XOR U21910 ( .A(n20779), .B(n20780), .Z(n20773) );
  AND U21911 ( .A(n20781), .B(n20782), .Z(n20779) );
  XOR U21912 ( .A(n20780), .B(n12816), .Z(n20782) );
  XNOR U21913 ( .A(n20783), .B(n20784), .Z(n12816) );
  XNOR U21914 ( .A(n[105]), .B(n20785), .Z(n20781) );
  IV U21915 ( .A(n20780), .Z(n20785) );
  XOR U21916 ( .A(n20786), .B(n20787), .Z(n20780) );
  AND U21917 ( .A(n20788), .B(n20789), .Z(n20786) );
  XOR U21918 ( .A(n20787), .B(n12821), .Z(n20789) );
  XNOR U21919 ( .A(n20790), .B(n20791), .Z(n12821) );
  XNOR U21920 ( .A(n[104]), .B(n20792), .Z(n20788) );
  IV U21921 ( .A(n20787), .Z(n20792) );
  XOR U21922 ( .A(n20793), .B(n20794), .Z(n20787) );
  AND U21923 ( .A(n20795), .B(n20796), .Z(n20793) );
  XOR U21924 ( .A(n20794), .B(n12826), .Z(n20796) );
  XNOR U21925 ( .A(n20797), .B(n20798), .Z(n12826) );
  XNOR U21926 ( .A(n[103]), .B(n20799), .Z(n20795) );
  IV U21927 ( .A(n20794), .Z(n20799) );
  XOR U21928 ( .A(n20800), .B(n20801), .Z(n20794) );
  AND U21929 ( .A(n20802), .B(n20803), .Z(n20800) );
  XOR U21930 ( .A(n20801), .B(n12831), .Z(n20803) );
  XNOR U21931 ( .A(n20804), .B(n20805), .Z(n12831) );
  XNOR U21932 ( .A(n[102]), .B(n20806), .Z(n20802) );
  IV U21933 ( .A(n20801), .Z(n20806) );
  XOR U21934 ( .A(n20807), .B(n20808), .Z(n20801) );
  AND U21935 ( .A(n20809), .B(n20810), .Z(n20807) );
  XOR U21936 ( .A(n20808), .B(n12836), .Z(n20810) );
  XNOR U21937 ( .A(n20811), .B(n20812), .Z(n12836) );
  XNOR U21938 ( .A(n[101]), .B(n20813), .Z(n20809) );
  IV U21939 ( .A(n20808), .Z(n20813) );
  XOR U21940 ( .A(n20814), .B(n20815), .Z(n20808) );
  AND U21941 ( .A(n20816), .B(n20817), .Z(n20814) );
  XOR U21942 ( .A(n20815), .B(n12841), .Z(n20817) );
  XNOR U21943 ( .A(n20818), .B(n20819), .Z(n12841) );
  XNOR U21944 ( .A(n[100]), .B(n20820), .Z(n20816) );
  IV U21945 ( .A(n20815), .Z(n20820) );
  XOR U21946 ( .A(n20821), .B(n20822), .Z(n20815) );
  AND U21947 ( .A(n20823), .B(n20824), .Z(n20821) );
  XOR U21948 ( .A(n20822), .B(n12846), .Z(n20824) );
  XNOR U21949 ( .A(n20825), .B(n20826), .Z(n12846) );
  XNOR U21950 ( .A(n[99]), .B(n20827), .Z(n20823) );
  IV U21951 ( .A(n20822), .Z(n20827) );
  XOR U21952 ( .A(n20828), .B(n20829), .Z(n20822) );
  AND U21953 ( .A(n20830), .B(n20831), .Z(n20828) );
  XOR U21954 ( .A(n20829), .B(n12851), .Z(n20831) );
  XNOR U21955 ( .A(n20832), .B(n20833), .Z(n12851) );
  XNOR U21956 ( .A(n[98]), .B(n20834), .Z(n20830) );
  IV U21957 ( .A(n20829), .Z(n20834) );
  XOR U21958 ( .A(n20835), .B(n20836), .Z(n20829) );
  AND U21959 ( .A(n20837), .B(n20838), .Z(n20835) );
  XOR U21960 ( .A(n20836), .B(n12856), .Z(n20838) );
  XNOR U21961 ( .A(n20839), .B(n20840), .Z(n12856) );
  XNOR U21962 ( .A(n[97]), .B(n20841), .Z(n20837) );
  IV U21963 ( .A(n20836), .Z(n20841) );
  XOR U21964 ( .A(n20842), .B(n20843), .Z(n20836) );
  AND U21965 ( .A(n20844), .B(n20845), .Z(n20842) );
  XOR U21966 ( .A(n20843), .B(n12861), .Z(n20845) );
  XNOR U21967 ( .A(n20846), .B(n20847), .Z(n12861) );
  XNOR U21968 ( .A(n[96]), .B(n20848), .Z(n20844) );
  IV U21969 ( .A(n20843), .Z(n20848) );
  XOR U21970 ( .A(n20849), .B(n20850), .Z(n20843) );
  AND U21971 ( .A(n20851), .B(n20852), .Z(n20849) );
  XOR U21972 ( .A(n20850), .B(n12866), .Z(n20852) );
  XNOR U21973 ( .A(n20853), .B(n20854), .Z(n12866) );
  XNOR U21974 ( .A(n[95]), .B(n20855), .Z(n20851) );
  IV U21975 ( .A(n20850), .Z(n20855) );
  XOR U21976 ( .A(n20856), .B(n20857), .Z(n20850) );
  AND U21977 ( .A(n20858), .B(n20859), .Z(n20856) );
  XOR U21978 ( .A(n20857), .B(n12871), .Z(n20859) );
  XNOR U21979 ( .A(n20860), .B(n20861), .Z(n12871) );
  XNOR U21980 ( .A(n[94]), .B(n20862), .Z(n20858) );
  IV U21981 ( .A(n20857), .Z(n20862) );
  XOR U21982 ( .A(n20863), .B(n20864), .Z(n20857) );
  AND U21983 ( .A(n20865), .B(n20866), .Z(n20863) );
  XOR U21984 ( .A(n20864), .B(n12876), .Z(n20866) );
  XNOR U21985 ( .A(n20867), .B(n20868), .Z(n12876) );
  XNOR U21986 ( .A(n[93]), .B(n20869), .Z(n20865) );
  IV U21987 ( .A(n20864), .Z(n20869) );
  XOR U21988 ( .A(n20870), .B(n20871), .Z(n20864) );
  AND U21989 ( .A(n20872), .B(n20873), .Z(n20870) );
  XOR U21990 ( .A(n20871), .B(n12881), .Z(n20873) );
  XNOR U21991 ( .A(n20874), .B(n20875), .Z(n12881) );
  XNOR U21992 ( .A(n[92]), .B(n20876), .Z(n20872) );
  IV U21993 ( .A(n20871), .Z(n20876) );
  XOR U21994 ( .A(n20877), .B(n20878), .Z(n20871) );
  AND U21995 ( .A(n20879), .B(n20880), .Z(n20877) );
  XOR U21996 ( .A(n20878), .B(n12886), .Z(n20880) );
  XNOR U21997 ( .A(n20881), .B(n20882), .Z(n12886) );
  XNOR U21998 ( .A(n[91]), .B(n20883), .Z(n20879) );
  IV U21999 ( .A(n20878), .Z(n20883) );
  XOR U22000 ( .A(n20884), .B(n20885), .Z(n20878) );
  AND U22001 ( .A(n20886), .B(n20887), .Z(n20884) );
  XOR U22002 ( .A(n20885), .B(n12891), .Z(n20887) );
  XNOR U22003 ( .A(n20888), .B(n20889), .Z(n12891) );
  XNOR U22004 ( .A(n[90]), .B(n20890), .Z(n20886) );
  IV U22005 ( .A(n20885), .Z(n20890) );
  XOR U22006 ( .A(n20891), .B(n20892), .Z(n20885) );
  AND U22007 ( .A(n20893), .B(n20894), .Z(n20891) );
  XOR U22008 ( .A(n20892), .B(n12896), .Z(n20894) );
  XNOR U22009 ( .A(n20895), .B(n20896), .Z(n12896) );
  XNOR U22010 ( .A(n[89]), .B(n20897), .Z(n20893) );
  IV U22011 ( .A(n20892), .Z(n20897) );
  XOR U22012 ( .A(n20898), .B(n20899), .Z(n20892) );
  AND U22013 ( .A(n20900), .B(n20901), .Z(n20898) );
  XOR U22014 ( .A(n20899), .B(n12901), .Z(n20901) );
  XNOR U22015 ( .A(n20902), .B(n20903), .Z(n12901) );
  XNOR U22016 ( .A(n[88]), .B(n20904), .Z(n20900) );
  IV U22017 ( .A(n20899), .Z(n20904) );
  XOR U22018 ( .A(n20905), .B(n20906), .Z(n20899) );
  AND U22019 ( .A(n20907), .B(n20908), .Z(n20905) );
  XOR U22020 ( .A(n20906), .B(n12906), .Z(n20908) );
  XNOR U22021 ( .A(n20909), .B(n20910), .Z(n12906) );
  XNOR U22022 ( .A(n[87]), .B(n20911), .Z(n20907) );
  IV U22023 ( .A(n20906), .Z(n20911) );
  XOR U22024 ( .A(n20912), .B(n20913), .Z(n20906) );
  AND U22025 ( .A(n20914), .B(n20915), .Z(n20912) );
  XOR U22026 ( .A(n20913), .B(n12911), .Z(n20915) );
  XNOR U22027 ( .A(n20916), .B(n20917), .Z(n12911) );
  XNOR U22028 ( .A(n[86]), .B(n20918), .Z(n20914) );
  IV U22029 ( .A(n20913), .Z(n20918) );
  XOR U22030 ( .A(n20919), .B(n20920), .Z(n20913) );
  AND U22031 ( .A(n20921), .B(n20922), .Z(n20919) );
  XOR U22032 ( .A(n20920), .B(n12916), .Z(n20922) );
  XNOR U22033 ( .A(n20923), .B(n20924), .Z(n12916) );
  XNOR U22034 ( .A(n[85]), .B(n20925), .Z(n20921) );
  IV U22035 ( .A(n20920), .Z(n20925) );
  XOR U22036 ( .A(n20926), .B(n20927), .Z(n20920) );
  AND U22037 ( .A(n20928), .B(n20929), .Z(n20926) );
  XOR U22038 ( .A(n20927), .B(n12921), .Z(n20929) );
  XNOR U22039 ( .A(n20930), .B(n20931), .Z(n12921) );
  XNOR U22040 ( .A(n[84]), .B(n20932), .Z(n20928) );
  IV U22041 ( .A(n20927), .Z(n20932) );
  XOR U22042 ( .A(n20933), .B(n20934), .Z(n20927) );
  AND U22043 ( .A(n20935), .B(n20936), .Z(n20933) );
  XOR U22044 ( .A(n20934), .B(n12926), .Z(n20936) );
  XNOR U22045 ( .A(n20937), .B(n20938), .Z(n12926) );
  XNOR U22046 ( .A(n[83]), .B(n20939), .Z(n20935) );
  IV U22047 ( .A(n20934), .Z(n20939) );
  XOR U22048 ( .A(n20940), .B(n20941), .Z(n20934) );
  AND U22049 ( .A(n20942), .B(n20943), .Z(n20940) );
  XOR U22050 ( .A(n20941), .B(n12931), .Z(n20943) );
  XNOR U22051 ( .A(n20944), .B(n20945), .Z(n12931) );
  XNOR U22052 ( .A(n[82]), .B(n20946), .Z(n20942) );
  IV U22053 ( .A(n20941), .Z(n20946) );
  XOR U22054 ( .A(n20947), .B(n20948), .Z(n20941) );
  AND U22055 ( .A(n20949), .B(n20950), .Z(n20947) );
  XOR U22056 ( .A(n20948), .B(n12936), .Z(n20950) );
  XNOR U22057 ( .A(n20951), .B(n20952), .Z(n12936) );
  XNOR U22058 ( .A(n[81]), .B(n20953), .Z(n20949) );
  IV U22059 ( .A(n20948), .Z(n20953) );
  XOR U22060 ( .A(n20954), .B(n20955), .Z(n20948) );
  AND U22061 ( .A(n20956), .B(n20957), .Z(n20954) );
  XOR U22062 ( .A(n20955), .B(n12941), .Z(n20957) );
  XNOR U22063 ( .A(n20958), .B(n20959), .Z(n12941) );
  XNOR U22064 ( .A(n[80]), .B(n20960), .Z(n20956) );
  IV U22065 ( .A(n20955), .Z(n20960) );
  XOR U22066 ( .A(n20961), .B(n20962), .Z(n20955) );
  AND U22067 ( .A(n20963), .B(n20964), .Z(n20961) );
  XOR U22068 ( .A(n20962), .B(n12946), .Z(n20964) );
  XNOR U22069 ( .A(n20965), .B(n20966), .Z(n12946) );
  XNOR U22070 ( .A(n[79]), .B(n20967), .Z(n20963) );
  IV U22071 ( .A(n20962), .Z(n20967) );
  XOR U22072 ( .A(n20968), .B(n20969), .Z(n20962) );
  AND U22073 ( .A(n20970), .B(n20971), .Z(n20968) );
  XOR U22074 ( .A(n20969), .B(n12951), .Z(n20971) );
  XNOR U22075 ( .A(n20972), .B(n20973), .Z(n12951) );
  XNOR U22076 ( .A(n[78]), .B(n20974), .Z(n20970) );
  IV U22077 ( .A(n20969), .Z(n20974) );
  XOR U22078 ( .A(n20975), .B(n20976), .Z(n20969) );
  AND U22079 ( .A(n20977), .B(n20978), .Z(n20975) );
  XOR U22080 ( .A(n20976), .B(n12956), .Z(n20978) );
  XNOR U22081 ( .A(n20979), .B(n20980), .Z(n12956) );
  XNOR U22082 ( .A(n[77]), .B(n20981), .Z(n20977) );
  IV U22083 ( .A(n20976), .Z(n20981) );
  XOR U22084 ( .A(n20982), .B(n20983), .Z(n20976) );
  AND U22085 ( .A(n20984), .B(n20985), .Z(n20982) );
  XOR U22086 ( .A(n20983), .B(n12961), .Z(n20985) );
  XNOR U22087 ( .A(n20986), .B(n20987), .Z(n12961) );
  XNOR U22088 ( .A(n[76]), .B(n20988), .Z(n20984) );
  IV U22089 ( .A(n20983), .Z(n20988) );
  XOR U22090 ( .A(n20989), .B(n20990), .Z(n20983) );
  AND U22091 ( .A(n20991), .B(n20992), .Z(n20989) );
  XOR U22092 ( .A(n20990), .B(n12966), .Z(n20992) );
  XNOR U22093 ( .A(n20993), .B(n20994), .Z(n12966) );
  XNOR U22094 ( .A(n[75]), .B(n20995), .Z(n20991) );
  IV U22095 ( .A(n20990), .Z(n20995) );
  XOR U22096 ( .A(n20996), .B(n20997), .Z(n20990) );
  AND U22097 ( .A(n20998), .B(n20999), .Z(n20996) );
  XOR U22098 ( .A(n20997), .B(n12971), .Z(n20999) );
  XNOR U22099 ( .A(n21000), .B(n21001), .Z(n12971) );
  XNOR U22100 ( .A(n[74]), .B(n21002), .Z(n20998) );
  IV U22101 ( .A(n20997), .Z(n21002) );
  XOR U22102 ( .A(n21003), .B(n21004), .Z(n20997) );
  AND U22103 ( .A(n21005), .B(n21006), .Z(n21003) );
  XOR U22104 ( .A(n21004), .B(n12976), .Z(n21006) );
  XNOR U22105 ( .A(n21007), .B(n21008), .Z(n12976) );
  XNOR U22106 ( .A(n[73]), .B(n21009), .Z(n21005) );
  IV U22107 ( .A(n21004), .Z(n21009) );
  XOR U22108 ( .A(n21010), .B(n21011), .Z(n21004) );
  AND U22109 ( .A(n21012), .B(n21013), .Z(n21010) );
  XOR U22110 ( .A(n21011), .B(n12981), .Z(n21013) );
  XNOR U22111 ( .A(n21014), .B(n21015), .Z(n12981) );
  XNOR U22112 ( .A(n[72]), .B(n21016), .Z(n21012) );
  IV U22113 ( .A(n21011), .Z(n21016) );
  XOR U22114 ( .A(n21017), .B(n21018), .Z(n21011) );
  AND U22115 ( .A(n21019), .B(n21020), .Z(n21017) );
  XOR U22116 ( .A(n21018), .B(n12986), .Z(n21020) );
  XNOR U22117 ( .A(n21021), .B(n21022), .Z(n12986) );
  XNOR U22118 ( .A(n[71]), .B(n21023), .Z(n21019) );
  IV U22119 ( .A(n21018), .Z(n21023) );
  XOR U22120 ( .A(n21024), .B(n21025), .Z(n21018) );
  AND U22121 ( .A(n21026), .B(n21027), .Z(n21024) );
  XOR U22122 ( .A(n21025), .B(n12991), .Z(n21027) );
  XNOR U22123 ( .A(n21028), .B(n21029), .Z(n12991) );
  XNOR U22124 ( .A(n[70]), .B(n21030), .Z(n21026) );
  IV U22125 ( .A(n21025), .Z(n21030) );
  XOR U22126 ( .A(n21031), .B(n21032), .Z(n21025) );
  AND U22127 ( .A(n21033), .B(n21034), .Z(n21031) );
  XOR U22128 ( .A(n21032), .B(n12996), .Z(n21034) );
  XNOR U22129 ( .A(n21035), .B(n21036), .Z(n12996) );
  XNOR U22130 ( .A(n[69]), .B(n21037), .Z(n21033) );
  IV U22131 ( .A(n21032), .Z(n21037) );
  XOR U22132 ( .A(n21038), .B(n21039), .Z(n21032) );
  AND U22133 ( .A(n21040), .B(n21041), .Z(n21038) );
  XOR U22134 ( .A(n21039), .B(n13001), .Z(n21041) );
  XNOR U22135 ( .A(n21042), .B(n21043), .Z(n13001) );
  XNOR U22136 ( .A(n[68]), .B(n21044), .Z(n21040) );
  IV U22137 ( .A(n21039), .Z(n21044) );
  XOR U22138 ( .A(n21045), .B(n21046), .Z(n21039) );
  AND U22139 ( .A(n21047), .B(n21048), .Z(n21045) );
  XOR U22140 ( .A(n21046), .B(n13006), .Z(n21048) );
  XNOR U22141 ( .A(n21049), .B(n21050), .Z(n13006) );
  XNOR U22142 ( .A(n[67]), .B(n21051), .Z(n21047) );
  IV U22143 ( .A(n21046), .Z(n21051) );
  XOR U22144 ( .A(n21052), .B(n21053), .Z(n21046) );
  AND U22145 ( .A(n21054), .B(n21055), .Z(n21052) );
  XOR U22146 ( .A(n21053), .B(n13011), .Z(n21055) );
  XNOR U22147 ( .A(n21056), .B(n21057), .Z(n13011) );
  XNOR U22148 ( .A(n[66]), .B(n21058), .Z(n21054) );
  IV U22149 ( .A(n21053), .Z(n21058) );
  XOR U22150 ( .A(n21059), .B(n21060), .Z(n21053) );
  AND U22151 ( .A(n21061), .B(n21062), .Z(n21059) );
  XOR U22152 ( .A(n21060), .B(n13016), .Z(n21062) );
  XNOR U22153 ( .A(n21063), .B(n21064), .Z(n13016) );
  XNOR U22154 ( .A(n[65]), .B(n21065), .Z(n21061) );
  IV U22155 ( .A(n21060), .Z(n21065) );
  XOR U22156 ( .A(n21066), .B(n21067), .Z(n21060) );
  AND U22157 ( .A(n21068), .B(n21069), .Z(n21066) );
  XOR U22158 ( .A(n21067), .B(n13021), .Z(n21069) );
  XNOR U22159 ( .A(n21070), .B(n21071), .Z(n13021) );
  XNOR U22160 ( .A(n[64]), .B(n21072), .Z(n21068) );
  IV U22161 ( .A(n21067), .Z(n21072) );
  XOR U22162 ( .A(n21073), .B(n21074), .Z(n21067) );
  AND U22163 ( .A(n21075), .B(n21076), .Z(n21073) );
  XOR U22164 ( .A(n21074), .B(n13026), .Z(n21076) );
  XNOR U22165 ( .A(n21077), .B(n21078), .Z(n13026) );
  XNOR U22166 ( .A(n[63]), .B(n21079), .Z(n21075) );
  IV U22167 ( .A(n21074), .Z(n21079) );
  XOR U22168 ( .A(n21080), .B(n21081), .Z(n21074) );
  AND U22169 ( .A(n21082), .B(n21083), .Z(n21080) );
  XOR U22170 ( .A(n21081), .B(n13031), .Z(n21083) );
  XNOR U22171 ( .A(n21084), .B(n21085), .Z(n13031) );
  XNOR U22172 ( .A(n[62]), .B(n21086), .Z(n21082) );
  IV U22173 ( .A(n21081), .Z(n21086) );
  XOR U22174 ( .A(n21087), .B(n21088), .Z(n21081) );
  AND U22175 ( .A(n21089), .B(n21090), .Z(n21087) );
  XOR U22176 ( .A(n21088), .B(n13036), .Z(n21090) );
  XNOR U22177 ( .A(n21091), .B(n21092), .Z(n13036) );
  XNOR U22178 ( .A(n[61]), .B(n21093), .Z(n21089) );
  IV U22179 ( .A(n21088), .Z(n21093) );
  XOR U22180 ( .A(n21094), .B(n21095), .Z(n21088) );
  AND U22181 ( .A(n21096), .B(n21097), .Z(n21094) );
  XOR U22182 ( .A(n21095), .B(n13041), .Z(n21097) );
  XNOR U22183 ( .A(n21098), .B(n21099), .Z(n13041) );
  XNOR U22184 ( .A(n[60]), .B(n21100), .Z(n21096) );
  IV U22185 ( .A(n21095), .Z(n21100) );
  XOR U22186 ( .A(n21101), .B(n21102), .Z(n21095) );
  AND U22187 ( .A(n21103), .B(n21104), .Z(n21101) );
  XOR U22188 ( .A(n21102), .B(n13046), .Z(n21104) );
  XNOR U22189 ( .A(n21105), .B(n21106), .Z(n13046) );
  XNOR U22190 ( .A(n[59]), .B(n21107), .Z(n21103) );
  IV U22191 ( .A(n21102), .Z(n21107) );
  XOR U22192 ( .A(n21108), .B(n21109), .Z(n21102) );
  AND U22193 ( .A(n21110), .B(n21111), .Z(n21108) );
  XOR U22194 ( .A(n21109), .B(n13051), .Z(n21111) );
  XNOR U22195 ( .A(n21112), .B(n21113), .Z(n13051) );
  XNOR U22196 ( .A(n[58]), .B(n21114), .Z(n21110) );
  IV U22197 ( .A(n21109), .Z(n21114) );
  XOR U22198 ( .A(n21115), .B(n21116), .Z(n21109) );
  AND U22199 ( .A(n21117), .B(n21118), .Z(n21115) );
  XOR U22200 ( .A(n21116), .B(n13056), .Z(n21118) );
  XNOR U22201 ( .A(n21119), .B(n21120), .Z(n13056) );
  XNOR U22202 ( .A(n[57]), .B(n21121), .Z(n21117) );
  IV U22203 ( .A(n21116), .Z(n21121) );
  XOR U22204 ( .A(n21122), .B(n21123), .Z(n21116) );
  AND U22205 ( .A(n21124), .B(n21125), .Z(n21122) );
  XOR U22206 ( .A(n21123), .B(n13061), .Z(n21125) );
  XNOR U22207 ( .A(n21126), .B(n21127), .Z(n13061) );
  XNOR U22208 ( .A(n[56]), .B(n21128), .Z(n21124) );
  IV U22209 ( .A(n21123), .Z(n21128) );
  XOR U22210 ( .A(n21129), .B(n21130), .Z(n21123) );
  AND U22211 ( .A(n21131), .B(n21132), .Z(n21129) );
  XOR U22212 ( .A(n21130), .B(n13066), .Z(n21132) );
  XNOR U22213 ( .A(n21133), .B(n21134), .Z(n13066) );
  XNOR U22214 ( .A(n[55]), .B(n21135), .Z(n21131) );
  IV U22215 ( .A(n21130), .Z(n21135) );
  XOR U22216 ( .A(n21136), .B(n21137), .Z(n21130) );
  AND U22217 ( .A(n21138), .B(n21139), .Z(n21136) );
  XOR U22218 ( .A(n21137), .B(n13071), .Z(n21139) );
  XNOR U22219 ( .A(n21140), .B(n21141), .Z(n13071) );
  XNOR U22220 ( .A(n[54]), .B(n21142), .Z(n21138) );
  IV U22221 ( .A(n21137), .Z(n21142) );
  XOR U22222 ( .A(n21143), .B(n21144), .Z(n21137) );
  AND U22223 ( .A(n21145), .B(n21146), .Z(n21143) );
  XOR U22224 ( .A(n21144), .B(n13076), .Z(n21146) );
  XNOR U22225 ( .A(n21147), .B(n21148), .Z(n13076) );
  XNOR U22226 ( .A(n[53]), .B(n21149), .Z(n21145) );
  IV U22227 ( .A(n21144), .Z(n21149) );
  XOR U22228 ( .A(n21150), .B(n21151), .Z(n21144) );
  AND U22229 ( .A(n21152), .B(n21153), .Z(n21150) );
  XOR U22230 ( .A(n21151), .B(n13081), .Z(n21153) );
  XNOR U22231 ( .A(n21154), .B(n21155), .Z(n13081) );
  XNOR U22232 ( .A(n[52]), .B(n21156), .Z(n21152) );
  IV U22233 ( .A(n21151), .Z(n21156) );
  XOR U22234 ( .A(n21157), .B(n21158), .Z(n21151) );
  AND U22235 ( .A(n21159), .B(n21160), .Z(n21157) );
  XOR U22236 ( .A(n21158), .B(n13086), .Z(n21160) );
  XNOR U22237 ( .A(n21161), .B(n21162), .Z(n13086) );
  XNOR U22238 ( .A(n[51]), .B(n21163), .Z(n21159) );
  IV U22239 ( .A(n21158), .Z(n21163) );
  XOR U22240 ( .A(n21164), .B(n21165), .Z(n21158) );
  AND U22241 ( .A(n21166), .B(n21167), .Z(n21164) );
  XOR U22242 ( .A(n21165), .B(n13091), .Z(n21167) );
  XNOR U22243 ( .A(n21168), .B(n21169), .Z(n13091) );
  XNOR U22244 ( .A(n[50]), .B(n21170), .Z(n21166) );
  IV U22245 ( .A(n21165), .Z(n21170) );
  XOR U22246 ( .A(n21171), .B(n21172), .Z(n21165) );
  AND U22247 ( .A(n21173), .B(n21174), .Z(n21171) );
  XOR U22248 ( .A(n21172), .B(n13096), .Z(n21174) );
  XNOR U22249 ( .A(n21175), .B(n21176), .Z(n13096) );
  XNOR U22250 ( .A(n[49]), .B(n21177), .Z(n21173) );
  IV U22251 ( .A(n21172), .Z(n21177) );
  XOR U22252 ( .A(n21178), .B(n21179), .Z(n21172) );
  AND U22253 ( .A(n21180), .B(n21181), .Z(n21178) );
  XOR U22254 ( .A(n21179), .B(n13101), .Z(n21181) );
  XNOR U22255 ( .A(n21182), .B(n21183), .Z(n13101) );
  XNOR U22256 ( .A(n[48]), .B(n21184), .Z(n21180) );
  IV U22257 ( .A(n21179), .Z(n21184) );
  XOR U22258 ( .A(n21185), .B(n21186), .Z(n21179) );
  AND U22259 ( .A(n21187), .B(n21188), .Z(n21185) );
  XOR U22260 ( .A(n21186), .B(n13106), .Z(n21188) );
  XNOR U22261 ( .A(n21189), .B(n21190), .Z(n13106) );
  XNOR U22262 ( .A(n[47]), .B(n21191), .Z(n21187) );
  IV U22263 ( .A(n21186), .Z(n21191) );
  XOR U22264 ( .A(n21192), .B(n21193), .Z(n21186) );
  AND U22265 ( .A(n21194), .B(n21195), .Z(n21192) );
  XOR U22266 ( .A(n21193), .B(n13111), .Z(n21195) );
  XNOR U22267 ( .A(n21196), .B(n21197), .Z(n13111) );
  XNOR U22268 ( .A(n[46]), .B(n21198), .Z(n21194) );
  IV U22269 ( .A(n21193), .Z(n21198) );
  XOR U22270 ( .A(n21199), .B(n21200), .Z(n21193) );
  AND U22271 ( .A(n21201), .B(n21202), .Z(n21199) );
  XOR U22272 ( .A(n21200), .B(n13116), .Z(n21202) );
  XNOR U22273 ( .A(n21203), .B(n21204), .Z(n13116) );
  XNOR U22274 ( .A(n[45]), .B(n21205), .Z(n21201) );
  IV U22275 ( .A(n21200), .Z(n21205) );
  XOR U22276 ( .A(n21206), .B(n21207), .Z(n21200) );
  AND U22277 ( .A(n21208), .B(n21209), .Z(n21206) );
  XOR U22278 ( .A(n21207), .B(n13121), .Z(n21209) );
  XNOR U22279 ( .A(n21210), .B(n21211), .Z(n13121) );
  XNOR U22280 ( .A(n[44]), .B(n21212), .Z(n21208) );
  IV U22281 ( .A(n21207), .Z(n21212) );
  XOR U22282 ( .A(n21213), .B(n21214), .Z(n21207) );
  AND U22283 ( .A(n21215), .B(n21216), .Z(n21213) );
  XOR U22284 ( .A(n21214), .B(n13126), .Z(n21216) );
  XNOR U22285 ( .A(n21217), .B(n21218), .Z(n13126) );
  XNOR U22286 ( .A(n[43]), .B(n21219), .Z(n21215) );
  IV U22287 ( .A(n21214), .Z(n21219) );
  XOR U22288 ( .A(n21220), .B(n21221), .Z(n21214) );
  AND U22289 ( .A(n21222), .B(n21223), .Z(n21220) );
  XOR U22290 ( .A(n21221), .B(n13131), .Z(n21223) );
  XNOR U22291 ( .A(n21224), .B(n21225), .Z(n13131) );
  XNOR U22292 ( .A(n[42]), .B(n21226), .Z(n21222) );
  IV U22293 ( .A(n21221), .Z(n21226) );
  XOR U22294 ( .A(n21227), .B(n21228), .Z(n21221) );
  AND U22295 ( .A(n21229), .B(n21230), .Z(n21227) );
  XOR U22296 ( .A(n21228), .B(n13136), .Z(n21230) );
  XNOR U22297 ( .A(n21231), .B(n21232), .Z(n13136) );
  XNOR U22298 ( .A(n[41]), .B(n21233), .Z(n21229) );
  IV U22299 ( .A(n21228), .Z(n21233) );
  XOR U22300 ( .A(n21234), .B(n21235), .Z(n21228) );
  AND U22301 ( .A(n21236), .B(n21237), .Z(n21234) );
  XOR U22302 ( .A(n21235), .B(n13141), .Z(n21237) );
  XNOR U22303 ( .A(n21238), .B(n21239), .Z(n13141) );
  XNOR U22304 ( .A(n[40]), .B(n21240), .Z(n21236) );
  IV U22305 ( .A(n21235), .Z(n21240) );
  XOR U22306 ( .A(n21241), .B(n21242), .Z(n21235) );
  AND U22307 ( .A(n21243), .B(n21244), .Z(n21241) );
  XOR U22308 ( .A(n21242), .B(n13146), .Z(n21244) );
  XNOR U22309 ( .A(n21245), .B(n21246), .Z(n13146) );
  XNOR U22310 ( .A(n[39]), .B(n21247), .Z(n21243) );
  IV U22311 ( .A(n21242), .Z(n21247) );
  XOR U22312 ( .A(n21248), .B(n21249), .Z(n21242) );
  AND U22313 ( .A(n21250), .B(n21251), .Z(n21248) );
  XOR U22314 ( .A(n21249), .B(n13151), .Z(n21251) );
  XNOR U22315 ( .A(n21252), .B(n21253), .Z(n13151) );
  XNOR U22316 ( .A(n[38]), .B(n21254), .Z(n21250) );
  IV U22317 ( .A(n21249), .Z(n21254) );
  XOR U22318 ( .A(n21255), .B(n21256), .Z(n21249) );
  AND U22319 ( .A(n21257), .B(n21258), .Z(n21255) );
  XOR U22320 ( .A(n21256), .B(n13156), .Z(n21258) );
  XNOR U22321 ( .A(n21259), .B(n21260), .Z(n13156) );
  XNOR U22322 ( .A(n[37]), .B(n21261), .Z(n21257) );
  IV U22323 ( .A(n21256), .Z(n21261) );
  XOR U22324 ( .A(n21262), .B(n21263), .Z(n21256) );
  AND U22325 ( .A(n21264), .B(n21265), .Z(n21262) );
  XOR U22326 ( .A(n21263), .B(n13161), .Z(n21265) );
  XNOR U22327 ( .A(n21266), .B(n21267), .Z(n13161) );
  XNOR U22328 ( .A(n[36]), .B(n21268), .Z(n21264) );
  IV U22329 ( .A(n21263), .Z(n21268) );
  XOR U22330 ( .A(n21269), .B(n21270), .Z(n21263) );
  AND U22331 ( .A(n21271), .B(n21272), .Z(n21269) );
  XOR U22332 ( .A(n21270), .B(n13166), .Z(n21272) );
  XNOR U22333 ( .A(n21273), .B(n21274), .Z(n13166) );
  XNOR U22334 ( .A(n[35]), .B(n21275), .Z(n21271) );
  IV U22335 ( .A(n21270), .Z(n21275) );
  XOR U22336 ( .A(n21276), .B(n21277), .Z(n21270) );
  AND U22337 ( .A(n21278), .B(n21279), .Z(n21276) );
  XOR U22338 ( .A(n21277), .B(n13171), .Z(n21279) );
  XNOR U22339 ( .A(n21280), .B(n21281), .Z(n13171) );
  XNOR U22340 ( .A(n[34]), .B(n21282), .Z(n21278) );
  IV U22341 ( .A(n21277), .Z(n21282) );
  XOR U22342 ( .A(n21283), .B(n21284), .Z(n21277) );
  AND U22343 ( .A(n21285), .B(n21286), .Z(n21283) );
  XOR U22344 ( .A(n21284), .B(n13176), .Z(n21286) );
  XNOR U22345 ( .A(n21287), .B(n21288), .Z(n13176) );
  XNOR U22346 ( .A(n[33]), .B(n21289), .Z(n21285) );
  IV U22347 ( .A(n21284), .Z(n21289) );
  XOR U22348 ( .A(n21290), .B(n21291), .Z(n21284) );
  AND U22349 ( .A(n21292), .B(n21293), .Z(n21290) );
  XOR U22350 ( .A(n21291), .B(n13181), .Z(n21293) );
  XNOR U22351 ( .A(n21294), .B(n21295), .Z(n13181) );
  XNOR U22352 ( .A(n[32]), .B(n21296), .Z(n21292) );
  IV U22353 ( .A(n21291), .Z(n21296) );
  XOR U22354 ( .A(n21297), .B(n21298), .Z(n21291) );
  AND U22355 ( .A(n21299), .B(n21300), .Z(n21297) );
  XOR U22356 ( .A(n21298), .B(n13186), .Z(n21300) );
  XNOR U22357 ( .A(n21301), .B(n21302), .Z(n13186) );
  XNOR U22358 ( .A(n[31]), .B(n21303), .Z(n21299) );
  IV U22359 ( .A(n21298), .Z(n21303) );
  XOR U22360 ( .A(n21304), .B(n21305), .Z(n21298) );
  AND U22361 ( .A(n21306), .B(n21307), .Z(n21304) );
  XOR U22362 ( .A(n21305), .B(n13191), .Z(n21307) );
  XNOR U22363 ( .A(n21308), .B(n21309), .Z(n13191) );
  XNOR U22364 ( .A(n[30]), .B(n21310), .Z(n21306) );
  IV U22365 ( .A(n21305), .Z(n21310) );
  XOR U22366 ( .A(n21311), .B(n21312), .Z(n21305) );
  AND U22367 ( .A(n21313), .B(n21314), .Z(n21311) );
  XOR U22368 ( .A(n21312), .B(n13196), .Z(n21314) );
  XNOR U22369 ( .A(n21315), .B(n21316), .Z(n13196) );
  XNOR U22370 ( .A(n[29]), .B(n21317), .Z(n21313) );
  IV U22371 ( .A(n21312), .Z(n21317) );
  XOR U22372 ( .A(n21318), .B(n21319), .Z(n21312) );
  AND U22373 ( .A(n21320), .B(n21321), .Z(n21318) );
  XOR U22374 ( .A(n21319), .B(n13201), .Z(n21321) );
  XNOR U22375 ( .A(n21322), .B(n21323), .Z(n13201) );
  XNOR U22376 ( .A(n[28]), .B(n21324), .Z(n21320) );
  IV U22377 ( .A(n21319), .Z(n21324) );
  XOR U22378 ( .A(n21325), .B(n21326), .Z(n21319) );
  AND U22379 ( .A(n21327), .B(n21328), .Z(n21325) );
  XOR U22380 ( .A(n21326), .B(n13206), .Z(n21328) );
  XNOR U22381 ( .A(n21329), .B(n21330), .Z(n13206) );
  XNOR U22382 ( .A(n[27]), .B(n21331), .Z(n21327) );
  IV U22383 ( .A(n21326), .Z(n21331) );
  XOR U22384 ( .A(n21332), .B(n21333), .Z(n21326) );
  AND U22385 ( .A(n21334), .B(n21335), .Z(n21332) );
  XOR U22386 ( .A(n21333), .B(n13211), .Z(n21335) );
  XNOR U22387 ( .A(n21336), .B(n21337), .Z(n13211) );
  XNOR U22388 ( .A(n[26]), .B(n21338), .Z(n21334) );
  IV U22389 ( .A(n21333), .Z(n21338) );
  XOR U22390 ( .A(n21339), .B(n21340), .Z(n21333) );
  AND U22391 ( .A(n21341), .B(n21342), .Z(n21339) );
  XOR U22392 ( .A(n21340), .B(n13216), .Z(n21342) );
  XNOR U22393 ( .A(n21343), .B(n21344), .Z(n13216) );
  XNOR U22394 ( .A(n[25]), .B(n21345), .Z(n21341) );
  IV U22395 ( .A(n21340), .Z(n21345) );
  XOR U22396 ( .A(n21346), .B(n21347), .Z(n21340) );
  AND U22397 ( .A(n21348), .B(n21349), .Z(n21346) );
  XOR U22398 ( .A(n21347), .B(n13221), .Z(n21349) );
  XNOR U22399 ( .A(n21350), .B(n21351), .Z(n13221) );
  XNOR U22400 ( .A(n[24]), .B(n21352), .Z(n21348) );
  IV U22401 ( .A(n21347), .Z(n21352) );
  XOR U22402 ( .A(n21353), .B(n21354), .Z(n21347) );
  AND U22403 ( .A(n21355), .B(n21356), .Z(n21353) );
  XOR U22404 ( .A(n21354), .B(n13226), .Z(n21356) );
  XNOR U22405 ( .A(n21357), .B(n21358), .Z(n13226) );
  XNOR U22406 ( .A(n[23]), .B(n21359), .Z(n21355) );
  IV U22407 ( .A(n21354), .Z(n21359) );
  XOR U22408 ( .A(n21360), .B(n21361), .Z(n21354) );
  AND U22409 ( .A(n21362), .B(n21363), .Z(n21360) );
  XOR U22410 ( .A(n21361), .B(n13231), .Z(n21363) );
  XNOR U22411 ( .A(n21364), .B(n21365), .Z(n13231) );
  XNOR U22412 ( .A(n[22]), .B(n21366), .Z(n21362) );
  IV U22413 ( .A(n21361), .Z(n21366) );
  XOR U22414 ( .A(n21367), .B(n21368), .Z(n21361) );
  AND U22415 ( .A(n21369), .B(n21370), .Z(n21367) );
  XOR U22416 ( .A(n21368), .B(n13236), .Z(n21370) );
  XNOR U22417 ( .A(n21371), .B(n21372), .Z(n13236) );
  XNOR U22418 ( .A(n[21]), .B(n21373), .Z(n21369) );
  IV U22419 ( .A(n21368), .Z(n21373) );
  XOR U22420 ( .A(n21374), .B(n21375), .Z(n21368) );
  AND U22421 ( .A(n21376), .B(n21377), .Z(n21374) );
  XOR U22422 ( .A(n21375), .B(n13241), .Z(n21377) );
  XNOR U22423 ( .A(n21378), .B(n21379), .Z(n13241) );
  XNOR U22424 ( .A(n[20]), .B(n21380), .Z(n21376) );
  IV U22425 ( .A(n21375), .Z(n21380) );
  XOR U22426 ( .A(n21381), .B(n21382), .Z(n21375) );
  AND U22427 ( .A(n21383), .B(n21384), .Z(n21381) );
  XOR U22428 ( .A(n21382), .B(n13246), .Z(n21384) );
  XNOR U22429 ( .A(n21385), .B(n21386), .Z(n13246) );
  XNOR U22430 ( .A(n[19]), .B(n21387), .Z(n21383) );
  IV U22431 ( .A(n21382), .Z(n21387) );
  XOR U22432 ( .A(n21388), .B(n21389), .Z(n21382) );
  AND U22433 ( .A(n21390), .B(n21391), .Z(n21388) );
  XOR U22434 ( .A(n21389), .B(n13251), .Z(n21391) );
  XNOR U22435 ( .A(n21392), .B(n21393), .Z(n13251) );
  XNOR U22436 ( .A(n[18]), .B(n21394), .Z(n21390) );
  IV U22437 ( .A(n21389), .Z(n21394) );
  XOR U22438 ( .A(n21395), .B(n21396), .Z(n21389) );
  AND U22439 ( .A(n21397), .B(n21398), .Z(n21395) );
  XOR U22440 ( .A(n21396), .B(n13256), .Z(n21398) );
  XNOR U22441 ( .A(n21399), .B(n21400), .Z(n13256) );
  XNOR U22442 ( .A(n[17]), .B(n21401), .Z(n21397) );
  IV U22443 ( .A(n21396), .Z(n21401) );
  XOR U22444 ( .A(n21402), .B(n21403), .Z(n21396) );
  AND U22445 ( .A(n21404), .B(n21405), .Z(n21402) );
  XOR U22446 ( .A(n21403), .B(n13261), .Z(n21405) );
  XNOR U22447 ( .A(n21406), .B(n21407), .Z(n13261) );
  XNOR U22448 ( .A(n[16]), .B(n21408), .Z(n21404) );
  IV U22449 ( .A(n21403), .Z(n21408) );
  XOR U22450 ( .A(n21409), .B(n21410), .Z(n21403) );
  AND U22451 ( .A(n21411), .B(n21412), .Z(n21409) );
  XOR U22452 ( .A(n21410), .B(n13266), .Z(n21412) );
  XNOR U22453 ( .A(n21413), .B(n21414), .Z(n13266) );
  XNOR U22454 ( .A(n[15]), .B(n21415), .Z(n21411) );
  IV U22455 ( .A(n21410), .Z(n21415) );
  XOR U22456 ( .A(n21416), .B(n21417), .Z(n21410) );
  AND U22457 ( .A(n21418), .B(n21419), .Z(n21416) );
  XOR U22458 ( .A(n21417), .B(n13271), .Z(n21419) );
  XNOR U22459 ( .A(n21420), .B(n21421), .Z(n13271) );
  XNOR U22460 ( .A(n[14]), .B(n21422), .Z(n21418) );
  IV U22461 ( .A(n21417), .Z(n21422) );
  XOR U22462 ( .A(n21423), .B(n21424), .Z(n21417) );
  AND U22463 ( .A(n21425), .B(n21426), .Z(n21423) );
  XOR U22464 ( .A(n21424), .B(n13276), .Z(n21426) );
  XNOR U22465 ( .A(n21427), .B(n21428), .Z(n13276) );
  XNOR U22466 ( .A(n[13]), .B(n21429), .Z(n21425) );
  IV U22467 ( .A(n21424), .Z(n21429) );
  XOR U22468 ( .A(n21430), .B(n21431), .Z(n21424) );
  AND U22469 ( .A(n21432), .B(n21433), .Z(n21430) );
  XOR U22470 ( .A(n21431), .B(n13281), .Z(n21433) );
  XNOR U22471 ( .A(n21434), .B(n21435), .Z(n13281) );
  XNOR U22472 ( .A(n[12]), .B(n21436), .Z(n21432) );
  IV U22473 ( .A(n21431), .Z(n21436) );
  XOR U22474 ( .A(n21437), .B(n21438), .Z(n21431) );
  AND U22475 ( .A(n21439), .B(n21440), .Z(n21437) );
  XOR U22476 ( .A(n21438), .B(n13286), .Z(n21440) );
  XNOR U22477 ( .A(n21441), .B(n21442), .Z(n13286) );
  XNOR U22478 ( .A(n[11]), .B(n21443), .Z(n21439) );
  IV U22479 ( .A(n21438), .Z(n21443) );
  XOR U22480 ( .A(n21444), .B(n21445), .Z(n21438) );
  AND U22481 ( .A(n21446), .B(n21447), .Z(n21444) );
  XOR U22482 ( .A(n21445), .B(n13291), .Z(n21447) );
  XNOR U22483 ( .A(n21448), .B(n21449), .Z(n13291) );
  XNOR U22484 ( .A(n[10]), .B(n21450), .Z(n21446) );
  IV U22485 ( .A(n21445), .Z(n21450) );
  XOR U22486 ( .A(n21451), .B(n21452), .Z(n21445) );
  AND U22487 ( .A(n21453), .B(n21454), .Z(n21451) );
  XOR U22488 ( .A(n13296), .B(n21452), .Z(n21454) );
  XNOR U22489 ( .A(n21455), .B(n21456), .Z(n13296) );
  XNOR U22490 ( .A(n[9]), .B(n21457), .Z(n21453) );
  IV U22491 ( .A(n21452), .Z(n21457) );
  XOR U22492 ( .A(n21458), .B(n21459), .Z(n21452) );
  AND U22493 ( .A(n21460), .B(n21461), .Z(n21458) );
  XOR U22494 ( .A(n21459), .B(n13301), .Z(n21461) );
  XNOR U22495 ( .A(n21462), .B(n21463), .Z(n13301) );
  XNOR U22496 ( .A(n[8]), .B(n21464), .Z(n21460) );
  IV U22497 ( .A(n21459), .Z(n21464) );
  XOR U22498 ( .A(n21465), .B(n21466), .Z(n21459) );
  AND U22499 ( .A(n21467), .B(n21468), .Z(n21465) );
  XOR U22500 ( .A(n21466), .B(n13306), .Z(n21468) );
  XNOR U22501 ( .A(n21469), .B(n21470), .Z(n13306) );
  XNOR U22502 ( .A(n[7]), .B(n21471), .Z(n21467) );
  IV U22503 ( .A(n21466), .Z(n21471) );
  XOR U22504 ( .A(n21472), .B(n21473), .Z(n21466) );
  AND U22505 ( .A(n21474), .B(n21475), .Z(n21472) );
  XOR U22506 ( .A(n21473), .B(n13311), .Z(n21475) );
  XNOR U22507 ( .A(n21476), .B(n21477), .Z(n13311) );
  XNOR U22508 ( .A(n[6]), .B(n21478), .Z(n21474) );
  IV U22509 ( .A(n21473), .Z(n21478) );
  XOR U22510 ( .A(n21479), .B(n21480), .Z(n21473) );
  AND U22511 ( .A(n21481), .B(n21482), .Z(n21479) );
  XOR U22512 ( .A(n21480), .B(n13316), .Z(n21482) );
  XNOR U22513 ( .A(n21483), .B(n21484), .Z(n13316) );
  XNOR U22514 ( .A(n[5]), .B(n21485), .Z(n21481) );
  IV U22515 ( .A(n21480), .Z(n21485) );
  XOR U22516 ( .A(n21486), .B(n21487), .Z(n21480) );
  AND U22517 ( .A(n21488), .B(n21489), .Z(n21486) );
  XOR U22518 ( .A(n21487), .B(n13321), .Z(n21489) );
  XNOR U22519 ( .A(n21490), .B(n21491), .Z(n13321) );
  XNOR U22520 ( .A(n[4]), .B(n21492), .Z(n21488) );
  IV U22521 ( .A(n21487), .Z(n21492) );
  XOR U22522 ( .A(n21493), .B(n21494), .Z(n21487) );
  AND U22523 ( .A(n21495), .B(n21496), .Z(n21493) );
  XOR U22524 ( .A(n21494), .B(n13326), .Z(n21496) );
  XNOR U22525 ( .A(n21497), .B(n21498), .Z(n13326) );
  XNOR U22526 ( .A(n[3]), .B(n21499), .Z(n21495) );
  IV U22527 ( .A(n21494), .Z(n21499) );
  XOR U22528 ( .A(n21500), .B(n21501), .Z(n21494) );
  AND U22529 ( .A(n21502), .B(n21503), .Z(n21500) );
  XOR U22530 ( .A(n21501), .B(n13331), .Z(n21503) );
  XNOR U22531 ( .A(n21504), .B(n21505), .Z(n13331) );
  XOR U22532 ( .A(n[2]), .B(n21501), .Z(n21502) );
  XOR U22533 ( .A(n21506), .B(n21507), .Z(n21501) );
  NAND U22534 ( .A(n21508), .B(n21509), .Z(n21507) );
  XOR U22535 ( .A(n21506), .B(n13337), .Z(n21509) );
  XNOR U22536 ( .A(n21510), .B(n21511), .Z(n13337) );
  XNOR U22537 ( .A(n[1]), .B(n21506), .Z(n21508) );
  NOR U22538 ( .A(n[0]), .B(n13339), .Z(n21506) );
  XNOR U22539 ( .A(n21512), .B(n21513), .Z(n13339) );
  IV U22540 ( .A(n21514), .Z(n21513) );
  XNOR U22541 ( .A(n21515), .B(n21516), .Z(n14346) );
  ANDN U22542 ( .B(n21517), .A(n1038), .Z(n21515) );
  XOR U22543 ( .A(n21518), .B(n21517), .Z(n1038) );
  IV U22544 ( .A(n14348), .Z(n21517) );
  XNOR U22545 ( .A(n21519), .B(n21520), .Z(n14348) );
  AND U22546 ( .A(n14358), .B(n21521), .Z(n21519) );
  XNOR U22547 ( .A(n14357), .B(n21520), .Z(n21521) );
  NAND U22548 ( .A(n21522), .B(n[1023]), .Z(n14357) );
  NAND U22549 ( .A(n21523), .B(n[1023]), .Z(n21522) );
  XNOR U22550 ( .A(n21524), .B(n21520), .Z(n14358) );
  XOR U22551 ( .A(n21525), .B(n21526), .Z(n21520) );
  AND U22552 ( .A(n14365), .B(n21527), .Z(n21525) );
  XNOR U22553 ( .A(n14364), .B(n21526), .Z(n21527) );
  NAND U22554 ( .A(n21528), .B(n[1022]), .Z(n14364) );
  NAND U22555 ( .A(n21523), .B(n[1022]), .Z(n21528) );
  XNOR U22556 ( .A(n21529), .B(n21526), .Z(n14365) );
  XOR U22557 ( .A(n21530), .B(n21531), .Z(n21526) );
  AND U22558 ( .A(n14372), .B(n21532), .Z(n21530) );
  XNOR U22559 ( .A(n14371), .B(n21531), .Z(n21532) );
  NAND U22560 ( .A(n21533), .B(n[1021]), .Z(n14371) );
  NAND U22561 ( .A(n21523), .B(n[1021]), .Z(n21533) );
  XNOR U22562 ( .A(n21534), .B(n21531), .Z(n14372) );
  XOR U22563 ( .A(n21535), .B(n21536), .Z(n21531) );
  AND U22564 ( .A(n14379), .B(n21537), .Z(n21535) );
  XNOR U22565 ( .A(n14378), .B(n21536), .Z(n21537) );
  NAND U22566 ( .A(n21538), .B(n[1020]), .Z(n14378) );
  NAND U22567 ( .A(n21523), .B(n[1020]), .Z(n21538) );
  XNOR U22568 ( .A(n21539), .B(n21536), .Z(n14379) );
  XOR U22569 ( .A(n21540), .B(n21541), .Z(n21536) );
  AND U22570 ( .A(n14386), .B(n21542), .Z(n21540) );
  XNOR U22571 ( .A(n14385), .B(n21541), .Z(n21542) );
  NAND U22572 ( .A(n21543), .B(n[1019]), .Z(n14385) );
  NAND U22573 ( .A(n21523), .B(n[1019]), .Z(n21543) );
  XNOR U22574 ( .A(n21544), .B(n21541), .Z(n14386) );
  XOR U22575 ( .A(n21545), .B(n21546), .Z(n21541) );
  AND U22576 ( .A(n14393), .B(n21547), .Z(n21545) );
  XNOR U22577 ( .A(n14392), .B(n21546), .Z(n21547) );
  NAND U22578 ( .A(n21548), .B(n[1018]), .Z(n14392) );
  NAND U22579 ( .A(n21523), .B(n[1018]), .Z(n21548) );
  XNOR U22580 ( .A(n21549), .B(n21546), .Z(n14393) );
  XOR U22581 ( .A(n21550), .B(n21551), .Z(n21546) );
  AND U22582 ( .A(n14400), .B(n21552), .Z(n21550) );
  XNOR U22583 ( .A(n14399), .B(n21551), .Z(n21552) );
  NAND U22584 ( .A(n21553), .B(n[1017]), .Z(n14399) );
  NAND U22585 ( .A(n21523), .B(n[1017]), .Z(n21553) );
  XNOR U22586 ( .A(n21554), .B(n21551), .Z(n14400) );
  XOR U22587 ( .A(n21555), .B(n21556), .Z(n21551) );
  AND U22588 ( .A(n14407), .B(n21557), .Z(n21555) );
  XNOR U22589 ( .A(n14406), .B(n21556), .Z(n21557) );
  NAND U22590 ( .A(n21558), .B(n[1016]), .Z(n14406) );
  NAND U22591 ( .A(n21523), .B(n[1016]), .Z(n21558) );
  XNOR U22592 ( .A(n21559), .B(n21556), .Z(n14407) );
  XOR U22593 ( .A(n21560), .B(n21561), .Z(n21556) );
  AND U22594 ( .A(n14414), .B(n21562), .Z(n21560) );
  XNOR U22595 ( .A(n14413), .B(n21561), .Z(n21562) );
  NAND U22596 ( .A(n21563), .B(n[1015]), .Z(n14413) );
  NAND U22597 ( .A(n21523), .B(n[1015]), .Z(n21563) );
  XNOR U22598 ( .A(n21564), .B(n21561), .Z(n14414) );
  XOR U22599 ( .A(n21565), .B(n21566), .Z(n21561) );
  AND U22600 ( .A(n14421), .B(n21567), .Z(n21565) );
  XNOR U22601 ( .A(n14420), .B(n21566), .Z(n21567) );
  NAND U22602 ( .A(n21568), .B(n[1014]), .Z(n14420) );
  NAND U22603 ( .A(n21523), .B(n[1014]), .Z(n21568) );
  XNOR U22604 ( .A(n21569), .B(n21566), .Z(n14421) );
  XOR U22605 ( .A(n21570), .B(n21571), .Z(n21566) );
  AND U22606 ( .A(n14428), .B(n21572), .Z(n21570) );
  XNOR U22607 ( .A(n14427), .B(n21571), .Z(n21572) );
  NAND U22608 ( .A(n21573), .B(n[1013]), .Z(n14427) );
  NAND U22609 ( .A(n21523), .B(n[1013]), .Z(n21573) );
  XNOR U22610 ( .A(n21574), .B(n21571), .Z(n14428) );
  XOR U22611 ( .A(n21575), .B(n21576), .Z(n21571) );
  AND U22612 ( .A(n14435), .B(n21577), .Z(n21575) );
  XNOR U22613 ( .A(n14434), .B(n21576), .Z(n21577) );
  NAND U22614 ( .A(n21578), .B(n[1012]), .Z(n14434) );
  NAND U22615 ( .A(n21523), .B(n[1012]), .Z(n21578) );
  XNOR U22616 ( .A(n21579), .B(n21576), .Z(n14435) );
  XOR U22617 ( .A(n21580), .B(n21581), .Z(n21576) );
  AND U22618 ( .A(n14442), .B(n21582), .Z(n21580) );
  XNOR U22619 ( .A(n14441), .B(n21581), .Z(n21582) );
  NAND U22620 ( .A(n21583), .B(n[1011]), .Z(n14441) );
  NAND U22621 ( .A(n21523), .B(n[1011]), .Z(n21583) );
  XNOR U22622 ( .A(n21584), .B(n21581), .Z(n14442) );
  XOR U22623 ( .A(n21585), .B(n21586), .Z(n21581) );
  AND U22624 ( .A(n14449), .B(n21587), .Z(n21585) );
  XNOR U22625 ( .A(n14448), .B(n21586), .Z(n21587) );
  NAND U22626 ( .A(n21588), .B(n[1010]), .Z(n14448) );
  NAND U22627 ( .A(n21523), .B(n[1010]), .Z(n21588) );
  XNOR U22628 ( .A(n21589), .B(n21586), .Z(n14449) );
  XOR U22629 ( .A(n21590), .B(n21591), .Z(n21586) );
  AND U22630 ( .A(n14456), .B(n21592), .Z(n21590) );
  XNOR U22631 ( .A(n14455), .B(n21591), .Z(n21592) );
  NAND U22632 ( .A(n21593), .B(n[1009]), .Z(n14455) );
  NAND U22633 ( .A(n21523), .B(n[1009]), .Z(n21593) );
  XNOR U22634 ( .A(n21594), .B(n21591), .Z(n14456) );
  XOR U22635 ( .A(n21595), .B(n21596), .Z(n21591) );
  AND U22636 ( .A(n14463), .B(n21597), .Z(n21595) );
  XNOR U22637 ( .A(n14462), .B(n21596), .Z(n21597) );
  NAND U22638 ( .A(n21598), .B(n[1008]), .Z(n14462) );
  NAND U22639 ( .A(n21523), .B(n[1008]), .Z(n21598) );
  XNOR U22640 ( .A(n21599), .B(n21596), .Z(n14463) );
  XOR U22641 ( .A(n21600), .B(n21601), .Z(n21596) );
  AND U22642 ( .A(n14470), .B(n21602), .Z(n21600) );
  XNOR U22643 ( .A(n14469), .B(n21601), .Z(n21602) );
  NAND U22644 ( .A(n21603), .B(n[1007]), .Z(n14469) );
  NAND U22645 ( .A(n21523), .B(n[1007]), .Z(n21603) );
  XNOR U22646 ( .A(n21604), .B(n21601), .Z(n14470) );
  XOR U22647 ( .A(n21605), .B(n21606), .Z(n21601) );
  AND U22648 ( .A(n14477), .B(n21607), .Z(n21605) );
  XNOR U22649 ( .A(n14476), .B(n21606), .Z(n21607) );
  NAND U22650 ( .A(n21608), .B(n[1006]), .Z(n14476) );
  NAND U22651 ( .A(n21523), .B(n[1006]), .Z(n21608) );
  XNOR U22652 ( .A(n21609), .B(n21606), .Z(n14477) );
  XOR U22653 ( .A(n21610), .B(n21611), .Z(n21606) );
  AND U22654 ( .A(n14484), .B(n21612), .Z(n21610) );
  XNOR U22655 ( .A(n14483), .B(n21611), .Z(n21612) );
  NAND U22656 ( .A(n21613), .B(n[1005]), .Z(n14483) );
  NAND U22657 ( .A(n21523), .B(n[1005]), .Z(n21613) );
  XNOR U22658 ( .A(n21614), .B(n21611), .Z(n14484) );
  XOR U22659 ( .A(n21615), .B(n21616), .Z(n21611) );
  AND U22660 ( .A(n14491), .B(n21617), .Z(n21615) );
  XNOR U22661 ( .A(n14490), .B(n21616), .Z(n21617) );
  NAND U22662 ( .A(n21618), .B(n[1004]), .Z(n14490) );
  NAND U22663 ( .A(n21523), .B(n[1004]), .Z(n21618) );
  XNOR U22664 ( .A(n21619), .B(n21616), .Z(n14491) );
  XOR U22665 ( .A(n21620), .B(n21621), .Z(n21616) );
  AND U22666 ( .A(n14498), .B(n21622), .Z(n21620) );
  XNOR U22667 ( .A(n14497), .B(n21621), .Z(n21622) );
  NAND U22668 ( .A(n21623), .B(n[1003]), .Z(n14497) );
  NAND U22669 ( .A(n21523), .B(n[1003]), .Z(n21623) );
  XNOR U22670 ( .A(n21624), .B(n21621), .Z(n14498) );
  XOR U22671 ( .A(n21625), .B(n21626), .Z(n21621) );
  AND U22672 ( .A(n14505), .B(n21627), .Z(n21625) );
  XNOR U22673 ( .A(n14504), .B(n21626), .Z(n21627) );
  NAND U22674 ( .A(n21628), .B(n[1002]), .Z(n14504) );
  NAND U22675 ( .A(n21523), .B(n[1002]), .Z(n21628) );
  XNOR U22676 ( .A(n21629), .B(n21626), .Z(n14505) );
  XOR U22677 ( .A(n21630), .B(n21631), .Z(n21626) );
  AND U22678 ( .A(n14512), .B(n21632), .Z(n21630) );
  XNOR U22679 ( .A(n14511), .B(n21631), .Z(n21632) );
  NAND U22680 ( .A(n21633), .B(n[1001]), .Z(n14511) );
  NAND U22681 ( .A(n21523), .B(n[1001]), .Z(n21633) );
  XNOR U22682 ( .A(n21634), .B(n21631), .Z(n14512) );
  XOR U22683 ( .A(n21635), .B(n21636), .Z(n21631) );
  AND U22684 ( .A(n14519), .B(n21637), .Z(n21635) );
  XNOR U22685 ( .A(n14518), .B(n21636), .Z(n21637) );
  NAND U22686 ( .A(n21638), .B(n[1000]), .Z(n14518) );
  NAND U22687 ( .A(n21523), .B(n[1000]), .Z(n21638) );
  XNOR U22688 ( .A(n21639), .B(n21636), .Z(n14519) );
  XOR U22689 ( .A(n21640), .B(n21641), .Z(n21636) );
  AND U22690 ( .A(n14526), .B(n21642), .Z(n21640) );
  XNOR U22691 ( .A(n14525), .B(n21641), .Z(n21642) );
  NAND U22692 ( .A(n21643), .B(n[999]), .Z(n14525) );
  NAND U22693 ( .A(n21523), .B(n[999]), .Z(n21643) );
  XNOR U22694 ( .A(n21644), .B(n21641), .Z(n14526) );
  XOR U22695 ( .A(n21645), .B(n21646), .Z(n21641) );
  AND U22696 ( .A(n14533), .B(n21647), .Z(n21645) );
  XNOR U22697 ( .A(n14532), .B(n21646), .Z(n21647) );
  NAND U22698 ( .A(n21648), .B(n[998]), .Z(n14532) );
  NAND U22699 ( .A(n21523), .B(n[998]), .Z(n21648) );
  XNOR U22700 ( .A(n21649), .B(n21646), .Z(n14533) );
  XOR U22701 ( .A(n21650), .B(n21651), .Z(n21646) );
  AND U22702 ( .A(n14540), .B(n21652), .Z(n21650) );
  XNOR U22703 ( .A(n14539), .B(n21651), .Z(n21652) );
  NAND U22704 ( .A(n21653), .B(n[997]), .Z(n14539) );
  NAND U22705 ( .A(n21523), .B(n[997]), .Z(n21653) );
  XNOR U22706 ( .A(n21654), .B(n21651), .Z(n14540) );
  XOR U22707 ( .A(n21655), .B(n21656), .Z(n21651) );
  AND U22708 ( .A(n14547), .B(n21657), .Z(n21655) );
  XNOR U22709 ( .A(n14546), .B(n21656), .Z(n21657) );
  NAND U22710 ( .A(n21658), .B(n[996]), .Z(n14546) );
  NAND U22711 ( .A(n21523), .B(n[996]), .Z(n21658) );
  XNOR U22712 ( .A(n21659), .B(n21656), .Z(n14547) );
  XOR U22713 ( .A(n21660), .B(n21661), .Z(n21656) );
  AND U22714 ( .A(n14554), .B(n21662), .Z(n21660) );
  XNOR U22715 ( .A(n14553), .B(n21661), .Z(n21662) );
  NAND U22716 ( .A(n21663), .B(n[995]), .Z(n14553) );
  NAND U22717 ( .A(n21523), .B(n[995]), .Z(n21663) );
  XNOR U22718 ( .A(n21664), .B(n21661), .Z(n14554) );
  XOR U22719 ( .A(n21665), .B(n21666), .Z(n21661) );
  AND U22720 ( .A(n14561), .B(n21667), .Z(n21665) );
  XNOR U22721 ( .A(n14560), .B(n21666), .Z(n21667) );
  NAND U22722 ( .A(n21668), .B(n[994]), .Z(n14560) );
  NAND U22723 ( .A(n21523), .B(n[994]), .Z(n21668) );
  XNOR U22724 ( .A(n21669), .B(n21666), .Z(n14561) );
  XOR U22725 ( .A(n21670), .B(n21671), .Z(n21666) );
  AND U22726 ( .A(n14568), .B(n21672), .Z(n21670) );
  XNOR U22727 ( .A(n14567), .B(n21671), .Z(n21672) );
  NAND U22728 ( .A(n21673), .B(n[993]), .Z(n14567) );
  NAND U22729 ( .A(n21523), .B(n[993]), .Z(n21673) );
  XNOR U22730 ( .A(n21674), .B(n21671), .Z(n14568) );
  XOR U22731 ( .A(n21675), .B(n21676), .Z(n21671) );
  AND U22732 ( .A(n14575), .B(n21677), .Z(n21675) );
  XNOR U22733 ( .A(n14574), .B(n21676), .Z(n21677) );
  NAND U22734 ( .A(n21678), .B(n[992]), .Z(n14574) );
  NAND U22735 ( .A(n21523), .B(n[992]), .Z(n21678) );
  XNOR U22736 ( .A(n21679), .B(n21676), .Z(n14575) );
  XOR U22737 ( .A(n21680), .B(n21681), .Z(n21676) );
  AND U22738 ( .A(n14582), .B(n21682), .Z(n21680) );
  XNOR U22739 ( .A(n14581), .B(n21681), .Z(n21682) );
  NAND U22740 ( .A(n21683), .B(n[991]), .Z(n14581) );
  NAND U22741 ( .A(n21523), .B(n[991]), .Z(n21683) );
  XNOR U22742 ( .A(n21684), .B(n21681), .Z(n14582) );
  XOR U22743 ( .A(n21685), .B(n21686), .Z(n21681) );
  AND U22744 ( .A(n14589), .B(n21687), .Z(n21685) );
  XNOR U22745 ( .A(n14588), .B(n21686), .Z(n21687) );
  NAND U22746 ( .A(n21688), .B(n[990]), .Z(n14588) );
  NAND U22747 ( .A(n21523), .B(n[990]), .Z(n21688) );
  XNOR U22748 ( .A(n21689), .B(n21686), .Z(n14589) );
  XOR U22749 ( .A(n21690), .B(n21691), .Z(n21686) );
  AND U22750 ( .A(n14596), .B(n21692), .Z(n21690) );
  XNOR U22751 ( .A(n14595), .B(n21691), .Z(n21692) );
  NAND U22752 ( .A(n21693), .B(n[989]), .Z(n14595) );
  NAND U22753 ( .A(n21523), .B(n[989]), .Z(n21693) );
  XNOR U22754 ( .A(n21694), .B(n21691), .Z(n14596) );
  XOR U22755 ( .A(n21695), .B(n21696), .Z(n21691) );
  AND U22756 ( .A(n14603), .B(n21697), .Z(n21695) );
  XNOR U22757 ( .A(n14602), .B(n21696), .Z(n21697) );
  NAND U22758 ( .A(n21698), .B(n[988]), .Z(n14602) );
  NAND U22759 ( .A(n21523), .B(n[988]), .Z(n21698) );
  XNOR U22760 ( .A(n21699), .B(n21696), .Z(n14603) );
  XOR U22761 ( .A(n21700), .B(n21701), .Z(n21696) );
  AND U22762 ( .A(n14610), .B(n21702), .Z(n21700) );
  XNOR U22763 ( .A(n14609), .B(n21701), .Z(n21702) );
  NAND U22764 ( .A(n21703), .B(n[987]), .Z(n14609) );
  NAND U22765 ( .A(n21523), .B(n[987]), .Z(n21703) );
  XNOR U22766 ( .A(n21704), .B(n21701), .Z(n14610) );
  XOR U22767 ( .A(n21705), .B(n21706), .Z(n21701) );
  AND U22768 ( .A(n14617), .B(n21707), .Z(n21705) );
  XNOR U22769 ( .A(n14616), .B(n21706), .Z(n21707) );
  NAND U22770 ( .A(n21708), .B(n[986]), .Z(n14616) );
  NAND U22771 ( .A(n21523), .B(n[986]), .Z(n21708) );
  XNOR U22772 ( .A(n21709), .B(n21706), .Z(n14617) );
  XOR U22773 ( .A(n21710), .B(n21711), .Z(n21706) );
  AND U22774 ( .A(n14624), .B(n21712), .Z(n21710) );
  XNOR U22775 ( .A(n14623), .B(n21711), .Z(n21712) );
  NAND U22776 ( .A(n21713), .B(n[985]), .Z(n14623) );
  NAND U22777 ( .A(n21523), .B(n[985]), .Z(n21713) );
  XNOR U22778 ( .A(n21714), .B(n21711), .Z(n14624) );
  XOR U22779 ( .A(n21715), .B(n21716), .Z(n21711) );
  AND U22780 ( .A(n14631), .B(n21717), .Z(n21715) );
  XNOR U22781 ( .A(n14630), .B(n21716), .Z(n21717) );
  NAND U22782 ( .A(n21718), .B(n[984]), .Z(n14630) );
  NAND U22783 ( .A(n21523), .B(n[984]), .Z(n21718) );
  XNOR U22784 ( .A(n21719), .B(n21716), .Z(n14631) );
  XOR U22785 ( .A(n21720), .B(n21721), .Z(n21716) );
  AND U22786 ( .A(n14638), .B(n21722), .Z(n21720) );
  XNOR U22787 ( .A(n14637), .B(n21721), .Z(n21722) );
  NAND U22788 ( .A(n21723), .B(n[983]), .Z(n14637) );
  NAND U22789 ( .A(n21523), .B(n[983]), .Z(n21723) );
  XNOR U22790 ( .A(n21724), .B(n21721), .Z(n14638) );
  XOR U22791 ( .A(n21725), .B(n21726), .Z(n21721) );
  AND U22792 ( .A(n14645), .B(n21727), .Z(n21725) );
  XNOR U22793 ( .A(n14644), .B(n21726), .Z(n21727) );
  NAND U22794 ( .A(n21728), .B(n[982]), .Z(n14644) );
  NAND U22795 ( .A(n21523), .B(n[982]), .Z(n21728) );
  XNOR U22796 ( .A(n21729), .B(n21726), .Z(n14645) );
  XOR U22797 ( .A(n21730), .B(n21731), .Z(n21726) );
  AND U22798 ( .A(n14652), .B(n21732), .Z(n21730) );
  XNOR U22799 ( .A(n14651), .B(n21731), .Z(n21732) );
  NAND U22800 ( .A(n21733), .B(n[981]), .Z(n14651) );
  NAND U22801 ( .A(n21523), .B(n[981]), .Z(n21733) );
  XNOR U22802 ( .A(n21734), .B(n21731), .Z(n14652) );
  XOR U22803 ( .A(n21735), .B(n21736), .Z(n21731) );
  AND U22804 ( .A(n14659), .B(n21737), .Z(n21735) );
  XNOR U22805 ( .A(n14658), .B(n21736), .Z(n21737) );
  NAND U22806 ( .A(n21738), .B(n[980]), .Z(n14658) );
  NAND U22807 ( .A(n21523), .B(n[980]), .Z(n21738) );
  XNOR U22808 ( .A(n21739), .B(n21736), .Z(n14659) );
  XOR U22809 ( .A(n21740), .B(n21741), .Z(n21736) );
  AND U22810 ( .A(n14666), .B(n21742), .Z(n21740) );
  XNOR U22811 ( .A(n14665), .B(n21741), .Z(n21742) );
  NAND U22812 ( .A(n21743), .B(n[979]), .Z(n14665) );
  NAND U22813 ( .A(n21523), .B(n[979]), .Z(n21743) );
  XNOR U22814 ( .A(n21744), .B(n21741), .Z(n14666) );
  XOR U22815 ( .A(n21745), .B(n21746), .Z(n21741) );
  AND U22816 ( .A(n14673), .B(n21747), .Z(n21745) );
  XNOR U22817 ( .A(n14672), .B(n21746), .Z(n21747) );
  NAND U22818 ( .A(n21748), .B(n[978]), .Z(n14672) );
  NAND U22819 ( .A(n21523), .B(n[978]), .Z(n21748) );
  XNOR U22820 ( .A(n21749), .B(n21746), .Z(n14673) );
  XOR U22821 ( .A(n21750), .B(n21751), .Z(n21746) );
  AND U22822 ( .A(n14680), .B(n21752), .Z(n21750) );
  XNOR U22823 ( .A(n14679), .B(n21751), .Z(n21752) );
  NAND U22824 ( .A(n21753), .B(n[977]), .Z(n14679) );
  NAND U22825 ( .A(n21523), .B(n[977]), .Z(n21753) );
  XNOR U22826 ( .A(n21754), .B(n21751), .Z(n14680) );
  XOR U22827 ( .A(n21755), .B(n21756), .Z(n21751) );
  AND U22828 ( .A(n14687), .B(n21757), .Z(n21755) );
  XNOR U22829 ( .A(n14686), .B(n21756), .Z(n21757) );
  NAND U22830 ( .A(n21758), .B(n[976]), .Z(n14686) );
  NAND U22831 ( .A(n21523), .B(n[976]), .Z(n21758) );
  XNOR U22832 ( .A(n21759), .B(n21756), .Z(n14687) );
  XOR U22833 ( .A(n21760), .B(n21761), .Z(n21756) );
  AND U22834 ( .A(n14694), .B(n21762), .Z(n21760) );
  XNOR U22835 ( .A(n14693), .B(n21761), .Z(n21762) );
  NAND U22836 ( .A(n21763), .B(n[975]), .Z(n14693) );
  NAND U22837 ( .A(n21523), .B(n[975]), .Z(n21763) );
  XNOR U22838 ( .A(n21764), .B(n21761), .Z(n14694) );
  XOR U22839 ( .A(n21765), .B(n21766), .Z(n21761) );
  AND U22840 ( .A(n14701), .B(n21767), .Z(n21765) );
  XNOR U22841 ( .A(n14700), .B(n21766), .Z(n21767) );
  NAND U22842 ( .A(n21768), .B(n[974]), .Z(n14700) );
  NAND U22843 ( .A(n21523), .B(n[974]), .Z(n21768) );
  XNOR U22844 ( .A(n21769), .B(n21766), .Z(n14701) );
  XOR U22845 ( .A(n21770), .B(n21771), .Z(n21766) );
  AND U22846 ( .A(n14708), .B(n21772), .Z(n21770) );
  XNOR U22847 ( .A(n14707), .B(n21771), .Z(n21772) );
  NAND U22848 ( .A(n21773), .B(n[973]), .Z(n14707) );
  NAND U22849 ( .A(n21523), .B(n[973]), .Z(n21773) );
  XNOR U22850 ( .A(n21774), .B(n21771), .Z(n14708) );
  XOR U22851 ( .A(n21775), .B(n21776), .Z(n21771) );
  AND U22852 ( .A(n14715), .B(n21777), .Z(n21775) );
  XNOR U22853 ( .A(n14714), .B(n21776), .Z(n21777) );
  NAND U22854 ( .A(n21778), .B(n[972]), .Z(n14714) );
  NAND U22855 ( .A(n21523), .B(n[972]), .Z(n21778) );
  XNOR U22856 ( .A(n21779), .B(n21776), .Z(n14715) );
  XOR U22857 ( .A(n21780), .B(n21781), .Z(n21776) );
  AND U22858 ( .A(n14722), .B(n21782), .Z(n21780) );
  XNOR U22859 ( .A(n14721), .B(n21781), .Z(n21782) );
  NAND U22860 ( .A(n21783), .B(n[971]), .Z(n14721) );
  NAND U22861 ( .A(n21523), .B(n[971]), .Z(n21783) );
  XNOR U22862 ( .A(n21784), .B(n21781), .Z(n14722) );
  XOR U22863 ( .A(n21785), .B(n21786), .Z(n21781) );
  AND U22864 ( .A(n14729), .B(n21787), .Z(n21785) );
  XNOR U22865 ( .A(n14728), .B(n21786), .Z(n21787) );
  NAND U22866 ( .A(n21788), .B(n[970]), .Z(n14728) );
  NAND U22867 ( .A(n21523), .B(n[970]), .Z(n21788) );
  XNOR U22868 ( .A(n21789), .B(n21786), .Z(n14729) );
  XOR U22869 ( .A(n21790), .B(n21791), .Z(n21786) );
  AND U22870 ( .A(n14736), .B(n21792), .Z(n21790) );
  XNOR U22871 ( .A(n14735), .B(n21791), .Z(n21792) );
  NAND U22872 ( .A(n21793), .B(n[969]), .Z(n14735) );
  NAND U22873 ( .A(n21523), .B(n[969]), .Z(n21793) );
  XNOR U22874 ( .A(n21794), .B(n21791), .Z(n14736) );
  XOR U22875 ( .A(n21795), .B(n21796), .Z(n21791) );
  AND U22876 ( .A(n14743), .B(n21797), .Z(n21795) );
  XNOR U22877 ( .A(n14742), .B(n21796), .Z(n21797) );
  NAND U22878 ( .A(n21798), .B(n[968]), .Z(n14742) );
  NAND U22879 ( .A(n21523), .B(n[968]), .Z(n21798) );
  XNOR U22880 ( .A(n21799), .B(n21796), .Z(n14743) );
  XOR U22881 ( .A(n21800), .B(n21801), .Z(n21796) );
  AND U22882 ( .A(n14750), .B(n21802), .Z(n21800) );
  XNOR U22883 ( .A(n14749), .B(n21801), .Z(n21802) );
  NAND U22884 ( .A(n21803), .B(n[967]), .Z(n14749) );
  NAND U22885 ( .A(n21523), .B(n[967]), .Z(n21803) );
  XNOR U22886 ( .A(n21804), .B(n21801), .Z(n14750) );
  XOR U22887 ( .A(n21805), .B(n21806), .Z(n21801) );
  AND U22888 ( .A(n14757), .B(n21807), .Z(n21805) );
  XNOR U22889 ( .A(n14756), .B(n21806), .Z(n21807) );
  NAND U22890 ( .A(n21808), .B(n[966]), .Z(n14756) );
  NAND U22891 ( .A(n21523), .B(n[966]), .Z(n21808) );
  XNOR U22892 ( .A(n21809), .B(n21806), .Z(n14757) );
  XOR U22893 ( .A(n21810), .B(n21811), .Z(n21806) );
  AND U22894 ( .A(n14764), .B(n21812), .Z(n21810) );
  XNOR U22895 ( .A(n14763), .B(n21811), .Z(n21812) );
  NAND U22896 ( .A(n21813), .B(n[965]), .Z(n14763) );
  NAND U22897 ( .A(n21523), .B(n[965]), .Z(n21813) );
  XNOR U22898 ( .A(n21814), .B(n21811), .Z(n14764) );
  XOR U22899 ( .A(n21815), .B(n21816), .Z(n21811) );
  AND U22900 ( .A(n14771), .B(n21817), .Z(n21815) );
  XNOR U22901 ( .A(n14770), .B(n21816), .Z(n21817) );
  NAND U22902 ( .A(n21818), .B(n[964]), .Z(n14770) );
  NAND U22903 ( .A(n21523), .B(n[964]), .Z(n21818) );
  XNOR U22904 ( .A(n21819), .B(n21816), .Z(n14771) );
  XOR U22905 ( .A(n21820), .B(n21821), .Z(n21816) );
  AND U22906 ( .A(n14778), .B(n21822), .Z(n21820) );
  XNOR U22907 ( .A(n14777), .B(n21821), .Z(n21822) );
  NAND U22908 ( .A(n21823), .B(n[963]), .Z(n14777) );
  NAND U22909 ( .A(n21523), .B(n[963]), .Z(n21823) );
  XNOR U22910 ( .A(n21824), .B(n21821), .Z(n14778) );
  XOR U22911 ( .A(n21825), .B(n21826), .Z(n21821) );
  AND U22912 ( .A(n14785), .B(n21827), .Z(n21825) );
  XNOR U22913 ( .A(n14784), .B(n21826), .Z(n21827) );
  NAND U22914 ( .A(n21828), .B(n[962]), .Z(n14784) );
  NAND U22915 ( .A(n21523), .B(n[962]), .Z(n21828) );
  XNOR U22916 ( .A(n21829), .B(n21826), .Z(n14785) );
  XOR U22917 ( .A(n21830), .B(n21831), .Z(n21826) );
  AND U22918 ( .A(n14792), .B(n21832), .Z(n21830) );
  XNOR U22919 ( .A(n14791), .B(n21831), .Z(n21832) );
  NAND U22920 ( .A(n21833), .B(n[961]), .Z(n14791) );
  NAND U22921 ( .A(n21523), .B(n[961]), .Z(n21833) );
  XNOR U22922 ( .A(n21834), .B(n21831), .Z(n14792) );
  XOR U22923 ( .A(n21835), .B(n21836), .Z(n21831) );
  AND U22924 ( .A(n14799), .B(n21837), .Z(n21835) );
  XNOR U22925 ( .A(n14798), .B(n21836), .Z(n21837) );
  NAND U22926 ( .A(n21838), .B(n[960]), .Z(n14798) );
  NAND U22927 ( .A(n21523), .B(n[960]), .Z(n21838) );
  XNOR U22928 ( .A(n21839), .B(n21836), .Z(n14799) );
  XOR U22929 ( .A(n21840), .B(n21841), .Z(n21836) );
  AND U22930 ( .A(n14806), .B(n21842), .Z(n21840) );
  XNOR U22931 ( .A(n14805), .B(n21841), .Z(n21842) );
  NAND U22932 ( .A(n21843), .B(n[959]), .Z(n14805) );
  NAND U22933 ( .A(n21523), .B(n[959]), .Z(n21843) );
  XNOR U22934 ( .A(n21844), .B(n21841), .Z(n14806) );
  XOR U22935 ( .A(n21845), .B(n21846), .Z(n21841) );
  AND U22936 ( .A(n14813), .B(n21847), .Z(n21845) );
  XNOR U22937 ( .A(n14812), .B(n21846), .Z(n21847) );
  NAND U22938 ( .A(n21848), .B(n[958]), .Z(n14812) );
  NAND U22939 ( .A(n21523), .B(n[958]), .Z(n21848) );
  XNOR U22940 ( .A(n21849), .B(n21846), .Z(n14813) );
  XOR U22941 ( .A(n21850), .B(n21851), .Z(n21846) );
  AND U22942 ( .A(n14820), .B(n21852), .Z(n21850) );
  XNOR U22943 ( .A(n14819), .B(n21851), .Z(n21852) );
  NAND U22944 ( .A(n21853), .B(n[957]), .Z(n14819) );
  NAND U22945 ( .A(n21523), .B(n[957]), .Z(n21853) );
  XNOR U22946 ( .A(n21854), .B(n21851), .Z(n14820) );
  XOR U22947 ( .A(n21855), .B(n21856), .Z(n21851) );
  AND U22948 ( .A(n14827), .B(n21857), .Z(n21855) );
  XNOR U22949 ( .A(n14826), .B(n21856), .Z(n21857) );
  NAND U22950 ( .A(n21858), .B(n[956]), .Z(n14826) );
  NAND U22951 ( .A(n21523), .B(n[956]), .Z(n21858) );
  XNOR U22952 ( .A(n21859), .B(n21856), .Z(n14827) );
  XOR U22953 ( .A(n21860), .B(n21861), .Z(n21856) );
  AND U22954 ( .A(n14834), .B(n21862), .Z(n21860) );
  XNOR U22955 ( .A(n14833), .B(n21861), .Z(n21862) );
  NAND U22956 ( .A(n21863), .B(n[955]), .Z(n14833) );
  NAND U22957 ( .A(n21523), .B(n[955]), .Z(n21863) );
  XNOR U22958 ( .A(n21864), .B(n21861), .Z(n14834) );
  XOR U22959 ( .A(n21865), .B(n21866), .Z(n21861) );
  AND U22960 ( .A(n14841), .B(n21867), .Z(n21865) );
  XNOR U22961 ( .A(n14840), .B(n21866), .Z(n21867) );
  NAND U22962 ( .A(n21868), .B(n[954]), .Z(n14840) );
  NAND U22963 ( .A(n21523), .B(n[954]), .Z(n21868) );
  XNOR U22964 ( .A(n21869), .B(n21866), .Z(n14841) );
  XOR U22965 ( .A(n21870), .B(n21871), .Z(n21866) );
  AND U22966 ( .A(n14848), .B(n21872), .Z(n21870) );
  XNOR U22967 ( .A(n14847), .B(n21871), .Z(n21872) );
  NAND U22968 ( .A(n21873), .B(n[953]), .Z(n14847) );
  NAND U22969 ( .A(n21523), .B(n[953]), .Z(n21873) );
  XNOR U22970 ( .A(n21874), .B(n21871), .Z(n14848) );
  XOR U22971 ( .A(n21875), .B(n21876), .Z(n21871) );
  AND U22972 ( .A(n14855), .B(n21877), .Z(n21875) );
  XNOR U22973 ( .A(n14854), .B(n21876), .Z(n21877) );
  NAND U22974 ( .A(n21878), .B(n[952]), .Z(n14854) );
  NAND U22975 ( .A(n21523), .B(n[952]), .Z(n21878) );
  XNOR U22976 ( .A(n21879), .B(n21876), .Z(n14855) );
  XOR U22977 ( .A(n21880), .B(n21881), .Z(n21876) );
  AND U22978 ( .A(n14862), .B(n21882), .Z(n21880) );
  XNOR U22979 ( .A(n14861), .B(n21881), .Z(n21882) );
  NAND U22980 ( .A(n21883), .B(n[951]), .Z(n14861) );
  NAND U22981 ( .A(n21523), .B(n[951]), .Z(n21883) );
  XNOR U22982 ( .A(n21884), .B(n21881), .Z(n14862) );
  XOR U22983 ( .A(n21885), .B(n21886), .Z(n21881) );
  AND U22984 ( .A(n14869), .B(n21887), .Z(n21885) );
  XNOR U22985 ( .A(n14868), .B(n21886), .Z(n21887) );
  NAND U22986 ( .A(n21888), .B(n[950]), .Z(n14868) );
  NAND U22987 ( .A(n21523), .B(n[950]), .Z(n21888) );
  XNOR U22988 ( .A(n21889), .B(n21886), .Z(n14869) );
  XOR U22989 ( .A(n21890), .B(n21891), .Z(n21886) );
  AND U22990 ( .A(n14876), .B(n21892), .Z(n21890) );
  XNOR U22991 ( .A(n14875), .B(n21891), .Z(n21892) );
  NAND U22992 ( .A(n21893), .B(n[949]), .Z(n14875) );
  NAND U22993 ( .A(n21523), .B(n[949]), .Z(n21893) );
  XNOR U22994 ( .A(n21894), .B(n21891), .Z(n14876) );
  XOR U22995 ( .A(n21895), .B(n21896), .Z(n21891) );
  AND U22996 ( .A(n14883), .B(n21897), .Z(n21895) );
  XNOR U22997 ( .A(n14882), .B(n21896), .Z(n21897) );
  NAND U22998 ( .A(n21898), .B(n[948]), .Z(n14882) );
  NAND U22999 ( .A(n21523), .B(n[948]), .Z(n21898) );
  XNOR U23000 ( .A(n21899), .B(n21896), .Z(n14883) );
  XOR U23001 ( .A(n21900), .B(n21901), .Z(n21896) );
  AND U23002 ( .A(n14890), .B(n21902), .Z(n21900) );
  XNOR U23003 ( .A(n14889), .B(n21901), .Z(n21902) );
  NAND U23004 ( .A(n21903), .B(n[947]), .Z(n14889) );
  NAND U23005 ( .A(n21523), .B(n[947]), .Z(n21903) );
  XNOR U23006 ( .A(n21904), .B(n21901), .Z(n14890) );
  XOR U23007 ( .A(n21905), .B(n21906), .Z(n21901) );
  AND U23008 ( .A(n14897), .B(n21907), .Z(n21905) );
  XNOR U23009 ( .A(n14896), .B(n21906), .Z(n21907) );
  NAND U23010 ( .A(n21908), .B(n[946]), .Z(n14896) );
  NAND U23011 ( .A(n21523), .B(n[946]), .Z(n21908) );
  XNOR U23012 ( .A(n21909), .B(n21906), .Z(n14897) );
  XOR U23013 ( .A(n21910), .B(n21911), .Z(n21906) );
  AND U23014 ( .A(n14904), .B(n21912), .Z(n21910) );
  XNOR U23015 ( .A(n14903), .B(n21911), .Z(n21912) );
  NAND U23016 ( .A(n21913), .B(n[945]), .Z(n14903) );
  NAND U23017 ( .A(n21523), .B(n[945]), .Z(n21913) );
  XNOR U23018 ( .A(n21914), .B(n21911), .Z(n14904) );
  XOR U23019 ( .A(n21915), .B(n21916), .Z(n21911) );
  AND U23020 ( .A(n14911), .B(n21917), .Z(n21915) );
  XNOR U23021 ( .A(n14910), .B(n21916), .Z(n21917) );
  NAND U23022 ( .A(n21918), .B(n[944]), .Z(n14910) );
  NAND U23023 ( .A(n21523), .B(n[944]), .Z(n21918) );
  XNOR U23024 ( .A(n21919), .B(n21916), .Z(n14911) );
  XOR U23025 ( .A(n21920), .B(n21921), .Z(n21916) );
  AND U23026 ( .A(n14918), .B(n21922), .Z(n21920) );
  XNOR U23027 ( .A(n14917), .B(n21921), .Z(n21922) );
  NAND U23028 ( .A(n21923), .B(n[943]), .Z(n14917) );
  NAND U23029 ( .A(n21523), .B(n[943]), .Z(n21923) );
  XNOR U23030 ( .A(n21924), .B(n21921), .Z(n14918) );
  XOR U23031 ( .A(n21925), .B(n21926), .Z(n21921) );
  AND U23032 ( .A(n14925), .B(n21927), .Z(n21925) );
  XNOR U23033 ( .A(n14924), .B(n21926), .Z(n21927) );
  NAND U23034 ( .A(n21928), .B(n[942]), .Z(n14924) );
  NAND U23035 ( .A(n21523), .B(n[942]), .Z(n21928) );
  XNOR U23036 ( .A(n21929), .B(n21926), .Z(n14925) );
  XOR U23037 ( .A(n21930), .B(n21931), .Z(n21926) );
  AND U23038 ( .A(n14932), .B(n21932), .Z(n21930) );
  XNOR U23039 ( .A(n14931), .B(n21931), .Z(n21932) );
  NAND U23040 ( .A(n21933), .B(n[941]), .Z(n14931) );
  NAND U23041 ( .A(n21523), .B(n[941]), .Z(n21933) );
  XNOR U23042 ( .A(n21934), .B(n21931), .Z(n14932) );
  XOR U23043 ( .A(n21935), .B(n21936), .Z(n21931) );
  AND U23044 ( .A(n14939), .B(n21937), .Z(n21935) );
  XNOR U23045 ( .A(n14938), .B(n21936), .Z(n21937) );
  NAND U23046 ( .A(n21938), .B(n[940]), .Z(n14938) );
  NAND U23047 ( .A(n21523), .B(n[940]), .Z(n21938) );
  XNOR U23048 ( .A(n21939), .B(n21936), .Z(n14939) );
  XOR U23049 ( .A(n21940), .B(n21941), .Z(n21936) );
  AND U23050 ( .A(n14946), .B(n21942), .Z(n21940) );
  XNOR U23051 ( .A(n14945), .B(n21941), .Z(n21942) );
  NAND U23052 ( .A(n21943), .B(n[939]), .Z(n14945) );
  NAND U23053 ( .A(n21523), .B(n[939]), .Z(n21943) );
  XNOR U23054 ( .A(n21944), .B(n21941), .Z(n14946) );
  XOR U23055 ( .A(n21945), .B(n21946), .Z(n21941) );
  AND U23056 ( .A(n14953), .B(n21947), .Z(n21945) );
  XNOR U23057 ( .A(n14952), .B(n21946), .Z(n21947) );
  NAND U23058 ( .A(n21948), .B(n[938]), .Z(n14952) );
  NAND U23059 ( .A(n21523), .B(n[938]), .Z(n21948) );
  XNOR U23060 ( .A(n21949), .B(n21946), .Z(n14953) );
  XOR U23061 ( .A(n21950), .B(n21951), .Z(n21946) );
  AND U23062 ( .A(n14960), .B(n21952), .Z(n21950) );
  XNOR U23063 ( .A(n14959), .B(n21951), .Z(n21952) );
  NAND U23064 ( .A(n21953), .B(n[937]), .Z(n14959) );
  NAND U23065 ( .A(n21523), .B(n[937]), .Z(n21953) );
  XNOR U23066 ( .A(n21954), .B(n21951), .Z(n14960) );
  XOR U23067 ( .A(n21955), .B(n21956), .Z(n21951) );
  AND U23068 ( .A(n14967), .B(n21957), .Z(n21955) );
  XNOR U23069 ( .A(n14966), .B(n21956), .Z(n21957) );
  NAND U23070 ( .A(n21958), .B(n[936]), .Z(n14966) );
  NAND U23071 ( .A(n21523), .B(n[936]), .Z(n21958) );
  XNOR U23072 ( .A(n21959), .B(n21956), .Z(n14967) );
  XOR U23073 ( .A(n21960), .B(n21961), .Z(n21956) );
  AND U23074 ( .A(n14974), .B(n21962), .Z(n21960) );
  XNOR U23075 ( .A(n14973), .B(n21961), .Z(n21962) );
  NAND U23076 ( .A(n21963), .B(n[935]), .Z(n14973) );
  NAND U23077 ( .A(n21523), .B(n[935]), .Z(n21963) );
  XNOR U23078 ( .A(n21964), .B(n21961), .Z(n14974) );
  XOR U23079 ( .A(n21965), .B(n21966), .Z(n21961) );
  AND U23080 ( .A(n14981), .B(n21967), .Z(n21965) );
  XNOR U23081 ( .A(n14980), .B(n21966), .Z(n21967) );
  NAND U23082 ( .A(n21968), .B(n[934]), .Z(n14980) );
  NAND U23083 ( .A(n21523), .B(n[934]), .Z(n21968) );
  XNOR U23084 ( .A(n21969), .B(n21966), .Z(n14981) );
  XOR U23085 ( .A(n21970), .B(n21971), .Z(n21966) );
  AND U23086 ( .A(n14988), .B(n21972), .Z(n21970) );
  XNOR U23087 ( .A(n14987), .B(n21971), .Z(n21972) );
  NAND U23088 ( .A(n21973), .B(n[933]), .Z(n14987) );
  NAND U23089 ( .A(n21523), .B(n[933]), .Z(n21973) );
  XNOR U23090 ( .A(n21974), .B(n21971), .Z(n14988) );
  XOR U23091 ( .A(n21975), .B(n21976), .Z(n21971) );
  AND U23092 ( .A(n14995), .B(n21977), .Z(n21975) );
  XNOR U23093 ( .A(n14994), .B(n21976), .Z(n21977) );
  NAND U23094 ( .A(n21978), .B(n[932]), .Z(n14994) );
  NAND U23095 ( .A(n21523), .B(n[932]), .Z(n21978) );
  XNOR U23096 ( .A(n21979), .B(n21976), .Z(n14995) );
  XOR U23097 ( .A(n21980), .B(n21981), .Z(n21976) );
  AND U23098 ( .A(n15002), .B(n21982), .Z(n21980) );
  XNOR U23099 ( .A(n15001), .B(n21981), .Z(n21982) );
  NAND U23100 ( .A(n21983), .B(n[931]), .Z(n15001) );
  NAND U23101 ( .A(n21523), .B(n[931]), .Z(n21983) );
  XNOR U23102 ( .A(n21984), .B(n21981), .Z(n15002) );
  XOR U23103 ( .A(n21985), .B(n21986), .Z(n21981) );
  AND U23104 ( .A(n15009), .B(n21987), .Z(n21985) );
  XNOR U23105 ( .A(n15008), .B(n21986), .Z(n21987) );
  NAND U23106 ( .A(n21988), .B(n[930]), .Z(n15008) );
  NAND U23107 ( .A(n21523), .B(n[930]), .Z(n21988) );
  XNOR U23108 ( .A(n21989), .B(n21986), .Z(n15009) );
  XOR U23109 ( .A(n21990), .B(n21991), .Z(n21986) );
  AND U23110 ( .A(n15016), .B(n21992), .Z(n21990) );
  XNOR U23111 ( .A(n15015), .B(n21991), .Z(n21992) );
  NAND U23112 ( .A(n21993), .B(n[929]), .Z(n15015) );
  NAND U23113 ( .A(n21523), .B(n[929]), .Z(n21993) );
  XNOR U23114 ( .A(n21994), .B(n21991), .Z(n15016) );
  XOR U23115 ( .A(n21995), .B(n21996), .Z(n21991) );
  AND U23116 ( .A(n15023), .B(n21997), .Z(n21995) );
  XNOR U23117 ( .A(n15022), .B(n21996), .Z(n21997) );
  NAND U23118 ( .A(n21998), .B(n[928]), .Z(n15022) );
  NAND U23119 ( .A(n21523), .B(n[928]), .Z(n21998) );
  XNOR U23120 ( .A(n21999), .B(n21996), .Z(n15023) );
  XOR U23121 ( .A(n22000), .B(n22001), .Z(n21996) );
  AND U23122 ( .A(n15030), .B(n22002), .Z(n22000) );
  XNOR U23123 ( .A(n15029), .B(n22001), .Z(n22002) );
  NAND U23124 ( .A(n22003), .B(n[927]), .Z(n15029) );
  NAND U23125 ( .A(n21523), .B(n[927]), .Z(n22003) );
  XNOR U23126 ( .A(n22004), .B(n22001), .Z(n15030) );
  XOR U23127 ( .A(n22005), .B(n22006), .Z(n22001) );
  AND U23128 ( .A(n15037), .B(n22007), .Z(n22005) );
  XNOR U23129 ( .A(n15036), .B(n22006), .Z(n22007) );
  NAND U23130 ( .A(n22008), .B(n[926]), .Z(n15036) );
  NAND U23131 ( .A(n21523), .B(n[926]), .Z(n22008) );
  XNOR U23132 ( .A(n22009), .B(n22006), .Z(n15037) );
  XOR U23133 ( .A(n22010), .B(n22011), .Z(n22006) );
  AND U23134 ( .A(n15044), .B(n22012), .Z(n22010) );
  XNOR U23135 ( .A(n15043), .B(n22011), .Z(n22012) );
  NAND U23136 ( .A(n22013), .B(n[925]), .Z(n15043) );
  NAND U23137 ( .A(n21523), .B(n[925]), .Z(n22013) );
  XNOR U23138 ( .A(n22014), .B(n22011), .Z(n15044) );
  XOR U23139 ( .A(n22015), .B(n22016), .Z(n22011) );
  AND U23140 ( .A(n15051), .B(n22017), .Z(n22015) );
  XNOR U23141 ( .A(n15050), .B(n22016), .Z(n22017) );
  NAND U23142 ( .A(n22018), .B(n[924]), .Z(n15050) );
  NAND U23143 ( .A(n21523), .B(n[924]), .Z(n22018) );
  XNOR U23144 ( .A(n22019), .B(n22016), .Z(n15051) );
  XOR U23145 ( .A(n22020), .B(n22021), .Z(n22016) );
  AND U23146 ( .A(n15058), .B(n22022), .Z(n22020) );
  XNOR U23147 ( .A(n15057), .B(n22021), .Z(n22022) );
  NAND U23148 ( .A(n22023), .B(n[923]), .Z(n15057) );
  NAND U23149 ( .A(n21523), .B(n[923]), .Z(n22023) );
  XNOR U23150 ( .A(n22024), .B(n22021), .Z(n15058) );
  XOR U23151 ( .A(n22025), .B(n22026), .Z(n22021) );
  AND U23152 ( .A(n15065), .B(n22027), .Z(n22025) );
  XNOR U23153 ( .A(n15064), .B(n22026), .Z(n22027) );
  NAND U23154 ( .A(n22028), .B(n[922]), .Z(n15064) );
  NAND U23155 ( .A(n21523), .B(n[922]), .Z(n22028) );
  XNOR U23156 ( .A(n22029), .B(n22026), .Z(n15065) );
  XOR U23157 ( .A(n22030), .B(n22031), .Z(n22026) );
  AND U23158 ( .A(n15072), .B(n22032), .Z(n22030) );
  XNOR U23159 ( .A(n15071), .B(n22031), .Z(n22032) );
  NAND U23160 ( .A(n22033), .B(n[921]), .Z(n15071) );
  NAND U23161 ( .A(n21523), .B(n[921]), .Z(n22033) );
  XNOR U23162 ( .A(n22034), .B(n22031), .Z(n15072) );
  XOR U23163 ( .A(n22035), .B(n22036), .Z(n22031) );
  AND U23164 ( .A(n15079), .B(n22037), .Z(n22035) );
  XNOR U23165 ( .A(n15078), .B(n22036), .Z(n22037) );
  NAND U23166 ( .A(n22038), .B(n[920]), .Z(n15078) );
  NAND U23167 ( .A(n21523), .B(n[920]), .Z(n22038) );
  XNOR U23168 ( .A(n22039), .B(n22036), .Z(n15079) );
  XOR U23169 ( .A(n22040), .B(n22041), .Z(n22036) );
  AND U23170 ( .A(n15086), .B(n22042), .Z(n22040) );
  XNOR U23171 ( .A(n15085), .B(n22041), .Z(n22042) );
  NAND U23172 ( .A(n22043), .B(n[919]), .Z(n15085) );
  NAND U23173 ( .A(n21523), .B(n[919]), .Z(n22043) );
  XNOR U23174 ( .A(n22044), .B(n22041), .Z(n15086) );
  XOR U23175 ( .A(n22045), .B(n22046), .Z(n22041) );
  AND U23176 ( .A(n15093), .B(n22047), .Z(n22045) );
  XNOR U23177 ( .A(n15092), .B(n22046), .Z(n22047) );
  NAND U23178 ( .A(n22048), .B(n[918]), .Z(n15092) );
  NAND U23179 ( .A(n21523), .B(n[918]), .Z(n22048) );
  XNOR U23180 ( .A(n22049), .B(n22046), .Z(n15093) );
  XOR U23181 ( .A(n22050), .B(n22051), .Z(n22046) );
  AND U23182 ( .A(n15100), .B(n22052), .Z(n22050) );
  XNOR U23183 ( .A(n15099), .B(n22051), .Z(n22052) );
  NAND U23184 ( .A(n22053), .B(n[917]), .Z(n15099) );
  NAND U23185 ( .A(n21523), .B(n[917]), .Z(n22053) );
  XNOR U23186 ( .A(n22054), .B(n22051), .Z(n15100) );
  XOR U23187 ( .A(n22055), .B(n22056), .Z(n22051) );
  AND U23188 ( .A(n15107), .B(n22057), .Z(n22055) );
  XNOR U23189 ( .A(n15106), .B(n22056), .Z(n22057) );
  NAND U23190 ( .A(n22058), .B(n[916]), .Z(n15106) );
  NAND U23191 ( .A(n21523), .B(n[916]), .Z(n22058) );
  XNOR U23192 ( .A(n22059), .B(n22056), .Z(n15107) );
  XOR U23193 ( .A(n22060), .B(n22061), .Z(n22056) );
  AND U23194 ( .A(n15114), .B(n22062), .Z(n22060) );
  XNOR U23195 ( .A(n15113), .B(n22061), .Z(n22062) );
  NAND U23196 ( .A(n22063), .B(n[915]), .Z(n15113) );
  NAND U23197 ( .A(n21523), .B(n[915]), .Z(n22063) );
  XNOR U23198 ( .A(n22064), .B(n22061), .Z(n15114) );
  XOR U23199 ( .A(n22065), .B(n22066), .Z(n22061) );
  AND U23200 ( .A(n15121), .B(n22067), .Z(n22065) );
  XNOR U23201 ( .A(n15120), .B(n22066), .Z(n22067) );
  NAND U23202 ( .A(n22068), .B(n[914]), .Z(n15120) );
  NAND U23203 ( .A(n21523), .B(n[914]), .Z(n22068) );
  XNOR U23204 ( .A(n22069), .B(n22066), .Z(n15121) );
  XOR U23205 ( .A(n22070), .B(n22071), .Z(n22066) );
  AND U23206 ( .A(n15128), .B(n22072), .Z(n22070) );
  XNOR U23207 ( .A(n15127), .B(n22071), .Z(n22072) );
  NAND U23208 ( .A(n22073), .B(n[913]), .Z(n15127) );
  NAND U23209 ( .A(n21523), .B(n[913]), .Z(n22073) );
  XNOR U23210 ( .A(n22074), .B(n22071), .Z(n15128) );
  XOR U23211 ( .A(n22075), .B(n22076), .Z(n22071) );
  AND U23212 ( .A(n15135), .B(n22077), .Z(n22075) );
  XNOR U23213 ( .A(n15134), .B(n22076), .Z(n22077) );
  NAND U23214 ( .A(n22078), .B(n[912]), .Z(n15134) );
  NAND U23215 ( .A(n21523), .B(n[912]), .Z(n22078) );
  XNOR U23216 ( .A(n22079), .B(n22076), .Z(n15135) );
  XOR U23217 ( .A(n22080), .B(n22081), .Z(n22076) );
  AND U23218 ( .A(n15142), .B(n22082), .Z(n22080) );
  XNOR U23219 ( .A(n15141), .B(n22081), .Z(n22082) );
  NAND U23220 ( .A(n22083), .B(n[911]), .Z(n15141) );
  NAND U23221 ( .A(n21523), .B(n[911]), .Z(n22083) );
  XNOR U23222 ( .A(n22084), .B(n22081), .Z(n15142) );
  XOR U23223 ( .A(n22085), .B(n22086), .Z(n22081) );
  AND U23224 ( .A(n15149), .B(n22087), .Z(n22085) );
  XNOR U23225 ( .A(n15148), .B(n22086), .Z(n22087) );
  NAND U23226 ( .A(n22088), .B(n[910]), .Z(n15148) );
  NAND U23227 ( .A(n21523), .B(n[910]), .Z(n22088) );
  XNOR U23228 ( .A(n22089), .B(n22086), .Z(n15149) );
  XOR U23229 ( .A(n22090), .B(n22091), .Z(n22086) );
  AND U23230 ( .A(n15156), .B(n22092), .Z(n22090) );
  XNOR U23231 ( .A(n15155), .B(n22091), .Z(n22092) );
  NAND U23232 ( .A(n22093), .B(n[909]), .Z(n15155) );
  NAND U23233 ( .A(n21523), .B(n[909]), .Z(n22093) );
  XNOR U23234 ( .A(n22094), .B(n22091), .Z(n15156) );
  XOR U23235 ( .A(n22095), .B(n22096), .Z(n22091) );
  AND U23236 ( .A(n15163), .B(n22097), .Z(n22095) );
  XNOR U23237 ( .A(n15162), .B(n22096), .Z(n22097) );
  NAND U23238 ( .A(n22098), .B(n[908]), .Z(n15162) );
  NAND U23239 ( .A(n21523), .B(n[908]), .Z(n22098) );
  XNOR U23240 ( .A(n22099), .B(n22096), .Z(n15163) );
  XOR U23241 ( .A(n22100), .B(n22101), .Z(n22096) );
  AND U23242 ( .A(n15170), .B(n22102), .Z(n22100) );
  XNOR U23243 ( .A(n15169), .B(n22101), .Z(n22102) );
  NAND U23244 ( .A(n22103), .B(n[907]), .Z(n15169) );
  NAND U23245 ( .A(n21523), .B(n[907]), .Z(n22103) );
  XNOR U23246 ( .A(n22104), .B(n22101), .Z(n15170) );
  XOR U23247 ( .A(n22105), .B(n22106), .Z(n22101) );
  AND U23248 ( .A(n15177), .B(n22107), .Z(n22105) );
  XNOR U23249 ( .A(n15176), .B(n22106), .Z(n22107) );
  NAND U23250 ( .A(n22108), .B(n[906]), .Z(n15176) );
  NAND U23251 ( .A(n21523), .B(n[906]), .Z(n22108) );
  XNOR U23252 ( .A(n22109), .B(n22106), .Z(n15177) );
  XOR U23253 ( .A(n22110), .B(n22111), .Z(n22106) );
  AND U23254 ( .A(n15184), .B(n22112), .Z(n22110) );
  XNOR U23255 ( .A(n15183), .B(n22111), .Z(n22112) );
  NAND U23256 ( .A(n22113), .B(n[905]), .Z(n15183) );
  NAND U23257 ( .A(n21523), .B(n[905]), .Z(n22113) );
  XNOR U23258 ( .A(n22114), .B(n22111), .Z(n15184) );
  XOR U23259 ( .A(n22115), .B(n22116), .Z(n22111) );
  AND U23260 ( .A(n15191), .B(n22117), .Z(n22115) );
  XNOR U23261 ( .A(n15190), .B(n22116), .Z(n22117) );
  NAND U23262 ( .A(n22118), .B(n[904]), .Z(n15190) );
  NAND U23263 ( .A(n21523), .B(n[904]), .Z(n22118) );
  XNOR U23264 ( .A(n22119), .B(n22116), .Z(n15191) );
  XOR U23265 ( .A(n22120), .B(n22121), .Z(n22116) );
  AND U23266 ( .A(n15198), .B(n22122), .Z(n22120) );
  XNOR U23267 ( .A(n15197), .B(n22121), .Z(n22122) );
  NAND U23268 ( .A(n22123), .B(n[903]), .Z(n15197) );
  NAND U23269 ( .A(n21523), .B(n[903]), .Z(n22123) );
  XNOR U23270 ( .A(n22124), .B(n22121), .Z(n15198) );
  XOR U23271 ( .A(n22125), .B(n22126), .Z(n22121) );
  AND U23272 ( .A(n15205), .B(n22127), .Z(n22125) );
  XNOR U23273 ( .A(n15204), .B(n22126), .Z(n22127) );
  NAND U23274 ( .A(n22128), .B(n[902]), .Z(n15204) );
  NAND U23275 ( .A(n21523), .B(n[902]), .Z(n22128) );
  XNOR U23276 ( .A(n22129), .B(n22126), .Z(n15205) );
  XOR U23277 ( .A(n22130), .B(n22131), .Z(n22126) );
  AND U23278 ( .A(n15212), .B(n22132), .Z(n22130) );
  XNOR U23279 ( .A(n15211), .B(n22131), .Z(n22132) );
  NAND U23280 ( .A(n22133), .B(n[901]), .Z(n15211) );
  NAND U23281 ( .A(n21523), .B(n[901]), .Z(n22133) );
  XNOR U23282 ( .A(n22134), .B(n22131), .Z(n15212) );
  XOR U23283 ( .A(n22135), .B(n22136), .Z(n22131) );
  AND U23284 ( .A(n15219), .B(n22137), .Z(n22135) );
  XNOR U23285 ( .A(n15218), .B(n22136), .Z(n22137) );
  NAND U23286 ( .A(n22138), .B(n[900]), .Z(n15218) );
  NAND U23287 ( .A(n21523), .B(n[900]), .Z(n22138) );
  XNOR U23288 ( .A(n22139), .B(n22136), .Z(n15219) );
  XOR U23289 ( .A(n22140), .B(n22141), .Z(n22136) );
  AND U23290 ( .A(n15226), .B(n22142), .Z(n22140) );
  XNOR U23291 ( .A(n15225), .B(n22141), .Z(n22142) );
  NAND U23292 ( .A(n22143), .B(n[899]), .Z(n15225) );
  NAND U23293 ( .A(n21523), .B(n[899]), .Z(n22143) );
  XNOR U23294 ( .A(n22144), .B(n22141), .Z(n15226) );
  XOR U23295 ( .A(n22145), .B(n22146), .Z(n22141) );
  AND U23296 ( .A(n15233), .B(n22147), .Z(n22145) );
  XNOR U23297 ( .A(n15232), .B(n22146), .Z(n22147) );
  NAND U23298 ( .A(n22148), .B(n[898]), .Z(n15232) );
  NAND U23299 ( .A(n21523), .B(n[898]), .Z(n22148) );
  XNOR U23300 ( .A(n22149), .B(n22146), .Z(n15233) );
  XOR U23301 ( .A(n22150), .B(n22151), .Z(n22146) );
  AND U23302 ( .A(n15240), .B(n22152), .Z(n22150) );
  XNOR U23303 ( .A(n15239), .B(n22151), .Z(n22152) );
  NAND U23304 ( .A(n22153), .B(n[897]), .Z(n15239) );
  NAND U23305 ( .A(n21523), .B(n[897]), .Z(n22153) );
  XNOR U23306 ( .A(n22154), .B(n22151), .Z(n15240) );
  XOR U23307 ( .A(n22155), .B(n22156), .Z(n22151) );
  AND U23308 ( .A(n15247), .B(n22157), .Z(n22155) );
  XNOR U23309 ( .A(n15246), .B(n22156), .Z(n22157) );
  NAND U23310 ( .A(n22158), .B(n[896]), .Z(n15246) );
  NAND U23311 ( .A(n21523), .B(n[896]), .Z(n22158) );
  XNOR U23312 ( .A(n22159), .B(n22156), .Z(n15247) );
  XOR U23313 ( .A(n22160), .B(n22161), .Z(n22156) );
  AND U23314 ( .A(n15254), .B(n22162), .Z(n22160) );
  XNOR U23315 ( .A(n15253), .B(n22161), .Z(n22162) );
  NAND U23316 ( .A(n22163), .B(n[895]), .Z(n15253) );
  NAND U23317 ( .A(n21523), .B(n[895]), .Z(n22163) );
  XNOR U23318 ( .A(n22164), .B(n22161), .Z(n15254) );
  XOR U23319 ( .A(n22165), .B(n22166), .Z(n22161) );
  AND U23320 ( .A(n15261), .B(n22167), .Z(n22165) );
  XNOR U23321 ( .A(n15260), .B(n22166), .Z(n22167) );
  NAND U23322 ( .A(n22168), .B(n[894]), .Z(n15260) );
  NAND U23323 ( .A(n21523), .B(n[894]), .Z(n22168) );
  XNOR U23324 ( .A(n22169), .B(n22166), .Z(n15261) );
  XOR U23325 ( .A(n22170), .B(n22171), .Z(n22166) );
  AND U23326 ( .A(n15268), .B(n22172), .Z(n22170) );
  XNOR U23327 ( .A(n15267), .B(n22171), .Z(n22172) );
  NAND U23328 ( .A(n22173), .B(n[893]), .Z(n15267) );
  NAND U23329 ( .A(n21523), .B(n[893]), .Z(n22173) );
  XNOR U23330 ( .A(n22174), .B(n22171), .Z(n15268) );
  XOR U23331 ( .A(n22175), .B(n22176), .Z(n22171) );
  AND U23332 ( .A(n15275), .B(n22177), .Z(n22175) );
  XNOR U23333 ( .A(n15274), .B(n22176), .Z(n22177) );
  NAND U23334 ( .A(n22178), .B(n[892]), .Z(n15274) );
  NAND U23335 ( .A(n21523), .B(n[892]), .Z(n22178) );
  XNOR U23336 ( .A(n22179), .B(n22176), .Z(n15275) );
  XOR U23337 ( .A(n22180), .B(n22181), .Z(n22176) );
  AND U23338 ( .A(n15282), .B(n22182), .Z(n22180) );
  XNOR U23339 ( .A(n15281), .B(n22181), .Z(n22182) );
  NAND U23340 ( .A(n22183), .B(n[891]), .Z(n15281) );
  NAND U23341 ( .A(n21523), .B(n[891]), .Z(n22183) );
  XNOR U23342 ( .A(n22184), .B(n22181), .Z(n15282) );
  XOR U23343 ( .A(n22185), .B(n22186), .Z(n22181) );
  AND U23344 ( .A(n15289), .B(n22187), .Z(n22185) );
  XNOR U23345 ( .A(n15288), .B(n22186), .Z(n22187) );
  NAND U23346 ( .A(n22188), .B(n[890]), .Z(n15288) );
  NAND U23347 ( .A(n21523), .B(n[890]), .Z(n22188) );
  XNOR U23348 ( .A(n22189), .B(n22186), .Z(n15289) );
  XOR U23349 ( .A(n22190), .B(n22191), .Z(n22186) );
  AND U23350 ( .A(n15296), .B(n22192), .Z(n22190) );
  XNOR U23351 ( .A(n15295), .B(n22191), .Z(n22192) );
  NAND U23352 ( .A(n22193), .B(n[889]), .Z(n15295) );
  NAND U23353 ( .A(n21523), .B(n[889]), .Z(n22193) );
  XNOR U23354 ( .A(n22194), .B(n22191), .Z(n15296) );
  XOR U23355 ( .A(n22195), .B(n22196), .Z(n22191) );
  AND U23356 ( .A(n15303), .B(n22197), .Z(n22195) );
  XNOR U23357 ( .A(n15302), .B(n22196), .Z(n22197) );
  NAND U23358 ( .A(n22198), .B(n[888]), .Z(n15302) );
  NAND U23359 ( .A(n21523), .B(n[888]), .Z(n22198) );
  XNOR U23360 ( .A(n22199), .B(n22196), .Z(n15303) );
  XOR U23361 ( .A(n22200), .B(n22201), .Z(n22196) );
  AND U23362 ( .A(n15310), .B(n22202), .Z(n22200) );
  XNOR U23363 ( .A(n15309), .B(n22201), .Z(n22202) );
  NAND U23364 ( .A(n22203), .B(n[887]), .Z(n15309) );
  NAND U23365 ( .A(n21523), .B(n[887]), .Z(n22203) );
  XNOR U23366 ( .A(n22204), .B(n22201), .Z(n15310) );
  XOR U23367 ( .A(n22205), .B(n22206), .Z(n22201) );
  AND U23368 ( .A(n15317), .B(n22207), .Z(n22205) );
  XNOR U23369 ( .A(n15316), .B(n22206), .Z(n22207) );
  NAND U23370 ( .A(n22208), .B(n[886]), .Z(n15316) );
  NAND U23371 ( .A(n21523), .B(n[886]), .Z(n22208) );
  XNOR U23372 ( .A(n22209), .B(n22206), .Z(n15317) );
  XOR U23373 ( .A(n22210), .B(n22211), .Z(n22206) );
  AND U23374 ( .A(n15324), .B(n22212), .Z(n22210) );
  XNOR U23375 ( .A(n15323), .B(n22211), .Z(n22212) );
  NAND U23376 ( .A(n22213), .B(n[885]), .Z(n15323) );
  NAND U23377 ( .A(n21523), .B(n[885]), .Z(n22213) );
  XNOR U23378 ( .A(n22214), .B(n22211), .Z(n15324) );
  XOR U23379 ( .A(n22215), .B(n22216), .Z(n22211) );
  AND U23380 ( .A(n15331), .B(n22217), .Z(n22215) );
  XNOR U23381 ( .A(n15330), .B(n22216), .Z(n22217) );
  NAND U23382 ( .A(n22218), .B(n[884]), .Z(n15330) );
  NAND U23383 ( .A(n21523), .B(n[884]), .Z(n22218) );
  XNOR U23384 ( .A(n22219), .B(n22216), .Z(n15331) );
  XOR U23385 ( .A(n22220), .B(n22221), .Z(n22216) );
  AND U23386 ( .A(n15338), .B(n22222), .Z(n22220) );
  XNOR U23387 ( .A(n15337), .B(n22221), .Z(n22222) );
  NAND U23388 ( .A(n22223), .B(n[883]), .Z(n15337) );
  NAND U23389 ( .A(n21523), .B(n[883]), .Z(n22223) );
  XNOR U23390 ( .A(n22224), .B(n22221), .Z(n15338) );
  XOR U23391 ( .A(n22225), .B(n22226), .Z(n22221) );
  AND U23392 ( .A(n15345), .B(n22227), .Z(n22225) );
  XNOR U23393 ( .A(n15344), .B(n22226), .Z(n22227) );
  NAND U23394 ( .A(n22228), .B(n[882]), .Z(n15344) );
  NAND U23395 ( .A(n21523), .B(n[882]), .Z(n22228) );
  XNOR U23396 ( .A(n22229), .B(n22226), .Z(n15345) );
  XOR U23397 ( .A(n22230), .B(n22231), .Z(n22226) );
  AND U23398 ( .A(n15352), .B(n22232), .Z(n22230) );
  XNOR U23399 ( .A(n15351), .B(n22231), .Z(n22232) );
  NAND U23400 ( .A(n22233), .B(n[881]), .Z(n15351) );
  NAND U23401 ( .A(n21523), .B(n[881]), .Z(n22233) );
  XNOR U23402 ( .A(n22234), .B(n22231), .Z(n15352) );
  XOR U23403 ( .A(n22235), .B(n22236), .Z(n22231) );
  AND U23404 ( .A(n15359), .B(n22237), .Z(n22235) );
  XNOR U23405 ( .A(n15358), .B(n22236), .Z(n22237) );
  NAND U23406 ( .A(n22238), .B(n[880]), .Z(n15358) );
  NAND U23407 ( .A(n21523), .B(n[880]), .Z(n22238) );
  XNOR U23408 ( .A(n22239), .B(n22236), .Z(n15359) );
  XOR U23409 ( .A(n22240), .B(n22241), .Z(n22236) );
  AND U23410 ( .A(n15366), .B(n22242), .Z(n22240) );
  XNOR U23411 ( .A(n15365), .B(n22241), .Z(n22242) );
  NAND U23412 ( .A(n22243), .B(n[879]), .Z(n15365) );
  NAND U23413 ( .A(n21523), .B(n[879]), .Z(n22243) );
  XNOR U23414 ( .A(n22244), .B(n22241), .Z(n15366) );
  XOR U23415 ( .A(n22245), .B(n22246), .Z(n22241) );
  AND U23416 ( .A(n15373), .B(n22247), .Z(n22245) );
  XNOR U23417 ( .A(n15372), .B(n22246), .Z(n22247) );
  NAND U23418 ( .A(n22248), .B(n[878]), .Z(n15372) );
  NAND U23419 ( .A(n21523), .B(n[878]), .Z(n22248) );
  XNOR U23420 ( .A(n22249), .B(n22246), .Z(n15373) );
  XOR U23421 ( .A(n22250), .B(n22251), .Z(n22246) );
  AND U23422 ( .A(n15380), .B(n22252), .Z(n22250) );
  XNOR U23423 ( .A(n15379), .B(n22251), .Z(n22252) );
  NAND U23424 ( .A(n22253), .B(n[877]), .Z(n15379) );
  NAND U23425 ( .A(n21523), .B(n[877]), .Z(n22253) );
  XNOR U23426 ( .A(n22254), .B(n22251), .Z(n15380) );
  XOR U23427 ( .A(n22255), .B(n22256), .Z(n22251) );
  AND U23428 ( .A(n15387), .B(n22257), .Z(n22255) );
  XNOR U23429 ( .A(n15386), .B(n22256), .Z(n22257) );
  NAND U23430 ( .A(n22258), .B(n[876]), .Z(n15386) );
  NAND U23431 ( .A(n21523), .B(n[876]), .Z(n22258) );
  XNOR U23432 ( .A(n22259), .B(n22256), .Z(n15387) );
  XOR U23433 ( .A(n22260), .B(n22261), .Z(n22256) );
  AND U23434 ( .A(n15394), .B(n22262), .Z(n22260) );
  XNOR U23435 ( .A(n15393), .B(n22261), .Z(n22262) );
  NAND U23436 ( .A(n22263), .B(n[875]), .Z(n15393) );
  NAND U23437 ( .A(n21523), .B(n[875]), .Z(n22263) );
  XNOR U23438 ( .A(n22264), .B(n22261), .Z(n15394) );
  XOR U23439 ( .A(n22265), .B(n22266), .Z(n22261) );
  AND U23440 ( .A(n15401), .B(n22267), .Z(n22265) );
  XNOR U23441 ( .A(n15400), .B(n22266), .Z(n22267) );
  NAND U23442 ( .A(n22268), .B(n[874]), .Z(n15400) );
  NAND U23443 ( .A(n21523), .B(n[874]), .Z(n22268) );
  XNOR U23444 ( .A(n22269), .B(n22266), .Z(n15401) );
  XOR U23445 ( .A(n22270), .B(n22271), .Z(n22266) );
  AND U23446 ( .A(n15408), .B(n22272), .Z(n22270) );
  XNOR U23447 ( .A(n15407), .B(n22271), .Z(n22272) );
  NAND U23448 ( .A(n22273), .B(n[873]), .Z(n15407) );
  NAND U23449 ( .A(n21523), .B(n[873]), .Z(n22273) );
  XNOR U23450 ( .A(n22274), .B(n22271), .Z(n15408) );
  XOR U23451 ( .A(n22275), .B(n22276), .Z(n22271) );
  AND U23452 ( .A(n15415), .B(n22277), .Z(n22275) );
  XNOR U23453 ( .A(n15414), .B(n22276), .Z(n22277) );
  NAND U23454 ( .A(n22278), .B(n[872]), .Z(n15414) );
  NAND U23455 ( .A(n21523), .B(n[872]), .Z(n22278) );
  XNOR U23456 ( .A(n22279), .B(n22276), .Z(n15415) );
  XOR U23457 ( .A(n22280), .B(n22281), .Z(n22276) );
  AND U23458 ( .A(n15422), .B(n22282), .Z(n22280) );
  XNOR U23459 ( .A(n15421), .B(n22281), .Z(n22282) );
  NAND U23460 ( .A(n22283), .B(n[871]), .Z(n15421) );
  NAND U23461 ( .A(n21523), .B(n[871]), .Z(n22283) );
  XNOR U23462 ( .A(n22284), .B(n22281), .Z(n15422) );
  XOR U23463 ( .A(n22285), .B(n22286), .Z(n22281) );
  AND U23464 ( .A(n15429), .B(n22287), .Z(n22285) );
  XNOR U23465 ( .A(n15428), .B(n22286), .Z(n22287) );
  NAND U23466 ( .A(n22288), .B(n[870]), .Z(n15428) );
  NAND U23467 ( .A(n21523), .B(n[870]), .Z(n22288) );
  XNOR U23468 ( .A(n22289), .B(n22286), .Z(n15429) );
  XOR U23469 ( .A(n22290), .B(n22291), .Z(n22286) );
  AND U23470 ( .A(n15436), .B(n22292), .Z(n22290) );
  XNOR U23471 ( .A(n15435), .B(n22291), .Z(n22292) );
  NAND U23472 ( .A(n22293), .B(n[869]), .Z(n15435) );
  NAND U23473 ( .A(n21523), .B(n[869]), .Z(n22293) );
  XNOR U23474 ( .A(n22294), .B(n22291), .Z(n15436) );
  XOR U23475 ( .A(n22295), .B(n22296), .Z(n22291) );
  AND U23476 ( .A(n15443), .B(n22297), .Z(n22295) );
  XNOR U23477 ( .A(n15442), .B(n22296), .Z(n22297) );
  NAND U23478 ( .A(n22298), .B(n[868]), .Z(n15442) );
  NAND U23479 ( .A(n21523), .B(n[868]), .Z(n22298) );
  XNOR U23480 ( .A(n22299), .B(n22296), .Z(n15443) );
  XOR U23481 ( .A(n22300), .B(n22301), .Z(n22296) );
  AND U23482 ( .A(n15450), .B(n22302), .Z(n22300) );
  XNOR U23483 ( .A(n15449), .B(n22301), .Z(n22302) );
  NAND U23484 ( .A(n22303), .B(n[867]), .Z(n15449) );
  NAND U23485 ( .A(n21523), .B(n[867]), .Z(n22303) );
  XNOR U23486 ( .A(n22304), .B(n22301), .Z(n15450) );
  XOR U23487 ( .A(n22305), .B(n22306), .Z(n22301) );
  AND U23488 ( .A(n15457), .B(n22307), .Z(n22305) );
  XNOR U23489 ( .A(n15456), .B(n22306), .Z(n22307) );
  NAND U23490 ( .A(n22308), .B(n[866]), .Z(n15456) );
  NAND U23491 ( .A(n21523), .B(n[866]), .Z(n22308) );
  XNOR U23492 ( .A(n22309), .B(n22306), .Z(n15457) );
  XOR U23493 ( .A(n22310), .B(n22311), .Z(n22306) );
  AND U23494 ( .A(n15464), .B(n22312), .Z(n22310) );
  XNOR U23495 ( .A(n15463), .B(n22311), .Z(n22312) );
  NAND U23496 ( .A(n22313), .B(n[865]), .Z(n15463) );
  NAND U23497 ( .A(n21523), .B(n[865]), .Z(n22313) );
  XNOR U23498 ( .A(n22314), .B(n22311), .Z(n15464) );
  XOR U23499 ( .A(n22315), .B(n22316), .Z(n22311) );
  AND U23500 ( .A(n15471), .B(n22317), .Z(n22315) );
  XNOR U23501 ( .A(n15470), .B(n22316), .Z(n22317) );
  NAND U23502 ( .A(n22318), .B(n[864]), .Z(n15470) );
  NAND U23503 ( .A(n21523), .B(n[864]), .Z(n22318) );
  XNOR U23504 ( .A(n22319), .B(n22316), .Z(n15471) );
  XOR U23505 ( .A(n22320), .B(n22321), .Z(n22316) );
  AND U23506 ( .A(n15478), .B(n22322), .Z(n22320) );
  XNOR U23507 ( .A(n15477), .B(n22321), .Z(n22322) );
  NAND U23508 ( .A(n22323), .B(n[863]), .Z(n15477) );
  NAND U23509 ( .A(n21523), .B(n[863]), .Z(n22323) );
  XNOR U23510 ( .A(n22324), .B(n22321), .Z(n15478) );
  XOR U23511 ( .A(n22325), .B(n22326), .Z(n22321) );
  AND U23512 ( .A(n15485), .B(n22327), .Z(n22325) );
  XNOR U23513 ( .A(n15484), .B(n22326), .Z(n22327) );
  NAND U23514 ( .A(n22328), .B(n[862]), .Z(n15484) );
  NAND U23515 ( .A(n21523), .B(n[862]), .Z(n22328) );
  XNOR U23516 ( .A(n22329), .B(n22326), .Z(n15485) );
  XOR U23517 ( .A(n22330), .B(n22331), .Z(n22326) );
  AND U23518 ( .A(n15492), .B(n22332), .Z(n22330) );
  XNOR U23519 ( .A(n15491), .B(n22331), .Z(n22332) );
  NAND U23520 ( .A(n22333), .B(n[861]), .Z(n15491) );
  NAND U23521 ( .A(n21523), .B(n[861]), .Z(n22333) );
  XNOR U23522 ( .A(n22334), .B(n22331), .Z(n15492) );
  XOR U23523 ( .A(n22335), .B(n22336), .Z(n22331) );
  AND U23524 ( .A(n15499), .B(n22337), .Z(n22335) );
  XNOR U23525 ( .A(n15498), .B(n22336), .Z(n22337) );
  NAND U23526 ( .A(n22338), .B(n[860]), .Z(n15498) );
  NAND U23527 ( .A(n21523), .B(n[860]), .Z(n22338) );
  XNOR U23528 ( .A(n22339), .B(n22336), .Z(n15499) );
  XOR U23529 ( .A(n22340), .B(n22341), .Z(n22336) );
  AND U23530 ( .A(n15506), .B(n22342), .Z(n22340) );
  XNOR U23531 ( .A(n15505), .B(n22341), .Z(n22342) );
  NAND U23532 ( .A(n22343), .B(n[859]), .Z(n15505) );
  NAND U23533 ( .A(n21523), .B(n[859]), .Z(n22343) );
  XNOR U23534 ( .A(n22344), .B(n22341), .Z(n15506) );
  XOR U23535 ( .A(n22345), .B(n22346), .Z(n22341) );
  AND U23536 ( .A(n15513), .B(n22347), .Z(n22345) );
  XNOR U23537 ( .A(n15512), .B(n22346), .Z(n22347) );
  NAND U23538 ( .A(n22348), .B(n[858]), .Z(n15512) );
  NAND U23539 ( .A(n21523), .B(n[858]), .Z(n22348) );
  XNOR U23540 ( .A(n22349), .B(n22346), .Z(n15513) );
  XOR U23541 ( .A(n22350), .B(n22351), .Z(n22346) );
  AND U23542 ( .A(n15520), .B(n22352), .Z(n22350) );
  XNOR U23543 ( .A(n15519), .B(n22351), .Z(n22352) );
  NAND U23544 ( .A(n22353), .B(n[857]), .Z(n15519) );
  NAND U23545 ( .A(n21523), .B(n[857]), .Z(n22353) );
  XNOR U23546 ( .A(n22354), .B(n22351), .Z(n15520) );
  XOR U23547 ( .A(n22355), .B(n22356), .Z(n22351) );
  AND U23548 ( .A(n15527), .B(n22357), .Z(n22355) );
  XNOR U23549 ( .A(n15526), .B(n22356), .Z(n22357) );
  NAND U23550 ( .A(n22358), .B(n[856]), .Z(n15526) );
  NAND U23551 ( .A(n21523), .B(n[856]), .Z(n22358) );
  XNOR U23552 ( .A(n22359), .B(n22356), .Z(n15527) );
  XOR U23553 ( .A(n22360), .B(n22361), .Z(n22356) );
  AND U23554 ( .A(n15534), .B(n22362), .Z(n22360) );
  XNOR U23555 ( .A(n15533), .B(n22361), .Z(n22362) );
  NAND U23556 ( .A(n22363), .B(n[855]), .Z(n15533) );
  NAND U23557 ( .A(n21523), .B(n[855]), .Z(n22363) );
  XNOR U23558 ( .A(n22364), .B(n22361), .Z(n15534) );
  XOR U23559 ( .A(n22365), .B(n22366), .Z(n22361) );
  AND U23560 ( .A(n15541), .B(n22367), .Z(n22365) );
  XNOR U23561 ( .A(n15540), .B(n22366), .Z(n22367) );
  NAND U23562 ( .A(n22368), .B(n[854]), .Z(n15540) );
  NAND U23563 ( .A(n21523), .B(n[854]), .Z(n22368) );
  XNOR U23564 ( .A(n22369), .B(n22366), .Z(n15541) );
  XOR U23565 ( .A(n22370), .B(n22371), .Z(n22366) );
  AND U23566 ( .A(n15548), .B(n22372), .Z(n22370) );
  XNOR U23567 ( .A(n15547), .B(n22371), .Z(n22372) );
  NAND U23568 ( .A(n22373), .B(n[853]), .Z(n15547) );
  NAND U23569 ( .A(n21523), .B(n[853]), .Z(n22373) );
  XNOR U23570 ( .A(n22374), .B(n22371), .Z(n15548) );
  XOR U23571 ( .A(n22375), .B(n22376), .Z(n22371) );
  AND U23572 ( .A(n15555), .B(n22377), .Z(n22375) );
  XNOR U23573 ( .A(n15554), .B(n22376), .Z(n22377) );
  NAND U23574 ( .A(n22378), .B(n[852]), .Z(n15554) );
  NAND U23575 ( .A(n21523), .B(n[852]), .Z(n22378) );
  XNOR U23576 ( .A(n22379), .B(n22376), .Z(n15555) );
  XOR U23577 ( .A(n22380), .B(n22381), .Z(n22376) );
  AND U23578 ( .A(n15562), .B(n22382), .Z(n22380) );
  XNOR U23579 ( .A(n15561), .B(n22381), .Z(n22382) );
  NAND U23580 ( .A(n22383), .B(n[851]), .Z(n15561) );
  NAND U23581 ( .A(n21523), .B(n[851]), .Z(n22383) );
  XNOR U23582 ( .A(n22384), .B(n22381), .Z(n15562) );
  XOR U23583 ( .A(n22385), .B(n22386), .Z(n22381) );
  AND U23584 ( .A(n15569), .B(n22387), .Z(n22385) );
  XNOR U23585 ( .A(n15568), .B(n22386), .Z(n22387) );
  NAND U23586 ( .A(n22388), .B(n[850]), .Z(n15568) );
  NAND U23587 ( .A(n21523), .B(n[850]), .Z(n22388) );
  XNOR U23588 ( .A(n22389), .B(n22386), .Z(n15569) );
  XOR U23589 ( .A(n22390), .B(n22391), .Z(n22386) );
  AND U23590 ( .A(n15576), .B(n22392), .Z(n22390) );
  XNOR U23591 ( .A(n15575), .B(n22391), .Z(n22392) );
  NAND U23592 ( .A(n22393), .B(n[849]), .Z(n15575) );
  NAND U23593 ( .A(n21523), .B(n[849]), .Z(n22393) );
  XNOR U23594 ( .A(n22394), .B(n22391), .Z(n15576) );
  XOR U23595 ( .A(n22395), .B(n22396), .Z(n22391) );
  AND U23596 ( .A(n15583), .B(n22397), .Z(n22395) );
  XNOR U23597 ( .A(n15582), .B(n22396), .Z(n22397) );
  NAND U23598 ( .A(n22398), .B(n[848]), .Z(n15582) );
  NAND U23599 ( .A(n21523), .B(n[848]), .Z(n22398) );
  XNOR U23600 ( .A(n22399), .B(n22396), .Z(n15583) );
  XOR U23601 ( .A(n22400), .B(n22401), .Z(n22396) );
  AND U23602 ( .A(n15590), .B(n22402), .Z(n22400) );
  XNOR U23603 ( .A(n15589), .B(n22401), .Z(n22402) );
  NAND U23604 ( .A(n22403), .B(n[847]), .Z(n15589) );
  NAND U23605 ( .A(n21523), .B(n[847]), .Z(n22403) );
  XNOR U23606 ( .A(n22404), .B(n22401), .Z(n15590) );
  XOR U23607 ( .A(n22405), .B(n22406), .Z(n22401) );
  AND U23608 ( .A(n15597), .B(n22407), .Z(n22405) );
  XNOR U23609 ( .A(n15596), .B(n22406), .Z(n22407) );
  NAND U23610 ( .A(n22408), .B(n[846]), .Z(n15596) );
  NAND U23611 ( .A(n21523), .B(n[846]), .Z(n22408) );
  XNOR U23612 ( .A(n22409), .B(n22406), .Z(n15597) );
  XOR U23613 ( .A(n22410), .B(n22411), .Z(n22406) );
  AND U23614 ( .A(n15604), .B(n22412), .Z(n22410) );
  XNOR U23615 ( .A(n15603), .B(n22411), .Z(n22412) );
  NAND U23616 ( .A(n22413), .B(n[845]), .Z(n15603) );
  NAND U23617 ( .A(n21523), .B(n[845]), .Z(n22413) );
  XNOR U23618 ( .A(n22414), .B(n22411), .Z(n15604) );
  XOR U23619 ( .A(n22415), .B(n22416), .Z(n22411) );
  AND U23620 ( .A(n15611), .B(n22417), .Z(n22415) );
  XNOR U23621 ( .A(n15610), .B(n22416), .Z(n22417) );
  NAND U23622 ( .A(n22418), .B(n[844]), .Z(n15610) );
  NAND U23623 ( .A(n21523), .B(n[844]), .Z(n22418) );
  XNOR U23624 ( .A(n22419), .B(n22416), .Z(n15611) );
  XOR U23625 ( .A(n22420), .B(n22421), .Z(n22416) );
  AND U23626 ( .A(n15618), .B(n22422), .Z(n22420) );
  XNOR U23627 ( .A(n15617), .B(n22421), .Z(n22422) );
  NAND U23628 ( .A(n22423), .B(n[843]), .Z(n15617) );
  NAND U23629 ( .A(n21523), .B(n[843]), .Z(n22423) );
  XNOR U23630 ( .A(n22424), .B(n22421), .Z(n15618) );
  XOR U23631 ( .A(n22425), .B(n22426), .Z(n22421) );
  AND U23632 ( .A(n15625), .B(n22427), .Z(n22425) );
  XNOR U23633 ( .A(n15624), .B(n22426), .Z(n22427) );
  NAND U23634 ( .A(n22428), .B(n[842]), .Z(n15624) );
  NAND U23635 ( .A(n21523), .B(n[842]), .Z(n22428) );
  XNOR U23636 ( .A(n22429), .B(n22426), .Z(n15625) );
  XOR U23637 ( .A(n22430), .B(n22431), .Z(n22426) );
  AND U23638 ( .A(n15632), .B(n22432), .Z(n22430) );
  XNOR U23639 ( .A(n15631), .B(n22431), .Z(n22432) );
  NAND U23640 ( .A(n22433), .B(n[841]), .Z(n15631) );
  NAND U23641 ( .A(n21523), .B(n[841]), .Z(n22433) );
  XNOR U23642 ( .A(n22434), .B(n22431), .Z(n15632) );
  XOR U23643 ( .A(n22435), .B(n22436), .Z(n22431) );
  AND U23644 ( .A(n15639), .B(n22437), .Z(n22435) );
  XNOR U23645 ( .A(n15638), .B(n22436), .Z(n22437) );
  NAND U23646 ( .A(n22438), .B(n[840]), .Z(n15638) );
  NAND U23647 ( .A(n21523), .B(n[840]), .Z(n22438) );
  XNOR U23648 ( .A(n22439), .B(n22436), .Z(n15639) );
  XOR U23649 ( .A(n22440), .B(n22441), .Z(n22436) );
  AND U23650 ( .A(n15646), .B(n22442), .Z(n22440) );
  XNOR U23651 ( .A(n15645), .B(n22441), .Z(n22442) );
  NAND U23652 ( .A(n22443), .B(n[839]), .Z(n15645) );
  NAND U23653 ( .A(n21523), .B(n[839]), .Z(n22443) );
  XNOR U23654 ( .A(n22444), .B(n22441), .Z(n15646) );
  XOR U23655 ( .A(n22445), .B(n22446), .Z(n22441) );
  AND U23656 ( .A(n15653), .B(n22447), .Z(n22445) );
  XNOR U23657 ( .A(n15652), .B(n22446), .Z(n22447) );
  NAND U23658 ( .A(n22448), .B(n[838]), .Z(n15652) );
  NAND U23659 ( .A(n21523), .B(n[838]), .Z(n22448) );
  XNOR U23660 ( .A(n22449), .B(n22446), .Z(n15653) );
  XOR U23661 ( .A(n22450), .B(n22451), .Z(n22446) );
  AND U23662 ( .A(n15660), .B(n22452), .Z(n22450) );
  XNOR U23663 ( .A(n15659), .B(n22451), .Z(n22452) );
  NAND U23664 ( .A(n22453), .B(n[837]), .Z(n15659) );
  NAND U23665 ( .A(n21523), .B(n[837]), .Z(n22453) );
  XNOR U23666 ( .A(n22454), .B(n22451), .Z(n15660) );
  XOR U23667 ( .A(n22455), .B(n22456), .Z(n22451) );
  AND U23668 ( .A(n15667), .B(n22457), .Z(n22455) );
  XNOR U23669 ( .A(n15666), .B(n22456), .Z(n22457) );
  NAND U23670 ( .A(n22458), .B(n[836]), .Z(n15666) );
  NAND U23671 ( .A(n21523), .B(n[836]), .Z(n22458) );
  XNOR U23672 ( .A(n22459), .B(n22456), .Z(n15667) );
  XOR U23673 ( .A(n22460), .B(n22461), .Z(n22456) );
  AND U23674 ( .A(n15674), .B(n22462), .Z(n22460) );
  XNOR U23675 ( .A(n15673), .B(n22461), .Z(n22462) );
  NAND U23676 ( .A(n22463), .B(n[835]), .Z(n15673) );
  NAND U23677 ( .A(n21523), .B(n[835]), .Z(n22463) );
  XNOR U23678 ( .A(n22464), .B(n22461), .Z(n15674) );
  XOR U23679 ( .A(n22465), .B(n22466), .Z(n22461) );
  AND U23680 ( .A(n15681), .B(n22467), .Z(n22465) );
  XNOR U23681 ( .A(n15680), .B(n22466), .Z(n22467) );
  NAND U23682 ( .A(n22468), .B(n[834]), .Z(n15680) );
  NAND U23683 ( .A(n21523), .B(n[834]), .Z(n22468) );
  XNOR U23684 ( .A(n22469), .B(n22466), .Z(n15681) );
  XOR U23685 ( .A(n22470), .B(n22471), .Z(n22466) );
  AND U23686 ( .A(n15688), .B(n22472), .Z(n22470) );
  XNOR U23687 ( .A(n15687), .B(n22471), .Z(n22472) );
  NAND U23688 ( .A(n22473), .B(n[833]), .Z(n15687) );
  NAND U23689 ( .A(n21523), .B(n[833]), .Z(n22473) );
  XNOR U23690 ( .A(n22474), .B(n22471), .Z(n15688) );
  XOR U23691 ( .A(n22475), .B(n22476), .Z(n22471) );
  AND U23692 ( .A(n15695), .B(n22477), .Z(n22475) );
  XNOR U23693 ( .A(n15694), .B(n22476), .Z(n22477) );
  NAND U23694 ( .A(n22478), .B(n[832]), .Z(n15694) );
  NAND U23695 ( .A(n21523), .B(n[832]), .Z(n22478) );
  XNOR U23696 ( .A(n22479), .B(n22476), .Z(n15695) );
  XOR U23697 ( .A(n22480), .B(n22481), .Z(n22476) );
  AND U23698 ( .A(n15702), .B(n22482), .Z(n22480) );
  XNOR U23699 ( .A(n15701), .B(n22481), .Z(n22482) );
  NAND U23700 ( .A(n22483), .B(n[831]), .Z(n15701) );
  NAND U23701 ( .A(n21523), .B(n[831]), .Z(n22483) );
  XNOR U23702 ( .A(n22484), .B(n22481), .Z(n15702) );
  XOR U23703 ( .A(n22485), .B(n22486), .Z(n22481) );
  AND U23704 ( .A(n15709), .B(n22487), .Z(n22485) );
  XNOR U23705 ( .A(n15708), .B(n22486), .Z(n22487) );
  NAND U23706 ( .A(n22488), .B(n[830]), .Z(n15708) );
  NAND U23707 ( .A(n21523), .B(n[830]), .Z(n22488) );
  XNOR U23708 ( .A(n22489), .B(n22486), .Z(n15709) );
  XOR U23709 ( .A(n22490), .B(n22491), .Z(n22486) );
  AND U23710 ( .A(n15716), .B(n22492), .Z(n22490) );
  XNOR U23711 ( .A(n15715), .B(n22491), .Z(n22492) );
  NAND U23712 ( .A(n22493), .B(n[829]), .Z(n15715) );
  NAND U23713 ( .A(n21523), .B(n[829]), .Z(n22493) );
  XNOR U23714 ( .A(n22494), .B(n22491), .Z(n15716) );
  XOR U23715 ( .A(n22495), .B(n22496), .Z(n22491) );
  AND U23716 ( .A(n15723), .B(n22497), .Z(n22495) );
  XNOR U23717 ( .A(n15722), .B(n22496), .Z(n22497) );
  NAND U23718 ( .A(n22498), .B(n[828]), .Z(n15722) );
  NAND U23719 ( .A(n21523), .B(n[828]), .Z(n22498) );
  XNOR U23720 ( .A(n22499), .B(n22496), .Z(n15723) );
  XOR U23721 ( .A(n22500), .B(n22501), .Z(n22496) );
  AND U23722 ( .A(n15730), .B(n22502), .Z(n22500) );
  XNOR U23723 ( .A(n15729), .B(n22501), .Z(n22502) );
  NAND U23724 ( .A(n22503), .B(n[827]), .Z(n15729) );
  NAND U23725 ( .A(n21523), .B(n[827]), .Z(n22503) );
  XNOR U23726 ( .A(n22504), .B(n22501), .Z(n15730) );
  XOR U23727 ( .A(n22505), .B(n22506), .Z(n22501) );
  AND U23728 ( .A(n15737), .B(n22507), .Z(n22505) );
  XNOR U23729 ( .A(n15736), .B(n22506), .Z(n22507) );
  NAND U23730 ( .A(n22508), .B(n[826]), .Z(n15736) );
  NAND U23731 ( .A(n21523), .B(n[826]), .Z(n22508) );
  XNOR U23732 ( .A(n22509), .B(n22506), .Z(n15737) );
  XOR U23733 ( .A(n22510), .B(n22511), .Z(n22506) );
  AND U23734 ( .A(n15744), .B(n22512), .Z(n22510) );
  XNOR U23735 ( .A(n15743), .B(n22511), .Z(n22512) );
  NAND U23736 ( .A(n22513), .B(n[825]), .Z(n15743) );
  NAND U23737 ( .A(n21523), .B(n[825]), .Z(n22513) );
  XNOR U23738 ( .A(n22514), .B(n22511), .Z(n15744) );
  XOR U23739 ( .A(n22515), .B(n22516), .Z(n22511) );
  AND U23740 ( .A(n15751), .B(n22517), .Z(n22515) );
  XNOR U23741 ( .A(n15750), .B(n22516), .Z(n22517) );
  NAND U23742 ( .A(n22518), .B(n[824]), .Z(n15750) );
  NAND U23743 ( .A(n21523), .B(n[824]), .Z(n22518) );
  XNOR U23744 ( .A(n22519), .B(n22516), .Z(n15751) );
  XOR U23745 ( .A(n22520), .B(n22521), .Z(n22516) );
  AND U23746 ( .A(n15758), .B(n22522), .Z(n22520) );
  XNOR U23747 ( .A(n15757), .B(n22521), .Z(n22522) );
  NAND U23748 ( .A(n22523), .B(n[823]), .Z(n15757) );
  NAND U23749 ( .A(n21523), .B(n[823]), .Z(n22523) );
  XNOR U23750 ( .A(n22524), .B(n22521), .Z(n15758) );
  XOR U23751 ( .A(n22525), .B(n22526), .Z(n22521) );
  AND U23752 ( .A(n15765), .B(n22527), .Z(n22525) );
  XNOR U23753 ( .A(n15764), .B(n22526), .Z(n22527) );
  NAND U23754 ( .A(n22528), .B(n[822]), .Z(n15764) );
  NAND U23755 ( .A(n21523), .B(n[822]), .Z(n22528) );
  XNOR U23756 ( .A(n22529), .B(n22526), .Z(n15765) );
  XOR U23757 ( .A(n22530), .B(n22531), .Z(n22526) );
  AND U23758 ( .A(n15772), .B(n22532), .Z(n22530) );
  XNOR U23759 ( .A(n15771), .B(n22531), .Z(n22532) );
  NAND U23760 ( .A(n22533), .B(n[821]), .Z(n15771) );
  NAND U23761 ( .A(n21523), .B(n[821]), .Z(n22533) );
  XNOR U23762 ( .A(n22534), .B(n22531), .Z(n15772) );
  XOR U23763 ( .A(n22535), .B(n22536), .Z(n22531) );
  AND U23764 ( .A(n15779), .B(n22537), .Z(n22535) );
  XNOR U23765 ( .A(n15778), .B(n22536), .Z(n22537) );
  NAND U23766 ( .A(n22538), .B(n[820]), .Z(n15778) );
  NAND U23767 ( .A(n21523), .B(n[820]), .Z(n22538) );
  XNOR U23768 ( .A(n22539), .B(n22536), .Z(n15779) );
  XOR U23769 ( .A(n22540), .B(n22541), .Z(n22536) );
  AND U23770 ( .A(n15786), .B(n22542), .Z(n22540) );
  XNOR U23771 ( .A(n15785), .B(n22541), .Z(n22542) );
  NAND U23772 ( .A(n22543), .B(n[819]), .Z(n15785) );
  NAND U23773 ( .A(n21523), .B(n[819]), .Z(n22543) );
  XNOR U23774 ( .A(n22544), .B(n22541), .Z(n15786) );
  XOR U23775 ( .A(n22545), .B(n22546), .Z(n22541) );
  AND U23776 ( .A(n15793), .B(n22547), .Z(n22545) );
  XNOR U23777 ( .A(n15792), .B(n22546), .Z(n22547) );
  NAND U23778 ( .A(n22548), .B(n[818]), .Z(n15792) );
  NAND U23779 ( .A(n21523), .B(n[818]), .Z(n22548) );
  XNOR U23780 ( .A(n22549), .B(n22546), .Z(n15793) );
  XOR U23781 ( .A(n22550), .B(n22551), .Z(n22546) );
  AND U23782 ( .A(n15800), .B(n22552), .Z(n22550) );
  XNOR U23783 ( .A(n15799), .B(n22551), .Z(n22552) );
  NAND U23784 ( .A(n22553), .B(n[817]), .Z(n15799) );
  NAND U23785 ( .A(n21523), .B(n[817]), .Z(n22553) );
  XNOR U23786 ( .A(n22554), .B(n22551), .Z(n15800) );
  XOR U23787 ( .A(n22555), .B(n22556), .Z(n22551) );
  AND U23788 ( .A(n15807), .B(n22557), .Z(n22555) );
  XNOR U23789 ( .A(n15806), .B(n22556), .Z(n22557) );
  NAND U23790 ( .A(n22558), .B(n[816]), .Z(n15806) );
  NAND U23791 ( .A(n21523), .B(n[816]), .Z(n22558) );
  XNOR U23792 ( .A(n22559), .B(n22556), .Z(n15807) );
  XOR U23793 ( .A(n22560), .B(n22561), .Z(n22556) );
  AND U23794 ( .A(n15814), .B(n22562), .Z(n22560) );
  XNOR U23795 ( .A(n15813), .B(n22561), .Z(n22562) );
  NAND U23796 ( .A(n22563), .B(n[815]), .Z(n15813) );
  NAND U23797 ( .A(n21523), .B(n[815]), .Z(n22563) );
  XNOR U23798 ( .A(n22564), .B(n22561), .Z(n15814) );
  XOR U23799 ( .A(n22565), .B(n22566), .Z(n22561) );
  AND U23800 ( .A(n15821), .B(n22567), .Z(n22565) );
  XNOR U23801 ( .A(n15820), .B(n22566), .Z(n22567) );
  NAND U23802 ( .A(n22568), .B(n[814]), .Z(n15820) );
  NAND U23803 ( .A(n21523), .B(n[814]), .Z(n22568) );
  XNOR U23804 ( .A(n22569), .B(n22566), .Z(n15821) );
  XOR U23805 ( .A(n22570), .B(n22571), .Z(n22566) );
  AND U23806 ( .A(n15828), .B(n22572), .Z(n22570) );
  XNOR U23807 ( .A(n15827), .B(n22571), .Z(n22572) );
  NAND U23808 ( .A(n22573), .B(n[813]), .Z(n15827) );
  NAND U23809 ( .A(n21523), .B(n[813]), .Z(n22573) );
  XNOR U23810 ( .A(n22574), .B(n22571), .Z(n15828) );
  XOR U23811 ( .A(n22575), .B(n22576), .Z(n22571) );
  AND U23812 ( .A(n15835), .B(n22577), .Z(n22575) );
  XNOR U23813 ( .A(n15834), .B(n22576), .Z(n22577) );
  NAND U23814 ( .A(n22578), .B(n[812]), .Z(n15834) );
  NAND U23815 ( .A(n21523), .B(n[812]), .Z(n22578) );
  XNOR U23816 ( .A(n22579), .B(n22576), .Z(n15835) );
  XOR U23817 ( .A(n22580), .B(n22581), .Z(n22576) );
  AND U23818 ( .A(n15842), .B(n22582), .Z(n22580) );
  XNOR U23819 ( .A(n15841), .B(n22581), .Z(n22582) );
  NAND U23820 ( .A(n22583), .B(n[811]), .Z(n15841) );
  NAND U23821 ( .A(n21523), .B(n[811]), .Z(n22583) );
  XNOR U23822 ( .A(n22584), .B(n22581), .Z(n15842) );
  XOR U23823 ( .A(n22585), .B(n22586), .Z(n22581) );
  AND U23824 ( .A(n15849), .B(n22587), .Z(n22585) );
  XNOR U23825 ( .A(n15848), .B(n22586), .Z(n22587) );
  NAND U23826 ( .A(n22588), .B(n[810]), .Z(n15848) );
  NAND U23827 ( .A(n21523), .B(n[810]), .Z(n22588) );
  XNOR U23828 ( .A(n22589), .B(n22586), .Z(n15849) );
  XOR U23829 ( .A(n22590), .B(n22591), .Z(n22586) );
  AND U23830 ( .A(n15856), .B(n22592), .Z(n22590) );
  XNOR U23831 ( .A(n15855), .B(n22591), .Z(n22592) );
  NAND U23832 ( .A(n22593), .B(n[809]), .Z(n15855) );
  NAND U23833 ( .A(n21523), .B(n[809]), .Z(n22593) );
  XNOR U23834 ( .A(n22594), .B(n22591), .Z(n15856) );
  XOR U23835 ( .A(n22595), .B(n22596), .Z(n22591) );
  AND U23836 ( .A(n15863), .B(n22597), .Z(n22595) );
  XNOR U23837 ( .A(n15862), .B(n22596), .Z(n22597) );
  NAND U23838 ( .A(n22598), .B(n[808]), .Z(n15862) );
  NAND U23839 ( .A(n21523), .B(n[808]), .Z(n22598) );
  XNOR U23840 ( .A(n22599), .B(n22596), .Z(n15863) );
  XOR U23841 ( .A(n22600), .B(n22601), .Z(n22596) );
  AND U23842 ( .A(n15870), .B(n22602), .Z(n22600) );
  XNOR U23843 ( .A(n15869), .B(n22601), .Z(n22602) );
  NAND U23844 ( .A(n22603), .B(n[807]), .Z(n15869) );
  NAND U23845 ( .A(n21523), .B(n[807]), .Z(n22603) );
  XNOR U23846 ( .A(n22604), .B(n22601), .Z(n15870) );
  XOR U23847 ( .A(n22605), .B(n22606), .Z(n22601) );
  AND U23848 ( .A(n15877), .B(n22607), .Z(n22605) );
  XNOR U23849 ( .A(n15876), .B(n22606), .Z(n22607) );
  NAND U23850 ( .A(n22608), .B(n[806]), .Z(n15876) );
  NAND U23851 ( .A(n21523), .B(n[806]), .Z(n22608) );
  XNOR U23852 ( .A(n22609), .B(n22606), .Z(n15877) );
  XOR U23853 ( .A(n22610), .B(n22611), .Z(n22606) );
  AND U23854 ( .A(n15884), .B(n22612), .Z(n22610) );
  XNOR U23855 ( .A(n15883), .B(n22611), .Z(n22612) );
  NAND U23856 ( .A(n22613), .B(n[805]), .Z(n15883) );
  NAND U23857 ( .A(n21523), .B(n[805]), .Z(n22613) );
  XNOR U23858 ( .A(n22614), .B(n22611), .Z(n15884) );
  XOR U23859 ( .A(n22615), .B(n22616), .Z(n22611) );
  AND U23860 ( .A(n15891), .B(n22617), .Z(n22615) );
  XNOR U23861 ( .A(n15890), .B(n22616), .Z(n22617) );
  NAND U23862 ( .A(n22618), .B(n[804]), .Z(n15890) );
  NAND U23863 ( .A(n21523), .B(n[804]), .Z(n22618) );
  XNOR U23864 ( .A(n22619), .B(n22616), .Z(n15891) );
  XOR U23865 ( .A(n22620), .B(n22621), .Z(n22616) );
  AND U23866 ( .A(n15898), .B(n22622), .Z(n22620) );
  XNOR U23867 ( .A(n15897), .B(n22621), .Z(n22622) );
  NAND U23868 ( .A(n22623), .B(n[803]), .Z(n15897) );
  NAND U23869 ( .A(n21523), .B(n[803]), .Z(n22623) );
  XNOR U23870 ( .A(n22624), .B(n22621), .Z(n15898) );
  XOR U23871 ( .A(n22625), .B(n22626), .Z(n22621) );
  AND U23872 ( .A(n15905), .B(n22627), .Z(n22625) );
  XNOR U23873 ( .A(n15904), .B(n22626), .Z(n22627) );
  NAND U23874 ( .A(n22628), .B(n[802]), .Z(n15904) );
  NAND U23875 ( .A(n21523), .B(n[802]), .Z(n22628) );
  XNOR U23876 ( .A(n22629), .B(n22626), .Z(n15905) );
  XOR U23877 ( .A(n22630), .B(n22631), .Z(n22626) );
  AND U23878 ( .A(n15912), .B(n22632), .Z(n22630) );
  XNOR U23879 ( .A(n15911), .B(n22631), .Z(n22632) );
  NAND U23880 ( .A(n22633), .B(n[801]), .Z(n15911) );
  NAND U23881 ( .A(n21523), .B(n[801]), .Z(n22633) );
  XNOR U23882 ( .A(n22634), .B(n22631), .Z(n15912) );
  XOR U23883 ( .A(n22635), .B(n22636), .Z(n22631) );
  AND U23884 ( .A(n15919), .B(n22637), .Z(n22635) );
  XNOR U23885 ( .A(n15918), .B(n22636), .Z(n22637) );
  NAND U23886 ( .A(n22638), .B(n[800]), .Z(n15918) );
  NAND U23887 ( .A(n21523), .B(n[800]), .Z(n22638) );
  XNOR U23888 ( .A(n22639), .B(n22636), .Z(n15919) );
  XOR U23889 ( .A(n22640), .B(n22641), .Z(n22636) );
  AND U23890 ( .A(n15926), .B(n22642), .Z(n22640) );
  XNOR U23891 ( .A(n15925), .B(n22641), .Z(n22642) );
  NAND U23892 ( .A(n22643), .B(n[799]), .Z(n15925) );
  NAND U23893 ( .A(n21523), .B(n[799]), .Z(n22643) );
  XNOR U23894 ( .A(n22644), .B(n22641), .Z(n15926) );
  XOR U23895 ( .A(n22645), .B(n22646), .Z(n22641) );
  AND U23896 ( .A(n15933), .B(n22647), .Z(n22645) );
  XNOR U23897 ( .A(n15932), .B(n22646), .Z(n22647) );
  NAND U23898 ( .A(n22648), .B(n[798]), .Z(n15932) );
  NAND U23899 ( .A(n21523), .B(n[798]), .Z(n22648) );
  XNOR U23900 ( .A(n22649), .B(n22646), .Z(n15933) );
  XOR U23901 ( .A(n22650), .B(n22651), .Z(n22646) );
  AND U23902 ( .A(n15940), .B(n22652), .Z(n22650) );
  XNOR U23903 ( .A(n15939), .B(n22651), .Z(n22652) );
  NAND U23904 ( .A(n22653), .B(n[797]), .Z(n15939) );
  NAND U23905 ( .A(n21523), .B(n[797]), .Z(n22653) );
  XNOR U23906 ( .A(n22654), .B(n22651), .Z(n15940) );
  XOR U23907 ( .A(n22655), .B(n22656), .Z(n22651) );
  AND U23908 ( .A(n15947), .B(n22657), .Z(n22655) );
  XNOR U23909 ( .A(n15946), .B(n22656), .Z(n22657) );
  NAND U23910 ( .A(n22658), .B(n[796]), .Z(n15946) );
  NAND U23911 ( .A(n21523), .B(n[796]), .Z(n22658) );
  XNOR U23912 ( .A(n22659), .B(n22656), .Z(n15947) );
  XOR U23913 ( .A(n22660), .B(n22661), .Z(n22656) );
  AND U23914 ( .A(n15954), .B(n22662), .Z(n22660) );
  XNOR U23915 ( .A(n15953), .B(n22661), .Z(n22662) );
  NAND U23916 ( .A(n22663), .B(n[795]), .Z(n15953) );
  NAND U23917 ( .A(n21523), .B(n[795]), .Z(n22663) );
  XNOR U23918 ( .A(n22664), .B(n22661), .Z(n15954) );
  XOR U23919 ( .A(n22665), .B(n22666), .Z(n22661) );
  AND U23920 ( .A(n15961), .B(n22667), .Z(n22665) );
  XNOR U23921 ( .A(n15960), .B(n22666), .Z(n22667) );
  NAND U23922 ( .A(n22668), .B(n[794]), .Z(n15960) );
  NAND U23923 ( .A(n21523), .B(n[794]), .Z(n22668) );
  XNOR U23924 ( .A(n22669), .B(n22666), .Z(n15961) );
  XOR U23925 ( .A(n22670), .B(n22671), .Z(n22666) );
  AND U23926 ( .A(n15968), .B(n22672), .Z(n22670) );
  XNOR U23927 ( .A(n15967), .B(n22671), .Z(n22672) );
  NAND U23928 ( .A(n22673), .B(n[793]), .Z(n15967) );
  NAND U23929 ( .A(n21523), .B(n[793]), .Z(n22673) );
  XNOR U23930 ( .A(n22674), .B(n22671), .Z(n15968) );
  XOR U23931 ( .A(n22675), .B(n22676), .Z(n22671) );
  AND U23932 ( .A(n15975), .B(n22677), .Z(n22675) );
  XNOR U23933 ( .A(n15974), .B(n22676), .Z(n22677) );
  NAND U23934 ( .A(n22678), .B(n[792]), .Z(n15974) );
  NAND U23935 ( .A(n21523), .B(n[792]), .Z(n22678) );
  XNOR U23936 ( .A(n22679), .B(n22676), .Z(n15975) );
  XOR U23937 ( .A(n22680), .B(n22681), .Z(n22676) );
  AND U23938 ( .A(n15982), .B(n22682), .Z(n22680) );
  XNOR U23939 ( .A(n15981), .B(n22681), .Z(n22682) );
  NAND U23940 ( .A(n22683), .B(n[791]), .Z(n15981) );
  NAND U23941 ( .A(n21523), .B(n[791]), .Z(n22683) );
  XNOR U23942 ( .A(n22684), .B(n22681), .Z(n15982) );
  XOR U23943 ( .A(n22685), .B(n22686), .Z(n22681) );
  AND U23944 ( .A(n15989), .B(n22687), .Z(n22685) );
  XNOR U23945 ( .A(n15988), .B(n22686), .Z(n22687) );
  NAND U23946 ( .A(n22688), .B(n[790]), .Z(n15988) );
  NAND U23947 ( .A(n21523), .B(n[790]), .Z(n22688) );
  XNOR U23948 ( .A(n22689), .B(n22686), .Z(n15989) );
  XOR U23949 ( .A(n22690), .B(n22691), .Z(n22686) );
  AND U23950 ( .A(n15996), .B(n22692), .Z(n22690) );
  XNOR U23951 ( .A(n15995), .B(n22691), .Z(n22692) );
  NAND U23952 ( .A(n22693), .B(n[789]), .Z(n15995) );
  NAND U23953 ( .A(n21523), .B(n[789]), .Z(n22693) );
  XNOR U23954 ( .A(n22694), .B(n22691), .Z(n15996) );
  XOR U23955 ( .A(n22695), .B(n22696), .Z(n22691) );
  AND U23956 ( .A(n16003), .B(n22697), .Z(n22695) );
  XNOR U23957 ( .A(n16002), .B(n22696), .Z(n22697) );
  NAND U23958 ( .A(n22698), .B(n[788]), .Z(n16002) );
  NAND U23959 ( .A(n21523), .B(n[788]), .Z(n22698) );
  XNOR U23960 ( .A(n22699), .B(n22696), .Z(n16003) );
  XOR U23961 ( .A(n22700), .B(n22701), .Z(n22696) );
  AND U23962 ( .A(n16010), .B(n22702), .Z(n22700) );
  XNOR U23963 ( .A(n16009), .B(n22701), .Z(n22702) );
  NAND U23964 ( .A(n22703), .B(n[787]), .Z(n16009) );
  NAND U23965 ( .A(n21523), .B(n[787]), .Z(n22703) );
  XNOR U23966 ( .A(n22704), .B(n22701), .Z(n16010) );
  XOR U23967 ( .A(n22705), .B(n22706), .Z(n22701) );
  AND U23968 ( .A(n16017), .B(n22707), .Z(n22705) );
  XNOR U23969 ( .A(n16016), .B(n22706), .Z(n22707) );
  NAND U23970 ( .A(n22708), .B(n[786]), .Z(n16016) );
  NAND U23971 ( .A(n21523), .B(n[786]), .Z(n22708) );
  XNOR U23972 ( .A(n22709), .B(n22706), .Z(n16017) );
  XOR U23973 ( .A(n22710), .B(n22711), .Z(n22706) );
  AND U23974 ( .A(n16024), .B(n22712), .Z(n22710) );
  XNOR U23975 ( .A(n16023), .B(n22711), .Z(n22712) );
  NAND U23976 ( .A(n22713), .B(n[785]), .Z(n16023) );
  NAND U23977 ( .A(n21523), .B(n[785]), .Z(n22713) );
  XNOR U23978 ( .A(n22714), .B(n22711), .Z(n16024) );
  XOR U23979 ( .A(n22715), .B(n22716), .Z(n22711) );
  AND U23980 ( .A(n16031), .B(n22717), .Z(n22715) );
  XNOR U23981 ( .A(n16030), .B(n22716), .Z(n22717) );
  NAND U23982 ( .A(n22718), .B(n[784]), .Z(n16030) );
  NAND U23983 ( .A(n21523), .B(n[784]), .Z(n22718) );
  XNOR U23984 ( .A(n22719), .B(n22716), .Z(n16031) );
  XOR U23985 ( .A(n22720), .B(n22721), .Z(n22716) );
  AND U23986 ( .A(n16038), .B(n22722), .Z(n22720) );
  XNOR U23987 ( .A(n16037), .B(n22721), .Z(n22722) );
  NAND U23988 ( .A(n22723), .B(n[783]), .Z(n16037) );
  NAND U23989 ( .A(n21523), .B(n[783]), .Z(n22723) );
  XNOR U23990 ( .A(n22724), .B(n22721), .Z(n16038) );
  XOR U23991 ( .A(n22725), .B(n22726), .Z(n22721) );
  AND U23992 ( .A(n16045), .B(n22727), .Z(n22725) );
  XNOR U23993 ( .A(n16044), .B(n22726), .Z(n22727) );
  NAND U23994 ( .A(n22728), .B(n[782]), .Z(n16044) );
  NAND U23995 ( .A(n21523), .B(n[782]), .Z(n22728) );
  XNOR U23996 ( .A(n22729), .B(n22726), .Z(n16045) );
  XOR U23997 ( .A(n22730), .B(n22731), .Z(n22726) );
  AND U23998 ( .A(n16052), .B(n22732), .Z(n22730) );
  XNOR U23999 ( .A(n16051), .B(n22731), .Z(n22732) );
  NAND U24000 ( .A(n22733), .B(n[781]), .Z(n16051) );
  NAND U24001 ( .A(n21523), .B(n[781]), .Z(n22733) );
  XNOR U24002 ( .A(n22734), .B(n22731), .Z(n16052) );
  XOR U24003 ( .A(n22735), .B(n22736), .Z(n22731) );
  AND U24004 ( .A(n16059), .B(n22737), .Z(n22735) );
  XNOR U24005 ( .A(n16058), .B(n22736), .Z(n22737) );
  NAND U24006 ( .A(n22738), .B(n[780]), .Z(n16058) );
  NAND U24007 ( .A(n21523), .B(n[780]), .Z(n22738) );
  XNOR U24008 ( .A(n22739), .B(n22736), .Z(n16059) );
  XOR U24009 ( .A(n22740), .B(n22741), .Z(n22736) );
  AND U24010 ( .A(n16066), .B(n22742), .Z(n22740) );
  XNOR U24011 ( .A(n16065), .B(n22741), .Z(n22742) );
  NAND U24012 ( .A(n22743), .B(n[779]), .Z(n16065) );
  NAND U24013 ( .A(n21523), .B(n[779]), .Z(n22743) );
  XNOR U24014 ( .A(n22744), .B(n22741), .Z(n16066) );
  XOR U24015 ( .A(n22745), .B(n22746), .Z(n22741) );
  AND U24016 ( .A(n16073), .B(n22747), .Z(n22745) );
  XNOR U24017 ( .A(n16072), .B(n22746), .Z(n22747) );
  NAND U24018 ( .A(n22748), .B(n[778]), .Z(n16072) );
  NAND U24019 ( .A(n21523), .B(n[778]), .Z(n22748) );
  XNOR U24020 ( .A(n22749), .B(n22746), .Z(n16073) );
  XOR U24021 ( .A(n22750), .B(n22751), .Z(n22746) );
  AND U24022 ( .A(n16080), .B(n22752), .Z(n22750) );
  XNOR U24023 ( .A(n16079), .B(n22751), .Z(n22752) );
  NAND U24024 ( .A(n22753), .B(n[777]), .Z(n16079) );
  NAND U24025 ( .A(n21523), .B(n[777]), .Z(n22753) );
  XNOR U24026 ( .A(n22754), .B(n22751), .Z(n16080) );
  XOR U24027 ( .A(n22755), .B(n22756), .Z(n22751) );
  AND U24028 ( .A(n16087), .B(n22757), .Z(n22755) );
  XNOR U24029 ( .A(n16086), .B(n22756), .Z(n22757) );
  NAND U24030 ( .A(n22758), .B(n[776]), .Z(n16086) );
  NAND U24031 ( .A(n21523), .B(n[776]), .Z(n22758) );
  XNOR U24032 ( .A(n22759), .B(n22756), .Z(n16087) );
  XOR U24033 ( .A(n22760), .B(n22761), .Z(n22756) );
  AND U24034 ( .A(n16094), .B(n22762), .Z(n22760) );
  XNOR U24035 ( .A(n16093), .B(n22761), .Z(n22762) );
  NAND U24036 ( .A(n22763), .B(n[775]), .Z(n16093) );
  NAND U24037 ( .A(n21523), .B(n[775]), .Z(n22763) );
  XNOR U24038 ( .A(n22764), .B(n22761), .Z(n16094) );
  XOR U24039 ( .A(n22765), .B(n22766), .Z(n22761) );
  AND U24040 ( .A(n16101), .B(n22767), .Z(n22765) );
  XNOR U24041 ( .A(n16100), .B(n22766), .Z(n22767) );
  NAND U24042 ( .A(n22768), .B(n[774]), .Z(n16100) );
  NAND U24043 ( .A(n21523), .B(n[774]), .Z(n22768) );
  XNOR U24044 ( .A(n22769), .B(n22766), .Z(n16101) );
  XOR U24045 ( .A(n22770), .B(n22771), .Z(n22766) );
  AND U24046 ( .A(n16108), .B(n22772), .Z(n22770) );
  XNOR U24047 ( .A(n16107), .B(n22771), .Z(n22772) );
  NAND U24048 ( .A(n22773), .B(n[773]), .Z(n16107) );
  NAND U24049 ( .A(n21523), .B(n[773]), .Z(n22773) );
  XNOR U24050 ( .A(n22774), .B(n22771), .Z(n16108) );
  XOR U24051 ( .A(n22775), .B(n22776), .Z(n22771) );
  AND U24052 ( .A(n16115), .B(n22777), .Z(n22775) );
  XNOR U24053 ( .A(n16114), .B(n22776), .Z(n22777) );
  NAND U24054 ( .A(n22778), .B(n[772]), .Z(n16114) );
  NAND U24055 ( .A(n21523), .B(n[772]), .Z(n22778) );
  XNOR U24056 ( .A(n22779), .B(n22776), .Z(n16115) );
  XOR U24057 ( .A(n22780), .B(n22781), .Z(n22776) );
  AND U24058 ( .A(n16122), .B(n22782), .Z(n22780) );
  XNOR U24059 ( .A(n16121), .B(n22781), .Z(n22782) );
  NAND U24060 ( .A(n22783), .B(n[771]), .Z(n16121) );
  NAND U24061 ( .A(n21523), .B(n[771]), .Z(n22783) );
  XNOR U24062 ( .A(n22784), .B(n22781), .Z(n16122) );
  XOR U24063 ( .A(n22785), .B(n22786), .Z(n22781) );
  AND U24064 ( .A(n16129), .B(n22787), .Z(n22785) );
  XNOR U24065 ( .A(n16128), .B(n22786), .Z(n22787) );
  NAND U24066 ( .A(n22788), .B(n[770]), .Z(n16128) );
  NAND U24067 ( .A(n21523), .B(n[770]), .Z(n22788) );
  XNOR U24068 ( .A(n22789), .B(n22786), .Z(n16129) );
  XOR U24069 ( .A(n22790), .B(n22791), .Z(n22786) );
  AND U24070 ( .A(n16136), .B(n22792), .Z(n22790) );
  XNOR U24071 ( .A(n16135), .B(n22791), .Z(n22792) );
  NAND U24072 ( .A(n22793), .B(n[769]), .Z(n16135) );
  NAND U24073 ( .A(n21523), .B(n[769]), .Z(n22793) );
  XNOR U24074 ( .A(n22794), .B(n22791), .Z(n16136) );
  XOR U24075 ( .A(n22795), .B(n22796), .Z(n22791) );
  AND U24076 ( .A(n16143), .B(n22797), .Z(n22795) );
  XNOR U24077 ( .A(n16142), .B(n22796), .Z(n22797) );
  NAND U24078 ( .A(n22798), .B(n[768]), .Z(n16142) );
  NAND U24079 ( .A(n21523), .B(n[768]), .Z(n22798) );
  XNOR U24080 ( .A(n22799), .B(n22796), .Z(n16143) );
  XOR U24081 ( .A(n22800), .B(n22801), .Z(n22796) );
  AND U24082 ( .A(n16150), .B(n22802), .Z(n22800) );
  XNOR U24083 ( .A(n16149), .B(n22801), .Z(n22802) );
  NAND U24084 ( .A(n22803), .B(n[767]), .Z(n16149) );
  NAND U24085 ( .A(n21523), .B(n[767]), .Z(n22803) );
  XNOR U24086 ( .A(n22804), .B(n22801), .Z(n16150) );
  XOR U24087 ( .A(n22805), .B(n22806), .Z(n22801) );
  AND U24088 ( .A(n16157), .B(n22807), .Z(n22805) );
  XNOR U24089 ( .A(n16156), .B(n22806), .Z(n22807) );
  NAND U24090 ( .A(n22808), .B(n[766]), .Z(n16156) );
  NAND U24091 ( .A(n21523), .B(n[766]), .Z(n22808) );
  XNOR U24092 ( .A(n22809), .B(n22806), .Z(n16157) );
  XOR U24093 ( .A(n22810), .B(n22811), .Z(n22806) );
  AND U24094 ( .A(n16164), .B(n22812), .Z(n22810) );
  XNOR U24095 ( .A(n16163), .B(n22811), .Z(n22812) );
  NAND U24096 ( .A(n22813), .B(n[765]), .Z(n16163) );
  NAND U24097 ( .A(n21523), .B(n[765]), .Z(n22813) );
  XNOR U24098 ( .A(n22814), .B(n22811), .Z(n16164) );
  XOR U24099 ( .A(n22815), .B(n22816), .Z(n22811) );
  AND U24100 ( .A(n16171), .B(n22817), .Z(n22815) );
  XNOR U24101 ( .A(n16170), .B(n22816), .Z(n22817) );
  NAND U24102 ( .A(n22818), .B(n[764]), .Z(n16170) );
  NAND U24103 ( .A(n21523), .B(n[764]), .Z(n22818) );
  XNOR U24104 ( .A(n22819), .B(n22816), .Z(n16171) );
  XOR U24105 ( .A(n22820), .B(n22821), .Z(n22816) );
  AND U24106 ( .A(n16178), .B(n22822), .Z(n22820) );
  XNOR U24107 ( .A(n16177), .B(n22821), .Z(n22822) );
  NAND U24108 ( .A(n22823), .B(n[763]), .Z(n16177) );
  NAND U24109 ( .A(n21523), .B(n[763]), .Z(n22823) );
  XNOR U24110 ( .A(n22824), .B(n22821), .Z(n16178) );
  XOR U24111 ( .A(n22825), .B(n22826), .Z(n22821) );
  AND U24112 ( .A(n16185), .B(n22827), .Z(n22825) );
  XNOR U24113 ( .A(n16184), .B(n22826), .Z(n22827) );
  NAND U24114 ( .A(n22828), .B(n[762]), .Z(n16184) );
  NAND U24115 ( .A(n21523), .B(n[762]), .Z(n22828) );
  XNOR U24116 ( .A(n22829), .B(n22826), .Z(n16185) );
  XOR U24117 ( .A(n22830), .B(n22831), .Z(n22826) );
  AND U24118 ( .A(n16192), .B(n22832), .Z(n22830) );
  XNOR U24119 ( .A(n16191), .B(n22831), .Z(n22832) );
  NAND U24120 ( .A(n22833), .B(n[761]), .Z(n16191) );
  NAND U24121 ( .A(n21523), .B(n[761]), .Z(n22833) );
  XNOR U24122 ( .A(n22834), .B(n22831), .Z(n16192) );
  XOR U24123 ( .A(n22835), .B(n22836), .Z(n22831) );
  AND U24124 ( .A(n16199), .B(n22837), .Z(n22835) );
  XNOR U24125 ( .A(n16198), .B(n22836), .Z(n22837) );
  NAND U24126 ( .A(n22838), .B(n[760]), .Z(n16198) );
  NAND U24127 ( .A(n21523), .B(n[760]), .Z(n22838) );
  XNOR U24128 ( .A(n22839), .B(n22836), .Z(n16199) );
  XOR U24129 ( .A(n22840), .B(n22841), .Z(n22836) );
  AND U24130 ( .A(n16206), .B(n22842), .Z(n22840) );
  XNOR U24131 ( .A(n16205), .B(n22841), .Z(n22842) );
  NAND U24132 ( .A(n22843), .B(n[759]), .Z(n16205) );
  NAND U24133 ( .A(n21523), .B(n[759]), .Z(n22843) );
  XNOR U24134 ( .A(n22844), .B(n22841), .Z(n16206) );
  XOR U24135 ( .A(n22845), .B(n22846), .Z(n22841) );
  AND U24136 ( .A(n16213), .B(n22847), .Z(n22845) );
  XNOR U24137 ( .A(n16212), .B(n22846), .Z(n22847) );
  NAND U24138 ( .A(n22848), .B(n[758]), .Z(n16212) );
  NAND U24139 ( .A(n21523), .B(n[758]), .Z(n22848) );
  XNOR U24140 ( .A(n22849), .B(n22846), .Z(n16213) );
  XOR U24141 ( .A(n22850), .B(n22851), .Z(n22846) );
  AND U24142 ( .A(n16220), .B(n22852), .Z(n22850) );
  XNOR U24143 ( .A(n16219), .B(n22851), .Z(n22852) );
  NAND U24144 ( .A(n22853), .B(n[757]), .Z(n16219) );
  NAND U24145 ( .A(n21523), .B(n[757]), .Z(n22853) );
  XNOR U24146 ( .A(n22854), .B(n22851), .Z(n16220) );
  XOR U24147 ( .A(n22855), .B(n22856), .Z(n22851) );
  AND U24148 ( .A(n16227), .B(n22857), .Z(n22855) );
  XNOR U24149 ( .A(n16226), .B(n22856), .Z(n22857) );
  NAND U24150 ( .A(n22858), .B(n[756]), .Z(n16226) );
  NAND U24151 ( .A(n21523), .B(n[756]), .Z(n22858) );
  XNOR U24152 ( .A(n22859), .B(n22856), .Z(n16227) );
  XOR U24153 ( .A(n22860), .B(n22861), .Z(n22856) );
  AND U24154 ( .A(n16234), .B(n22862), .Z(n22860) );
  XNOR U24155 ( .A(n16233), .B(n22861), .Z(n22862) );
  NAND U24156 ( .A(n22863), .B(n[755]), .Z(n16233) );
  NAND U24157 ( .A(n21523), .B(n[755]), .Z(n22863) );
  XNOR U24158 ( .A(n22864), .B(n22861), .Z(n16234) );
  XOR U24159 ( .A(n22865), .B(n22866), .Z(n22861) );
  AND U24160 ( .A(n16241), .B(n22867), .Z(n22865) );
  XNOR U24161 ( .A(n16240), .B(n22866), .Z(n22867) );
  NAND U24162 ( .A(n22868), .B(n[754]), .Z(n16240) );
  NAND U24163 ( .A(n21523), .B(n[754]), .Z(n22868) );
  XNOR U24164 ( .A(n22869), .B(n22866), .Z(n16241) );
  XOR U24165 ( .A(n22870), .B(n22871), .Z(n22866) );
  AND U24166 ( .A(n16248), .B(n22872), .Z(n22870) );
  XNOR U24167 ( .A(n16247), .B(n22871), .Z(n22872) );
  NAND U24168 ( .A(n22873), .B(n[753]), .Z(n16247) );
  NAND U24169 ( .A(n21523), .B(n[753]), .Z(n22873) );
  XNOR U24170 ( .A(n22874), .B(n22871), .Z(n16248) );
  XOR U24171 ( .A(n22875), .B(n22876), .Z(n22871) );
  AND U24172 ( .A(n16255), .B(n22877), .Z(n22875) );
  XNOR U24173 ( .A(n16254), .B(n22876), .Z(n22877) );
  NAND U24174 ( .A(n22878), .B(n[752]), .Z(n16254) );
  NAND U24175 ( .A(n21523), .B(n[752]), .Z(n22878) );
  XNOR U24176 ( .A(n22879), .B(n22876), .Z(n16255) );
  XOR U24177 ( .A(n22880), .B(n22881), .Z(n22876) );
  AND U24178 ( .A(n16262), .B(n22882), .Z(n22880) );
  XNOR U24179 ( .A(n16261), .B(n22881), .Z(n22882) );
  NAND U24180 ( .A(n22883), .B(n[751]), .Z(n16261) );
  NAND U24181 ( .A(n21523), .B(n[751]), .Z(n22883) );
  XNOR U24182 ( .A(n22884), .B(n22881), .Z(n16262) );
  XOR U24183 ( .A(n22885), .B(n22886), .Z(n22881) );
  AND U24184 ( .A(n16269), .B(n22887), .Z(n22885) );
  XNOR U24185 ( .A(n16268), .B(n22886), .Z(n22887) );
  NAND U24186 ( .A(n22888), .B(n[750]), .Z(n16268) );
  NAND U24187 ( .A(n21523), .B(n[750]), .Z(n22888) );
  XNOR U24188 ( .A(n22889), .B(n22886), .Z(n16269) );
  XOR U24189 ( .A(n22890), .B(n22891), .Z(n22886) );
  AND U24190 ( .A(n16276), .B(n22892), .Z(n22890) );
  XNOR U24191 ( .A(n16275), .B(n22891), .Z(n22892) );
  NAND U24192 ( .A(n22893), .B(n[749]), .Z(n16275) );
  NAND U24193 ( .A(n21523), .B(n[749]), .Z(n22893) );
  XNOR U24194 ( .A(n22894), .B(n22891), .Z(n16276) );
  XOR U24195 ( .A(n22895), .B(n22896), .Z(n22891) );
  AND U24196 ( .A(n16283), .B(n22897), .Z(n22895) );
  XNOR U24197 ( .A(n16282), .B(n22896), .Z(n22897) );
  NAND U24198 ( .A(n22898), .B(n[748]), .Z(n16282) );
  NAND U24199 ( .A(n21523), .B(n[748]), .Z(n22898) );
  XNOR U24200 ( .A(n22899), .B(n22896), .Z(n16283) );
  XOR U24201 ( .A(n22900), .B(n22901), .Z(n22896) );
  AND U24202 ( .A(n16290), .B(n22902), .Z(n22900) );
  XNOR U24203 ( .A(n16289), .B(n22901), .Z(n22902) );
  NAND U24204 ( .A(n22903), .B(n[747]), .Z(n16289) );
  NAND U24205 ( .A(n21523), .B(n[747]), .Z(n22903) );
  XNOR U24206 ( .A(n22904), .B(n22901), .Z(n16290) );
  XOR U24207 ( .A(n22905), .B(n22906), .Z(n22901) );
  AND U24208 ( .A(n16297), .B(n22907), .Z(n22905) );
  XNOR U24209 ( .A(n16296), .B(n22906), .Z(n22907) );
  NAND U24210 ( .A(n22908), .B(n[746]), .Z(n16296) );
  NAND U24211 ( .A(n21523), .B(n[746]), .Z(n22908) );
  XNOR U24212 ( .A(n22909), .B(n22906), .Z(n16297) );
  XOR U24213 ( .A(n22910), .B(n22911), .Z(n22906) );
  AND U24214 ( .A(n16304), .B(n22912), .Z(n22910) );
  XNOR U24215 ( .A(n16303), .B(n22911), .Z(n22912) );
  NAND U24216 ( .A(n22913), .B(n[745]), .Z(n16303) );
  NAND U24217 ( .A(n21523), .B(n[745]), .Z(n22913) );
  XNOR U24218 ( .A(n22914), .B(n22911), .Z(n16304) );
  XOR U24219 ( .A(n22915), .B(n22916), .Z(n22911) );
  AND U24220 ( .A(n16311), .B(n22917), .Z(n22915) );
  XNOR U24221 ( .A(n16310), .B(n22916), .Z(n22917) );
  NAND U24222 ( .A(n22918), .B(n[744]), .Z(n16310) );
  NAND U24223 ( .A(n21523), .B(n[744]), .Z(n22918) );
  XNOR U24224 ( .A(n22919), .B(n22916), .Z(n16311) );
  XOR U24225 ( .A(n22920), .B(n22921), .Z(n22916) );
  AND U24226 ( .A(n16318), .B(n22922), .Z(n22920) );
  XNOR U24227 ( .A(n16317), .B(n22921), .Z(n22922) );
  NAND U24228 ( .A(n22923), .B(n[743]), .Z(n16317) );
  NAND U24229 ( .A(n21523), .B(n[743]), .Z(n22923) );
  XNOR U24230 ( .A(n22924), .B(n22921), .Z(n16318) );
  XOR U24231 ( .A(n22925), .B(n22926), .Z(n22921) );
  AND U24232 ( .A(n16325), .B(n22927), .Z(n22925) );
  XNOR U24233 ( .A(n16324), .B(n22926), .Z(n22927) );
  NAND U24234 ( .A(n22928), .B(n[742]), .Z(n16324) );
  NAND U24235 ( .A(n21523), .B(n[742]), .Z(n22928) );
  XNOR U24236 ( .A(n22929), .B(n22926), .Z(n16325) );
  XOR U24237 ( .A(n22930), .B(n22931), .Z(n22926) );
  AND U24238 ( .A(n16332), .B(n22932), .Z(n22930) );
  XNOR U24239 ( .A(n16331), .B(n22931), .Z(n22932) );
  NAND U24240 ( .A(n22933), .B(n[741]), .Z(n16331) );
  NAND U24241 ( .A(n21523), .B(n[741]), .Z(n22933) );
  XNOR U24242 ( .A(n22934), .B(n22931), .Z(n16332) );
  XOR U24243 ( .A(n22935), .B(n22936), .Z(n22931) );
  AND U24244 ( .A(n16339), .B(n22937), .Z(n22935) );
  XNOR U24245 ( .A(n16338), .B(n22936), .Z(n22937) );
  NAND U24246 ( .A(n22938), .B(n[740]), .Z(n16338) );
  NAND U24247 ( .A(n21523), .B(n[740]), .Z(n22938) );
  XNOR U24248 ( .A(n22939), .B(n22936), .Z(n16339) );
  XOR U24249 ( .A(n22940), .B(n22941), .Z(n22936) );
  AND U24250 ( .A(n16346), .B(n22942), .Z(n22940) );
  XNOR U24251 ( .A(n16345), .B(n22941), .Z(n22942) );
  NAND U24252 ( .A(n22943), .B(n[739]), .Z(n16345) );
  NAND U24253 ( .A(n21523), .B(n[739]), .Z(n22943) );
  XNOR U24254 ( .A(n22944), .B(n22941), .Z(n16346) );
  XOR U24255 ( .A(n22945), .B(n22946), .Z(n22941) );
  AND U24256 ( .A(n16353), .B(n22947), .Z(n22945) );
  XNOR U24257 ( .A(n16352), .B(n22946), .Z(n22947) );
  NAND U24258 ( .A(n22948), .B(n[738]), .Z(n16352) );
  NAND U24259 ( .A(n21523), .B(n[738]), .Z(n22948) );
  XNOR U24260 ( .A(n22949), .B(n22946), .Z(n16353) );
  XOR U24261 ( .A(n22950), .B(n22951), .Z(n22946) );
  AND U24262 ( .A(n16360), .B(n22952), .Z(n22950) );
  XNOR U24263 ( .A(n16359), .B(n22951), .Z(n22952) );
  NAND U24264 ( .A(n22953), .B(n[737]), .Z(n16359) );
  NAND U24265 ( .A(n21523), .B(n[737]), .Z(n22953) );
  XNOR U24266 ( .A(n22954), .B(n22951), .Z(n16360) );
  XOR U24267 ( .A(n22955), .B(n22956), .Z(n22951) );
  AND U24268 ( .A(n16367), .B(n22957), .Z(n22955) );
  XNOR U24269 ( .A(n16366), .B(n22956), .Z(n22957) );
  NAND U24270 ( .A(n22958), .B(n[736]), .Z(n16366) );
  NAND U24271 ( .A(n21523), .B(n[736]), .Z(n22958) );
  XNOR U24272 ( .A(n22959), .B(n22956), .Z(n16367) );
  XOR U24273 ( .A(n22960), .B(n22961), .Z(n22956) );
  AND U24274 ( .A(n16374), .B(n22962), .Z(n22960) );
  XNOR U24275 ( .A(n16373), .B(n22961), .Z(n22962) );
  NAND U24276 ( .A(n22963), .B(n[735]), .Z(n16373) );
  NAND U24277 ( .A(n21523), .B(n[735]), .Z(n22963) );
  XNOR U24278 ( .A(n22964), .B(n22961), .Z(n16374) );
  XOR U24279 ( .A(n22965), .B(n22966), .Z(n22961) );
  AND U24280 ( .A(n16381), .B(n22967), .Z(n22965) );
  XNOR U24281 ( .A(n16380), .B(n22966), .Z(n22967) );
  NAND U24282 ( .A(n22968), .B(n[734]), .Z(n16380) );
  NAND U24283 ( .A(n21523), .B(n[734]), .Z(n22968) );
  XNOR U24284 ( .A(n22969), .B(n22966), .Z(n16381) );
  XOR U24285 ( .A(n22970), .B(n22971), .Z(n22966) );
  AND U24286 ( .A(n16388), .B(n22972), .Z(n22970) );
  XNOR U24287 ( .A(n16387), .B(n22971), .Z(n22972) );
  NAND U24288 ( .A(n22973), .B(n[733]), .Z(n16387) );
  NAND U24289 ( .A(n21523), .B(n[733]), .Z(n22973) );
  XNOR U24290 ( .A(n22974), .B(n22971), .Z(n16388) );
  XOR U24291 ( .A(n22975), .B(n22976), .Z(n22971) );
  AND U24292 ( .A(n16395), .B(n22977), .Z(n22975) );
  XNOR U24293 ( .A(n16394), .B(n22976), .Z(n22977) );
  NAND U24294 ( .A(n22978), .B(n[732]), .Z(n16394) );
  NAND U24295 ( .A(n21523), .B(n[732]), .Z(n22978) );
  XNOR U24296 ( .A(n22979), .B(n22976), .Z(n16395) );
  XOR U24297 ( .A(n22980), .B(n22981), .Z(n22976) );
  AND U24298 ( .A(n16402), .B(n22982), .Z(n22980) );
  XNOR U24299 ( .A(n16401), .B(n22981), .Z(n22982) );
  NAND U24300 ( .A(n22983), .B(n[731]), .Z(n16401) );
  NAND U24301 ( .A(n21523), .B(n[731]), .Z(n22983) );
  XNOR U24302 ( .A(n22984), .B(n22981), .Z(n16402) );
  XOR U24303 ( .A(n22985), .B(n22986), .Z(n22981) );
  AND U24304 ( .A(n16409), .B(n22987), .Z(n22985) );
  XNOR U24305 ( .A(n16408), .B(n22986), .Z(n22987) );
  NAND U24306 ( .A(n22988), .B(n[730]), .Z(n16408) );
  NAND U24307 ( .A(n21523), .B(n[730]), .Z(n22988) );
  XNOR U24308 ( .A(n22989), .B(n22986), .Z(n16409) );
  XOR U24309 ( .A(n22990), .B(n22991), .Z(n22986) );
  AND U24310 ( .A(n16416), .B(n22992), .Z(n22990) );
  XNOR U24311 ( .A(n16415), .B(n22991), .Z(n22992) );
  NAND U24312 ( .A(n22993), .B(n[729]), .Z(n16415) );
  NAND U24313 ( .A(n21523), .B(n[729]), .Z(n22993) );
  XNOR U24314 ( .A(n22994), .B(n22991), .Z(n16416) );
  XOR U24315 ( .A(n22995), .B(n22996), .Z(n22991) );
  AND U24316 ( .A(n16423), .B(n22997), .Z(n22995) );
  XNOR U24317 ( .A(n16422), .B(n22996), .Z(n22997) );
  NAND U24318 ( .A(n22998), .B(n[728]), .Z(n16422) );
  NAND U24319 ( .A(n21523), .B(n[728]), .Z(n22998) );
  XNOR U24320 ( .A(n22999), .B(n22996), .Z(n16423) );
  XOR U24321 ( .A(n23000), .B(n23001), .Z(n22996) );
  AND U24322 ( .A(n16430), .B(n23002), .Z(n23000) );
  XNOR U24323 ( .A(n16429), .B(n23001), .Z(n23002) );
  NAND U24324 ( .A(n23003), .B(n[727]), .Z(n16429) );
  NAND U24325 ( .A(n21523), .B(n[727]), .Z(n23003) );
  XNOR U24326 ( .A(n23004), .B(n23001), .Z(n16430) );
  XOR U24327 ( .A(n23005), .B(n23006), .Z(n23001) );
  AND U24328 ( .A(n16437), .B(n23007), .Z(n23005) );
  XNOR U24329 ( .A(n16436), .B(n23006), .Z(n23007) );
  NAND U24330 ( .A(n23008), .B(n[726]), .Z(n16436) );
  NAND U24331 ( .A(n21523), .B(n[726]), .Z(n23008) );
  XNOR U24332 ( .A(n23009), .B(n23006), .Z(n16437) );
  XOR U24333 ( .A(n23010), .B(n23011), .Z(n23006) );
  AND U24334 ( .A(n16444), .B(n23012), .Z(n23010) );
  XNOR U24335 ( .A(n16443), .B(n23011), .Z(n23012) );
  NAND U24336 ( .A(n23013), .B(n[725]), .Z(n16443) );
  NAND U24337 ( .A(n21523), .B(n[725]), .Z(n23013) );
  XNOR U24338 ( .A(n23014), .B(n23011), .Z(n16444) );
  XOR U24339 ( .A(n23015), .B(n23016), .Z(n23011) );
  AND U24340 ( .A(n16451), .B(n23017), .Z(n23015) );
  XNOR U24341 ( .A(n16450), .B(n23016), .Z(n23017) );
  NAND U24342 ( .A(n23018), .B(n[724]), .Z(n16450) );
  NAND U24343 ( .A(n21523), .B(n[724]), .Z(n23018) );
  XNOR U24344 ( .A(n23019), .B(n23016), .Z(n16451) );
  XOR U24345 ( .A(n23020), .B(n23021), .Z(n23016) );
  AND U24346 ( .A(n16458), .B(n23022), .Z(n23020) );
  XNOR U24347 ( .A(n16457), .B(n23021), .Z(n23022) );
  NAND U24348 ( .A(n23023), .B(n[723]), .Z(n16457) );
  NAND U24349 ( .A(n21523), .B(n[723]), .Z(n23023) );
  XNOR U24350 ( .A(n23024), .B(n23021), .Z(n16458) );
  XOR U24351 ( .A(n23025), .B(n23026), .Z(n23021) );
  AND U24352 ( .A(n16465), .B(n23027), .Z(n23025) );
  XNOR U24353 ( .A(n16464), .B(n23026), .Z(n23027) );
  NAND U24354 ( .A(n23028), .B(n[722]), .Z(n16464) );
  NAND U24355 ( .A(n21523), .B(n[722]), .Z(n23028) );
  XNOR U24356 ( .A(n23029), .B(n23026), .Z(n16465) );
  XOR U24357 ( .A(n23030), .B(n23031), .Z(n23026) );
  AND U24358 ( .A(n16472), .B(n23032), .Z(n23030) );
  XNOR U24359 ( .A(n16471), .B(n23031), .Z(n23032) );
  NAND U24360 ( .A(n23033), .B(n[721]), .Z(n16471) );
  NAND U24361 ( .A(n21523), .B(n[721]), .Z(n23033) );
  XNOR U24362 ( .A(n23034), .B(n23031), .Z(n16472) );
  XOR U24363 ( .A(n23035), .B(n23036), .Z(n23031) );
  AND U24364 ( .A(n16479), .B(n23037), .Z(n23035) );
  XNOR U24365 ( .A(n16478), .B(n23036), .Z(n23037) );
  NAND U24366 ( .A(n23038), .B(n[720]), .Z(n16478) );
  NAND U24367 ( .A(n21523), .B(n[720]), .Z(n23038) );
  XNOR U24368 ( .A(n23039), .B(n23036), .Z(n16479) );
  XOR U24369 ( .A(n23040), .B(n23041), .Z(n23036) );
  AND U24370 ( .A(n16486), .B(n23042), .Z(n23040) );
  XNOR U24371 ( .A(n16485), .B(n23041), .Z(n23042) );
  NAND U24372 ( .A(n23043), .B(n[719]), .Z(n16485) );
  NAND U24373 ( .A(n21523), .B(n[719]), .Z(n23043) );
  XNOR U24374 ( .A(n23044), .B(n23041), .Z(n16486) );
  XOR U24375 ( .A(n23045), .B(n23046), .Z(n23041) );
  AND U24376 ( .A(n16493), .B(n23047), .Z(n23045) );
  XNOR U24377 ( .A(n16492), .B(n23046), .Z(n23047) );
  NAND U24378 ( .A(n23048), .B(n[718]), .Z(n16492) );
  NAND U24379 ( .A(n21523), .B(n[718]), .Z(n23048) );
  XNOR U24380 ( .A(n23049), .B(n23046), .Z(n16493) );
  XOR U24381 ( .A(n23050), .B(n23051), .Z(n23046) );
  AND U24382 ( .A(n16500), .B(n23052), .Z(n23050) );
  XNOR U24383 ( .A(n16499), .B(n23051), .Z(n23052) );
  NAND U24384 ( .A(n23053), .B(n[717]), .Z(n16499) );
  NAND U24385 ( .A(n21523), .B(n[717]), .Z(n23053) );
  XNOR U24386 ( .A(n23054), .B(n23051), .Z(n16500) );
  XOR U24387 ( .A(n23055), .B(n23056), .Z(n23051) );
  AND U24388 ( .A(n16507), .B(n23057), .Z(n23055) );
  XNOR U24389 ( .A(n16506), .B(n23056), .Z(n23057) );
  NAND U24390 ( .A(n23058), .B(n[716]), .Z(n16506) );
  NAND U24391 ( .A(n21523), .B(n[716]), .Z(n23058) );
  XNOR U24392 ( .A(n23059), .B(n23056), .Z(n16507) );
  XOR U24393 ( .A(n23060), .B(n23061), .Z(n23056) );
  AND U24394 ( .A(n16514), .B(n23062), .Z(n23060) );
  XNOR U24395 ( .A(n16513), .B(n23061), .Z(n23062) );
  NAND U24396 ( .A(n23063), .B(n[715]), .Z(n16513) );
  NAND U24397 ( .A(n21523), .B(n[715]), .Z(n23063) );
  XNOR U24398 ( .A(n23064), .B(n23061), .Z(n16514) );
  XOR U24399 ( .A(n23065), .B(n23066), .Z(n23061) );
  AND U24400 ( .A(n16521), .B(n23067), .Z(n23065) );
  XNOR U24401 ( .A(n16520), .B(n23066), .Z(n23067) );
  NAND U24402 ( .A(n23068), .B(n[714]), .Z(n16520) );
  NAND U24403 ( .A(n21523), .B(n[714]), .Z(n23068) );
  XNOR U24404 ( .A(n23069), .B(n23066), .Z(n16521) );
  XOR U24405 ( .A(n23070), .B(n23071), .Z(n23066) );
  AND U24406 ( .A(n16528), .B(n23072), .Z(n23070) );
  XNOR U24407 ( .A(n16527), .B(n23071), .Z(n23072) );
  NAND U24408 ( .A(n23073), .B(n[713]), .Z(n16527) );
  NAND U24409 ( .A(n21523), .B(n[713]), .Z(n23073) );
  XNOR U24410 ( .A(n23074), .B(n23071), .Z(n16528) );
  XOR U24411 ( .A(n23075), .B(n23076), .Z(n23071) );
  AND U24412 ( .A(n16535), .B(n23077), .Z(n23075) );
  XNOR U24413 ( .A(n16534), .B(n23076), .Z(n23077) );
  NAND U24414 ( .A(n23078), .B(n[712]), .Z(n16534) );
  NAND U24415 ( .A(n21523), .B(n[712]), .Z(n23078) );
  XNOR U24416 ( .A(n23079), .B(n23076), .Z(n16535) );
  XOR U24417 ( .A(n23080), .B(n23081), .Z(n23076) );
  AND U24418 ( .A(n16542), .B(n23082), .Z(n23080) );
  XNOR U24419 ( .A(n16541), .B(n23081), .Z(n23082) );
  NAND U24420 ( .A(n23083), .B(n[711]), .Z(n16541) );
  NAND U24421 ( .A(n21523), .B(n[711]), .Z(n23083) );
  XNOR U24422 ( .A(n23084), .B(n23081), .Z(n16542) );
  XOR U24423 ( .A(n23085), .B(n23086), .Z(n23081) );
  AND U24424 ( .A(n16549), .B(n23087), .Z(n23085) );
  XNOR U24425 ( .A(n16548), .B(n23086), .Z(n23087) );
  NAND U24426 ( .A(n23088), .B(n[710]), .Z(n16548) );
  NAND U24427 ( .A(n21523), .B(n[710]), .Z(n23088) );
  XNOR U24428 ( .A(n23089), .B(n23086), .Z(n16549) );
  XOR U24429 ( .A(n23090), .B(n23091), .Z(n23086) );
  AND U24430 ( .A(n16556), .B(n23092), .Z(n23090) );
  XNOR U24431 ( .A(n16555), .B(n23091), .Z(n23092) );
  NAND U24432 ( .A(n23093), .B(n[709]), .Z(n16555) );
  NAND U24433 ( .A(n21523), .B(n[709]), .Z(n23093) );
  XNOR U24434 ( .A(n23094), .B(n23091), .Z(n16556) );
  XOR U24435 ( .A(n23095), .B(n23096), .Z(n23091) );
  AND U24436 ( .A(n16563), .B(n23097), .Z(n23095) );
  XNOR U24437 ( .A(n16562), .B(n23096), .Z(n23097) );
  NAND U24438 ( .A(n23098), .B(n[708]), .Z(n16562) );
  NAND U24439 ( .A(n21523), .B(n[708]), .Z(n23098) );
  XNOR U24440 ( .A(n23099), .B(n23096), .Z(n16563) );
  XOR U24441 ( .A(n23100), .B(n23101), .Z(n23096) );
  AND U24442 ( .A(n16570), .B(n23102), .Z(n23100) );
  XNOR U24443 ( .A(n16569), .B(n23101), .Z(n23102) );
  NAND U24444 ( .A(n23103), .B(n[707]), .Z(n16569) );
  NAND U24445 ( .A(n21523), .B(n[707]), .Z(n23103) );
  XNOR U24446 ( .A(n23104), .B(n23101), .Z(n16570) );
  XOR U24447 ( .A(n23105), .B(n23106), .Z(n23101) );
  AND U24448 ( .A(n16577), .B(n23107), .Z(n23105) );
  XNOR U24449 ( .A(n16576), .B(n23106), .Z(n23107) );
  NAND U24450 ( .A(n23108), .B(n[706]), .Z(n16576) );
  NAND U24451 ( .A(n21523), .B(n[706]), .Z(n23108) );
  XNOR U24452 ( .A(n23109), .B(n23106), .Z(n16577) );
  XOR U24453 ( .A(n23110), .B(n23111), .Z(n23106) );
  AND U24454 ( .A(n16584), .B(n23112), .Z(n23110) );
  XNOR U24455 ( .A(n16583), .B(n23111), .Z(n23112) );
  NAND U24456 ( .A(n23113), .B(n[705]), .Z(n16583) );
  NAND U24457 ( .A(n21523), .B(n[705]), .Z(n23113) );
  XNOR U24458 ( .A(n23114), .B(n23111), .Z(n16584) );
  XOR U24459 ( .A(n23115), .B(n23116), .Z(n23111) );
  AND U24460 ( .A(n16591), .B(n23117), .Z(n23115) );
  XNOR U24461 ( .A(n16590), .B(n23116), .Z(n23117) );
  NAND U24462 ( .A(n23118), .B(n[704]), .Z(n16590) );
  NAND U24463 ( .A(n21523), .B(n[704]), .Z(n23118) );
  XNOR U24464 ( .A(n23119), .B(n23116), .Z(n16591) );
  XOR U24465 ( .A(n23120), .B(n23121), .Z(n23116) );
  AND U24466 ( .A(n16598), .B(n23122), .Z(n23120) );
  XNOR U24467 ( .A(n16597), .B(n23121), .Z(n23122) );
  NAND U24468 ( .A(n23123), .B(n[703]), .Z(n16597) );
  NAND U24469 ( .A(n21523), .B(n[703]), .Z(n23123) );
  XNOR U24470 ( .A(n23124), .B(n23121), .Z(n16598) );
  XOR U24471 ( .A(n23125), .B(n23126), .Z(n23121) );
  AND U24472 ( .A(n16605), .B(n23127), .Z(n23125) );
  XNOR U24473 ( .A(n16604), .B(n23126), .Z(n23127) );
  NAND U24474 ( .A(n23128), .B(n[702]), .Z(n16604) );
  NAND U24475 ( .A(n21523), .B(n[702]), .Z(n23128) );
  XNOR U24476 ( .A(n23129), .B(n23126), .Z(n16605) );
  XOR U24477 ( .A(n23130), .B(n23131), .Z(n23126) );
  AND U24478 ( .A(n16612), .B(n23132), .Z(n23130) );
  XNOR U24479 ( .A(n16611), .B(n23131), .Z(n23132) );
  NAND U24480 ( .A(n23133), .B(n[701]), .Z(n16611) );
  NAND U24481 ( .A(n21523), .B(n[701]), .Z(n23133) );
  XNOR U24482 ( .A(n23134), .B(n23131), .Z(n16612) );
  XOR U24483 ( .A(n23135), .B(n23136), .Z(n23131) );
  AND U24484 ( .A(n16619), .B(n23137), .Z(n23135) );
  XNOR U24485 ( .A(n16618), .B(n23136), .Z(n23137) );
  NAND U24486 ( .A(n23138), .B(n[700]), .Z(n16618) );
  NAND U24487 ( .A(n21523), .B(n[700]), .Z(n23138) );
  XNOR U24488 ( .A(n23139), .B(n23136), .Z(n16619) );
  XOR U24489 ( .A(n23140), .B(n23141), .Z(n23136) );
  AND U24490 ( .A(n16626), .B(n23142), .Z(n23140) );
  XNOR U24491 ( .A(n16625), .B(n23141), .Z(n23142) );
  NAND U24492 ( .A(n23143), .B(n[699]), .Z(n16625) );
  NAND U24493 ( .A(n21523), .B(n[699]), .Z(n23143) );
  XNOR U24494 ( .A(n23144), .B(n23141), .Z(n16626) );
  XOR U24495 ( .A(n23145), .B(n23146), .Z(n23141) );
  AND U24496 ( .A(n16633), .B(n23147), .Z(n23145) );
  XNOR U24497 ( .A(n16632), .B(n23146), .Z(n23147) );
  NAND U24498 ( .A(n23148), .B(n[698]), .Z(n16632) );
  NAND U24499 ( .A(n21523), .B(n[698]), .Z(n23148) );
  XNOR U24500 ( .A(n23149), .B(n23146), .Z(n16633) );
  XOR U24501 ( .A(n23150), .B(n23151), .Z(n23146) );
  AND U24502 ( .A(n16640), .B(n23152), .Z(n23150) );
  XNOR U24503 ( .A(n16639), .B(n23151), .Z(n23152) );
  NAND U24504 ( .A(n23153), .B(n[697]), .Z(n16639) );
  NAND U24505 ( .A(n21523), .B(n[697]), .Z(n23153) );
  XNOR U24506 ( .A(n23154), .B(n23151), .Z(n16640) );
  XOR U24507 ( .A(n23155), .B(n23156), .Z(n23151) );
  AND U24508 ( .A(n16647), .B(n23157), .Z(n23155) );
  XNOR U24509 ( .A(n16646), .B(n23156), .Z(n23157) );
  NAND U24510 ( .A(n23158), .B(n[696]), .Z(n16646) );
  NAND U24511 ( .A(n21523), .B(n[696]), .Z(n23158) );
  XNOR U24512 ( .A(n23159), .B(n23156), .Z(n16647) );
  XOR U24513 ( .A(n23160), .B(n23161), .Z(n23156) );
  AND U24514 ( .A(n16654), .B(n23162), .Z(n23160) );
  XNOR U24515 ( .A(n16653), .B(n23161), .Z(n23162) );
  NAND U24516 ( .A(n23163), .B(n[695]), .Z(n16653) );
  NAND U24517 ( .A(n21523), .B(n[695]), .Z(n23163) );
  XNOR U24518 ( .A(n23164), .B(n23161), .Z(n16654) );
  XOR U24519 ( .A(n23165), .B(n23166), .Z(n23161) );
  AND U24520 ( .A(n16661), .B(n23167), .Z(n23165) );
  XNOR U24521 ( .A(n16660), .B(n23166), .Z(n23167) );
  NAND U24522 ( .A(n23168), .B(n[694]), .Z(n16660) );
  NAND U24523 ( .A(n21523), .B(n[694]), .Z(n23168) );
  XNOR U24524 ( .A(n23169), .B(n23166), .Z(n16661) );
  XOR U24525 ( .A(n23170), .B(n23171), .Z(n23166) );
  AND U24526 ( .A(n16668), .B(n23172), .Z(n23170) );
  XNOR U24527 ( .A(n16667), .B(n23171), .Z(n23172) );
  NAND U24528 ( .A(n23173), .B(n[693]), .Z(n16667) );
  NAND U24529 ( .A(n21523), .B(n[693]), .Z(n23173) );
  XNOR U24530 ( .A(n23174), .B(n23171), .Z(n16668) );
  XOR U24531 ( .A(n23175), .B(n23176), .Z(n23171) );
  AND U24532 ( .A(n16675), .B(n23177), .Z(n23175) );
  XNOR U24533 ( .A(n16674), .B(n23176), .Z(n23177) );
  NAND U24534 ( .A(n23178), .B(n[692]), .Z(n16674) );
  NAND U24535 ( .A(n21523), .B(n[692]), .Z(n23178) );
  XNOR U24536 ( .A(n23179), .B(n23176), .Z(n16675) );
  XOR U24537 ( .A(n23180), .B(n23181), .Z(n23176) );
  AND U24538 ( .A(n16682), .B(n23182), .Z(n23180) );
  XNOR U24539 ( .A(n16681), .B(n23181), .Z(n23182) );
  NAND U24540 ( .A(n23183), .B(n[691]), .Z(n16681) );
  NAND U24541 ( .A(n21523), .B(n[691]), .Z(n23183) );
  XNOR U24542 ( .A(n23184), .B(n23181), .Z(n16682) );
  XOR U24543 ( .A(n23185), .B(n23186), .Z(n23181) );
  AND U24544 ( .A(n16689), .B(n23187), .Z(n23185) );
  XNOR U24545 ( .A(n16688), .B(n23186), .Z(n23187) );
  NAND U24546 ( .A(n23188), .B(n[690]), .Z(n16688) );
  NAND U24547 ( .A(n21523), .B(n[690]), .Z(n23188) );
  XNOR U24548 ( .A(n23189), .B(n23186), .Z(n16689) );
  XOR U24549 ( .A(n23190), .B(n23191), .Z(n23186) );
  AND U24550 ( .A(n16696), .B(n23192), .Z(n23190) );
  XNOR U24551 ( .A(n16695), .B(n23191), .Z(n23192) );
  NAND U24552 ( .A(n23193), .B(n[689]), .Z(n16695) );
  NAND U24553 ( .A(n21523), .B(n[689]), .Z(n23193) );
  XNOR U24554 ( .A(n23194), .B(n23191), .Z(n16696) );
  XOR U24555 ( .A(n23195), .B(n23196), .Z(n23191) );
  AND U24556 ( .A(n16703), .B(n23197), .Z(n23195) );
  XNOR U24557 ( .A(n16702), .B(n23196), .Z(n23197) );
  NAND U24558 ( .A(n23198), .B(n[688]), .Z(n16702) );
  NAND U24559 ( .A(n21523), .B(n[688]), .Z(n23198) );
  XNOR U24560 ( .A(n23199), .B(n23196), .Z(n16703) );
  XOR U24561 ( .A(n23200), .B(n23201), .Z(n23196) );
  AND U24562 ( .A(n16710), .B(n23202), .Z(n23200) );
  XNOR U24563 ( .A(n16709), .B(n23201), .Z(n23202) );
  NAND U24564 ( .A(n23203), .B(n[687]), .Z(n16709) );
  NAND U24565 ( .A(n21523), .B(n[687]), .Z(n23203) );
  XNOR U24566 ( .A(n23204), .B(n23201), .Z(n16710) );
  XOR U24567 ( .A(n23205), .B(n23206), .Z(n23201) );
  AND U24568 ( .A(n16717), .B(n23207), .Z(n23205) );
  XNOR U24569 ( .A(n16716), .B(n23206), .Z(n23207) );
  NAND U24570 ( .A(n23208), .B(n[686]), .Z(n16716) );
  NAND U24571 ( .A(n21523), .B(n[686]), .Z(n23208) );
  XNOR U24572 ( .A(n23209), .B(n23206), .Z(n16717) );
  XOR U24573 ( .A(n23210), .B(n23211), .Z(n23206) );
  AND U24574 ( .A(n16724), .B(n23212), .Z(n23210) );
  XNOR U24575 ( .A(n16723), .B(n23211), .Z(n23212) );
  NAND U24576 ( .A(n23213), .B(n[685]), .Z(n16723) );
  NAND U24577 ( .A(n21523), .B(n[685]), .Z(n23213) );
  XNOR U24578 ( .A(n23214), .B(n23211), .Z(n16724) );
  XOR U24579 ( .A(n23215), .B(n23216), .Z(n23211) );
  AND U24580 ( .A(n16731), .B(n23217), .Z(n23215) );
  XNOR U24581 ( .A(n16730), .B(n23216), .Z(n23217) );
  NAND U24582 ( .A(n23218), .B(n[684]), .Z(n16730) );
  NAND U24583 ( .A(n21523), .B(n[684]), .Z(n23218) );
  XNOR U24584 ( .A(n23219), .B(n23216), .Z(n16731) );
  XOR U24585 ( .A(n23220), .B(n23221), .Z(n23216) );
  AND U24586 ( .A(n16738), .B(n23222), .Z(n23220) );
  XNOR U24587 ( .A(n16737), .B(n23221), .Z(n23222) );
  NAND U24588 ( .A(n23223), .B(n[683]), .Z(n16737) );
  NAND U24589 ( .A(n21523), .B(n[683]), .Z(n23223) );
  XNOR U24590 ( .A(n23224), .B(n23221), .Z(n16738) );
  XOR U24591 ( .A(n23225), .B(n23226), .Z(n23221) );
  AND U24592 ( .A(n16745), .B(n23227), .Z(n23225) );
  XNOR U24593 ( .A(n16744), .B(n23226), .Z(n23227) );
  NAND U24594 ( .A(n23228), .B(n[682]), .Z(n16744) );
  NAND U24595 ( .A(n21523), .B(n[682]), .Z(n23228) );
  XNOR U24596 ( .A(n23229), .B(n23226), .Z(n16745) );
  XOR U24597 ( .A(n23230), .B(n23231), .Z(n23226) );
  AND U24598 ( .A(n16752), .B(n23232), .Z(n23230) );
  XNOR U24599 ( .A(n16751), .B(n23231), .Z(n23232) );
  NAND U24600 ( .A(n23233), .B(n[681]), .Z(n16751) );
  NAND U24601 ( .A(n21523), .B(n[681]), .Z(n23233) );
  XNOR U24602 ( .A(n23234), .B(n23231), .Z(n16752) );
  XOR U24603 ( .A(n23235), .B(n23236), .Z(n23231) );
  AND U24604 ( .A(n16759), .B(n23237), .Z(n23235) );
  XNOR U24605 ( .A(n16758), .B(n23236), .Z(n23237) );
  NAND U24606 ( .A(n23238), .B(n[680]), .Z(n16758) );
  NAND U24607 ( .A(n21523), .B(n[680]), .Z(n23238) );
  XNOR U24608 ( .A(n23239), .B(n23236), .Z(n16759) );
  XOR U24609 ( .A(n23240), .B(n23241), .Z(n23236) );
  AND U24610 ( .A(n16766), .B(n23242), .Z(n23240) );
  XNOR U24611 ( .A(n16765), .B(n23241), .Z(n23242) );
  NAND U24612 ( .A(n23243), .B(n[679]), .Z(n16765) );
  NAND U24613 ( .A(n21523), .B(n[679]), .Z(n23243) );
  XNOR U24614 ( .A(n23244), .B(n23241), .Z(n16766) );
  XOR U24615 ( .A(n23245), .B(n23246), .Z(n23241) );
  AND U24616 ( .A(n16773), .B(n23247), .Z(n23245) );
  XNOR U24617 ( .A(n16772), .B(n23246), .Z(n23247) );
  NAND U24618 ( .A(n23248), .B(n[678]), .Z(n16772) );
  NAND U24619 ( .A(n21523), .B(n[678]), .Z(n23248) );
  XNOR U24620 ( .A(n23249), .B(n23246), .Z(n16773) );
  XOR U24621 ( .A(n23250), .B(n23251), .Z(n23246) );
  AND U24622 ( .A(n16780), .B(n23252), .Z(n23250) );
  XNOR U24623 ( .A(n16779), .B(n23251), .Z(n23252) );
  NAND U24624 ( .A(n23253), .B(n[677]), .Z(n16779) );
  NAND U24625 ( .A(n21523), .B(n[677]), .Z(n23253) );
  XNOR U24626 ( .A(n23254), .B(n23251), .Z(n16780) );
  XOR U24627 ( .A(n23255), .B(n23256), .Z(n23251) );
  AND U24628 ( .A(n16787), .B(n23257), .Z(n23255) );
  XNOR U24629 ( .A(n16786), .B(n23256), .Z(n23257) );
  NAND U24630 ( .A(n23258), .B(n[676]), .Z(n16786) );
  NAND U24631 ( .A(n21523), .B(n[676]), .Z(n23258) );
  XNOR U24632 ( .A(n23259), .B(n23256), .Z(n16787) );
  XOR U24633 ( .A(n23260), .B(n23261), .Z(n23256) );
  AND U24634 ( .A(n16794), .B(n23262), .Z(n23260) );
  XNOR U24635 ( .A(n16793), .B(n23261), .Z(n23262) );
  NAND U24636 ( .A(n23263), .B(n[675]), .Z(n16793) );
  NAND U24637 ( .A(n21523), .B(n[675]), .Z(n23263) );
  XNOR U24638 ( .A(n23264), .B(n23261), .Z(n16794) );
  XOR U24639 ( .A(n23265), .B(n23266), .Z(n23261) );
  AND U24640 ( .A(n16801), .B(n23267), .Z(n23265) );
  XNOR U24641 ( .A(n16800), .B(n23266), .Z(n23267) );
  NAND U24642 ( .A(n23268), .B(n[674]), .Z(n16800) );
  NAND U24643 ( .A(n21523), .B(n[674]), .Z(n23268) );
  XNOR U24644 ( .A(n23269), .B(n23266), .Z(n16801) );
  XOR U24645 ( .A(n23270), .B(n23271), .Z(n23266) );
  AND U24646 ( .A(n16808), .B(n23272), .Z(n23270) );
  XNOR U24647 ( .A(n16807), .B(n23271), .Z(n23272) );
  NAND U24648 ( .A(n23273), .B(n[673]), .Z(n16807) );
  NAND U24649 ( .A(n21523), .B(n[673]), .Z(n23273) );
  XNOR U24650 ( .A(n23274), .B(n23271), .Z(n16808) );
  XOR U24651 ( .A(n23275), .B(n23276), .Z(n23271) );
  AND U24652 ( .A(n16815), .B(n23277), .Z(n23275) );
  XNOR U24653 ( .A(n16814), .B(n23276), .Z(n23277) );
  NAND U24654 ( .A(n23278), .B(n[672]), .Z(n16814) );
  NAND U24655 ( .A(n21523), .B(n[672]), .Z(n23278) );
  XNOR U24656 ( .A(n23279), .B(n23276), .Z(n16815) );
  XOR U24657 ( .A(n23280), .B(n23281), .Z(n23276) );
  AND U24658 ( .A(n16822), .B(n23282), .Z(n23280) );
  XNOR U24659 ( .A(n16821), .B(n23281), .Z(n23282) );
  NAND U24660 ( .A(n23283), .B(n[671]), .Z(n16821) );
  NAND U24661 ( .A(n21523), .B(n[671]), .Z(n23283) );
  XNOR U24662 ( .A(n23284), .B(n23281), .Z(n16822) );
  XOR U24663 ( .A(n23285), .B(n23286), .Z(n23281) );
  AND U24664 ( .A(n16829), .B(n23287), .Z(n23285) );
  XNOR U24665 ( .A(n16828), .B(n23286), .Z(n23287) );
  NAND U24666 ( .A(n23288), .B(n[670]), .Z(n16828) );
  NAND U24667 ( .A(n21523), .B(n[670]), .Z(n23288) );
  XNOR U24668 ( .A(n23289), .B(n23286), .Z(n16829) );
  XOR U24669 ( .A(n23290), .B(n23291), .Z(n23286) );
  AND U24670 ( .A(n16836), .B(n23292), .Z(n23290) );
  XNOR U24671 ( .A(n16835), .B(n23291), .Z(n23292) );
  NAND U24672 ( .A(n23293), .B(n[669]), .Z(n16835) );
  NAND U24673 ( .A(n21523), .B(n[669]), .Z(n23293) );
  XNOR U24674 ( .A(n23294), .B(n23291), .Z(n16836) );
  XOR U24675 ( .A(n23295), .B(n23296), .Z(n23291) );
  AND U24676 ( .A(n16843), .B(n23297), .Z(n23295) );
  XNOR U24677 ( .A(n16842), .B(n23296), .Z(n23297) );
  NAND U24678 ( .A(n23298), .B(n[668]), .Z(n16842) );
  NAND U24679 ( .A(n21523), .B(n[668]), .Z(n23298) );
  XNOR U24680 ( .A(n23299), .B(n23296), .Z(n16843) );
  XOR U24681 ( .A(n23300), .B(n23301), .Z(n23296) );
  AND U24682 ( .A(n16850), .B(n23302), .Z(n23300) );
  XNOR U24683 ( .A(n16849), .B(n23301), .Z(n23302) );
  NAND U24684 ( .A(n23303), .B(n[667]), .Z(n16849) );
  NAND U24685 ( .A(n21523), .B(n[667]), .Z(n23303) );
  XNOR U24686 ( .A(n23304), .B(n23301), .Z(n16850) );
  XOR U24687 ( .A(n23305), .B(n23306), .Z(n23301) );
  AND U24688 ( .A(n16857), .B(n23307), .Z(n23305) );
  XNOR U24689 ( .A(n16856), .B(n23306), .Z(n23307) );
  NAND U24690 ( .A(n23308), .B(n[666]), .Z(n16856) );
  NAND U24691 ( .A(n21523), .B(n[666]), .Z(n23308) );
  XNOR U24692 ( .A(n23309), .B(n23306), .Z(n16857) );
  XOR U24693 ( .A(n23310), .B(n23311), .Z(n23306) );
  AND U24694 ( .A(n16864), .B(n23312), .Z(n23310) );
  XNOR U24695 ( .A(n16863), .B(n23311), .Z(n23312) );
  NAND U24696 ( .A(n23313), .B(n[665]), .Z(n16863) );
  NAND U24697 ( .A(n21523), .B(n[665]), .Z(n23313) );
  XNOR U24698 ( .A(n23314), .B(n23311), .Z(n16864) );
  XOR U24699 ( .A(n23315), .B(n23316), .Z(n23311) );
  AND U24700 ( .A(n16871), .B(n23317), .Z(n23315) );
  XNOR U24701 ( .A(n16870), .B(n23316), .Z(n23317) );
  NAND U24702 ( .A(n23318), .B(n[664]), .Z(n16870) );
  NAND U24703 ( .A(n21523), .B(n[664]), .Z(n23318) );
  XNOR U24704 ( .A(n23319), .B(n23316), .Z(n16871) );
  XOR U24705 ( .A(n23320), .B(n23321), .Z(n23316) );
  AND U24706 ( .A(n16878), .B(n23322), .Z(n23320) );
  XNOR U24707 ( .A(n16877), .B(n23321), .Z(n23322) );
  NAND U24708 ( .A(n23323), .B(n[663]), .Z(n16877) );
  NAND U24709 ( .A(n21523), .B(n[663]), .Z(n23323) );
  XNOR U24710 ( .A(n23324), .B(n23321), .Z(n16878) );
  XOR U24711 ( .A(n23325), .B(n23326), .Z(n23321) );
  AND U24712 ( .A(n16885), .B(n23327), .Z(n23325) );
  XNOR U24713 ( .A(n16884), .B(n23326), .Z(n23327) );
  NAND U24714 ( .A(n23328), .B(n[662]), .Z(n16884) );
  NAND U24715 ( .A(n21523), .B(n[662]), .Z(n23328) );
  XNOR U24716 ( .A(n23329), .B(n23326), .Z(n16885) );
  XOR U24717 ( .A(n23330), .B(n23331), .Z(n23326) );
  AND U24718 ( .A(n16892), .B(n23332), .Z(n23330) );
  XNOR U24719 ( .A(n16891), .B(n23331), .Z(n23332) );
  NAND U24720 ( .A(n23333), .B(n[661]), .Z(n16891) );
  NAND U24721 ( .A(n21523), .B(n[661]), .Z(n23333) );
  XNOR U24722 ( .A(n23334), .B(n23331), .Z(n16892) );
  XOR U24723 ( .A(n23335), .B(n23336), .Z(n23331) );
  AND U24724 ( .A(n16899), .B(n23337), .Z(n23335) );
  XNOR U24725 ( .A(n16898), .B(n23336), .Z(n23337) );
  NAND U24726 ( .A(n23338), .B(n[660]), .Z(n16898) );
  NAND U24727 ( .A(n21523), .B(n[660]), .Z(n23338) );
  XNOR U24728 ( .A(n23339), .B(n23336), .Z(n16899) );
  XOR U24729 ( .A(n23340), .B(n23341), .Z(n23336) );
  AND U24730 ( .A(n16906), .B(n23342), .Z(n23340) );
  XNOR U24731 ( .A(n16905), .B(n23341), .Z(n23342) );
  NAND U24732 ( .A(n23343), .B(n[659]), .Z(n16905) );
  NAND U24733 ( .A(n21523), .B(n[659]), .Z(n23343) );
  XNOR U24734 ( .A(n23344), .B(n23341), .Z(n16906) );
  XOR U24735 ( .A(n23345), .B(n23346), .Z(n23341) );
  AND U24736 ( .A(n16913), .B(n23347), .Z(n23345) );
  XNOR U24737 ( .A(n16912), .B(n23346), .Z(n23347) );
  NAND U24738 ( .A(n23348), .B(n[658]), .Z(n16912) );
  NAND U24739 ( .A(n21523), .B(n[658]), .Z(n23348) );
  XNOR U24740 ( .A(n23349), .B(n23346), .Z(n16913) );
  XOR U24741 ( .A(n23350), .B(n23351), .Z(n23346) );
  AND U24742 ( .A(n16920), .B(n23352), .Z(n23350) );
  XNOR U24743 ( .A(n16919), .B(n23351), .Z(n23352) );
  NAND U24744 ( .A(n23353), .B(n[657]), .Z(n16919) );
  NAND U24745 ( .A(n21523), .B(n[657]), .Z(n23353) );
  XNOR U24746 ( .A(n23354), .B(n23351), .Z(n16920) );
  XOR U24747 ( .A(n23355), .B(n23356), .Z(n23351) );
  AND U24748 ( .A(n16927), .B(n23357), .Z(n23355) );
  XNOR U24749 ( .A(n16926), .B(n23356), .Z(n23357) );
  NAND U24750 ( .A(n23358), .B(n[656]), .Z(n16926) );
  NAND U24751 ( .A(n21523), .B(n[656]), .Z(n23358) );
  XNOR U24752 ( .A(n23359), .B(n23356), .Z(n16927) );
  XOR U24753 ( .A(n23360), .B(n23361), .Z(n23356) );
  AND U24754 ( .A(n16934), .B(n23362), .Z(n23360) );
  XNOR U24755 ( .A(n16933), .B(n23361), .Z(n23362) );
  NAND U24756 ( .A(n23363), .B(n[655]), .Z(n16933) );
  NAND U24757 ( .A(n21523), .B(n[655]), .Z(n23363) );
  XNOR U24758 ( .A(n23364), .B(n23361), .Z(n16934) );
  XOR U24759 ( .A(n23365), .B(n23366), .Z(n23361) );
  AND U24760 ( .A(n16941), .B(n23367), .Z(n23365) );
  XNOR U24761 ( .A(n16940), .B(n23366), .Z(n23367) );
  NAND U24762 ( .A(n23368), .B(n[654]), .Z(n16940) );
  NAND U24763 ( .A(n21523), .B(n[654]), .Z(n23368) );
  XNOR U24764 ( .A(n23369), .B(n23366), .Z(n16941) );
  XOR U24765 ( .A(n23370), .B(n23371), .Z(n23366) );
  AND U24766 ( .A(n16948), .B(n23372), .Z(n23370) );
  XNOR U24767 ( .A(n16947), .B(n23371), .Z(n23372) );
  NAND U24768 ( .A(n23373), .B(n[653]), .Z(n16947) );
  NAND U24769 ( .A(n21523), .B(n[653]), .Z(n23373) );
  XNOR U24770 ( .A(n23374), .B(n23371), .Z(n16948) );
  XOR U24771 ( .A(n23375), .B(n23376), .Z(n23371) );
  AND U24772 ( .A(n16955), .B(n23377), .Z(n23375) );
  XNOR U24773 ( .A(n16954), .B(n23376), .Z(n23377) );
  NAND U24774 ( .A(n23378), .B(n[652]), .Z(n16954) );
  NAND U24775 ( .A(n21523), .B(n[652]), .Z(n23378) );
  XNOR U24776 ( .A(n23379), .B(n23376), .Z(n16955) );
  XOR U24777 ( .A(n23380), .B(n23381), .Z(n23376) );
  AND U24778 ( .A(n16962), .B(n23382), .Z(n23380) );
  XNOR U24779 ( .A(n16961), .B(n23381), .Z(n23382) );
  NAND U24780 ( .A(n23383), .B(n[651]), .Z(n16961) );
  NAND U24781 ( .A(n21523), .B(n[651]), .Z(n23383) );
  XNOR U24782 ( .A(n23384), .B(n23381), .Z(n16962) );
  XOR U24783 ( .A(n23385), .B(n23386), .Z(n23381) );
  AND U24784 ( .A(n16969), .B(n23387), .Z(n23385) );
  XNOR U24785 ( .A(n16968), .B(n23386), .Z(n23387) );
  NAND U24786 ( .A(n23388), .B(n[650]), .Z(n16968) );
  NAND U24787 ( .A(n21523), .B(n[650]), .Z(n23388) );
  XNOR U24788 ( .A(n23389), .B(n23386), .Z(n16969) );
  XOR U24789 ( .A(n23390), .B(n23391), .Z(n23386) );
  AND U24790 ( .A(n16976), .B(n23392), .Z(n23390) );
  XNOR U24791 ( .A(n16975), .B(n23391), .Z(n23392) );
  NAND U24792 ( .A(n23393), .B(n[649]), .Z(n16975) );
  NAND U24793 ( .A(n21523), .B(n[649]), .Z(n23393) );
  XNOR U24794 ( .A(n23394), .B(n23391), .Z(n16976) );
  XOR U24795 ( .A(n23395), .B(n23396), .Z(n23391) );
  AND U24796 ( .A(n16983), .B(n23397), .Z(n23395) );
  XNOR U24797 ( .A(n16982), .B(n23396), .Z(n23397) );
  NAND U24798 ( .A(n23398), .B(n[648]), .Z(n16982) );
  NAND U24799 ( .A(n21523), .B(n[648]), .Z(n23398) );
  XNOR U24800 ( .A(n23399), .B(n23396), .Z(n16983) );
  XOR U24801 ( .A(n23400), .B(n23401), .Z(n23396) );
  AND U24802 ( .A(n16990), .B(n23402), .Z(n23400) );
  XNOR U24803 ( .A(n16989), .B(n23401), .Z(n23402) );
  NAND U24804 ( .A(n23403), .B(n[647]), .Z(n16989) );
  NAND U24805 ( .A(n21523), .B(n[647]), .Z(n23403) );
  XNOR U24806 ( .A(n23404), .B(n23401), .Z(n16990) );
  XOR U24807 ( .A(n23405), .B(n23406), .Z(n23401) );
  AND U24808 ( .A(n16997), .B(n23407), .Z(n23405) );
  XNOR U24809 ( .A(n16996), .B(n23406), .Z(n23407) );
  NAND U24810 ( .A(n23408), .B(n[646]), .Z(n16996) );
  NAND U24811 ( .A(n21523), .B(n[646]), .Z(n23408) );
  XNOR U24812 ( .A(n23409), .B(n23406), .Z(n16997) );
  XOR U24813 ( .A(n23410), .B(n23411), .Z(n23406) );
  AND U24814 ( .A(n17004), .B(n23412), .Z(n23410) );
  XNOR U24815 ( .A(n17003), .B(n23411), .Z(n23412) );
  NAND U24816 ( .A(n23413), .B(n[645]), .Z(n17003) );
  NAND U24817 ( .A(n21523), .B(n[645]), .Z(n23413) );
  XNOR U24818 ( .A(n23414), .B(n23411), .Z(n17004) );
  XOR U24819 ( .A(n23415), .B(n23416), .Z(n23411) );
  AND U24820 ( .A(n17011), .B(n23417), .Z(n23415) );
  XNOR U24821 ( .A(n17010), .B(n23416), .Z(n23417) );
  NAND U24822 ( .A(n23418), .B(n[644]), .Z(n17010) );
  NAND U24823 ( .A(n21523), .B(n[644]), .Z(n23418) );
  XNOR U24824 ( .A(n23419), .B(n23416), .Z(n17011) );
  XOR U24825 ( .A(n23420), .B(n23421), .Z(n23416) );
  AND U24826 ( .A(n17018), .B(n23422), .Z(n23420) );
  XNOR U24827 ( .A(n17017), .B(n23421), .Z(n23422) );
  NAND U24828 ( .A(n23423), .B(n[643]), .Z(n17017) );
  NAND U24829 ( .A(n21523), .B(n[643]), .Z(n23423) );
  XNOR U24830 ( .A(n23424), .B(n23421), .Z(n17018) );
  XOR U24831 ( .A(n23425), .B(n23426), .Z(n23421) );
  AND U24832 ( .A(n17025), .B(n23427), .Z(n23425) );
  XNOR U24833 ( .A(n17024), .B(n23426), .Z(n23427) );
  NAND U24834 ( .A(n23428), .B(n[642]), .Z(n17024) );
  NAND U24835 ( .A(n21523), .B(n[642]), .Z(n23428) );
  XNOR U24836 ( .A(n23429), .B(n23426), .Z(n17025) );
  XOR U24837 ( .A(n23430), .B(n23431), .Z(n23426) );
  AND U24838 ( .A(n17032), .B(n23432), .Z(n23430) );
  XNOR U24839 ( .A(n17031), .B(n23431), .Z(n23432) );
  NAND U24840 ( .A(n23433), .B(n[641]), .Z(n17031) );
  NAND U24841 ( .A(n21523), .B(n[641]), .Z(n23433) );
  XNOR U24842 ( .A(n23434), .B(n23431), .Z(n17032) );
  XOR U24843 ( .A(n23435), .B(n23436), .Z(n23431) );
  AND U24844 ( .A(n17039), .B(n23437), .Z(n23435) );
  XNOR U24845 ( .A(n17038), .B(n23436), .Z(n23437) );
  NAND U24846 ( .A(n23438), .B(n[640]), .Z(n17038) );
  NAND U24847 ( .A(n21523), .B(n[640]), .Z(n23438) );
  XNOR U24848 ( .A(n23439), .B(n23436), .Z(n17039) );
  XOR U24849 ( .A(n23440), .B(n23441), .Z(n23436) );
  AND U24850 ( .A(n17046), .B(n23442), .Z(n23440) );
  XNOR U24851 ( .A(n17045), .B(n23441), .Z(n23442) );
  NAND U24852 ( .A(n23443), .B(n[639]), .Z(n17045) );
  NAND U24853 ( .A(n21523), .B(n[639]), .Z(n23443) );
  XNOR U24854 ( .A(n23444), .B(n23441), .Z(n17046) );
  XOR U24855 ( .A(n23445), .B(n23446), .Z(n23441) );
  AND U24856 ( .A(n17053), .B(n23447), .Z(n23445) );
  XNOR U24857 ( .A(n17052), .B(n23446), .Z(n23447) );
  NAND U24858 ( .A(n23448), .B(n[638]), .Z(n17052) );
  NAND U24859 ( .A(n21523), .B(n[638]), .Z(n23448) );
  XNOR U24860 ( .A(n23449), .B(n23446), .Z(n17053) );
  XOR U24861 ( .A(n23450), .B(n23451), .Z(n23446) );
  AND U24862 ( .A(n17060), .B(n23452), .Z(n23450) );
  XNOR U24863 ( .A(n17059), .B(n23451), .Z(n23452) );
  NAND U24864 ( .A(n23453), .B(n[637]), .Z(n17059) );
  NAND U24865 ( .A(n21523), .B(n[637]), .Z(n23453) );
  XNOR U24866 ( .A(n23454), .B(n23451), .Z(n17060) );
  XOR U24867 ( .A(n23455), .B(n23456), .Z(n23451) );
  AND U24868 ( .A(n17067), .B(n23457), .Z(n23455) );
  XNOR U24869 ( .A(n17066), .B(n23456), .Z(n23457) );
  NAND U24870 ( .A(n23458), .B(n[636]), .Z(n17066) );
  NAND U24871 ( .A(n21523), .B(n[636]), .Z(n23458) );
  XNOR U24872 ( .A(n23459), .B(n23456), .Z(n17067) );
  XOR U24873 ( .A(n23460), .B(n23461), .Z(n23456) );
  AND U24874 ( .A(n17074), .B(n23462), .Z(n23460) );
  XNOR U24875 ( .A(n17073), .B(n23461), .Z(n23462) );
  NAND U24876 ( .A(n23463), .B(n[635]), .Z(n17073) );
  NAND U24877 ( .A(n21523), .B(n[635]), .Z(n23463) );
  XNOR U24878 ( .A(n23464), .B(n23461), .Z(n17074) );
  XOR U24879 ( .A(n23465), .B(n23466), .Z(n23461) );
  AND U24880 ( .A(n17081), .B(n23467), .Z(n23465) );
  XNOR U24881 ( .A(n17080), .B(n23466), .Z(n23467) );
  NAND U24882 ( .A(n23468), .B(n[634]), .Z(n17080) );
  NAND U24883 ( .A(n21523), .B(n[634]), .Z(n23468) );
  XNOR U24884 ( .A(n23469), .B(n23466), .Z(n17081) );
  XOR U24885 ( .A(n23470), .B(n23471), .Z(n23466) );
  AND U24886 ( .A(n17088), .B(n23472), .Z(n23470) );
  XNOR U24887 ( .A(n17087), .B(n23471), .Z(n23472) );
  NAND U24888 ( .A(n23473), .B(n[633]), .Z(n17087) );
  NAND U24889 ( .A(n21523), .B(n[633]), .Z(n23473) );
  XNOR U24890 ( .A(n23474), .B(n23471), .Z(n17088) );
  XOR U24891 ( .A(n23475), .B(n23476), .Z(n23471) );
  AND U24892 ( .A(n17095), .B(n23477), .Z(n23475) );
  XNOR U24893 ( .A(n17094), .B(n23476), .Z(n23477) );
  NAND U24894 ( .A(n23478), .B(n[632]), .Z(n17094) );
  NAND U24895 ( .A(n21523), .B(n[632]), .Z(n23478) );
  XNOR U24896 ( .A(n23479), .B(n23476), .Z(n17095) );
  XOR U24897 ( .A(n23480), .B(n23481), .Z(n23476) );
  AND U24898 ( .A(n17102), .B(n23482), .Z(n23480) );
  XNOR U24899 ( .A(n17101), .B(n23481), .Z(n23482) );
  NAND U24900 ( .A(n23483), .B(n[631]), .Z(n17101) );
  NAND U24901 ( .A(n21523), .B(n[631]), .Z(n23483) );
  XNOR U24902 ( .A(n23484), .B(n23481), .Z(n17102) );
  XOR U24903 ( .A(n23485), .B(n23486), .Z(n23481) );
  AND U24904 ( .A(n17109), .B(n23487), .Z(n23485) );
  XNOR U24905 ( .A(n17108), .B(n23486), .Z(n23487) );
  NAND U24906 ( .A(n23488), .B(n[630]), .Z(n17108) );
  NAND U24907 ( .A(n21523), .B(n[630]), .Z(n23488) );
  XNOR U24908 ( .A(n23489), .B(n23486), .Z(n17109) );
  XOR U24909 ( .A(n23490), .B(n23491), .Z(n23486) );
  AND U24910 ( .A(n17116), .B(n23492), .Z(n23490) );
  XNOR U24911 ( .A(n17115), .B(n23491), .Z(n23492) );
  NAND U24912 ( .A(n23493), .B(n[629]), .Z(n17115) );
  NAND U24913 ( .A(n21523), .B(n[629]), .Z(n23493) );
  XNOR U24914 ( .A(n23494), .B(n23491), .Z(n17116) );
  XOR U24915 ( .A(n23495), .B(n23496), .Z(n23491) );
  AND U24916 ( .A(n17123), .B(n23497), .Z(n23495) );
  XNOR U24917 ( .A(n17122), .B(n23496), .Z(n23497) );
  NAND U24918 ( .A(n23498), .B(n[628]), .Z(n17122) );
  NAND U24919 ( .A(n21523), .B(n[628]), .Z(n23498) );
  XNOR U24920 ( .A(n23499), .B(n23496), .Z(n17123) );
  XOR U24921 ( .A(n23500), .B(n23501), .Z(n23496) );
  AND U24922 ( .A(n17130), .B(n23502), .Z(n23500) );
  XNOR U24923 ( .A(n17129), .B(n23501), .Z(n23502) );
  NAND U24924 ( .A(n23503), .B(n[627]), .Z(n17129) );
  NAND U24925 ( .A(n21523), .B(n[627]), .Z(n23503) );
  XNOR U24926 ( .A(n23504), .B(n23501), .Z(n17130) );
  XOR U24927 ( .A(n23505), .B(n23506), .Z(n23501) );
  AND U24928 ( .A(n17137), .B(n23507), .Z(n23505) );
  XNOR U24929 ( .A(n17136), .B(n23506), .Z(n23507) );
  NAND U24930 ( .A(n23508), .B(n[626]), .Z(n17136) );
  NAND U24931 ( .A(n21523), .B(n[626]), .Z(n23508) );
  XNOR U24932 ( .A(n23509), .B(n23506), .Z(n17137) );
  XOR U24933 ( .A(n23510), .B(n23511), .Z(n23506) );
  AND U24934 ( .A(n17144), .B(n23512), .Z(n23510) );
  XNOR U24935 ( .A(n17143), .B(n23511), .Z(n23512) );
  NAND U24936 ( .A(n23513), .B(n[625]), .Z(n17143) );
  NAND U24937 ( .A(n21523), .B(n[625]), .Z(n23513) );
  XNOR U24938 ( .A(n23514), .B(n23511), .Z(n17144) );
  XOR U24939 ( .A(n23515), .B(n23516), .Z(n23511) );
  AND U24940 ( .A(n17151), .B(n23517), .Z(n23515) );
  XNOR U24941 ( .A(n17150), .B(n23516), .Z(n23517) );
  NAND U24942 ( .A(n23518), .B(n[624]), .Z(n17150) );
  NAND U24943 ( .A(n21523), .B(n[624]), .Z(n23518) );
  XNOR U24944 ( .A(n23519), .B(n23516), .Z(n17151) );
  XOR U24945 ( .A(n23520), .B(n23521), .Z(n23516) );
  AND U24946 ( .A(n17158), .B(n23522), .Z(n23520) );
  XNOR U24947 ( .A(n17157), .B(n23521), .Z(n23522) );
  NAND U24948 ( .A(n23523), .B(n[623]), .Z(n17157) );
  NAND U24949 ( .A(n21523), .B(n[623]), .Z(n23523) );
  XNOR U24950 ( .A(n23524), .B(n23521), .Z(n17158) );
  XOR U24951 ( .A(n23525), .B(n23526), .Z(n23521) );
  AND U24952 ( .A(n17165), .B(n23527), .Z(n23525) );
  XNOR U24953 ( .A(n17164), .B(n23526), .Z(n23527) );
  NAND U24954 ( .A(n23528), .B(n[622]), .Z(n17164) );
  NAND U24955 ( .A(n21523), .B(n[622]), .Z(n23528) );
  XNOR U24956 ( .A(n23529), .B(n23526), .Z(n17165) );
  XOR U24957 ( .A(n23530), .B(n23531), .Z(n23526) );
  AND U24958 ( .A(n17172), .B(n23532), .Z(n23530) );
  XNOR U24959 ( .A(n17171), .B(n23531), .Z(n23532) );
  NAND U24960 ( .A(n23533), .B(n[621]), .Z(n17171) );
  NAND U24961 ( .A(n21523), .B(n[621]), .Z(n23533) );
  XNOR U24962 ( .A(n23534), .B(n23531), .Z(n17172) );
  XOR U24963 ( .A(n23535), .B(n23536), .Z(n23531) );
  AND U24964 ( .A(n17179), .B(n23537), .Z(n23535) );
  XNOR U24965 ( .A(n17178), .B(n23536), .Z(n23537) );
  NAND U24966 ( .A(n23538), .B(n[620]), .Z(n17178) );
  NAND U24967 ( .A(n21523), .B(n[620]), .Z(n23538) );
  XNOR U24968 ( .A(n23539), .B(n23536), .Z(n17179) );
  XOR U24969 ( .A(n23540), .B(n23541), .Z(n23536) );
  AND U24970 ( .A(n17186), .B(n23542), .Z(n23540) );
  XNOR U24971 ( .A(n17185), .B(n23541), .Z(n23542) );
  NAND U24972 ( .A(n23543), .B(n[619]), .Z(n17185) );
  NAND U24973 ( .A(n21523), .B(n[619]), .Z(n23543) );
  XNOR U24974 ( .A(n23544), .B(n23541), .Z(n17186) );
  XOR U24975 ( .A(n23545), .B(n23546), .Z(n23541) );
  AND U24976 ( .A(n17193), .B(n23547), .Z(n23545) );
  XNOR U24977 ( .A(n17192), .B(n23546), .Z(n23547) );
  NAND U24978 ( .A(n23548), .B(n[618]), .Z(n17192) );
  NAND U24979 ( .A(n21523), .B(n[618]), .Z(n23548) );
  XNOR U24980 ( .A(n23549), .B(n23546), .Z(n17193) );
  XOR U24981 ( .A(n23550), .B(n23551), .Z(n23546) );
  AND U24982 ( .A(n17200), .B(n23552), .Z(n23550) );
  XNOR U24983 ( .A(n17199), .B(n23551), .Z(n23552) );
  NAND U24984 ( .A(n23553), .B(n[617]), .Z(n17199) );
  NAND U24985 ( .A(n21523), .B(n[617]), .Z(n23553) );
  XNOR U24986 ( .A(n23554), .B(n23551), .Z(n17200) );
  XOR U24987 ( .A(n23555), .B(n23556), .Z(n23551) );
  AND U24988 ( .A(n17207), .B(n23557), .Z(n23555) );
  XNOR U24989 ( .A(n17206), .B(n23556), .Z(n23557) );
  NAND U24990 ( .A(n23558), .B(n[616]), .Z(n17206) );
  NAND U24991 ( .A(n21523), .B(n[616]), .Z(n23558) );
  XNOR U24992 ( .A(n23559), .B(n23556), .Z(n17207) );
  XOR U24993 ( .A(n23560), .B(n23561), .Z(n23556) );
  AND U24994 ( .A(n17214), .B(n23562), .Z(n23560) );
  XNOR U24995 ( .A(n17213), .B(n23561), .Z(n23562) );
  NAND U24996 ( .A(n23563), .B(n[615]), .Z(n17213) );
  NAND U24997 ( .A(n21523), .B(n[615]), .Z(n23563) );
  XNOR U24998 ( .A(n23564), .B(n23561), .Z(n17214) );
  XOR U24999 ( .A(n23565), .B(n23566), .Z(n23561) );
  AND U25000 ( .A(n17221), .B(n23567), .Z(n23565) );
  XNOR U25001 ( .A(n17220), .B(n23566), .Z(n23567) );
  NAND U25002 ( .A(n23568), .B(n[614]), .Z(n17220) );
  NAND U25003 ( .A(n21523), .B(n[614]), .Z(n23568) );
  XNOR U25004 ( .A(n23569), .B(n23566), .Z(n17221) );
  XOR U25005 ( .A(n23570), .B(n23571), .Z(n23566) );
  AND U25006 ( .A(n17228), .B(n23572), .Z(n23570) );
  XNOR U25007 ( .A(n17227), .B(n23571), .Z(n23572) );
  NAND U25008 ( .A(n23573), .B(n[613]), .Z(n17227) );
  NAND U25009 ( .A(n21523), .B(n[613]), .Z(n23573) );
  XNOR U25010 ( .A(n23574), .B(n23571), .Z(n17228) );
  XOR U25011 ( .A(n23575), .B(n23576), .Z(n23571) );
  AND U25012 ( .A(n17235), .B(n23577), .Z(n23575) );
  XNOR U25013 ( .A(n17234), .B(n23576), .Z(n23577) );
  NAND U25014 ( .A(n23578), .B(n[612]), .Z(n17234) );
  NAND U25015 ( .A(n21523), .B(n[612]), .Z(n23578) );
  XNOR U25016 ( .A(n23579), .B(n23576), .Z(n17235) );
  XOR U25017 ( .A(n23580), .B(n23581), .Z(n23576) );
  AND U25018 ( .A(n17242), .B(n23582), .Z(n23580) );
  XNOR U25019 ( .A(n17241), .B(n23581), .Z(n23582) );
  NAND U25020 ( .A(n23583), .B(n[611]), .Z(n17241) );
  NAND U25021 ( .A(n21523), .B(n[611]), .Z(n23583) );
  XNOR U25022 ( .A(n23584), .B(n23581), .Z(n17242) );
  XOR U25023 ( .A(n23585), .B(n23586), .Z(n23581) );
  AND U25024 ( .A(n17249), .B(n23587), .Z(n23585) );
  XNOR U25025 ( .A(n17248), .B(n23586), .Z(n23587) );
  NAND U25026 ( .A(n23588), .B(n[610]), .Z(n17248) );
  NAND U25027 ( .A(n21523), .B(n[610]), .Z(n23588) );
  XNOR U25028 ( .A(n23589), .B(n23586), .Z(n17249) );
  XOR U25029 ( .A(n23590), .B(n23591), .Z(n23586) );
  AND U25030 ( .A(n17256), .B(n23592), .Z(n23590) );
  XNOR U25031 ( .A(n17255), .B(n23591), .Z(n23592) );
  NAND U25032 ( .A(n23593), .B(n[609]), .Z(n17255) );
  NAND U25033 ( .A(n21523), .B(n[609]), .Z(n23593) );
  XNOR U25034 ( .A(n23594), .B(n23591), .Z(n17256) );
  XOR U25035 ( .A(n23595), .B(n23596), .Z(n23591) );
  AND U25036 ( .A(n17263), .B(n23597), .Z(n23595) );
  XNOR U25037 ( .A(n17262), .B(n23596), .Z(n23597) );
  NAND U25038 ( .A(n23598), .B(n[608]), .Z(n17262) );
  NAND U25039 ( .A(n21523), .B(n[608]), .Z(n23598) );
  XNOR U25040 ( .A(n23599), .B(n23596), .Z(n17263) );
  XOR U25041 ( .A(n23600), .B(n23601), .Z(n23596) );
  AND U25042 ( .A(n17270), .B(n23602), .Z(n23600) );
  XNOR U25043 ( .A(n17269), .B(n23601), .Z(n23602) );
  NAND U25044 ( .A(n23603), .B(n[607]), .Z(n17269) );
  NAND U25045 ( .A(n21523), .B(n[607]), .Z(n23603) );
  XNOR U25046 ( .A(n23604), .B(n23601), .Z(n17270) );
  XOR U25047 ( .A(n23605), .B(n23606), .Z(n23601) );
  AND U25048 ( .A(n17277), .B(n23607), .Z(n23605) );
  XNOR U25049 ( .A(n17276), .B(n23606), .Z(n23607) );
  NAND U25050 ( .A(n23608), .B(n[606]), .Z(n17276) );
  NAND U25051 ( .A(n21523), .B(n[606]), .Z(n23608) );
  XNOR U25052 ( .A(n23609), .B(n23606), .Z(n17277) );
  XOR U25053 ( .A(n23610), .B(n23611), .Z(n23606) );
  AND U25054 ( .A(n17284), .B(n23612), .Z(n23610) );
  XNOR U25055 ( .A(n17283), .B(n23611), .Z(n23612) );
  NAND U25056 ( .A(n23613), .B(n[605]), .Z(n17283) );
  NAND U25057 ( .A(n21523), .B(n[605]), .Z(n23613) );
  XNOR U25058 ( .A(n23614), .B(n23611), .Z(n17284) );
  XOR U25059 ( .A(n23615), .B(n23616), .Z(n23611) );
  AND U25060 ( .A(n17291), .B(n23617), .Z(n23615) );
  XNOR U25061 ( .A(n17290), .B(n23616), .Z(n23617) );
  NAND U25062 ( .A(n23618), .B(n[604]), .Z(n17290) );
  NAND U25063 ( .A(n21523), .B(n[604]), .Z(n23618) );
  XNOR U25064 ( .A(n23619), .B(n23616), .Z(n17291) );
  XOR U25065 ( .A(n23620), .B(n23621), .Z(n23616) );
  AND U25066 ( .A(n17298), .B(n23622), .Z(n23620) );
  XNOR U25067 ( .A(n17297), .B(n23621), .Z(n23622) );
  NAND U25068 ( .A(n23623), .B(n[603]), .Z(n17297) );
  NAND U25069 ( .A(n21523), .B(n[603]), .Z(n23623) );
  XNOR U25070 ( .A(n23624), .B(n23621), .Z(n17298) );
  XOR U25071 ( .A(n23625), .B(n23626), .Z(n23621) );
  AND U25072 ( .A(n17305), .B(n23627), .Z(n23625) );
  XNOR U25073 ( .A(n17304), .B(n23626), .Z(n23627) );
  NAND U25074 ( .A(n23628), .B(n[602]), .Z(n17304) );
  NAND U25075 ( .A(n21523), .B(n[602]), .Z(n23628) );
  XNOR U25076 ( .A(n23629), .B(n23626), .Z(n17305) );
  XOR U25077 ( .A(n23630), .B(n23631), .Z(n23626) );
  AND U25078 ( .A(n17312), .B(n23632), .Z(n23630) );
  XNOR U25079 ( .A(n17311), .B(n23631), .Z(n23632) );
  NAND U25080 ( .A(n23633), .B(n[601]), .Z(n17311) );
  NAND U25081 ( .A(n21523), .B(n[601]), .Z(n23633) );
  XNOR U25082 ( .A(n23634), .B(n23631), .Z(n17312) );
  XOR U25083 ( .A(n23635), .B(n23636), .Z(n23631) );
  AND U25084 ( .A(n17319), .B(n23637), .Z(n23635) );
  XNOR U25085 ( .A(n17318), .B(n23636), .Z(n23637) );
  NAND U25086 ( .A(n23638), .B(n[600]), .Z(n17318) );
  NAND U25087 ( .A(n21523), .B(n[600]), .Z(n23638) );
  XNOR U25088 ( .A(n23639), .B(n23636), .Z(n17319) );
  XOR U25089 ( .A(n23640), .B(n23641), .Z(n23636) );
  AND U25090 ( .A(n17326), .B(n23642), .Z(n23640) );
  XNOR U25091 ( .A(n17325), .B(n23641), .Z(n23642) );
  NAND U25092 ( .A(n23643), .B(n[599]), .Z(n17325) );
  NAND U25093 ( .A(n21523), .B(n[599]), .Z(n23643) );
  XNOR U25094 ( .A(n23644), .B(n23641), .Z(n17326) );
  XOR U25095 ( .A(n23645), .B(n23646), .Z(n23641) );
  AND U25096 ( .A(n17333), .B(n23647), .Z(n23645) );
  XNOR U25097 ( .A(n17332), .B(n23646), .Z(n23647) );
  NAND U25098 ( .A(n23648), .B(n[598]), .Z(n17332) );
  NAND U25099 ( .A(n21523), .B(n[598]), .Z(n23648) );
  XNOR U25100 ( .A(n23649), .B(n23646), .Z(n17333) );
  XOR U25101 ( .A(n23650), .B(n23651), .Z(n23646) );
  AND U25102 ( .A(n17340), .B(n23652), .Z(n23650) );
  XNOR U25103 ( .A(n17339), .B(n23651), .Z(n23652) );
  NAND U25104 ( .A(n23653), .B(n[597]), .Z(n17339) );
  NAND U25105 ( .A(n21523), .B(n[597]), .Z(n23653) );
  XNOR U25106 ( .A(n23654), .B(n23651), .Z(n17340) );
  XOR U25107 ( .A(n23655), .B(n23656), .Z(n23651) );
  AND U25108 ( .A(n17347), .B(n23657), .Z(n23655) );
  XNOR U25109 ( .A(n17346), .B(n23656), .Z(n23657) );
  NAND U25110 ( .A(n23658), .B(n[596]), .Z(n17346) );
  NAND U25111 ( .A(n21523), .B(n[596]), .Z(n23658) );
  XNOR U25112 ( .A(n23659), .B(n23656), .Z(n17347) );
  XOR U25113 ( .A(n23660), .B(n23661), .Z(n23656) );
  AND U25114 ( .A(n17354), .B(n23662), .Z(n23660) );
  XNOR U25115 ( .A(n17353), .B(n23661), .Z(n23662) );
  NAND U25116 ( .A(n23663), .B(n[595]), .Z(n17353) );
  NAND U25117 ( .A(n21523), .B(n[595]), .Z(n23663) );
  XNOR U25118 ( .A(n23664), .B(n23661), .Z(n17354) );
  XOR U25119 ( .A(n23665), .B(n23666), .Z(n23661) );
  AND U25120 ( .A(n17361), .B(n23667), .Z(n23665) );
  XNOR U25121 ( .A(n17360), .B(n23666), .Z(n23667) );
  NAND U25122 ( .A(n23668), .B(n[594]), .Z(n17360) );
  NAND U25123 ( .A(n21523), .B(n[594]), .Z(n23668) );
  XNOR U25124 ( .A(n23669), .B(n23666), .Z(n17361) );
  XOR U25125 ( .A(n23670), .B(n23671), .Z(n23666) );
  AND U25126 ( .A(n17368), .B(n23672), .Z(n23670) );
  XNOR U25127 ( .A(n17367), .B(n23671), .Z(n23672) );
  NAND U25128 ( .A(n23673), .B(n[593]), .Z(n17367) );
  NAND U25129 ( .A(n21523), .B(n[593]), .Z(n23673) );
  XNOR U25130 ( .A(n23674), .B(n23671), .Z(n17368) );
  XOR U25131 ( .A(n23675), .B(n23676), .Z(n23671) );
  AND U25132 ( .A(n17375), .B(n23677), .Z(n23675) );
  XNOR U25133 ( .A(n17374), .B(n23676), .Z(n23677) );
  NAND U25134 ( .A(n23678), .B(n[592]), .Z(n17374) );
  NAND U25135 ( .A(n21523), .B(n[592]), .Z(n23678) );
  XNOR U25136 ( .A(n23679), .B(n23676), .Z(n17375) );
  XOR U25137 ( .A(n23680), .B(n23681), .Z(n23676) );
  AND U25138 ( .A(n17382), .B(n23682), .Z(n23680) );
  XNOR U25139 ( .A(n17381), .B(n23681), .Z(n23682) );
  NAND U25140 ( .A(n23683), .B(n[591]), .Z(n17381) );
  NAND U25141 ( .A(n21523), .B(n[591]), .Z(n23683) );
  XNOR U25142 ( .A(n23684), .B(n23681), .Z(n17382) );
  XOR U25143 ( .A(n23685), .B(n23686), .Z(n23681) );
  AND U25144 ( .A(n17389), .B(n23687), .Z(n23685) );
  XNOR U25145 ( .A(n17388), .B(n23686), .Z(n23687) );
  NAND U25146 ( .A(n23688), .B(n[590]), .Z(n17388) );
  NAND U25147 ( .A(n21523), .B(n[590]), .Z(n23688) );
  XNOR U25148 ( .A(n23689), .B(n23686), .Z(n17389) );
  XOR U25149 ( .A(n23690), .B(n23691), .Z(n23686) );
  AND U25150 ( .A(n17396), .B(n23692), .Z(n23690) );
  XNOR U25151 ( .A(n17395), .B(n23691), .Z(n23692) );
  NAND U25152 ( .A(n23693), .B(n[589]), .Z(n17395) );
  NAND U25153 ( .A(n21523), .B(n[589]), .Z(n23693) );
  XNOR U25154 ( .A(n23694), .B(n23691), .Z(n17396) );
  XOR U25155 ( .A(n23695), .B(n23696), .Z(n23691) );
  AND U25156 ( .A(n17403), .B(n23697), .Z(n23695) );
  XNOR U25157 ( .A(n17402), .B(n23696), .Z(n23697) );
  NAND U25158 ( .A(n23698), .B(n[588]), .Z(n17402) );
  NAND U25159 ( .A(n21523), .B(n[588]), .Z(n23698) );
  XNOR U25160 ( .A(n23699), .B(n23696), .Z(n17403) );
  XOR U25161 ( .A(n23700), .B(n23701), .Z(n23696) );
  AND U25162 ( .A(n17410), .B(n23702), .Z(n23700) );
  XNOR U25163 ( .A(n17409), .B(n23701), .Z(n23702) );
  NAND U25164 ( .A(n23703), .B(n[587]), .Z(n17409) );
  NAND U25165 ( .A(n21523), .B(n[587]), .Z(n23703) );
  XNOR U25166 ( .A(n23704), .B(n23701), .Z(n17410) );
  XOR U25167 ( .A(n23705), .B(n23706), .Z(n23701) );
  AND U25168 ( .A(n17417), .B(n23707), .Z(n23705) );
  XNOR U25169 ( .A(n17416), .B(n23706), .Z(n23707) );
  NAND U25170 ( .A(n23708), .B(n[586]), .Z(n17416) );
  NAND U25171 ( .A(n21523), .B(n[586]), .Z(n23708) );
  XNOR U25172 ( .A(n23709), .B(n23706), .Z(n17417) );
  XOR U25173 ( .A(n23710), .B(n23711), .Z(n23706) );
  AND U25174 ( .A(n17424), .B(n23712), .Z(n23710) );
  XNOR U25175 ( .A(n17423), .B(n23711), .Z(n23712) );
  NAND U25176 ( .A(n23713), .B(n[585]), .Z(n17423) );
  NAND U25177 ( .A(n21523), .B(n[585]), .Z(n23713) );
  XNOR U25178 ( .A(n23714), .B(n23711), .Z(n17424) );
  XOR U25179 ( .A(n23715), .B(n23716), .Z(n23711) );
  AND U25180 ( .A(n17431), .B(n23717), .Z(n23715) );
  XNOR U25181 ( .A(n17430), .B(n23716), .Z(n23717) );
  NAND U25182 ( .A(n23718), .B(n[584]), .Z(n17430) );
  NAND U25183 ( .A(n21523), .B(n[584]), .Z(n23718) );
  XNOR U25184 ( .A(n23719), .B(n23716), .Z(n17431) );
  XOR U25185 ( .A(n23720), .B(n23721), .Z(n23716) );
  AND U25186 ( .A(n17438), .B(n23722), .Z(n23720) );
  XNOR U25187 ( .A(n17437), .B(n23721), .Z(n23722) );
  NAND U25188 ( .A(n23723), .B(n[583]), .Z(n17437) );
  NAND U25189 ( .A(n21523), .B(n[583]), .Z(n23723) );
  XNOR U25190 ( .A(n23724), .B(n23721), .Z(n17438) );
  XOR U25191 ( .A(n23725), .B(n23726), .Z(n23721) );
  AND U25192 ( .A(n17445), .B(n23727), .Z(n23725) );
  XNOR U25193 ( .A(n17444), .B(n23726), .Z(n23727) );
  NAND U25194 ( .A(n23728), .B(n[582]), .Z(n17444) );
  NAND U25195 ( .A(n21523), .B(n[582]), .Z(n23728) );
  XNOR U25196 ( .A(n23729), .B(n23726), .Z(n17445) );
  XOR U25197 ( .A(n23730), .B(n23731), .Z(n23726) );
  AND U25198 ( .A(n17452), .B(n23732), .Z(n23730) );
  XNOR U25199 ( .A(n17451), .B(n23731), .Z(n23732) );
  NAND U25200 ( .A(n23733), .B(n[581]), .Z(n17451) );
  NAND U25201 ( .A(n21523), .B(n[581]), .Z(n23733) );
  XNOR U25202 ( .A(n23734), .B(n23731), .Z(n17452) );
  XOR U25203 ( .A(n23735), .B(n23736), .Z(n23731) );
  AND U25204 ( .A(n17459), .B(n23737), .Z(n23735) );
  XNOR U25205 ( .A(n17458), .B(n23736), .Z(n23737) );
  NAND U25206 ( .A(n23738), .B(n[580]), .Z(n17458) );
  NAND U25207 ( .A(n21523), .B(n[580]), .Z(n23738) );
  XNOR U25208 ( .A(n23739), .B(n23736), .Z(n17459) );
  XOR U25209 ( .A(n23740), .B(n23741), .Z(n23736) );
  AND U25210 ( .A(n17466), .B(n23742), .Z(n23740) );
  XNOR U25211 ( .A(n17465), .B(n23741), .Z(n23742) );
  NAND U25212 ( .A(n23743), .B(n[579]), .Z(n17465) );
  NAND U25213 ( .A(n21523), .B(n[579]), .Z(n23743) );
  XNOR U25214 ( .A(n23744), .B(n23741), .Z(n17466) );
  XOR U25215 ( .A(n23745), .B(n23746), .Z(n23741) );
  AND U25216 ( .A(n17473), .B(n23747), .Z(n23745) );
  XNOR U25217 ( .A(n17472), .B(n23746), .Z(n23747) );
  NAND U25218 ( .A(n23748), .B(n[578]), .Z(n17472) );
  NAND U25219 ( .A(n21523), .B(n[578]), .Z(n23748) );
  XNOR U25220 ( .A(n23749), .B(n23746), .Z(n17473) );
  XOR U25221 ( .A(n23750), .B(n23751), .Z(n23746) );
  AND U25222 ( .A(n17480), .B(n23752), .Z(n23750) );
  XNOR U25223 ( .A(n17479), .B(n23751), .Z(n23752) );
  NAND U25224 ( .A(n23753), .B(n[577]), .Z(n17479) );
  NAND U25225 ( .A(n21523), .B(n[577]), .Z(n23753) );
  XNOR U25226 ( .A(n23754), .B(n23751), .Z(n17480) );
  XOR U25227 ( .A(n23755), .B(n23756), .Z(n23751) );
  AND U25228 ( .A(n17487), .B(n23757), .Z(n23755) );
  XNOR U25229 ( .A(n17486), .B(n23756), .Z(n23757) );
  NAND U25230 ( .A(n23758), .B(n[576]), .Z(n17486) );
  NAND U25231 ( .A(n21523), .B(n[576]), .Z(n23758) );
  XNOR U25232 ( .A(n23759), .B(n23756), .Z(n17487) );
  XOR U25233 ( .A(n23760), .B(n23761), .Z(n23756) );
  AND U25234 ( .A(n17494), .B(n23762), .Z(n23760) );
  XNOR U25235 ( .A(n17493), .B(n23761), .Z(n23762) );
  NAND U25236 ( .A(n23763), .B(n[575]), .Z(n17493) );
  NAND U25237 ( .A(n21523), .B(n[575]), .Z(n23763) );
  XNOR U25238 ( .A(n23764), .B(n23761), .Z(n17494) );
  XOR U25239 ( .A(n23765), .B(n23766), .Z(n23761) );
  AND U25240 ( .A(n17501), .B(n23767), .Z(n23765) );
  XNOR U25241 ( .A(n17500), .B(n23766), .Z(n23767) );
  NAND U25242 ( .A(n23768), .B(n[574]), .Z(n17500) );
  NAND U25243 ( .A(n21523), .B(n[574]), .Z(n23768) );
  XNOR U25244 ( .A(n23769), .B(n23766), .Z(n17501) );
  XOR U25245 ( .A(n23770), .B(n23771), .Z(n23766) );
  AND U25246 ( .A(n17508), .B(n23772), .Z(n23770) );
  XNOR U25247 ( .A(n17507), .B(n23771), .Z(n23772) );
  NAND U25248 ( .A(n23773), .B(n[573]), .Z(n17507) );
  NAND U25249 ( .A(n21523), .B(n[573]), .Z(n23773) );
  XNOR U25250 ( .A(n23774), .B(n23771), .Z(n17508) );
  XOR U25251 ( .A(n23775), .B(n23776), .Z(n23771) );
  AND U25252 ( .A(n17515), .B(n23777), .Z(n23775) );
  XNOR U25253 ( .A(n17514), .B(n23776), .Z(n23777) );
  NAND U25254 ( .A(n23778), .B(n[572]), .Z(n17514) );
  NAND U25255 ( .A(n21523), .B(n[572]), .Z(n23778) );
  XNOR U25256 ( .A(n23779), .B(n23776), .Z(n17515) );
  XOR U25257 ( .A(n23780), .B(n23781), .Z(n23776) );
  AND U25258 ( .A(n17522), .B(n23782), .Z(n23780) );
  XNOR U25259 ( .A(n17521), .B(n23781), .Z(n23782) );
  NAND U25260 ( .A(n23783), .B(n[571]), .Z(n17521) );
  NAND U25261 ( .A(n21523), .B(n[571]), .Z(n23783) );
  XNOR U25262 ( .A(n23784), .B(n23781), .Z(n17522) );
  XOR U25263 ( .A(n23785), .B(n23786), .Z(n23781) );
  AND U25264 ( .A(n17529), .B(n23787), .Z(n23785) );
  XNOR U25265 ( .A(n17528), .B(n23786), .Z(n23787) );
  NAND U25266 ( .A(n23788), .B(n[570]), .Z(n17528) );
  NAND U25267 ( .A(n21523), .B(n[570]), .Z(n23788) );
  XNOR U25268 ( .A(n23789), .B(n23786), .Z(n17529) );
  XOR U25269 ( .A(n23790), .B(n23791), .Z(n23786) );
  AND U25270 ( .A(n17536), .B(n23792), .Z(n23790) );
  XNOR U25271 ( .A(n17535), .B(n23791), .Z(n23792) );
  NAND U25272 ( .A(n23793), .B(n[569]), .Z(n17535) );
  NAND U25273 ( .A(n21523), .B(n[569]), .Z(n23793) );
  XNOR U25274 ( .A(n23794), .B(n23791), .Z(n17536) );
  XOR U25275 ( .A(n23795), .B(n23796), .Z(n23791) );
  AND U25276 ( .A(n17543), .B(n23797), .Z(n23795) );
  XNOR U25277 ( .A(n17542), .B(n23796), .Z(n23797) );
  NAND U25278 ( .A(n23798), .B(n[568]), .Z(n17542) );
  NAND U25279 ( .A(n21523), .B(n[568]), .Z(n23798) );
  XNOR U25280 ( .A(n23799), .B(n23796), .Z(n17543) );
  XOR U25281 ( .A(n23800), .B(n23801), .Z(n23796) );
  AND U25282 ( .A(n17550), .B(n23802), .Z(n23800) );
  XNOR U25283 ( .A(n17549), .B(n23801), .Z(n23802) );
  NAND U25284 ( .A(n23803), .B(n[567]), .Z(n17549) );
  NAND U25285 ( .A(n21523), .B(n[567]), .Z(n23803) );
  XNOR U25286 ( .A(n23804), .B(n23801), .Z(n17550) );
  XOR U25287 ( .A(n23805), .B(n23806), .Z(n23801) );
  AND U25288 ( .A(n17557), .B(n23807), .Z(n23805) );
  XNOR U25289 ( .A(n17556), .B(n23806), .Z(n23807) );
  NAND U25290 ( .A(n23808), .B(n[566]), .Z(n17556) );
  NAND U25291 ( .A(n21523), .B(n[566]), .Z(n23808) );
  XNOR U25292 ( .A(n23809), .B(n23806), .Z(n17557) );
  XOR U25293 ( .A(n23810), .B(n23811), .Z(n23806) );
  AND U25294 ( .A(n17564), .B(n23812), .Z(n23810) );
  XNOR U25295 ( .A(n17563), .B(n23811), .Z(n23812) );
  NAND U25296 ( .A(n23813), .B(n[565]), .Z(n17563) );
  NAND U25297 ( .A(n21523), .B(n[565]), .Z(n23813) );
  XNOR U25298 ( .A(n23814), .B(n23811), .Z(n17564) );
  XOR U25299 ( .A(n23815), .B(n23816), .Z(n23811) );
  AND U25300 ( .A(n17571), .B(n23817), .Z(n23815) );
  XNOR U25301 ( .A(n17570), .B(n23816), .Z(n23817) );
  NAND U25302 ( .A(n23818), .B(n[564]), .Z(n17570) );
  NAND U25303 ( .A(n21523), .B(n[564]), .Z(n23818) );
  XNOR U25304 ( .A(n23819), .B(n23816), .Z(n17571) );
  XOR U25305 ( .A(n23820), .B(n23821), .Z(n23816) );
  AND U25306 ( .A(n17578), .B(n23822), .Z(n23820) );
  XNOR U25307 ( .A(n17577), .B(n23821), .Z(n23822) );
  NAND U25308 ( .A(n23823), .B(n[563]), .Z(n17577) );
  NAND U25309 ( .A(n21523), .B(n[563]), .Z(n23823) );
  XNOR U25310 ( .A(n23824), .B(n23821), .Z(n17578) );
  XOR U25311 ( .A(n23825), .B(n23826), .Z(n23821) );
  AND U25312 ( .A(n17585), .B(n23827), .Z(n23825) );
  XNOR U25313 ( .A(n17584), .B(n23826), .Z(n23827) );
  NAND U25314 ( .A(n23828), .B(n[562]), .Z(n17584) );
  NAND U25315 ( .A(n21523), .B(n[562]), .Z(n23828) );
  XNOR U25316 ( .A(n23829), .B(n23826), .Z(n17585) );
  XOR U25317 ( .A(n23830), .B(n23831), .Z(n23826) );
  AND U25318 ( .A(n17592), .B(n23832), .Z(n23830) );
  XNOR U25319 ( .A(n17591), .B(n23831), .Z(n23832) );
  NAND U25320 ( .A(n23833), .B(n[561]), .Z(n17591) );
  NAND U25321 ( .A(n21523), .B(n[561]), .Z(n23833) );
  XNOR U25322 ( .A(n23834), .B(n23831), .Z(n17592) );
  XOR U25323 ( .A(n23835), .B(n23836), .Z(n23831) );
  AND U25324 ( .A(n17599), .B(n23837), .Z(n23835) );
  XNOR U25325 ( .A(n17598), .B(n23836), .Z(n23837) );
  NAND U25326 ( .A(n23838), .B(n[560]), .Z(n17598) );
  NAND U25327 ( .A(n21523), .B(n[560]), .Z(n23838) );
  XNOR U25328 ( .A(n23839), .B(n23836), .Z(n17599) );
  XOR U25329 ( .A(n23840), .B(n23841), .Z(n23836) );
  AND U25330 ( .A(n17606), .B(n23842), .Z(n23840) );
  XNOR U25331 ( .A(n17605), .B(n23841), .Z(n23842) );
  NAND U25332 ( .A(n23843), .B(n[559]), .Z(n17605) );
  NAND U25333 ( .A(n21523), .B(n[559]), .Z(n23843) );
  XNOR U25334 ( .A(n23844), .B(n23841), .Z(n17606) );
  XOR U25335 ( .A(n23845), .B(n23846), .Z(n23841) );
  AND U25336 ( .A(n17613), .B(n23847), .Z(n23845) );
  XNOR U25337 ( .A(n17612), .B(n23846), .Z(n23847) );
  NAND U25338 ( .A(n23848), .B(n[558]), .Z(n17612) );
  NAND U25339 ( .A(n21523), .B(n[558]), .Z(n23848) );
  XNOR U25340 ( .A(n23849), .B(n23846), .Z(n17613) );
  XOR U25341 ( .A(n23850), .B(n23851), .Z(n23846) );
  AND U25342 ( .A(n17620), .B(n23852), .Z(n23850) );
  XNOR U25343 ( .A(n17619), .B(n23851), .Z(n23852) );
  NAND U25344 ( .A(n23853), .B(n[557]), .Z(n17619) );
  NAND U25345 ( .A(n21523), .B(n[557]), .Z(n23853) );
  XNOR U25346 ( .A(n23854), .B(n23851), .Z(n17620) );
  XOR U25347 ( .A(n23855), .B(n23856), .Z(n23851) );
  AND U25348 ( .A(n17627), .B(n23857), .Z(n23855) );
  XNOR U25349 ( .A(n17626), .B(n23856), .Z(n23857) );
  NAND U25350 ( .A(n23858), .B(n[556]), .Z(n17626) );
  NAND U25351 ( .A(n21523), .B(n[556]), .Z(n23858) );
  XNOR U25352 ( .A(n23859), .B(n23856), .Z(n17627) );
  XOR U25353 ( .A(n23860), .B(n23861), .Z(n23856) );
  AND U25354 ( .A(n17634), .B(n23862), .Z(n23860) );
  XNOR U25355 ( .A(n17633), .B(n23861), .Z(n23862) );
  NAND U25356 ( .A(n23863), .B(n[555]), .Z(n17633) );
  NAND U25357 ( .A(n21523), .B(n[555]), .Z(n23863) );
  XNOR U25358 ( .A(n23864), .B(n23861), .Z(n17634) );
  XOR U25359 ( .A(n23865), .B(n23866), .Z(n23861) );
  AND U25360 ( .A(n17641), .B(n23867), .Z(n23865) );
  XNOR U25361 ( .A(n17640), .B(n23866), .Z(n23867) );
  NAND U25362 ( .A(n23868), .B(n[554]), .Z(n17640) );
  NAND U25363 ( .A(n21523), .B(n[554]), .Z(n23868) );
  XNOR U25364 ( .A(n23869), .B(n23866), .Z(n17641) );
  XOR U25365 ( .A(n23870), .B(n23871), .Z(n23866) );
  AND U25366 ( .A(n17648), .B(n23872), .Z(n23870) );
  XNOR U25367 ( .A(n17647), .B(n23871), .Z(n23872) );
  NAND U25368 ( .A(n23873), .B(n[553]), .Z(n17647) );
  NAND U25369 ( .A(n21523), .B(n[553]), .Z(n23873) );
  XNOR U25370 ( .A(n23874), .B(n23871), .Z(n17648) );
  XOR U25371 ( .A(n23875), .B(n23876), .Z(n23871) );
  AND U25372 ( .A(n17655), .B(n23877), .Z(n23875) );
  XNOR U25373 ( .A(n17654), .B(n23876), .Z(n23877) );
  NAND U25374 ( .A(n23878), .B(n[552]), .Z(n17654) );
  NAND U25375 ( .A(n21523), .B(n[552]), .Z(n23878) );
  XNOR U25376 ( .A(n23879), .B(n23876), .Z(n17655) );
  XOR U25377 ( .A(n23880), .B(n23881), .Z(n23876) );
  AND U25378 ( .A(n17662), .B(n23882), .Z(n23880) );
  XNOR U25379 ( .A(n17661), .B(n23881), .Z(n23882) );
  NAND U25380 ( .A(n23883), .B(n[551]), .Z(n17661) );
  NAND U25381 ( .A(n21523), .B(n[551]), .Z(n23883) );
  XNOR U25382 ( .A(n23884), .B(n23881), .Z(n17662) );
  XOR U25383 ( .A(n23885), .B(n23886), .Z(n23881) );
  AND U25384 ( .A(n17669), .B(n23887), .Z(n23885) );
  XNOR U25385 ( .A(n17668), .B(n23886), .Z(n23887) );
  NAND U25386 ( .A(n23888), .B(n[550]), .Z(n17668) );
  NAND U25387 ( .A(n21523), .B(n[550]), .Z(n23888) );
  XNOR U25388 ( .A(n23889), .B(n23886), .Z(n17669) );
  XOR U25389 ( .A(n23890), .B(n23891), .Z(n23886) );
  AND U25390 ( .A(n17676), .B(n23892), .Z(n23890) );
  XNOR U25391 ( .A(n17675), .B(n23891), .Z(n23892) );
  NAND U25392 ( .A(n23893), .B(n[549]), .Z(n17675) );
  NAND U25393 ( .A(n21523), .B(n[549]), .Z(n23893) );
  XNOR U25394 ( .A(n23894), .B(n23891), .Z(n17676) );
  XOR U25395 ( .A(n23895), .B(n23896), .Z(n23891) );
  AND U25396 ( .A(n17683), .B(n23897), .Z(n23895) );
  XNOR U25397 ( .A(n17682), .B(n23896), .Z(n23897) );
  NAND U25398 ( .A(n23898), .B(n[548]), .Z(n17682) );
  NAND U25399 ( .A(n21523), .B(n[548]), .Z(n23898) );
  XNOR U25400 ( .A(n23899), .B(n23896), .Z(n17683) );
  XOR U25401 ( .A(n23900), .B(n23901), .Z(n23896) );
  AND U25402 ( .A(n17690), .B(n23902), .Z(n23900) );
  XNOR U25403 ( .A(n17689), .B(n23901), .Z(n23902) );
  NAND U25404 ( .A(n23903), .B(n[547]), .Z(n17689) );
  NAND U25405 ( .A(n21523), .B(n[547]), .Z(n23903) );
  XNOR U25406 ( .A(n23904), .B(n23901), .Z(n17690) );
  XOR U25407 ( .A(n23905), .B(n23906), .Z(n23901) );
  AND U25408 ( .A(n17697), .B(n23907), .Z(n23905) );
  XNOR U25409 ( .A(n17696), .B(n23906), .Z(n23907) );
  NAND U25410 ( .A(n23908), .B(n[546]), .Z(n17696) );
  NAND U25411 ( .A(n21523), .B(n[546]), .Z(n23908) );
  XNOR U25412 ( .A(n23909), .B(n23906), .Z(n17697) );
  XOR U25413 ( .A(n23910), .B(n23911), .Z(n23906) );
  AND U25414 ( .A(n17704), .B(n23912), .Z(n23910) );
  XNOR U25415 ( .A(n17703), .B(n23911), .Z(n23912) );
  NAND U25416 ( .A(n23913), .B(n[545]), .Z(n17703) );
  NAND U25417 ( .A(n21523), .B(n[545]), .Z(n23913) );
  XNOR U25418 ( .A(n23914), .B(n23911), .Z(n17704) );
  XOR U25419 ( .A(n23915), .B(n23916), .Z(n23911) );
  AND U25420 ( .A(n17711), .B(n23917), .Z(n23915) );
  XNOR U25421 ( .A(n17710), .B(n23916), .Z(n23917) );
  NAND U25422 ( .A(n23918), .B(n[544]), .Z(n17710) );
  NAND U25423 ( .A(n21523), .B(n[544]), .Z(n23918) );
  XNOR U25424 ( .A(n23919), .B(n23916), .Z(n17711) );
  XOR U25425 ( .A(n23920), .B(n23921), .Z(n23916) );
  AND U25426 ( .A(n17718), .B(n23922), .Z(n23920) );
  XNOR U25427 ( .A(n17717), .B(n23921), .Z(n23922) );
  NAND U25428 ( .A(n23923), .B(n[543]), .Z(n17717) );
  NAND U25429 ( .A(n21523), .B(n[543]), .Z(n23923) );
  XNOR U25430 ( .A(n23924), .B(n23921), .Z(n17718) );
  XOR U25431 ( .A(n23925), .B(n23926), .Z(n23921) );
  AND U25432 ( .A(n17725), .B(n23927), .Z(n23925) );
  XNOR U25433 ( .A(n17724), .B(n23926), .Z(n23927) );
  NAND U25434 ( .A(n23928), .B(n[542]), .Z(n17724) );
  NAND U25435 ( .A(n21523), .B(n[542]), .Z(n23928) );
  XNOR U25436 ( .A(n23929), .B(n23926), .Z(n17725) );
  XOR U25437 ( .A(n23930), .B(n23931), .Z(n23926) );
  AND U25438 ( .A(n17732), .B(n23932), .Z(n23930) );
  XNOR U25439 ( .A(n17731), .B(n23931), .Z(n23932) );
  NAND U25440 ( .A(n23933), .B(n[541]), .Z(n17731) );
  NAND U25441 ( .A(n21523), .B(n[541]), .Z(n23933) );
  XNOR U25442 ( .A(n23934), .B(n23931), .Z(n17732) );
  XOR U25443 ( .A(n23935), .B(n23936), .Z(n23931) );
  AND U25444 ( .A(n17739), .B(n23937), .Z(n23935) );
  XNOR U25445 ( .A(n17738), .B(n23936), .Z(n23937) );
  NAND U25446 ( .A(n23938), .B(n[540]), .Z(n17738) );
  NAND U25447 ( .A(n21523), .B(n[540]), .Z(n23938) );
  XNOR U25448 ( .A(n23939), .B(n23936), .Z(n17739) );
  XOR U25449 ( .A(n23940), .B(n23941), .Z(n23936) );
  AND U25450 ( .A(n17746), .B(n23942), .Z(n23940) );
  XNOR U25451 ( .A(n17745), .B(n23941), .Z(n23942) );
  NAND U25452 ( .A(n23943), .B(n[539]), .Z(n17745) );
  NAND U25453 ( .A(n21523), .B(n[539]), .Z(n23943) );
  XNOR U25454 ( .A(n23944), .B(n23941), .Z(n17746) );
  XOR U25455 ( .A(n23945), .B(n23946), .Z(n23941) );
  AND U25456 ( .A(n17753), .B(n23947), .Z(n23945) );
  XNOR U25457 ( .A(n17752), .B(n23946), .Z(n23947) );
  NAND U25458 ( .A(n23948), .B(n[538]), .Z(n17752) );
  NAND U25459 ( .A(n21523), .B(n[538]), .Z(n23948) );
  XNOR U25460 ( .A(n23949), .B(n23946), .Z(n17753) );
  XOR U25461 ( .A(n23950), .B(n23951), .Z(n23946) );
  AND U25462 ( .A(n17760), .B(n23952), .Z(n23950) );
  XNOR U25463 ( .A(n17759), .B(n23951), .Z(n23952) );
  NAND U25464 ( .A(n23953), .B(n[537]), .Z(n17759) );
  NAND U25465 ( .A(n21523), .B(n[537]), .Z(n23953) );
  XNOR U25466 ( .A(n23954), .B(n23951), .Z(n17760) );
  XOR U25467 ( .A(n23955), .B(n23956), .Z(n23951) );
  AND U25468 ( .A(n17767), .B(n23957), .Z(n23955) );
  XNOR U25469 ( .A(n17766), .B(n23956), .Z(n23957) );
  NAND U25470 ( .A(n23958), .B(n[536]), .Z(n17766) );
  NAND U25471 ( .A(n21523), .B(n[536]), .Z(n23958) );
  XNOR U25472 ( .A(n23959), .B(n23956), .Z(n17767) );
  XOR U25473 ( .A(n23960), .B(n23961), .Z(n23956) );
  AND U25474 ( .A(n17774), .B(n23962), .Z(n23960) );
  XNOR U25475 ( .A(n17773), .B(n23961), .Z(n23962) );
  NAND U25476 ( .A(n23963), .B(n[535]), .Z(n17773) );
  NAND U25477 ( .A(n21523), .B(n[535]), .Z(n23963) );
  XNOR U25478 ( .A(n23964), .B(n23961), .Z(n17774) );
  XOR U25479 ( .A(n23965), .B(n23966), .Z(n23961) );
  AND U25480 ( .A(n17781), .B(n23967), .Z(n23965) );
  XNOR U25481 ( .A(n17780), .B(n23966), .Z(n23967) );
  NAND U25482 ( .A(n23968), .B(n[534]), .Z(n17780) );
  NAND U25483 ( .A(n21523), .B(n[534]), .Z(n23968) );
  XNOR U25484 ( .A(n23969), .B(n23966), .Z(n17781) );
  XOR U25485 ( .A(n23970), .B(n23971), .Z(n23966) );
  AND U25486 ( .A(n17788), .B(n23972), .Z(n23970) );
  XNOR U25487 ( .A(n17787), .B(n23971), .Z(n23972) );
  NAND U25488 ( .A(n23973), .B(n[533]), .Z(n17787) );
  NAND U25489 ( .A(n21523), .B(n[533]), .Z(n23973) );
  XNOR U25490 ( .A(n23974), .B(n23971), .Z(n17788) );
  XOR U25491 ( .A(n23975), .B(n23976), .Z(n23971) );
  AND U25492 ( .A(n17795), .B(n23977), .Z(n23975) );
  XNOR U25493 ( .A(n17794), .B(n23976), .Z(n23977) );
  NAND U25494 ( .A(n23978), .B(n[532]), .Z(n17794) );
  NAND U25495 ( .A(n21523), .B(n[532]), .Z(n23978) );
  XNOR U25496 ( .A(n23979), .B(n23976), .Z(n17795) );
  XOR U25497 ( .A(n23980), .B(n23981), .Z(n23976) );
  AND U25498 ( .A(n17802), .B(n23982), .Z(n23980) );
  XNOR U25499 ( .A(n17801), .B(n23981), .Z(n23982) );
  NAND U25500 ( .A(n23983), .B(n[531]), .Z(n17801) );
  NAND U25501 ( .A(n21523), .B(n[531]), .Z(n23983) );
  XNOR U25502 ( .A(n23984), .B(n23981), .Z(n17802) );
  XOR U25503 ( .A(n23985), .B(n23986), .Z(n23981) );
  AND U25504 ( .A(n17809), .B(n23987), .Z(n23985) );
  XNOR U25505 ( .A(n17808), .B(n23986), .Z(n23987) );
  NAND U25506 ( .A(n23988), .B(n[530]), .Z(n17808) );
  NAND U25507 ( .A(n21523), .B(n[530]), .Z(n23988) );
  XNOR U25508 ( .A(n23989), .B(n23986), .Z(n17809) );
  XOR U25509 ( .A(n23990), .B(n23991), .Z(n23986) );
  AND U25510 ( .A(n17816), .B(n23992), .Z(n23990) );
  XNOR U25511 ( .A(n17815), .B(n23991), .Z(n23992) );
  NAND U25512 ( .A(n23993), .B(n[529]), .Z(n17815) );
  NAND U25513 ( .A(n21523), .B(n[529]), .Z(n23993) );
  XNOR U25514 ( .A(n23994), .B(n23991), .Z(n17816) );
  XOR U25515 ( .A(n23995), .B(n23996), .Z(n23991) );
  AND U25516 ( .A(n17823), .B(n23997), .Z(n23995) );
  XNOR U25517 ( .A(n17822), .B(n23996), .Z(n23997) );
  NAND U25518 ( .A(n23998), .B(n[528]), .Z(n17822) );
  NAND U25519 ( .A(n21523), .B(n[528]), .Z(n23998) );
  XNOR U25520 ( .A(n23999), .B(n23996), .Z(n17823) );
  XOR U25521 ( .A(n24000), .B(n24001), .Z(n23996) );
  AND U25522 ( .A(n17830), .B(n24002), .Z(n24000) );
  XNOR U25523 ( .A(n17829), .B(n24001), .Z(n24002) );
  NAND U25524 ( .A(n24003), .B(n[527]), .Z(n17829) );
  NAND U25525 ( .A(n21523), .B(n[527]), .Z(n24003) );
  XNOR U25526 ( .A(n24004), .B(n24001), .Z(n17830) );
  XOR U25527 ( .A(n24005), .B(n24006), .Z(n24001) );
  AND U25528 ( .A(n17837), .B(n24007), .Z(n24005) );
  XNOR U25529 ( .A(n17836), .B(n24006), .Z(n24007) );
  NAND U25530 ( .A(n24008), .B(n[526]), .Z(n17836) );
  NAND U25531 ( .A(n21523), .B(n[526]), .Z(n24008) );
  XNOR U25532 ( .A(n24009), .B(n24006), .Z(n17837) );
  XOR U25533 ( .A(n24010), .B(n24011), .Z(n24006) );
  AND U25534 ( .A(n17844), .B(n24012), .Z(n24010) );
  XNOR U25535 ( .A(n17843), .B(n24011), .Z(n24012) );
  NAND U25536 ( .A(n24013), .B(n[525]), .Z(n17843) );
  NAND U25537 ( .A(n21523), .B(n[525]), .Z(n24013) );
  XNOR U25538 ( .A(n24014), .B(n24011), .Z(n17844) );
  XOR U25539 ( .A(n24015), .B(n24016), .Z(n24011) );
  AND U25540 ( .A(n17851), .B(n24017), .Z(n24015) );
  XNOR U25541 ( .A(n17850), .B(n24016), .Z(n24017) );
  NAND U25542 ( .A(n24018), .B(n[524]), .Z(n17850) );
  NAND U25543 ( .A(n21523), .B(n[524]), .Z(n24018) );
  XNOR U25544 ( .A(n24019), .B(n24016), .Z(n17851) );
  XOR U25545 ( .A(n24020), .B(n24021), .Z(n24016) );
  AND U25546 ( .A(n17858), .B(n24022), .Z(n24020) );
  XNOR U25547 ( .A(n17857), .B(n24021), .Z(n24022) );
  NAND U25548 ( .A(n24023), .B(n[523]), .Z(n17857) );
  NAND U25549 ( .A(n21523), .B(n[523]), .Z(n24023) );
  XNOR U25550 ( .A(n24024), .B(n24021), .Z(n17858) );
  XOR U25551 ( .A(n24025), .B(n24026), .Z(n24021) );
  AND U25552 ( .A(n17865), .B(n24027), .Z(n24025) );
  XNOR U25553 ( .A(n17864), .B(n24026), .Z(n24027) );
  NAND U25554 ( .A(n24028), .B(n[522]), .Z(n17864) );
  NAND U25555 ( .A(n21523), .B(n[522]), .Z(n24028) );
  XNOR U25556 ( .A(n24029), .B(n24026), .Z(n17865) );
  XOR U25557 ( .A(n24030), .B(n24031), .Z(n24026) );
  AND U25558 ( .A(n17872), .B(n24032), .Z(n24030) );
  XNOR U25559 ( .A(n17871), .B(n24031), .Z(n24032) );
  NAND U25560 ( .A(n24033), .B(n[521]), .Z(n17871) );
  NAND U25561 ( .A(n21523), .B(n[521]), .Z(n24033) );
  XNOR U25562 ( .A(n24034), .B(n24031), .Z(n17872) );
  XOR U25563 ( .A(n24035), .B(n24036), .Z(n24031) );
  AND U25564 ( .A(n17879), .B(n24037), .Z(n24035) );
  XNOR U25565 ( .A(n17878), .B(n24036), .Z(n24037) );
  NAND U25566 ( .A(n24038), .B(n[520]), .Z(n17878) );
  NAND U25567 ( .A(n21523), .B(n[520]), .Z(n24038) );
  XNOR U25568 ( .A(n24039), .B(n24036), .Z(n17879) );
  XOR U25569 ( .A(n24040), .B(n24041), .Z(n24036) );
  AND U25570 ( .A(n17886), .B(n24042), .Z(n24040) );
  XNOR U25571 ( .A(n17885), .B(n24041), .Z(n24042) );
  NAND U25572 ( .A(n24043), .B(n[519]), .Z(n17885) );
  NAND U25573 ( .A(n21523), .B(n[519]), .Z(n24043) );
  XNOR U25574 ( .A(n24044), .B(n24041), .Z(n17886) );
  XOR U25575 ( .A(n24045), .B(n24046), .Z(n24041) );
  AND U25576 ( .A(n17893), .B(n24047), .Z(n24045) );
  XNOR U25577 ( .A(n17892), .B(n24046), .Z(n24047) );
  NAND U25578 ( .A(n24048), .B(n[518]), .Z(n17892) );
  NAND U25579 ( .A(n21523), .B(n[518]), .Z(n24048) );
  XNOR U25580 ( .A(n24049), .B(n24046), .Z(n17893) );
  XOR U25581 ( .A(n24050), .B(n24051), .Z(n24046) );
  AND U25582 ( .A(n17900), .B(n24052), .Z(n24050) );
  XNOR U25583 ( .A(n17899), .B(n24051), .Z(n24052) );
  NAND U25584 ( .A(n24053), .B(n[517]), .Z(n17899) );
  NAND U25585 ( .A(n21523), .B(n[517]), .Z(n24053) );
  XNOR U25586 ( .A(n24054), .B(n24051), .Z(n17900) );
  XOR U25587 ( .A(n24055), .B(n24056), .Z(n24051) );
  AND U25588 ( .A(n17907), .B(n24057), .Z(n24055) );
  XNOR U25589 ( .A(n17906), .B(n24056), .Z(n24057) );
  NAND U25590 ( .A(n24058), .B(n[516]), .Z(n17906) );
  NAND U25591 ( .A(n21523), .B(n[516]), .Z(n24058) );
  XNOR U25592 ( .A(n24059), .B(n24056), .Z(n17907) );
  XOR U25593 ( .A(n24060), .B(n24061), .Z(n24056) );
  AND U25594 ( .A(n17914), .B(n24062), .Z(n24060) );
  XNOR U25595 ( .A(n17913), .B(n24061), .Z(n24062) );
  NAND U25596 ( .A(n24063), .B(n[515]), .Z(n17913) );
  NAND U25597 ( .A(n21523), .B(n[515]), .Z(n24063) );
  XNOR U25598 ( .A(n24064), .B(n24061), .Z(n17914) );
  XOR U25599 ( .A(n24065), .B(n24066), .Z(n24061) );
  AND U25600 ( .A(n17921), .B(n24067), .Z(n24065) );
  XNOR U25601 ( .A(n17920), .B(n24066), .Z(n24067) );
  NAND U25602 ( .A(n24068), .B(n[514]), .Z(n17920) );
  NAND U25603 ( .A(n21523), .B(n[514]), .Z(n24068) );
  XNOR U25604 ( .A(n24069), .B(n24066), .Z(n17921) );
  XOR U25605 ( .A(n24070), .B(n24071), .Z(n24066) );
  AND U25606 ( .A(n17928), .B(n24072), .Z(n24070) );
  XNOR U25607 ( .A(n17927), .B(n24071), .Z(n24072) );
  NAND U25608 ( .A(n24073), .B(n[513]), .Z(n17927) );
  NAND U25609 ( .A(n21523), .B(n[513]), .Z(n24073) );
  XNOR U25610 ( .A(n24074), .B(n24071), .Z(n17928) );
  XOR U25611 ( .A(n24075), .B(n24076), .Z(n24071) );
  AND U25612 ( .A(n17935), .B(n24077), .Z(n24075) );
  XNOR U25613 ( .A(n17934), .B(n24076), .Z(n24077) );
  NAND U25614 ( .A(n24078), .B(n[512]), .Z(n17934) );
  NAND U25615 ( .A(n21523), .B(n[512]), .Z(n24078) );
  XNOR U25616 ( .A(n24079), .B(n24076), .Z(n17935) );
  XOR U25617 ( .A(n24080), .B(n24081), .Z(n24076) );
  AND U25618 ( .A(n17942), .B(n24082), .Z(n24080) );
  XNOR U25619 ( .A(n17941), .B(n24081), .Z(n24082) );
  NAND U25620 ( .A(n24083), .B(n[511]), .Z(n17941) );
  NAND U25621 ( .A(n21523), .B(n[511]), .Z(n24083) );
  XNOR U25622 ( .A(n24084), .B(n24081), .Z(n17942) );
  XOR U25623 ( .A(n24085), .B(n24086), .Z(n24081) );
  AND U25624 ( .A(n17949), .B(n24087), .Z(n24085) );
  XNOR U25625 ( .A(n17948), .B(n24086), .Z(n24087) );
  NAND U25626 ( .A(n24088), .B(n[510]), .Z(n17948) );
  NAND U25627 ( .A(n21523), .B(n[510]), .Z(n24088) );
  XNOR U25628 ( .A(n24089), .B(n24086), .Z(n17949) );
  XOR U25629 ( .A(n24090), .B(n24091), .Z(n24086) );
  AND U25630 ( .A(n17956), .B(n24092), .Z(n24090) );
  XNOR U25631 ( .A(n17955), .B(n24091), .Z(n24092) );
  NAND U25632 ( .A(n24093), .B(n[509]), .Z(n17955) );
  NAND U25633 ( .A(n21523), .B(n[509]), .Z(n24093) );
  XNOR U25634 ( .A(n24094), .B(n24091), .Z(n17956) );
  XOR U25635 ( .A(n24095), .B(n24096), .Z(n24091) );
  AND U25636 ( .A(n17963), .B(n24097), .Z(n24095) );
  XNOR U25637 ( .A(n17962), .B(n24096), .Z(n24097) );
  NAND U25638 ( .A(n24098), .B(n[508]), .Z(n17962) );
  NAND U25639 ( .A(n21523), .B(n[508]), .Z(n24098) );
  XNOR U25640 ( .A(n24099), .B(n24096), .Z(n17963) );
  XOR U25641 ( .A(n24100), .B(n24101), .Z(n24096) );
  AND U25642 ( .A(n17970), .B(n24102), .Z(n24100) );
  XNOR U25643 ( .A(n17969), .B(n24101), .Z(n24102) );
  NAND U25644 ( .A(n24103), .B(n[507]), .Z(n17969) );
  NAND U25645 ( .A(n21523), .B(n[507]), .Z(n24103) );
  XNOR U25646 ( .A(n24104), .B(n24101), .Z(n17970) );
  XOR U25647 ( .A(n24105), .B(n24106), .Z(n24101) );
  AND U25648 ( .A(n17977), .B(n24107), .Z(n24105) );
  XNOR U25649 ( .A(n17976), .B(n24106), .Z(n24107) );
  NAND U25650 ( .A(n24108), .B(n[506]), .Z(n17976) );
  NAND U25651 ( .A(n21523), .B(n[506]), .Z(n24108) );
  XNOR U25652 ( .A(n24109), .B(n24106), .Z(n17977) );
  XOR U25653 ( .A(n24110), .B(n24111), .Z(n24106) );
  AND U25654 ( .A(n17984), .B(n24112), .Z(n24110) );
  XNOR U25655 ( .A(n17983), .B(n24111), .Z(n24112) );
  NAND U25656 ( .A(n24113), .B(n[505]), .Z(n17983) );
  NAND U25657 ( .A(n21523), .B(n[505]), .Z(n24113) );
  XNOR U25658 ( .A(n24114), .B(n24111), .Z(n17984) );
  XOR U25659 ( .A(n24115), .B(n24116), .Z(n24111) );
  AND U25660 ( .A(n17991), .B(n24117), .Z(n24115) );
  XNOR U25661 ( .A(n17990), .B(n24116), .Z(n24117) );
  NAND U25662 ( .A(n24118), .B(n[504]), .Z(n17990) );
  NAND U25663 ( .A(n21523), .B(n[504]), .Z(n24118) );
  XNOR U25664 ( .A(n24119), .B(n24116), .Z(n17991) );
  XOR U25665 ( .A(n24120), .B(n24121), .Z(n24116) );
  AND U25666 ( .A(n17998), .B(n24122), .Z(n24120) );
  XNOR U25667 ( .A(n17997), .B(n24121), .Z(n24122) );
  NAND U25668 ( .A(n24123), .B(n[503]), .Z(n17997) );
  NAND U25669 ( .A(n21523), .B(n[503]), .Z(n24123) );
  XNOR U25670 ( .A(n24124), .B(n24121), .Z(n17998) );
  XOR U25671 ( .A(n24125), .B(n24126), .Z(n24121) );
  AND U25672 ( .A(n18005), .B(n24127), .Z(n24125) );
  XNOR U25673 ( .A(n18004), .B(n24126), .Z(n24127) );
  NAND U25674 ( .A(n24128), .B(n[502]), .Z(n18004) );
  NAND U25675 ( .A(n21523), .B(n[502]), .Z(n24128) );
  XNOR U25676 ( .A(n24129), .B(n24126), .Z(n18005) );
  XOR U25677 ( .A(n24130), .B(n24131), .Z(n24126) );
  AND U25678 ( .A(n18012), .B(n24132), .Z(n24130) );
  XNOR U25679 ( .A(n18011), .B(n24131), .Z(n24132) );
  NAND U25680 ( .A(n24133), .B(n[501]), .Z(n18011) );
  NAND U25681 ( .A(n21523), .B(n[501]), .Z(n24133) );
  XNOR U25682 ( .A(n24134), .B(n24131), .Z(n18012) );
  XOR U25683 ( .A(n24135), .B(n24136), .Z(n24131) );
  AND U25684 ( .A(n18019), .B(n24137), .Z(n24135) );
  XNOR U25685 ( .A(n18018), .B(n24136), .Z(n24137) );
  NAND U25686 ( .A(n24138), .B(n[500]), .Z(n18018) );
  NAND U25687 ( .A(n21523), .B(n[500]), .Z(n24138) );
  XNOR U25688 ( .A(n24139), .B(n24136), .Z(n18019) );
  XOR U25689 ( .A(n24140), .B(n24141), .Z(n24136) );
  AND U25690 ( .A(n18026), .B(n24142), .Z(n24140) );
  XNOR U25691 ( .A(n18025), .B(n24141), .Z(n24142) );
  NAND U25692 ( .A(n24143), .B(n[499]), .Z(n18025) );
  NAND U25693 ( .A(n21523), .B(n[499]), .Z(n24143) );
  XNOR U25694 ( .A(n24144), .B(n24141), .Z(n18026) );
  XOR U25695 ( .A(n24145), .B(n24146), .Z(n24141) );
  AND U25696 ( .A(n18033), .B(n24147), .Z(n24145) );
  XNOR U25697 ( .A(n18032), .B(n24146), .Z(n24147) );
  NAND U25698 ( .A(n24148), .B(n[498]), .Z(n18032) );
  NAND U25699 ( .A(n21523), .B(n[498]), .Z(n24148) );
  XNOR U25700 ( .A(n24149), .B(n24146), .Z(n18033) );
  XOR U25701 ( .A(n24150), .B(n24151), .Z(n24146) );
  AND U25702 ( .A(n18040), .B(n24152), .Z(n24150) );
  XNOR U25703 ( .A(n18039), .B(n24151), .Z(n24152) );
  NAND U25704 ( .A(n24153), .B(n[497]), .Z(n18039) );
  NAND U25705 ( .A(n21523), .B(n[497]), .Z(n24153) );
  XNOR U25706 ( .A(n24154), .B(n24151), .Z(n18040) );
  XOR U25707 ( .A(n24155), .B(n24156), .Z(n24151) );
  AND U25708 ( .A(n18047), .B(n24157), .Z(n24155) );
  XNOR U25709 ( .A(n18046), .B(n24156), .Z(n24157) );
  NAND U25710 ( .A(n24158), .B(n[496]), .Z(n18046) );
  NAND U25711 ( .A(n21523), .B(n[496]), .Z(n24158) );
  XNOR U25712 ( .A(n24159), .B(n24156), .Z(n18047) );
  XOR U25713 ( .A(n24160), .B(n24161), .Z(n24156) );
  AND U25714 ( .A(n18054), .B(n24162), .Z(n24160) );
  XNOR U25715 ( .A(n18053), .B(n24161), .Z(n24162) );
  NAND U25716 ( .A(n24163), .B(n[495]), .Z(n18053) );
  NAND U25717 ( .A(n21523), .B(n[495]), .Z(n24163) );
  XNOR U25718 ( .A(n24164), .B(n24161), .Z(n18054) );
  XOR U25719 ( .A(n24165), .B(n24166), .Z(n24161) );
  AND U25720 ( .A(n18061), .B(n24167), .Z(n24165) );
  XNOR U25721 ( .A(n18060), .B(n24166), .Z(n24167) );
  NAND U25722 ( .A(n24168), .B(n[494]), .Z(n18060) );
  NAND U25723 ( .A(n21523), .B(n[494]), .Z(n24168) );
  XNOR U25724 ( .A(n24169), .B(n24166), .Z(n18061) );
  XOR U25725 ( .A(n24170), .B(n24171), .Z(n24166) );
  AND U25726 ( .A(n18068), .B(n24172), .Z(n24170) );
  XNOR U25727 ( .A(n18067), .B(n24171), .Z(n24172) );
  NAND U25728 ( .A(n24173), .B(n[493]), .Z(n18067) );
  NAND U25729 ( .A(n21523), .B(n[493]), .Z(n24173) );
  XNOR U25730 ( .A(n24174), .B(n24171), .Z(n18068) );
  XOR U25731 ( .A(n24175), .B(n24176), .Z(n24171) );
  AND U25732 ( .A(n18075), .B(n24177), .Z(n24175) );
  XNOR U25733 ( .A(n18074), .B(n24176), .Z(n24177) );
  NAND U25734 ( .A(n24178), .B(n[492]), .Z(n18074) );
  NAND U25735 ( .A(n21523), .B(n[492]), .Z(n24178) );
  XNOR U25736 ( .A(n24179), .B(n24176), .Z(n18075) );
  XOR U25737 ( .A(n24180), .B(n24181), .Z(n24176) );
  AND U25738 ( .A(n18082), .B(n24182), .Z(n24180) );
  XNOR U25739 ( .A(n18081), .B(n24181), .Z(n24182) );
  NAND U25740 ( .A(n24183), .B(n[491]), .Z(n18081) );
  NAND U25741 ( .A(n21523), .B(n[491]), .Z(n24183) );
  XNOR U25742 ( .A(n24184), .B(n24181), .Z(n18082) );
  XOR U25743 ( .A(n24185), .B(n24186), .Z(n24181) );
  AND U25744 ( .A(n18089), .B(n24187), .Z(n24185) );
  XNOR U25745 ( .A(n18088), .B(n24186), .Z(n24187) );
  NAND U25746 ( .A(n24188), .B(n[490]), .Z(n18088) );
  NAND U25747 ( .A(n21523), .B(n[490]), .Z(n24188) );
  XNOR U25748 ( .A(n24189), .B(n24186), .Z(n18089) );
  XOR U25749 ( .A(n24190), .B(n24191), .Z(n24186) );
  AND U25750 ( .A(n18096), .B(n24192), .Z(n24190) );
  XNOR U25751 ( .A(n18095), .B(n24191), .Z(n24192) );
  NAND U25752 ( .A(n24193), .B(n[489]), .Z(n18095) );
  NAND U25753 ( .A(n21523), .B(n[489]), .Z(n24193) );
  XNOR U25754 ( .A(n24194), .B(n24191), .Z(n18096) );
  XOR U25755 ( .A(n24195), .B(n24196), .Z(n24191) );
  AND U25756 ( .A(n18103), .B(n24197), .Z(n24195) );
  XNOR U25757 ( .A(n18102), .B(n24196), .Z(n24197) );
  NAND U25758 ( .A(n24198), .B(n[488]), .Z(n18102) );
  NAND U25759 ( .A(n21523), .B(n[488]), .Z(n24198) );
  XNOR U25760 ( .A(n24199), .B(n24196), .Z(n18103) );
  XOR U25761 ( .A(n24200), .B(n24201), .Z(n24196) );
  AND U25762 ( .A(n18110), .B(n24202), .Z(n24200) );
  XNOR U25763 ( .A(n18109), .B(n24201), .Z(n24202) );
  NAND U25764 ( .A(n24203), .B(n[487]), .Z(n18109) );
  NAND U25765 ( .A(n21523), .B(n[487]), .Z(n24203) );
  XNOR U25766 ( .A(n24204), .B(n24201), .Z(n18110) );
  XOR U25767 ( .A(n24205), .B(n24206), .Z(n24201) );
  AND U25768 ( .A(n18117), .B(n24207), .Z(n24205) );
  XNOR U25769 ( .A(n18116), .B(n24206), .Z(n24207) );
  NAND U25770 ( .A(n24208), .B(n[486]), .Z(n18116) );
  NAND U25771 ( .A(n21523), .B(n[486]), .Z(n24208) );
  XNOR U25772 ( .A(n24209), .B(n24206), .Z(n18117) );
  XOR U25773 ( .A(n24210), .B(n24211), .Z(n24206) );
  AND U25774 ( .A(n18124), .B(n24212), .Z(n24210) );
  XNOR U25775 ( .A(n18123), .B(n24211), .Z(n24212) );
  NAND U25776 ( .A(n24213), .B(n[485]), .Z(n18123) );
  NAND U25777 ( .A(n21523), .B(n[485]), .Z(n24213) );
  XNOR U25778 ( .A(n24214), .B(n24211), .Z(n18124) );
  XOR U25779 ( .A(n24215), .B(n24216), .Z(n24211) );
  AND U25780 ( .A(n18131), .B(n24217), .Z(n24215) );
  XNOR U25781 ( .A(n18130), .B(n24216), .Z(n24217) );
  NAND U25782 ( .A(n24218), .B(n[484]), .Z(n18130) );
  NAND U25783 ( .A(n21523), .B(n[484]), .Z(n24218) );
  XNOR U25784 ( .A(n24219), .B(n24216), .Z(n18131) );
  XOR U25785 ( .A(n24220), .B(n24221), .Z(n24216) );
  AND U25786 ( .A(n18138), .B(n24222), .Z(n24220) );
  XNOR U25787 ( .A(n18137), .B(n24221), .Z(n24222) );
  NAND U25788 ( .A(n24223), .B(n[483]), .Z(n18137) );
  NAND U25789 ( .A(n21523), .B(n[483]), .Z(n24223) );
  XNOR U25790 ( .A(n24224), .B(n24221), .Z(n18138) );
  XOR U25791 ( .A(n24225), .B(n24226), .Z(n24221) );
  AND U25792 ( .A(n18145), .B(n24227), .Z(n24225) );
  XNOR U25793 ( .A(n18144), .B(n24226), .Z(n24227) );
  NAND U25794 ( .A(n24228), .B(n[482]), .Z(n18144) );
  NAND U25795 ( .A(n21523), .B(n[482]), .Z(n24228) );
  XNOR U25796 ( .A(n24229), .B(n24226), .Z(n18145) );
  XOR U25797 ( .A(n24230), .B(n24231), .Z(n24226) );
  AND U25798 ( .A(n18152), .B(n24232), .Z(n24230) );
  XNOR U25799 ( .A(n18151), .B(n24231), .Z(n24232) );
  NAND U25800 ( .A(n24233), .B(n[481]), .Z(n18151) );
  NAND U25801 ( .A(n21523), .B(n[481]), .Z(n24233) );
  XNOR U25802 ( .A(n24234), .B(n24231), .Z(n18152) );
  XOR U25803 ( .A(n24235), .B(n24236), .Z(n24231) );
  AND U25804 ( .A(n18159), .B(n24237), .Z(n24235) );
  XNOR U25805 ( .A(n18158), .B(n24236), .Z(n24237) );
  NAND U25806 ( .A(n24238), .B(n[480]), .Z(n18158) );
  NAND U25807 ( .A(n21523), .B(n[480]), .Z(n24238) );
  XNOR U25808 ( .A(n24239), .B(n24236), .Z(n18159) );
  XOR U25809 ( .A(n24240), .B(n24241), .Z(n24236) );
  AND U25810 ( .A(n18166), .B(n24242), .Z(n24240) );
  XNOR U25811 ( .A(n18165), .B(n24241), .Z(n24242) );
  NAND U25812 ( .A(n24243), .B(n[479]), .Z(n18165) );
  NAND U25813 ( .A(n21523), .B(n[479]), .Z(n24243) );
  XNOR U25814 ( .A(n24244), .B(n24241), .Z(n18166) );
  XOR U25815 ( .A(n24245), .B(n24246), .Z(n24241) );
  AND U25816 ( .A(n18173), .B(n24247), .Z(n24245) );
  XNOR U25817 ( .A(n18172), .B(n24246), .Z(n24247) );
  NAND U25818 ( .A(n24248), .B(n[478]), .Z(n18172) );
  NAND U25819 ( .A(n21523), .B(n[478]), .Z(n24248) );
  XNOR U25820 ( .A(n24249), .B(n24246), .Z(n18173) );
  XOR U25821 ( .A(n24250), .B(n24251), .Z(n24246) );
  AND U25822 ( .A(n18180), .B(n24252), .Z(n24250) );
  XNOR U25823 ( .A(n18179), .B(n24251), .Z(n24252) );
  NAND U25824 ( .A(n24253), .B(n[477]), .Z(n18179) );
  NAND U25825 ( .A(n21523), .B(n[477]), .Z(n24253) );
  XNOR U25826 ( .A(n24254), .B(n24251), .Z(n18180) );
  XOR U25827 ( .A(n24255), .B(n24256), .Z(n24251) );
  AND U25828 ( .A(n18187), .B(n24257), .Z(n24255) );
  XNOR U25829 ( .A(n18186), .B(n24256), .Z(n24257) );
  NAND U25830 ( .A(n24258), .B(n[476]), .Z(n18186) );
  NAND U25831 ( .A(n21523), .B(n[476]), .Z(n24258) );
  XNOR U25832 ( .A(n24259), .B(n24256), .Z(n18187) );
  XOR U25833 ( .A(n24260), .B(n24261), .Z(n24256) );
  AND U25834 ( .A(n18194), .B(n24262), .Z(n24260) );
  XNOR U25835 ( .A(n18193), .B(n24261), .Z(n24262) );
  NAND U25836 ( .A(n24263), .B(n[475]), .Z(n18193) );
  NAND U25837 ( .A(n21523), .B(n[475]), .Z(n24263) );
  XNOR U25838 ( .A(n24264), .B(n24261), .Z(n18194) );
  XOR U25839 ( .A(n24265), .B(n24266), .Z(n24261) );
  AND U25840 ( .A(n18201), .B(n24267), .Z(n24265) );
  XNOR U25841 ( .A(n18200), .B(n24266), .Z(n24267) );
  NAND U25842 ( .A(n24268), .B(n[474]), .Z(n18200) );
  NAND U25843 ( .A(n21523), .B(n[474]), .Z(n24268) );
  XNOR U25844 ( .A(n24269), .B(n24266), .Z(n18201) );
  XOR U25845 ( .A(n24270), .B(n24271), .Z(n24266) );
  AND U25846 ( .A(n18208), .B(n24272), .Z(n24270) );
  XNOR U25847 ( .A(n18207), .B(n24271), .Z(n24272) );
  NAND U25848 ( .A(n24273), .B(n[473]), .Z(n18207) );
  NAND U25849 ( .A(n21523), .B(n[473]), .Z(n24273) );
  XNOR U25850 ( .A(n24274), .B(n24271), .Z(n18208) );
  XOR U25851 ( .A(n24275), .B(n24276), .Z(n24271) );
  AND U25852 ( .A(n18215), .B(n24277), .Z(n24275) );
  XNOR U25853 ( .A(n18214), .B(n24276), .Z(n24277) );
  NAND U25854 ( .A(n24278), .B(n[472]), .Z(n18214) );
  NAND U25855 ( .A(n21523), .B(n[472]), .Z(n24278) );
  XNOR U25856 ( .A(n24279), .B(n24276), .Z(n18215) );
  XOR U25857 ( .A(n24280), .B(n24281), .Z(n24276) );
  AND U25858 ( .A(n18222), .B(n24282), .Z(n24280) );
  XNOR U25859 ( .A(n18221), .B(n24281), .Z(n24282) );
  NAND U25860 ( .A(n24283), .B(n[471]), .Z(n18221) );
  NAND U25861 ( .A(n21523), .B(n[471]), .Z(n24283) );
  XNOR U25862 ( .A(n24284), .B(n24281), .Z(n18222) );
  XOR U25863 ( .A(n24285), .B(n24286), .Z(n24281) );
  AND U25864 ( .A(n18229), .B(n24287), .Z(n24285) );
  XNOR U25865 ( .A(n18228), .B(n24286), .Z(n24287) );
  NAND U25866 ( .A(n24288), .B(n[470]), .Z(n18228) );
  NAND U25867 ( .A(n21523), .B(n[470]), .Z(n24288) );
  XNOR U25868 ( .A(n24289), .B(n24286), .Z(n18229) );
  XOR U25869 ( .A(n24290), .B(n24291), .Z(n24286) );
  AND U25870 ( .A(n18236), .B(n24292), .Z(n24290) );
  XNOR U25871 ( .A(n18235), .B(n24291), .Z(n24292) );
  NAND U25872 ( .A(n24293), .B(n[469]), .Z(n18235) );
  NAND U25873 ( .A(n21523), .B(n[469]), .Z(n24293) );
  XNOR U25874 ( .A(n24294), .B(n24291), .Z(n18236) );
  XOR U25875 ( .A(n24295), .B(n24296), .Z(n24291) );
  AND U25876 ( .A(n18243), .B(n24297), .Z(n24295) );
  XNOR U25877 ( .A(n18242), .B(n24296), .Z(n24297) );
  NAND U25878 ( .A(n24298), .B(n[468]), .Z(n18242) );
  NAND U25879 ( .A(n21523), .B(n[468]), .Z(n24298) );
  XNOR U25880 ( .A(n24299), .B(n24296), .Z(n18243) );
  XOR U25881 ( .A(n24300), .B(n24301), .Z(n24296) );
  AND U25882 ( .A(n18250), .B(n24302), .Z(n24300) );
  XNOR U25883 ( .A(n18249), .B(n24301), .Z(n24302) );
  NAND U25884 ( .A(n24303), .B(n[467]), .Z(n18249) );
  NAND U25885 ( .A(n21523), .B(n[467]), .Z(n24303) );
  XNOR U25886 ( .A(n24304), .B(n24301), .Z(n18250) );
  XOR U25887 ( .A(n24305), .B(n24306), .Z(n24301) );
  AND U25888 ( .A(n18257), .B(n24307), .Z(n24305) );
  XNOR U25889 ( .A(n18256), .B(n24306), .Z(n24307) );
  NAND U25890 ( .A(n24308), .B(n[466]), .Z(n18256) );
  NAND U25891 ( .A(n21523), .B(n[466]), .Z(n24308) );
  XNOR U25892 ( .A(n24309), .B(n24306), .Z(n18257) );
  XOR U25893 ( .A(n24310), .B(n24311), .Z(n24306) );
  AND U25894 ( .A(n18264), .B(n24312), .Z(n24310) );
  XNOR U25895 ( .A(n18263), .B(n24311), .Z(n24312) );
  NAND U25896 ( .A(n24313), .B(n[465]), .Z(n18263) );
  NAND U25897 ( .A(n21523), .B(n[465]), .Z(n24313) );
  XNOR U25898 ( .A(n24314), .B(n24311), .Z(n18264) );
  XOR U25899 ( .A(n24315), .B(n24316), .Z(n24311) );
  AND U25900 ( .A(n18271), .B(n24317), .Z(n24315) );
  XNOR U25901 ( .A(n18270), .B(n24316), .Z(n24317) );
  NAND U25902 ( .A(n24318), .B(n[464]), .Z(n18270) );
  NAND U25903 ( .A(n21523), .B(n[464]), .Z(n24318) );
  XNOR U25904 ( .A(n24319), .B(n24316), .Z(n18271) );
  XOR U25905 ( .A(n24320), .B(n24321), .Z(n24316) );
  AND U25906 ( .A(n18278), .B(n24322), .Z(n24320) );
  XNOR U25907 ( .A(n18277), .B(n24321), .Z(n24322) );
  NAND U25908 ( .A(n24323), .B(n[463]), .Z(n18277) );
  NAND U25909 ( .A(n21523), .B(n[463]), .Z(n24323) );
  XNOR U25910 ( .A(n24324), .B(n24321), .Z(n18278) );
  XOR U25911 ( .A(n24325), .B(n24326), .Z(n24321) );
  AND U25912 ( .A(n18285), .B(n24327), .Z(n24325) );
  XNOR U25913 ( .A(n18284), .B(n24326), .Z(n24327) );
  NAND U25914 ( .A(n24328), .B(n[462]), .Z(n18284) );
  NAND U25915 ( .A(n21523), .B(n[462]), .Z(n24328) );
  XNOR U25916 ( .A(n24329), .B(n24326), .Z(n18285) );
  XOR U25917 ( .A(n24330), .B(n24331), .Z(n24326) );
  AND U25918 ( .A(n18292), .B(n24332), .Z(n24330) );
  XNOR U25919 ( .A(n18291), .B(n24331), .Z(n24332) );
  NAND U25920 ( .A(n24333), .B(n[461]), .Z(n18291) );
  NAND U25921 ( .A(n21523), .B(n[461]), .Z(n24333) );
  XNOR U25922 ( .A(n24334), .B(n24331), .Z(n18292) );
  XOR U25923 ( .A(n24335), .B(n24336), .Z(n24331) );
  AND U25924 ( .A(n18299), .B(n24337), .Z(n24335) );
  XNOR U25925 ( .A(n18298), .B(n24336), .Z(n24337) );
  NAND U25926 ( .A(n24338), .B(n[460]), .Z(n18298) );
  NAND U25927 ( .A(n21523), .B(n[460]), .Z(n24338) );
  XNOR U25928 ( .A(n24339), .B(n24336), .Z(n18299) );
  XOR U25929 ( .A(n24340), .B(n24341), .Z(n24336) );
  AND U25930 ( .A(n18306), .B(n24342), .Z(n24340) );
  XNOR U25931 ( .A(n18305), .B(n24341), .Z(n24342) );
  NAND U25932 ( .A(n24343), .B(n[459]), .Z(n18305) );
  NAND U25933 ( .A(n21523), .B(n[459]), .Z(n24343) );
  XNOR U25934 ( .A(n24344), .B(n24341), .Z(n18306) );
  XOR U25935 ( .A(n24345), .B(n24346), .Z(n24341) );
  AND U25936 ( .A(n18313), .B(n24347), .Z(n24345) );
  XNOR U25937 ( .A(n18312), .B(n24346), .Z(n24347) );
  NAND U25938 ( .A(n24348), .B(n[458]), .Z(n18312) );
  NAND U25939 ( .A(n21523), .B(n[458]), .Z(n24348) );
  XNOR U25940 ( .A(n24349), .B(n24346), .Z(n18313) );
  XOR U25941 ( .A(n24350), .B(n24351), .Z(n24346) );
  AND U25942 ( .A(n18320), .B(n24352), .Z(n24350) );
  XNOR U25943 ( .A(n18319), .B(n24351), .Z(n24352) );
  NAND U25944 ( .A(n24353), .B(n[457]), .Z(n18319) );
  NAND U25945 ( .A(n21523), .B(n[457]), .Z(n24353) );
  XNOR U25946 ( .A(n24354), .B(n24351), .Z(n18320) );
  XOR U25947 ( .A(n24355), .B(n24356), .Z(n24351) );
  AND U25948 ( .A(n18327), .B(n24357), .Z(n24355) );
  XNOR U25949 ( .A(n18326), .B(n24356), .Z(n24357) );
  NAND U25950 ( .A(n24358), .B(n[456]), .Z(n18326) );
  NAND U25951 ( .A(n21523), .B(n[456]), .Z(n24358) );
  XNOR U25952 ( .A(n24359), .B(n24356), .Z(n18327) );
  XOR U25953 ( .A(n24360), .B(n24361), .Z(n24356) );
  AND U25954 ( .A(n18334), .B(n24362), .Z(n24360) );
  XNOR U25955 ( .A(n18333), .B(n24361), .Z(n24362) );
  NAND U25956 ( .A(n24363), .B(n[455]), .Z(n18333) );
  NAND U25957 ( .A(n21523), .B(n[455]), .Z(n24363) );
  XNOR U25958 ( .A(n24364), .B(n24361), .Z(n18334) );
  XOR U25959 ( .A(n24365), .B(n24366), .Z(n24361) );
  AND U25960 ( .A(n18341), .B(n24367), .Z(n24365) );
  XNOR U25961 ( .A(n18340), .B(n24366), .Z(n24367) );
  NAND U25962 ( .A(n24368), .B(n[454]), .Z(n18340) );
  NAND U25963 ( .A(n21523), .B(n[454]), .Z(n24368) );
  XNOR U25964 ( .A(n24369), .B(n24366), .Z(n18341) );
  XOR U25965 ( .A(n24370), .B(n24371), .Z(n24366) );
  AND U25966 ( .A(n18348), .B(n24372), .Z(n24370) );
  XNOR U25967 ( .A(n18347), .B(n24371), .Z(n24372) );
  NAND U25968 ( .A(n24373), .B(n[453]), .Z(n18347) );
  NAND U25969 ( .A(n21523), .B(n[453]), .Z(n24373) );
  XNOR U25970 ( .A(n24374), .B(n24371), .Z(n18348) );
  XOR U25971 ( .A(n24375), .B(n24376), .Z(n24371) );
  AND U25972 ( .A(n18355), .B(n24377), .Z(n24375) );
  XNOR U25973 ( .A(n18354), .B(n24376), .Z(n24377) );
  NAND U25974 ( .A(n24378), .B(n[452]), .Z(n18354) );
  NAND U25975 ( .A(n21523), .B(n[452]), .Z(n24378) );
  XNOR U25976 ( .A(n24379), .B(n24376), .Z(n18355) );
  XOR U25977 ( .A(n24380), .B(n24381), .Z(n24376) );
  AND U25978 ( .A(n18362), .B(n24382), .Z(n24380) );
  XNOR U25979 ( .A(n18361), .B(n24381), .Z(n24382) );
  NAND U25980 ( .A(n24383), .B(n[451]), .Z(n18361) );
  NAND U25981 ( .A(n21523), .B(n[451]), .Z(n24383) );
  XNOR U25982 ( .A(n24384), .B(n24381), .Z(n18362) );
  XOR U25983 ( .A(n24385), .B(n24386), .Z(n24381) );
  AND U25984 ( .A(n18369), .B(n24387), .Z(n24385) );
  XNOR U25985 ( .A(n18368), .B(n24386), .Z(n24387) );
  NAND U25986 ( .A(n24388), .B(n[450]), .Z(n18368) );
  NAND U25987 ( .A(n21523), .B(n[450]), .Z(n24388) );
  XNOR U25988 ( .A(n24389), .B(n24386), .Z(n18369) );
  XOR U25989 ( .A(n24390), .B(n24391), .Z(n24386) );
  AND U25990 ( .A(n18376), .B(n24392), .Z(n24390) );
  XNOR U25991 ( .A(n18375), .B(n24391), .Z(n24392) );
  NAND U25992 ( .A(n24393), .B(n[449]), .Z(n18375) );
  NAND U25993 ( .A(n21523), .B(n[449]), .Z(n24393) );
  XNOR U25994 ( .A(n24394), .B(n24391), .Z(n18376) );
  XOR U25995 ( .A(n24395), .B(n24396), .Z(n24391) );
  AND U25996 ( .A(n18383), .B(n24397), .Z(n24395) );
  XNOR U25997 ( .A(n18382), .B(n24396), .Z(n24397) );
  NAND U25998 ( .A(n24398), .B(n[448]), .Z(n18382) );
  NAND U25999 ( .A(n21523), .B(n[448]), .Z(n24398) );
  XNOR U26000 ( .A(n24399), .B(n24396), .Z(n18383) );
  XOR U26001 ( .A(n24400), .B(n24401), .Z(n24396) );
  AND U26002 ( .A(n18390), .B(n24402), .Z(n24400) );
  XNOR U26003 ( .A(n18389), .B(n24401), .Z(n24402) );
  NAND U26004 ( .A(n24403), .B(n[447]), .Z(n18389) );
  NAND U26005 ( .A(n21523), .B(n[447]), .Z(n24403) );
  XNOR U26006 ( .A(n24404), .B(n24401), .Z(n18390) );
  XOR U26007 ( .A(n24405), .B(n24406), .Z(n24401) );
  AND U26008 ( .A(n18397), .B(n24407), .Z(n24405) );
  XNOR U26009 ( .A(n18396), .B(n24406), .Z(n24407) );
  NAND U26010 ( .A(n24408), .B(n[446]), .Z(n18396) );
  NAND U26011 ( .A(n21523), .B(n[446]), .Z(n24408) );
  XNOR U26012 ( .A(n24409), .B(n24406), .Z(n18397) );
  XOR U26013 ( .A(n24410), .B(n24411), .Z(n24406) );
  AND U26014 ( .A(n18404), .B(n24412), .Z(n24410) );
  XNOR U26015 ( .A(n18403), .B(n24411), .Z(n24412) );
  NAND U26016 ( .A(n24413), .B(n[445]), .Z(n18403) );
  NAND U26017 ( .A(n21523), .B(n[445]), .Z(n24413) );
  XNOR U26018 ( .A(n24414), .B(n24411), .Z(n18404) );
  XOR U26019 ( .A(n24415), .B(n24416), .Z(n24411) );
  AND U26020 ( .A(n18411), .B(n24417), .Z(n24415) );
  XNOR U26021 ( .A(n18410), .B(n24416), .Z(n24417) );
  NAND U26022 ( .A(n24418), .B(n[444]), .Z(n18410) );
  NAND U26023 ( .A(n21523), .B(n[444]), .Z(n24418) );
  XNOR U26024 ( .A(n24419), .B(n24416), .Z(n18411) );
  XOR U26025 ( .A(n24420), .B(n24421), .Z(n24416) );
  AND U26026 ( .A(n18418), .B(n24422), .Z(n24420) );
  XNOR U26027 ( .A(n18417), .B(n24421), .Z(n24422) );
  NAND U26028 ( .A(n24423), .B(n[443]), .Z(n18417) );
  NAND U26029 ( .A(n21523), .B(n[443]), .Z(n24423) );
  XNOR U26030 ( .A(n24424), .B(n24421), .Z(n18418) );
  XOR U26031 ( .A(n24425), .B(n24426), .Z(n24421) );
  AND U26032 ( .A(n18425), .B(n24427), .Z(n24425) );
  XNOR U26033 ( .A(n18424), .B(n24426), .Z(n24427) );
  NAND U26034 ( .A(n24428), .B(n[442]), .Z(n18424) );
  NAND U26035 ( .A(n21523), .B(n[442]), .Z(n24428) );
  XNOR U26036 ( .A(n24429), .B(n24426), .Z(n18425) );
  XOR U26037 ( .A(n24430), .B(n24431), .Z(n24426) );
  AND U26038 ( .A(n18432), .B(n24432), .Z(n24430) );
  XNOR U26039 ( .A(n18431), .B(n24431), .Z(n24432) );
  NAND U26040 ( .A(n24433), .B(n[441]), .Z(n18431) );
  NAND U26041 ( .A(n21523), .B(n[441]), .Z(n24433) );
  XNOR U26042 ( .A(n24434), .B(n24431), .Z(n18432) );
  XOR U26043 ( .A(n24435), .B(n24436), .Z(n24431) );
  AND U26044 ( .A(n18439), .B(n24437), .Z(n24435) );
  XNOR U26045 ( .A(n18438), .B(n24436), .Z(n24437) );
  NAND U26046 ( .A(n24438), .B(n[440]), .Z(n18438) );
  NAND U26047 ( .A(n21523), .B(n[440]), .Z(n24438) );
  XNOR U26048 ( .A(n24439), .B(n24436), .Z(n18439) );
  XOR U26049 ( .A(n24440), .B(n24441), .Z(n24436) );
  AND U26050 ( .A(n18446), .B(n24442), .Z(n24440) );
  XNOR U26051 ( .A(n18445), .B(n24441), .Z(n24442) );
  NAND U26052 ( .A(n24443), .B(n[439]), .Z(n18445) );
  NAND U26053 ( .A(n21523), .B(n[439]), .Z(n24443) );
  XNOR U26054 ( .A(n24444), .B(n24441), .Z(n18446) );
  XOR U26055 ( .A(n24445), .B(n24446), .Z(n24441) );
  AND U26056 ( .A(n18453), .B(n24447), .Z(n24445) );
  XNOR U26057 ( .A(n18452), .B(n24446), .Z(n24447) );
  NAND U26058 ( .A(n24448), .B(n[438]), .Z(n18452) );
  NAND U26059 ( .A(n21523), .B(n[438]), .Z(n24448) );
  XNOR U26060 ( .A(n24449), .B(n24446), .Z(n18453) );
  XOR U26061 ( .A(n24450), .B(n24451), .Z(n24446) );
  AND U26062 ( .A(n18460), .B(n24452), .Z(n24450) );
  XNOR U26063 ( .A(n18459), .B(n24451), .Z(n24452) );
  NAND U26064 ( .A(n24453), .B(n[437]), .Z(n18459) );
  NAND U26065 ( .A(n21523), .B(n[437]), .Z(n24453) );
  XNOR U26066 ( .A(n24454), .B(n24451), .Z(n18460) );
  XOR U26067 ( .A(n24455), .B(n24456), .Z(n24451) );
  AND U26068 ( .A(n18467), .B(n24457), .Z(n24455) );
  XNOR U26069 ( .A(n18466), .B(n24456), .Z(n24457) );
  NAND U26070 ( .A(n24458), .B(n[436]), .Z(n18466) );
  NAND U26071 ( .A(n21523), .B(n[436]), .Z(n24458) );
  XNOR U26072 ( .A(n24459), .B(n24456), .Z(n18467) );
  XOR U26073 ( .A(n24460), .B(n24461), .Z(n24456) );
  AND U26074 ( .A(n18474), .B(n24462), .Z(n24460) );
  XNOR U26075 ( .A(n18473), .B(n24461), .Z(n24462) );
  NAND U26076 ( .A(n24463), .B(n[435]), .Z(n18473) );
  NAND U26077 ( .A(n21523), .B(n[435]), .Z(n24463) );
  XNOR U26078 ( .A(n24464), .B(n24461), .Z(n18474) );
  XOR U26079 ( .A(n24465), .B(n24466), .Z(n24461) );
  AND U26080 ( .A(n18481), .B(n24467), .Z(n24465) );
  XNOR U26081 ( .A(n18480), .B(n24466), .Z(n24467) );
  NAND U26082 ( .A(n24468), .B(n[434]), .Z(n18480) );
  NAND U26083 ( .A(n21523), .B(n[434]), .Z(n24468) );
  XNOR U26084 ( .A(n24469), .B(n24466), .Z(n18481) );
  XOR U26085 ( .A(n24470), .B(n24471), .Z(n24466) );
  AND U26086 ( .A(n18488), .B(n24472), .Z(n24470) );
  XNOR U26087 ( .A(n18487), .B(n24471), .Z(n24472) );
  NAND U26088 ( .A(n24473), .B(n[433]), .Z(n18487) );
  NAND U26089 ( .A(n21523), .B(n[433]), .Z(n24473) );
  XNOR U26090 ( .A(n24474), .B(n24471), .Z(n18488) );
  XOR U26091 ( .A(n24475), .B(n24476), .Z(n24471) );
  AND U26092 ( .A(n18495), .B(n24477), .Z(n24475) );
  XNOR U26093 ( .A(n18494), .B(n24476), .Z(n24477) );
  NAND U26094 ( .A(n24478), .B(n[432]), .Z(n18494) );
  NAND U26095 ( .A(n21523), .B(n[432]), .Z(n24478) );
  XNOR U26096 ( .A(n24479), .B(n24476), .Z(n18495) );
  XOR U26097 ( .A(n24480), .B(n24481), .Z(n24476) );
  AND U26098 ( .A(n18502), .B(n24482), .Z(n24480) );
  XNOR U26099 ( .A(n18501), .B(n24481), .Z(n24482) );
  NAND U26100 ( .A(n24483), .B(n[431]), .Z(n18501) );
  NAND U26101 ( .A(n21523), .B(n[431]), .Z(n24483) );
  XNOR U26102 ( .A(n24484), .B(n24481), .Z(n18502) );
  XOR U26103 ( .A(n24485), .B(n24486), .Z(n24481) );
  AND U26104 ( .A(n18509), .B(n24487), .Z(n24485) );
  XNOR U26105 ( .A(n18508), .B(n24486), .Z(n24487) );
  NAND U26106 ( .A(n24488), .B(n[430]), .Z(n18508) );
  NAND U26107 ( .A(n21523), .B(n[430]), .Z(n24488) );
  XNOR U26108 ( .A(n24489), .B(n24486), .Z(n18509) );
  XOR U26109 ( .A(n24490), .B(n24491), .Z(n24486) );
  AND U26110 ( .A(n18516), .B(n24492), .Z(n24490) );
  XNOR U26111 ( .A(n18515), .B(n24491), .Z(n24492) );
  NAND U26112 ( .A(n24493), .B(n[429]), .Z(n18515) );
  NAND U26113 ( .A(n21523), .B(n[429]), .Z(n24493) );
  XNOR U26114 ( .A(n24494), .B(n24491), .Z(n18516) );
  XOR U26115 ( .A(n24495), .B(n24496), .Z(n24491) );
  AND U26116 ( .A(n18523), .B(n24497), .Z(n24495) );
  XNOR U26117 ( .A(n18522), .B(n24496), .Z(n24497) );
  NAND U26118 ( .A(n24498), .B(n[428]), .Z(n18522) );
  NAND U26119 ( .A(n21523), .B(n[428]), .Z(n24498) );
  XNOR U26120 ( .A(n24499), .B(n24496), .Z(n18523) );
  XOR U26121 ( .A(n24500), .B(n24501), .Z(n24496) );
  AND U26122 ( .A(n18530), .B(n24502), .Z(n24500) );
  XNOR U26123 ( .A(n18529), .B(n24501), .Z(n24502) );
  NAND U26124 ( .A(n24503), .B(n[427]), .Z(n18529) );
  NAND U26125 ( .A(n21523), .B(n[427]), .Z(n24503) );
  XNOR U26126 ( .A(n24504), .B(n24501), .Z(n18530) );
  XOR U26127 ( .A(n24505), .B(n24506), .Z(n24501) );
  AND U26128 ( .A(n18537), .B(n24507), .Z(n24505) );
  XNOR U26129 ( .A(n18536), .B(n24506), .Z(n24507) );
  NAND U26130 ( .A(n24508), .B(n[426]), .Z(n18536) );
  NAND U26131 ( .A(n21523), .B(n[426]), .Z(n24508) );
  XNOR U26132 ( .A(n24509), .B(n24506), .Z(n18537) );
  XOR U26133 ( .A(n24510), .B(n24511), .Z(n24506) );
  AND U26134 ( .A(n18544), .B(n24512), .Z(n24510) );
  XNOR U26135 ( .A(n18543), .B(n24511), .Z(n24512) );
  NAND U26136 ( .A(n24513), .B(n[425]), .Z(n18543) );
  NAND U26137 ( .A(n21523), .B(n[425]), .Z(n24513) );
  XNOR U26138 ( .A(n24514), .B(n24511), .Z(n18544) );
  XOR U26139 ( .A(n24515), .B(n24516), .Z(n24511) );
  AND U26140 ( .A(n18551), .B(n24517), .Z(n24515) );
  XNOR U26141 ( .A(n18550), .B(n24516), .Z(n24517) );
  NAND U26142 ( .A(n24518), .B(n[424]), .Z(n18550) );
  NAND U26143 ( .A(n21523), .B(n[424]), .Z(n24518) );
  XNOR U26144 ( .A(n24519), .B(n24516), .Z(n18551) );
  XOR U26145 ( .A(n24520), .B(n24521), .Z(n24516) );
  AND U26146 ( .A(n18558), .B(n24522), .Z(n24520) );
  XNOR U26147 ( .A(n18557), .B(n24521), .Z(n24522) );
  NAND U26148 ( .A(n24523), .B(n[423]), .Z(n18557) );
  NAND U26149 ( .A(n21523), .B(n[423]), .Z(n24523) );
  XNOR U26150 ( .A(n24524), .B(n24521), .Z(n18558) );
  XOR U26151 ( .A(n24525), .B(n24526), .Z(n24521) );
  AND U26152 ( .A(n18565), .B(n24527), .Z(n24525) );
  XNOR U26153 ( .A(n18564), .B(n24526), .Z(n24527) );
  NAND U26154 ( .A(n24528), .B(n[422]), .Z(n18564) );
  NAND U26155 ( .A(n21523), .B(n[422]), .Z(n24528) );
  XNOR U26156 ( .A(n24529), .B(n24526), .Z(n18565) );
  XOR U26157 ( .A(n24530), .B(n24531), .Z(n24526) );
  AND U26158 ( .A(n18572), .B(n24532), .Z(n24530) );
  XNOR U26159 ( .A(n18571), .B(n24531), .Z(n24532) );
  NAND U26160 ( .A(n24533), .B(n[421]), .Z(n18571) );
  NAND U26161 ( .A(n21523), .B(n[421]), .Z(n24533) );
  XNOR U26162 ( .A(n24534), .B(n24531), .Z(n18572) );
  XOR U26163 ( .A(n24535), .B(n24536), .Z(n24531) );
  AND U26164 ( .A(n18579), .B(n24537), .Z(n24535) );
  XNOR U26165 ( .A(n18578), .B(n24536), .Z(n24537) );
  NAND U26166 ( .A(n24538), .B(n[420]), .Z(n18578) );
  NAND U26167 ( .A(n21523), .B(n[420]), .Z(n24538) );
  XNOR U26168 ( .A(n24539), .B(n24536), .Z(n18579) );
  XOR U26169 ( .A(n24540), .B(n24541), .Z(n24536) );
  AND U26170 ( .A(n18586), .B(n24542), .Z(n24540) );
  XNOR U26171 ( .A(n18585), .B(n24541), .Z(n24542) );
  NAND U26172 ( .A(n24543), .B(n[419]), .Z(n18585) );
  NAND U26173 ( .A(n21523), .B(n[419]), .Z(n24543) );
  XNOR U26174 ( .A(n24544), .B(n24541), .Z(n18586) );
  XOR U26175 ( .A(n24545), .B(n24546), .Z(n24541) );
  AND U26176 ( .A(n18593), .B(n24547), .Z(n24545) );
  XNOR U26177 ( .A(n18592), .B(n24546), .Z(n24547) );
  NAND U26178 ( .A(n24548), .B(n[418]), .Z(n18592) );
  NAND U26179 ( .A(n21523), .B(n[418]), .Z(n24548) );
  XNOR U26180 ( .A(n24549), .B(n24546), .Z(n18593) );
  XOR U26181 ( .A(n24550), .B(n24551), .Z(n24546) );
  AND U26182 ( .A(n18600), .B(n24552), .Z(n24550) );
  XNOR U26183 ( .A(n18599), .B(n24551), .Z(n24552) );
  NAND U26184 ( .A(n24553), .B(n[417]), .Z(n18599) );
  NAND U26185 ( .A(n21523), .B(n[417]), .Z(n24553) );
  XNOR U26186 ( .A(n24554), .B(n24551), .Z(n18600) );
  XOR U26187 ( .A(n24555), .B(n24556), .Z(n24551) );
  AND U26188 ( .A(n18607), .B(n24557), .Z(n24555) );
  XNOR U26189 ( .A(n18606), .B(n24556), .Z(n24557) );
  NAND U26190 ( .A(n24558), .B(n[416]), .Z(n18606) );
  NAND U26191 ( .A(n21523), .B(n[416]), .Z(n24558) );
  XNOR U26192 ( .A(n24559), .B(n24556), .Z(n18607) );
  XOR U26193 ( .A(n24560), .B(n24561), .Z(n24556) );
  AND U26194 ( .A(n18614), .B(n24562), .Z(n24560) );
  XNOR U26195 ( .A(n18613), .B(n24561), .Z(n24562) );
  NAND U26196 ( .A(n24563), .B(n[415]), .Z(n18613) );
  NAND U26197 ( .A(n21523), .B(n[415]), .Z(n24563) );
  XNOR U26198 ( .A(n24564), .B(n24561), .Z(n18614) );
  XOR U26199 ( .A(n24565), .B(n24566), .Z(n24561) );
  AND U26200 ( .A(n18621), .B(n24567), .Z(n24565) );
  XNOR U26201 ( .A(n18620), .B(n24566), .Z(n24567) );
  NAND U26202 ( .A(n24568), .B(n[414]), .Z(n18620) );
  NAND U26203 ( .A(n21523), .B(n[414]), .Z(n24568) );
  XNOR U26204 ( .A(n24569), .B(n24566), .Z(n18621) );
  XOR U26205 ( .A(n24570), .B(n24571), .Z(n24566) );
  AND U26206 ( .A(n18628), .B(n24572), .Z(n24570) );
  XNOR U26207 ( .A(n18627), .B(n24571), .Z(n24572) );
  NAND U26208 ( .A(n24573), .B(n[413]), .Z(n18627) );
  NAND U26209 ( .A(n21523), .B(n[413]), .Z(n24573) );
  XNOR U26210 ( .A(n24574), .B(n24571), .Z(n18628) );
  XOR U26211 ( .A(n24575), .B(n24576), .Z(n24571) );
  AND U26212 ( .A(n18635), .B(n24577), .Z(n24575) );
  XNOR U26213 ( .A(n18634), .B(n24576), .Z(n24577) );
  NAND U26214 ( .A(n24578), .B(n[412]), .Z(n18634) );
  NAND U26215 ( .A(n21523), .B(n[412]), .Z(n24578) );
  XNOR U26216 ( .A(n24579), .B(n24576), .Z(n18635) );
  XOR U26217 ( .A(n24580), .B(n24581), .Z(n24576) );
  AND U26218 ( .A(n18642), .B(n24582), .Z(n24580) );
  XNOR U26219 ( .A(n18641), .B(n24581), .Z(n24582) );
  NAND U26220 ( .A(n24583), .B(n[411]), .Z(n18641) );
  NAND U26221 ( .A(n21523), .B(n[411]), .Z(n24583) );
  XNOR U26222 ( .A(n24584), .B(n24581), .Z(n18642) );
  XOR U26223 ( .A(n24585), .B(n24586), .Z(n24581) );
  AND U26224 ( .A(n18649), .B(n24587), .Z(n24585) );
  XNOR U26225 ( .A(n18648), .B(n24586), .Z(n24587) );
  NAND U26226 ( .A(n24588), .B(n[410]), .Z(n18648) );
  NAND U26227 ( .A(n21523), .B(n[410]), .Z(n24588) );
  XNOR U26228 ( .A(n24589), .B(n24586), .Z(n18649) );
  XOR U26229 ( .A(n24590), .B(n24591), .Z(n24586) );
  AND U26230 ( .A(n18656), .B(n24592), .Z(n24590) );
  XNOR U26231 ( .A(n18655), .B(n24591), .Z(n24592) );
  NAND U26232 ( .A(n24593), .B(n[409]), .Z(n18655) );
  NAND U26233 ( .A(n21523), .B(n[409]), .Z(n24593) );
  XNOR U26234 ( .A(n24594), .B(n24591), .Z(n18656) );
  XOR U26235 ( .A(n24595), .B(n24596), .Z(n24591) );
  AND U26236 ( .A(n18663), .B(n24597), .Z(n24595) );
  XNOR U26237 ( .A(n18662), .B(n24596), .Z(n24597) );
  NAND U26238 ( .A(n24598), .B(n[408]), .Z(n18662) );
  NAND U26239 ( .A(n21523), .B(n[408]), .Z(n24598) );
  XNOR U26240 ( .A(n24599), .B(n24596), .Z(n18663) );
  XOR U26241 ( .A(n24600), .B(n24601), .Z(n24596) );
  AND U26242 ( .A(n18670), .B(n24602), .Z(n24600) );
  XNOR U26243 ( .A(n18669), .B(n24601), .Z(n24602) );
  NAND U26244 ( .A(n24603), .B(n[407]), .Z(n18669) );
  NAND U26245 ( .A(n21523), .B(n[407]), .Z(n24603) );
  XNOR U26246 ( .A(n24604), .B(n24601), .Z(n18670) );
  XOR U26247 ( .A(n24605), .B(n24606), .Z(n24601) );
  AND U26248 ( .A(n18677), .B(n24607), .Z(n24605) );
  XNOR U26249 ( .A(n18676), .B(n24606), .Z(n24607) );
  NAND U26250 ( .A(n24608), .B(n[406]), .Z(n18676) );
  NAND U26251 ( .A(n21523), .B(n[406]), .Z(n24608) );
  XNOR U26252 ( .A(n24609), .B(n24606), .Z(n18677) );
  XOR U26253 ( .A(n24610), .B(n24611), .Z(n24606) );
  AND U26254 ( .A(n18684), .B(n24612), .Z(n24610) );
  XNOR U26255 ( .A(n18683), .B(n24611), .Z(n24612) );
  NAND U26256 ( .A(n24613), .B(n[405]), .Z(n18683) );
  NAND U26257 ( .A(n21523), .B(n[405]), .Z(n24613) );
  XNOR U26258 ( .A(n24614), .B(n24611), .Z(n18684) );
  XOR U26259 ( .A(n24615), .B(n24616), .Z(n24611) );
  AND U26260 ( .A(n18691), .B(n24617), .Z(n24615) );
  XNOR U26261 ( .A(n18690), .B(n24616), .Z(n24617) );
  NAND U26262 ( .A(n24618), .B(n[404]), .Z(n18690) );
  NAND U26263 ( .A(n21523), .B(n[404]), .Z(n24618) );
  XNOR U26264 ( .A(n24619), .B(n24616), .Z(n18691) );
  XOR U26265 ( .A(n24620), .B(n24621), .Z(n24616) );
  AND U26266 ( .A(n18698), .B(n24622), .Z(n24620) );
  XNOR U26267 ( .A(n18697), .B(n24621), .Z(n24622) );
  NAND U26268 ( .A(n24623), .B(n[403]), .Z(n18697) );
  NAND U26269 ( .A(n21523), .B(n[403]), .Z(n24623) );
  XNOR U26270 ( .A(n24624), .B(n24621), .Z(n18698) );
  XOR U26271 ( .A(n24625), .B(n24626), .Z(n24621) );
  AND U26272 ( .A(n18705), .B(n24627), .Z(n24625) );
  XNOR U26273 ( .A(n18704), .B(n24626), .Z(n24627) );
  NAND U26274 ( .A(n24628), .B(n[402]), .Z(n18704) );
  NAND U26275 ( .A(n21523), .B(n[402]), .Z(n24628) );
  XNOR U26276 ( .A(n24629), .B(n24626), .Z(n18705) );
  XOR U26277 ( .A(n24630), .B(n24631), .Z(n24626) );
  AND U26278 ( .A(n18712), .B(n24632), .Z(n24630) );
  XNOR U26279 ( .A(n18711), .B(n24631), .Z(n24632) );
  NAND U26280 ( .A(n24633), .B(n[401]), .Z(n18711) );
  NAND U26281 ( .A(n21523), .B(n[401]), .Z(n24633) );
  XNOR U26282 ( .A(n24634), .B(n24631), .Z(n18712) );
  XOR U26283 ( .A(n24635), .B(n24636), .Z(n24631) );
  AND U26284 ( .A(n18719), .B(n24637), .Z(n24635) );
  XNOR U26285 ( .A(n18718), .B(n24636), .Z(n24637) );
  NAND U26286 ( .A(n24638), .B(n[400]), .Z(n18718) );
  NAND U26287 ( .A(n21523), .B(n[400]), .Z(n24638) );
  XNOR U26288 ( .A(n24639), .B(n24636), .Z(n18719) );
  XOR U26289 ( .A(n24640), .B(n24641), .Z(n24636) );
  AND U26290 ( .A(n18726), .B(n24642), .Z(n24640) );
  XNOR U26291 ( .A(n18725), .B(n24641), .Z(n24642) );
  NAND U26292 ( .A(n24643), .B(n[399]), .Z(n18725) );
  NAND U26293 ( .A(n21523), .B(n[399]), .Z(n24643) );
  XNOR U26294 ( .A(n24644), .B(n24641), .Z(n18726) );
  XOR U26295 ( .A(n24645), .B(n24646), .Z(n24641) );
  AND U26296 ( .A(n18733), .B(n24647), .Z(n24645) );
  XNOR U26297 ( .A(n18732), .B(n24646), .Z(n24647) );
  NAND U26298 ( .A(n24648), .B(n[398]), .Z(n18732) );
  NAND U26299 ( .A(n21523), .B(n[398]), .Z(n24648) );
  XNOR U26300 ( .A(n24649), .B(n24646), .Z(n18733) );
  XOR U26301 ( .A(n24650), .B(n24651), .Z(n24646) );
  AND U26302 ( .A(n18740), .B(n24652), .Z(n24650) );
  XNOR U26303 ( .A(n18739), .B(n24651), .Z(n24652) );
  NAND U26304 ( .A(n24653), .B(n[397]), .Z(n18739) );
  NAND U26305 ( .A(n21523), .B(n[397]), .Z(n24653) );
  XNOR U26306 ( .A(n24654), .B(n24651), .Z(n18740) );
  XOR U26307 ( .A(n24655), .B(n24656), .Z(n24651) );
  AND U26308 ( .A(n18747), .B(n24657), .Z(n24655) );
  XNOR U26309 ( .A(n18746), .B(n24656), .Z(n24657) );
  NAND U26310 ( .A(n24658), .B(n[396]), .Z(n18746) );
  NAND U26311 ( .A(n21523), .B(n[396]), .Z(n24658) );
  XNOR U26312 ( .A(n24659), .B(n24656), .Z(n18747) );
  XOR U26313 ( .A(n24660), .B(n24661), .Z(n24656) );
  AND U26314 ( .A(n18754), .B(n24662), .Z(n24660) );
  XNOR U26315 ( .A(n18753), .B(n24661), .Z(n24662) );
  NAND U26316 ( .A(n24663), .B(n[395]), .Z(n18753) );
  NAND U26317 ( .A(n21523), .B(n[395]), .Z(n24663) );
  XNOR U26318 ( .A(n24664), .B(n24661), .Z(n18754) );
  XOR U26319 ( .A(n24665), .B(n24666), .Z(n24661) );
  AND U26320 ( .A(n18761), .B(n24667), .Z(n24665) );
  XNOR U26321 ( .A(n18760), .B(n24666), .Z(n24667) );
  NAND U26322 ( .A(n24668), .B(n[394]), .Z(n18760) );
  NAND U26323 ( .A(n21523), .B(n[394]), .Z(n24668) );
  XNOR U26324 ( .A(n24669), .B(n24666), .Z(n18761) );
  XOR U26325 ( .A(n24670), .B(n24671), .Z(n24666) );
  AND U26326 ( .A(n18768), .B(n24672), .Z(n24670) );
  XNOR U26327 ( .A(n18767), .B(n24671), .Z(n24672) );
  NAND U26328 ( .A(n24673), .B(n[393]), .Z(n18767) );
  NAND U26329 ( .A(n21523), .B(n[393]), .Z(n24673) );
  XNOR U26330 ( .A(n24674), .B(n24671), .Z(n18768) );
  XOR U26331 ( .A(n24675), .B(n24676), .Z(n24671) );
  AND U26332 ( .A(n18775), .B(n24677), .Z(n24675) );
  XNOR U26333 ( .A(n18774), .B(n24676), .Z(n24677) );
  NAND U26334 ( .A(n24678), .B(n[392]), .Z(n18774) );
  NAND U26335 ( .A(n21523), .B(n[392]), .Z(n24678) );
  XNOR U26336 ( .A(n24679), .B(n24676), .Z(n18775) );
  XOR U26337 ( .A(n24680), .B(n24681), .Z(n24676) );
  AND U26338 ( .A(n18782), .B(n24682), .Z(n24680) );
  XNOR U26339 ( .A(n18781), .B(n24681), .Z(n24682) );
  NAND U26340 ( .A(n24683), .B(n[391]), .Z(n18781) );
  NAND U26341 ( .A(n21523), .B(n[391]), .Z(n24683) );
  XNOR U26342 ( .A(n24684), .B(n24681), .Z(n18782) );
  XOR U26343 ( .A(n24685), .B(n24686), .Z(n24681) );
  AND U26344 ( .A(n18789), .B(n24687), .Z(n24685) );
  XNOR U26345 ( .A(n18788), .B(n24686), .Z(n24687) );
  NAND U26346 ( .A(n24688), .B(n[390]), .Z(n18788) );
  NAND U26347 ( .A(n21523), .B(n[390]), .Z(n24688) );
  XNOR U26348 ( .A(n24689), .B(n24686), .Z(n18789) );
  XOR U26349 ( .A(n24690), .B(n24691), .Z(n24686) );
  AND U26350 ( .A(n18796), .B(n24692), .Z(n24690) );
  XNOR U26351 ( .A(n18795), .B(n24691), .Z(n24692) );
  NAND U26352 ( .A(n24693), .B(n[389]), .Z(n18795) );
  NAND U26353 ( .A(n21523), .B(n[389]), .Z(n24693) );
  XNOR U26354 ( .A(n24694), .B(n24691), .Z(n18796) );
  XOR U26355 ( .A(n24695), .B(n24696), .Z(n24691) );
  AND U26356 ( .A(n18803), .B(n24697), .Z(n24695) );
  XNOR U26357 ( .A(n18802), .B(n24696), .Z(n24697) );
  NAND U26358 ( .A(n24698), .B(n[388]), .Z(n18802) );
  NAND U26359 ( .A(n21523), .B(n[388]), .Z(n24698) );
  XNOR U26360 ( .A(n24699), .B(n24696), .Z(n18803) );
  XOR U26361 ( .A(n24700), .B(n24701), .Z(n24696) );
  AND U26362 ( .A(n18810), .B(n24702), .Z(n24700) );
  XNOR U26363 ( .A(n18809), .B(n24701), .Z(n24702) );
  NAND U26364 ( .A(n24703), .B(n[387]), .Z(n18809) );
  NAND U26365 ( .A(n21523), .B(n[387]), .Z(n24703) );
  XNOR U26366 ( .A(n24704), .B(n24701), .Z(n18810) );
  XOR U26367 ( .A(n24705), .B(n24706), .Z(n24701) );
  AND U26368 ( .A(n18817), .B(n24707), .Z(n24705) );
  XNOR U26369 ( .A(n18816), .B(n24706), .Z(n24707) );
  NAND U26370 ( .A(n24708), .B(n[386]), .Z(n18816) );
  NAND U26371 ( .A(n21523), .B(n[386]), .Z(n24708) );
  XNOR U26372 ( .A(n24709), .B(n24706), .Z(n18817) );
  XOR U26373 ( .A(n24710), .B(n24711), .Z(n24706) );
  AND U26374 ( .A(n18824), .B(n24712), .Z(n24710) );
  XNOR U26375 ( .A(n18823), .B(n24711), .Z(n24712) );
  NAND U26376 ( .A(n24713), .B(n[385]), .Z(n18823) );
  NAND U26377 ( .A(n21523), .B(n[385]), .Z(n24713) );
  XNOR U26378 ( .A(n24714), .B(n24711), .Z(n18824) );
  XOR U26379 ( .A(n24715), .B(n24716), .Z(n24711) );
  AND U26380 ( .A(n18831), .B(n24717), .Z(n24715) );
  XNOR U26381 ( .A(n18830), .B(n24716), .Z(n24717) );
  NAND U26382 ( .A(n24718), .B(n[384]), .Z(n18830) );
  NAND U26383 ( .A(n21523), .B(n[384]), .Z(n24718) );
  XNOR U26384 ( .A(n24719), .B(n24716), .Z(n18831) );
  XOR U26385 ( .A(n24720), .B(n24721), .Z(n24716) );
  AND U26386 ( .A(n18838), .B(n24722), .Z(n24720) );
  XNOR U26387 ( .A(n18837), .B(n24721), .Z(n24722) );
  NAND U26388 ( .A(n24723), .B(n[383]), .Z(n18837) );
  NAND U26389 ( .A(n21523), .B(n[383]), .Z(n24723) );
  XNOR U26390 ( .A(n24724), .B(n24721), .Z(n18838) );
  XOR U26391 ( .A(n24725), .B(n24726), .Z(n24721) );
  AND U26392 ( .A(n18845), .B(n24727), .Z(n24725) );
  XNOR U26393 ( .A(n18844), .B(n24726), .Z(n24727) );
  NAND U26394 ( .A(n24728), .B(n[382]), .Z(n18844) );
  NAND U26395 ( .A(n21523), .B(n[382]), .Z(n24728) );
  XNOR U26396 ( .A(n24729), .B(n24726), .Z(n18845) );
  XOR U26397 ( .A(n24730), .B(n24731), .Z(n24726) );
  AND U26398 ( .A(n18852), .B(n24732), .Z(n24730) );
  XNOR U26399 ( .A(n18851), .B(n24731), .Z(n24732) );
  NAND U26400 ( .A(n24733), .B(n[381]), .Z(n18851) );
  NAND U26401 ( .A(n21523), .B(n[381]), .Z(n24733) );
  XNOR U26402 ( .A(n24734), .B(n24731), .Z(n18852) );
  XOR U26403 ( .A(n24735), .B(n24736), .Z(n24731) );
  AND U26404 ( .A(n18859), .B(n24737), .Z(n24735) );
  XNOR U26405 ( .A(n18858), .B(n24736), .Z(n24737) );
  NAND U26406 ( .A(n24738), .B(n[380]), .Z(n18858) );
  NAND U26407 ( .A(n21523), .B(n[380]), .Z(n24738) );
  XNOR U26408 ( .A(n24739), .B(n24736), .Z(n18859) );
  XOR U26409 ( .A(n24740), .B(n24741), .Z(n24736) );
  AND U26410 ( .A(n18866), .B(n24742), .Z(n24740) );
  XNOR U26411 ( .A(n18865), .B(n24741), .Z(n24742) );
  NAND U26412 ( .A(n24743), .B(n[379]), .Z(n18865) );
  NAND U26413 ( .A(n21523), .B(n[379]), .Z(n24743) );
  XNOR U26414 ( .A(n24744), .B(n24741), .Z(n18866) );
  XOR U26415 ( .A(n24745), .B(n24746), .Z(n24741) );
  AND U26416 ( .A(n18873), .B(n24747), .Z(n24745) );
  XNOR U26417 ( .A(n18872), .B(n24746), .Z(n24747) );
  NAND U26418 ( .A(n24748), .B(n[378]), .Z(n18872) );
  NAND U26419 ( .A(n21523), .B(n[378]), .Z(n24748) );
  XNOR U26420 ( .A(n24749), .B(n24746), .Z(n18873) );
  XOR U26421 ( .A(n24750), .B(n24751), .Z(n24746) );
  AND U26422 ( .A(n18880), .B(n24752), .Z(n24750) );
  XNOR U26423 ( .A(n18879), .B(n24751), .Z(n24752) );
  NAND U26424 ( .A(n24753), .B(n[377]), .Z(n18879) );
  NAND U26425 ( .A(n21523), .B(n[377]), .Z(n24753) );
  XNOR U26426 ( .A(n24754), .B(n24751), .Z(n18880) );
  XOR U26427 ( .A(n24755), .B(n24756), .Z(n24751) );
  AND U26428 ( .A(n18887), .B(n24757), .Z(n24755) );
  XNOR U26429 ( .A(n18886), .B(n24756), .Z(n24757) );
  NAND U26430 ( .A(n24758), .B(n[376]), .Z(n18886) );
  NAND U26431 ( .A(n21523), .B(n[376]), .Z(n24758) );
  XNOR U26432 ( .A(n24759), .B(n24756), .Z(n18887) );
  XOR U26433 ( .A(n24760), .B(n24761), .Z(n24756) );
  AND U26434 ( .A(n18894), .B(n24762), .Z(n24760) );
  XNOR U26435 ( .A(n18893), .B(n24761), .Z(n24762) );
  NAND U26436 ( .A(n24763), .B(n[375]), .Z(n18893) );
  NAND U26437 ( .A(n21523), .B(n[375]), .Z(n24763) );
  XNOR U26438 ( .A(n24764), .B(n24761), .Z(n18894) );
  XOR U26439 ( .A(n24765), .B(n24766), .Z(n24761) );
  AND U26440 ( .A(n18901), .B(n24767), .Z(n24765) );
  XNOR U26441 ( .A(n18900), .B(n24766), .Z(n24767) );
  NAND U26442 ( .A(n24768), .B(n[374]), .Z(n18900) );
  NAND U26443 ( .A(n21523), .B(n[374]), .Z(n24768) );
  XNOR U26444 ( .A(n24769), .B(n24766), .Z(n18901) );
  XOR U26445 ( .A(n24770), .B(n24771), .Z(n24766) );
  AND U26446 ( .A(n18908), .B(n24772), .Z(n24770) );
  XNOR U26447 ( .A(n18907), .B(n24771), .Z(n24772) );
  NAND U26448 ( .A(n24773), .B(n[373]), .Z(n18907) );
  NAND U26449 ( .A(n21523), .B(n[373]), .Z(n24773) );
  XNOR U26450 ( .A(n24774), .B(n24771), .Z(n18908) );
  XOR U26451 ( .A(n24775), .B(n24776), .Z(n24771) );
  AND U26452 ( .A(n18915), .B(n24777), .Z(n24775) );
  XNOR U26453 ( .A(n18914), .B(n24776), .Z(n24777) );
  NAND U26454 ( .A(n24778), .B(n[372]), .Z(n18914) );
  NAND U26455 ( .A(n21523), .B(n[372]), .Z(n24778) );
  XNOR U26456 ( .A(n24779), .B(n24776), .Z(n18915) );
  XOR U26457 ( .A(n24780), .B(n24781), .Z(n24776) );
  AND U26458 ( .A(n18922), .B(n24782), .Z(n24780) );
  XNOR U26459 ( .A(n18921), .B(n24781), .Z(n24782) );
  NAND U26460 ( .A(n24783), .B(n[371]), .Z(n18921) );
  NAND U26461 ( .A(n21523), .B(n[371]), .Z(n24783) );
  XNOR U26462 ( .A(n24784), .B(n24781), .Z(n18922) );
  XOR U26463 ( .A(n24785), .B(n24786), .Z(n24781) );
  AND U26464 ( .A(n18929), .B(n24787), .Z(n24785) );
  XNOR U26465 ( .A(n18928), .B(n24786), .Z(n24787) );
  NAND U26466 ( .A(n24788), .B(n[370]), .Z(n18928) );
  NAND U26467 ( .A(n21523), .B(n[370]), .Z(n24788) );
  XNOR U26468 ( .A(n24789), .B(n24786), .Z(n18929) );
  XOR U26469 ( .A(n24790), .B(n24791), .Z(n24786) );
  AND U26470 ( .A(n18936), .B(n24792), .Z(n24790) );
  XNOR U26471 ( .A(n18935), .B(n24791), .Z(n24792) );
  NAND U26472 ( .A(n24793), .B(n[369]), .Z(n18935) );
  NAND U26473 ( .A(n21523), .B(n[369]), .Z(n24793) );
  XNOR U26474 ( .A(n24794), .B(n24791), .Z(n18936) );
  XOR U26475 ( .A(n24795), .B(n24796), .Z(n24791) );
  AND U26476 ( .A(n18943), .B(n24797), .Z(n24795) );
  XNOR U26477 ( .A(n18942), .B(n24796), .Z(n24797) );
  NAND U26478 ( .A(n24798), .B(n[368]), .Z(n18942) );
  NAND U26479 ( .A(n21523), .B(n[368]), .Z(n24798) );
  XNOR U26480 ( .A(n24799), .B(n24796), .Z(n18943) );
  XOR U26481 ( .A(n24800), .B(n24801), .Z(n24796) );
  AND U26482 ( .A(n18950), .B(n24802), .Z(n24800) );
  XNOR U26483 ( .A(n18949), .B(n24801), .Z(n24802) );
  NAND U26484 ( .A(n24803), .B(n[367]), .Z(n18949) );
  NAND U26485 ( .A(n21523), .B(n[367]), .Z(n24803) );
  XNOR U26486 ( .A(n24804), .B(n24801), .Z(n18950) );
  XOR U26487 ( .A(n24805), .B(n24806), .Z(n24801) );
  AND U26488 ( .A(n18957), .B(n24807), .Z(n24805) );
  XNOR U26489 ( .A(n18956), .B(n24806), .Z(n24807) );
  NAND U26490 ( .A(n24808), .B(n[366]), .Z(n18956) );
  NAND U26491 ( .A(n21523), .B(n[366]), .Z(n24808) );
  XNOR U26492 ( .A(n24809), .B(n24806), .Z(n18957) );
  XOR U26493 ( .A(n24810), .B(n24811), .Z(n24806) );
  AND U26494 ( .A(n18964), .B(n24812), .Z(n24810) );
  XNOR U26495 ( .A(n18963), .B(n24811), .Z(n24812) );
  NAND U26496 ( .A(n24813), .B(n[365]), .Z(n18963) );
  NAND U26497 ( .A(n21523), .B(n[365]), .Z(n24813) );
  XNOR U26498 ( .A(n24814), .B(n24811), .Z(n18964) );
  XOR U26499 ( .A(n24815), .B(n24816), .Z(n24811) );
  AND U26500 ( .A(n18971), .B(n24817), .Z(n24815) );
  XNOR U26501 ( .A(n18970), .B(n24816), .Z(n24817) );
  NAND U26502 ( .A(n24818), .B(n[364]), .Z(n18970) );
  NAND U26503 ( .A(n21523), .B(n[364]), .Z(n24818) );
  XNOR U26504 ( .A(n24819), .B(n24816), .Z(n18971) );
  XOR U26505 ( .A(n24820), .B(n24821), .Z(n24816) );
  AND U26506 ( .A(n18978), .B(n24822), .Z(n24820) );
  XNOR U26507 ( .A(n18977), .B(n24821), .Z(n24822) );
  NAND U26508 ( .A(n24823), .B(n[363]), .Z(n18977) );
  NAND U26509 ( .A(n21523), .B(n[363]), .Z(n24823) );
  XNOR U26510 ( .A(n24824), .B(n24821), .Z(n18978) );
  XOR U26511 ( .A(n24825), .B(n24826), .Z(n24821) );
  AND U26512 ( .A(n18985), .B(n24827), .Z(n24825) );
  XNOR U26513 ( .A(n18984), .B(n24826), .Z(n24827) );
  NAND U26514 ( .A(n24828), .B(n[362]), .Z(n18984) );
  NAND U26515 ( .A(n21523), .B(n[362]), .Z(n24828) );
  XNOR U26516 ( .A(n24829), .B(n24826), .Z(n18985) );
  XOR U26517 ( .A(n24830), .B(n24831), .Z(n24826) );
  AND U26518 ( .A(n18992), .B(n24832), .Z(n24830) );
  XNOR U26519 ( .A(n18991), .B(n24831), .Z(n24832) );
  NAND U26520 ( .A(n24833), .B(n[361]), .Z(n18991) );
  NAND U26521 ( .A(n21523), .B(n[361]), .Z(n24833) );
  XNOR U26522 ( .A(n24834), .B(n24831), .Z(n18992) );
  XOR U26523 ( .A(n24835), .B(n24836), .Z(n24831) );
  AND U26524 ( .A(n18999), .B(n24837), .Z(n24835) );
  XNOR U26525 ( .A(n18998), .B(n24836), .Z(n24837) );
  NAND U26526 ( .A(n24838), .B(n[360]), .Z(n18998) );
  NAND U26527 ( .A(n21523), .B(n[360]), .Z(n24838) );
  XNOR U26528 ( .A(n24839), .B(n24836), .Z(n18999) );
  XOR U26529 ( .A(n24840), .B(n24841), .Z(n24836) );
  AND U26530 ( .A(n19006), .B(n24842), .Z(n24840) );
  XNOR U26531 ( .A(n19005), .B(n24841), .Z(n24842) );
  NAND U26532 ( .A(n24843), .B(n[359]), .Z(n19005) );
  NAND U26533 ( .A(n21523), .B(n[359]), .Z(n24843) );
  XNOR U26534 ( .A(n24844), .B(n24841), .Z(n19006) );
  XOR U26535 ( .A(n24845), .B(n24846), .Z(n24841) );
  AND U26536 ( .A(n19013), .B(n24847), .Z(n24845) );
  XNOR U26537 ( .A(n19012), .B(n24846), .Z(n24847) );
  NAND U26538 ( .A(n24848), .B(n[358]), .Z(n19012) );
  NAND U26539 ( .A(n21523), .B(n[358]), .Z(n24848) );
  XNOR U26540 ( .A(n24849), .B(n24846), .Z(n19013) );
  XOR U26541 ( .A(n24850), .B(n24851), .Z(n24846) );
  AND U26542 ( .A(n19020), .B(n24852), .Z(n24850) );
  XNOR U26543 ( .A(n19019), .B(n24851), .Z(n24852) );
  NAND U26544 ( .A(n24853), .B(n[357]), .Z(n19019) );
  NAND U26545 ( .A(n21523), .B(n[357]), .Z(n24853) );
  XNOR U26546 ( .A(n24854), .B(n24851), .Z(n19020) );
  XOR U26547 ( .A(n24855), .B(n24856), .Z(n24851) );
  AND U26548 ( .A(n19027), .B(n24857), .Z(n24855) );
  XNOR U26549 ( .A(n19026), .B(n24856), .Z(n24857) );
  NAND U26550 ( .A(n24858), .B(n[356]), .Z(n19026) );
  NAND U26551 ( .A(n21523), .B(n[356]), .Z(n24858) );
  XNOR U26552 ( .A(n24859), .B(n24856), .Z(n19027) );
  XOR U26553 ( .A(n24860), .B(n24861), .Z(n24856) );
  AND U26554 ( .A(n19034), .B(n24862), .Z(n24860) );
  XNOR U26555 ( .A(n19033), .B(n24861), .Z(n24862) );
  NAND U26556 ( .A(n24863), .B(n[355]), .Z(n19033) );
  NAND U26557 ( .A(n21523), .B(n[355]), .Z(n24863) );
  XNOR U26558 ( .A(n24864), .B(n24861), .Z(n19034) );
  XOR U26559 ( .A(n24865), .B(n24866), .Z(n24861) );
  AND U26560 ( .A(n19041), .B(n24867), .Z(n24865) );
  XNOR U26561 ( .A(n19040), .B(n24866), .Z(n24867) );
  NAND U26562 ( .A(n24868), .B(n[354]), .Z(n19040) );
  NAND U26563 ( .A(n21523), .B(n[354]), .Z(n24868) );
  XNOR U26564 ( .A(n24869), .B(n24866), .Z(n19041) );
  XOR U26565 ( .A(n24870), .B(n24871), .Z(n24866) );
  AND U26566 ( .A(n19048), .B(n24872), .Z(n24870) );
  XNOR U26567 ( .A(n19047), .B(n24871), .Z(n24872) );
  NAND U26568 ( .A(n24873), .B(n[353]), .Z(n19047) );
  NAND U26569 ( .A(n21523), .B(n[353]), .Z(n24873) );
  XNOR U26570 ( .A(n24874), .B(n24871), .Z(n19048) );
  XOR U26571 ( .A(n24875), .B(n24876), .Z(n24871) );
  AND U26572 ( .A(n19055), .B(n24877), .Z(n24875) );
  XNOR U26573 ( .A(n19054), .B(n24876), .Z(n24877) );
  NAND U26574 ( .A(n24878), .B(n[352]), .Z(n19054) );
  NAND U26575 ( .A(n21523), .B(n[352]), .Z(n24878) );
  XNOR U26576 ( .A(n24879), .B(n24876), .Z(n19055) );
  XOR U26577 ( .A(n24880), .B(n24881), .Z(n24876) );
  AND U26578 ( .A(n19062), .B(n24882), .Z(n24880) );
  XNOR U26579 ( .A(n19061), .B(n24881), .Z(n24882) );
  NAND U26580 ( .A(n24883), .B(n[351]), .Z(n19061) );
  NAND U26581 ( .A(n21523), .B(n[351]), .Z(n24883) );
  XNOR U26582 ( .A(n24884), .B(n24881), .Z(n19062) );
  XOR U26583 ( .A(n24885), .B(n24886), .Z(n24881) );
  AND U26584 ( .A(n19069), .B(n24887), .Z(n24885) );
  XNOR U26585 ( .A(n19068), .B(n24886), .Z(n24887) );
  NAND U26586 ( .A(n24888), .B(n[350]), .Z(n19068) );
  NAND U26587 ( .A(n21523), .B(n[350]), .Z(n24888) );
  XNOR U26588 ( .A(n24889), .B(n24886), .Z(n19069) );
  XOR U26589 ( .A(n24890), .B(n24891), .Z(n24886) );
  AND U26590 ( .A(n19076), .B(n24892), .Z(n24890) );
  XNOR U26591 ( .A(n19075), .B(n24891), .Z(n24892) );
  NAND U26592 ( .A(n24893), .B(n[349]), .Z(n19075) );
  NAND U26593 ( .A(n21523), .B(n[349]), .Z(n24893) );
  XNOR U26594 ( .A(n24894), .B(n24891), .Z(n19076) );
  XOR U26595 ( .A(n24895), .B(n24896), .Z(n24891) );
  AND U26596 ( .A(n19083), .B(n24897), .Z(n24895) );
  XNOR U26597 ( .A(n19082), .B(n24896), .Z(n24897) );
  NAND U26598 ( .A(n24898), .B(n[348]), .Z(n19082) );
  NAND U26599 ( .A(n21523), .B(n[348]), .Z(n24898) );
  XNOR U26600 ( .A(n24899), .B(n24896), .Z(n19083) );
  XOR U26601 ( .A(n24900), .B(n24901), .Z(n24896) );
  AND U26602 ( .A(n19090), .B(n24902), .Z(n24900) );
  XNOR U26603 ( .A(n19089), .B(n24901), .Z(n24902) );
  NAND U26604 ( .A(n24903), .B(n[347]), .Z(n19089) );
  NAND U26605 ( .A(n21523), .B(n[347]), .Z(n24903) );
  XNOR U26606 ( .A(n24904), .B(n24901), .Z(n19090) );
  XOR U26607 ( .A(n24905), .B(n24906), .Z(n24901) );
  AND U26608 ( .A(n19097), .B(n24907), .Z(n24905) );
  XNOR U26609 ( .A(n19096), .B(n24906), .Z(n24907) );
  NAND U26610 ( .A(n24908), .B(n[346]), .Z(n19096) );
  NAND U26611 ( .A(n21523), .B(n[346]), .Z(n24908) );
  XNOR U26612 ( .A(n24909), .B(n24906), .Z(n19097) );
  XOR U26613 ( .A(n24910), .B(n24911), .Z(n24906) );
  AND U26614 ( .A(n19104), .B(n24912), .Z(n24910) );
  XNOR U26615 ( .A(n19103), .B(n24911), .Z(n24912) );
  NAND U26616 ( .A(n24913), .B(n[345]), .Z(n19103) );
  NAND U26617 ( .A(n21523), .B(n[345]), .Z(n24913) );
  XNOR U26618 ( .A(n24914), .B(n24911), .Z(n19104) );
  XOR U26619 ( .A(n24915), .B(n24916), .Z(n24911) );
  AND U26620 ( .A(n19111), .B(n24917), .Z(n24915) );
  XNOR U26621 ( .A(n19110), .B(n24916), .Z(n24917) );
  NAND U26622 ( .A(n24918), .B(n[344]), .Z(n19110) );
  NAND U26623 ( .A(n21523), .B(n[344]), .Z(n24918) );
  XNOR U26624 ( .A(n24919), .B(n24916), .Z(n19111) );
  XOR U26625 ( .A(n24920), .B(n24921), .Z(n24916) );
  AND U26626 ( .A(n19118), .B(n24922), .Z(n24920) );
  XNOR U26627 ( .A(n19117), .B(n24921), .Z(n24922) );
  NAND U26628 ( .A(n24923), .B(n[343]), .Z(n19117) );
  NAND U26629 ( .A(n21523), .B(n[343]), .Z(n24923) );
  XNOR U26630 ( .A(n24924), .B(n24921), .Z(n19118) );
  XOR U26631 ( .A(n24925), .B(n24926), .Z(n24921) );
  AND U26632 ( .A(n19125), .B(n24927), .Z(n24925) );
  XNOR U26633 ( .A(n19124), .B(n24926), .Z(n24927) );
  NAND U26634 ( .A(n24928), .B(n[342]), .Z(n19124) );
  NAND U26635 ( .A(n21523), .B(n[342]), .Z(n24928) );
  XNOR U26636 ( .A(n24929), .B(n24926), .Z(n19125) );
  XOR U26637 ( .A(n24930), .B(n24931), .Z(n24926) );
  AND U26638 ( .A(n19132), .B(n24932), .Z(n24930) );
  XNOR U26639 ( .A(n19131), .B(n24931), .Z(n24932) );
  NAND U26640 ( .A(n24933), .B(n[341]), .Z(n19131) );
  NAND U26641 ( .A(n21523), .B(n[341]), .Z(n24933) );
  XNOR U26642 ( .A(n24934), .B(n24931), .Z(n19132) );
  XOR U26643 ( .A(n24935), .B(n24936), .Z(n24931) );
  AND U26644 ( .A(n19139), .B(n24937), .Z(n24935) );
  XNOR U26645 ( .A(n19138), .B(n24936), .Z(n24937) );
  NAND U26646 ( .A(n24938), .B(n[340]), .Z(n19138) );
  NAND U26647 ( .A(n21523), .B(n[340]), .Z(n24938) );
  XNOR U26648 ( .A(n24939), .B(n24936), .Z(n19139) );
  XOR U26649 ( .A(n24940), .B(n24941), .Z(n24936) );
  AND U26650 ( .A(n19146), .B(n24942), .Z(n24940) );
  XNOR U26651 ( .A(n19145), .B(n24941), .Z(n24942) );
  NAND U26652 ( .A(n24943), .B(n[339]), .Z(n19145) );
  NAND U26653 ( .A(n21523), .B(n[339]), .Z(n24943) );
  XNOR U26654 ( .A(n24944), .B(n24941), .Z(n19146) );
  XOR U26655 ( .A(n24945), .B(n24946), .Z(n24941) );
  AND U26656 ( .A(n19153), .B(n24947), .Z(n24945) );
  XNOR U26657 ( .A(n19152), .B(n24946), .Z(n24947) );
  NAND U26658 ( .A(n24948), .B(n[338]), .Z(n19152) );
  NAND U26659 ( .A(n21523), .B(n[338]), .Z(n24948) );
  XNOR U26660 ( .A(n24949), .B(n24946), .Z(n19153) );
  XOR U26661 ( .A(n24950), .B(n24951), .Z(n24946) );
  AND U26662 ( .A(n19160), .B(n24952), .Z(n24950) );
  XNOR U26663 ( .A(n19159), .B(n24951), .Z(n24952) );
  NAND U26664 ( .A(n24953), .B(n[337]), .Z(n19159) );
  NAND U26665 ( .A(n21523), .B(n[337]), .Z(n24953) );
  XNOR U26666 ( .A(n24954), .B(n24951), .Z(n19160) );
  XOR U26667 ( .A(n24955), .B(n24956), .Z(n24951) );
  AND U26668 ( .A(n19167), .B(n24957), .Z(n24955) );
  XNOR U26669 ( .A(n19166), .B(n24956), .Z(n24957) );
  NAND U26670 ( .A(n24958), .B(n[336]), .Z(n19166) );
  NAND U26671 ( .A(n21523), .B(n[336]), .Z(n24958) );
  XNOR U26672 ( .A(n24959), .B(n24956), .Z(n19167) );
  XOR U26673 ( .A(n24960), .B(n24961), .Z(n24956) );
  AND U26674 ( .A(n19174), .B(n24962), .Z(n24960) );
  XNOR U26675 ( .A(n19173), .B(n24961), .Z(n24962) );
  NAND U26676 ( .A(n24963), .B(n[335]), .Z(n19173) );
  NAND U26677 ( .A(n21523), .B(n[335]), .Z(n24963) );
  XNOR U26678 ( .A(n24964), .B(n24961), .Z(n19174) );
  XOR U26679 ( .A(n24965), .B(n24966), .Z(n24961) );
  AND U26680 ( .A(n19181), .B(n24967), .Z(n24965) );
  XNOR U26681 ( .A(n19180), .B(n24966), .Z(n24967) );
  NAND U26682 ( .A(n24968), .B(n[334]), .Z(n19180) );
  NAND U26683 ( .A(n21523), .B(n[334]), .Z(n24968) );
  XNOR U26684 ( .A(n24969), .B(n24966), .Z(n19181) );
  XOR U26685 ( .A(n24970), .B(n24971), .Z(n24966) );
  AND U26686 ( .A(n19188), .B(n24972), .Z(n24970) );
  XNOR U26687 ( .A(n19187), .B(n24971), .Z(n24972) );
  NAND U26688 ( .A(n24973), .B(n[333]), .Z(n19187) );
  NAND U26689 ( .A(n21523), .B(n[333]), .Z(n24973) );
  XNOR U26690 ( .A(n24974), .B(n24971), .Z(n19188) );
  XOR U26691 ( .A(n24975), .B(n24976), .Z(n24971) );
  AND U26692 ( .A(n19195), .B(n24977), .Z(n24975) );
  XNOR U26693 ( .A(n19194), .B(n24976), .Z(n24977) );
  NAND U26694 ( .A(n24978), .B(n[332]), .Z(n19194) );
  NAND U26695 ( .A(n21523), .B(n[332]), .Z(n24978) );
  XNOR U26696 ( .A(n24979), .B(n24976), .Z(n19195) );
  XOR U26697 ( .A(n24980), .B(n24981), .Z(n24976) );
  AND U26698 ( .A(n19202), .B(n24982), .Z(n24980) );
  XNOR U26699 ( .A(n19201), .B(n24981), .Z(n24982) );
  NAND U26700 ( .A(n24983), .B(n[331]), .Z(n19201) );
  NAND U26701 ( .A(n21523), .B(n[331]), .Z(n24983) );
  XNOR U26702 ( .A(n24984), .B(n24981), .Z(n19202) );
  XOR U26703 ( .A(n24985), .B(n24986), .Z(n24981) );
  AND U26704 ( .A(n19209), .B(n24987), .Z(n24985) );
  XNOR U26705 ( .A(n19208), .B(n24986), .Z(n24987) );
  NAND U26706 ( .A(n24988), .B(n[330]), .Z(n19208) );
  NAND U26707 ( .A(n21523), .B(n[330]), .Z(n24988) );
  XNOR U26708 ( .A(n24989), .B(n24986), .Z(n19209) );
  XOR U26709 ( .A(n24990), .B(n24991), .Z(n24986) );
  AND U26710 ( .A(n19216), .B(n24992), .Z(n24990) );
  XNOR U26711 ( .A(n19215), .B(n24991), .Z(n24992) );
  NAND U26712 ( .A(n24993), .B(n[329]), .Z(n19215) );
  NAND U26713 ( .A(n21523), .B(n[329]), .Z(n24993) );
  XNOR U26714 ( .A(n24994), .B(n24991), .Z(n19216) );
  XOR U26715 ( .A(n24995), .B(n24996), .Z(n24991) );
  AND U26716 ( .A(n19223), .B(n24997), .Z(n24995) );
  XNOR U26717 ( .A(n19222), .B(n24996), .Z(n24997) );
  NAND U26718 ( .A(n24998), .B(n[328]), .Z(n19222) );
  NAND U26719 ( .A(n21523), .B(n[328]), .Z(n24998) );
  XNOR U26720 ( .A(n24999), .B(n24996), .Z(n19223) );
  XOR U26721 ( .A(n25000), .B(n25001), .Z(n24996) );
  AND U26722 ( .A(n19230), .B(n25002), .Z(n25000) );
  XNOR U26723 ( .A(n19229), .B(n25001), .Z(n25002) );
  NAND U26724 ( .A(n25003), .B(n[327]), .Z(n19229) );
  NAND U26725 ( .A(n21523), .B(n[327]), .Z(n25003) );
  XNOR U26726 ( .A(n25004), .B(n25001), .Z(n19230) );
  XOR U26727 ( .A(n25005), .B(n25006), .Z(n25001) );
  AND U26728 ( .A(n19237), .B(n25007), .Z(n25005) );
  XNOR U26729 ( .A(n19236), .B(n25006), .Z(n25007) );
  NAND U26730 ( .A(n25008), .B(n[326]), .Z(n19236) );
  NAND U26731 ( .A(n21523), .B(n[326]), .Z(n25008) );
  XNOR U26732 ( .A(n25009), .B(n25006), .Z(n19237) );
  XOR U26733 ( .A(n25010), .B(n25011), .Z(n25006) );
  AND U26734 ( .A(n19244), .B(n25012), .Z(n25010) );
  XNOR U26735 ( .A(n19243), .B(n25011), .Z(n25012) );
  NAND U26736 ( .A(n25013), .B(n[325]), .Z(n19243) );
  NAND U26737 ( .A(n21523), .B(n[325]), .Z(n25013) );
  XNOR U26738 ( .A(n25014), .B(n25011), .Z(n19244) );
  XOR U26739 ( .A(n25015), .B(n25016), .Z(n25011) );
  AND U26740 ( .A(n19251), .B(n25017), .Z(n25015) );
  XNOR U26741 ( .A(n19250), .B(n25016), .Z(n25017) );
  NAND U26742 ( .A(n25018), .B(n[324]), .Z(n19250) );
  NAND U26743 ( .A(n21523), .B(n[324]), .Z(n25018) );
  XNOR U26744 ( .A(n25019), .B(n25016), .Z(n19251) );
  XOR U26745 ( .A(n25020), .B(n25021), .Z(n25016) );
  AND U26746 ( .A(n19258), .B(n25022), .Z(n25020) );
  XNOR U26747 ( .A(n19257), .B(n25021), .Z(n25022) );
  NAND U26748 ( .A(n25023), .B(n[323]), .Z(n19257) );
  NAND U26749 ( .A(n21523), .B(n[323]), .Z(n25023) );
  XNOR U26750 ( .A(n25024), .B(n25021), .Z(n19258) );
  XOR U26751 ( .A(n25025), .B(n25026), .Z(n25021) );
  AND U26752 ( .A(n19265), .B(n25027), .Z(n25025) );
  XNOR U26753 ( .A(n19264), .B(n25026), .Z(n25027) );
  NAND U26754 ( .A(n25028), .B(n[322]), .Z(n19264) );
  NAND U26755 ( .A(n21523), .B(n[322]), .Z(n25028) );
  XNOR U26756 ( .A(n25029), .B(n25026), .Z(n19265) );
  XOR U26757 ( .A(n25030), .B(n25031), .Z(n25026) );
  AND U26758 ( .A(n19272), .B(n25032), .Z(n25030) );
  XNOR U26759 ( .A(n19271), .B(n25031), .Z(n25032) );
  NAND U26760 ( .A(n25033), .B(n[321]), .Z(n19271) );
  NAND U26761 ( .A(n21523), .B(n[321]), .Z(n25033) );
  XNOR U26762 ( .A(n25034), .B(n25031), .Z(n19272) );
  XOR U26763 ( .A(n25035), .B(n25036), .Z(n25031) );
  AND U26764 ( .A(n19279), .B(n25037), .Z(n25035) );
  XNOR U26765 ( .A(n19278), .B(n25036), .Z(n25037) );
  NAND U26766 ( .A(n25038), .B(n[320]), .Z(n19278) );
  NAND U26767 ( .A(n21523), .B(n[320]), .Z(n25038) );
  XNOR U26768 ( .A(n25039), .B(n25036), .Z(n19279) );
  XOR U26769 ( .A(n25040), .B(n25041), .Z(n25036) );
  AND U26770 ( .A(n19286), .B(n25042), .Z(n25040) );
  XNOR U26771 ( .A(n19285), .B(n25041), .Z(n25042) );
  NAND U26772 ( .A(n25043), .B(n[319]), .Z(n19285) );
  NAND U26773 ( .A(n21523), .B(n[319]), .Z(n25043) );
  XNOR U26774 ( .A(n25044), .B(n25041), .Z(n19286) );
  XOR U26775 ( .A(n25045), .B(n25046), .Z(n25041) );
  AND U26776 ( .A(n19293), .B(n25047), .Z(n25045) );
  XNOR U26777 ( .A(n19292), .B(n25046), .Z(n25047) );
  NAND U26778 ( .A(n25048), .B(n[318]), .Z(n19292) );
  NAND U26779 ( .A(n21523), .B(n[318]), .Z(n25048) );
  XNOR U26780 ( .A(n25049), .B(n25046), .Z(n19293) );
  XOR U26781 ( .A(n25050), .B(n25051), .Z(n25046) );
  AND U26782 ( .A(n19300), .B(n25052), .Z(n25050) );
  XNOR U26783 ( .A(n19299), .B(n25051), .Z(n25052) );
  NAND U26784 ( .A(n25053), .B(n[317]), .Z(n19299) );
  NAND U26785 ( .A(n21523), .B(n[317]), .Z(n25053) );
  XNOR U26786 ( .A(n25054), .B(n25051), .Z(n19300) );
  XOR U26787 ( .A(n25055), .B(n25056), .Z(n25051) );
  AND U26788 ( .A(n19307), .B(n25057), .Z(n25055) );
  XNOR U26789 ( .A(n19306), .B(n25056), .Z(n25057) );
  NAND U26790 ( .A(n25058), .B(n[316]), .Z(n19306) );
  NAND U26791 ( .A(n21523), .B(n[316]), .Z(n25058) );
  XNOR U26792 ( .A(n25059), .B(n25056), .Z(n19307) );
  XOR U26793 ( .A(n25060), .B(n25061), .Z(n25056) );
  AND U26794 ( .A(n19314), .B(n25062), .Z(n25060) );
  XNOR U26795 ( .A(n19313), .B(n25061), .Z(n25062) );
  NAND U26796 ( .A(n25063), .B(n[315]), .Z(n19313) );
  NAND U26797 ( .A(n21523), .B(n[315]), .Z(n25063) );
  XNOR U26798 ( .A(n25064), .B(n25061), .Z(n19314) );
  XOR U26799 ( .A(n25065), .B(n25066), .Z(n25061) );
  AND U26800 ( .A(n19321), .B(n25067), .Z(n25065) );
  XNOR U26801 ( .A(n19320), .B(n25066), .Z(n25067) );
  NAND U26802 ( .A(n25068), .B(n[314]), .Z(n19320) );
  NAND U26803 ( .A(n21523), .B(n[314]), .Z(n25068) );
  XNOR U26804 ( .A(n25069), .B(n25066), .Z(n19321) );
  XOR U26805 ( .A(n25070), .B(n25071), .Z(n25066) );
  AND U26806 ( .A(n19328), .B(n25072), .Z(n25070) );
  XNOR U26807 ( .A(n19327), .B(n25071), .Z(n25072) );
  NAND U26808 ( .A(n25073), .B(n[313]), .Z(n19327) );
  NAND U26809 ( .A(n21523), .B(n[313]), .Z(n25073) );
  XNOR U26810 ( .A(n25074), .B(n25071), .Z(n19328) );
  XOR U26811 ( .A(n25075), .B(n25076), .Z(n25071) );
  AND U26812 ( .A(n19335), .B(n25077), .Z(n25075) );
  XNOR U26813 ( .A(n19334), .B(n25076), .Z(n25077) );
  NAND U26814 ( .A(n25078), .B(n[312]), .Z(n19334) );
  NAND U26815 ( .A(n21523), .B(n[312]), .Z(n25078) );
  XNOR U26816 ( .A(n25079), .B(n25076), .Z(n19335) );
  XOR U26817 ( .A(n25080), .B(n25081), .Z(n25076) );
  AND U26818 ( .A(n19342), .B(n25082), .Z(n25080) );
  XNOR U26819 ( .A(n19341), .B(n25081), .Z(n25082) );
  NAND U26820 ( .A(n25083), .B(n[311]), .Z(n19341) );
  NAND U26821 ( .A(n21523), .B(n[311]), .Z(n25083) );
  XNOR U26822 ( .A(n25084), .B(n25081), .Z(n19342) );
  XOR U26823 ( .A(n25085), .B(n25086), .Z(n25081) );
  AND U26824 ( .A(n19349), .B(n25087), .Z(n25085) );
  XNOR U26825 ( .A(n19348), .B(n25086), .Z(n25087) );
  NAND U26826 ( .A(n25088), .B(n[310]), .Z(n19348) );
  NAND U26827 ( .A(n21523), .B(n[310]), .Z(n25088) );
  XNOR U26828 ( .A(n25089), .B(n25086), .Z(n19349) );
  XOR U26829 ( .A(n25090), .B(n25091), .Z(n25086) );
  AND U26830 ( .A(n19356), .B(n25092), .Z(n25090) );
  XNOR U26831 ( .A(n19355), .B(n25091), .Z(n25092) );
  NAND U26832 ( .A(n25093), .B(n[309]), .Z(n19355) );
  NAND U26833 ( .A(n21523), .B(n[309]), .Z(n25093) );
  XNOR U26834 ( .A(n25094), .B(n25091), .Z(n19356) );
  XOR U26835 ( .A(n25095), .B(n25096), .Z(n25091) );
  AND U26836 ( .A(n19363), .B(n25097), .Z(n25095) );
  XNOR U26837 ( .A(n19362), .B(n25096), .Z(n25097) );
  NAND U26838 ( .A(n25098), .B(n[308]), .Z(n19362) );
  NAND U26839 ( .A(n21523), .B(n[308]), .Z(n25098) );
  XNOR U26840 ( .A(n25099), .B(n25096), .Z(n19363) );
  XOR U26841 ( .A(n25100), .B(n25101), .Z(n25096) );
  AND U26842 ( .A(n19370), .B(n25102), .Z(n25100) );
  XNOR U26843 ( .A(n19369), .B(n25101), .Z(n25102) );
  NAND U26844 ( .A(n25103), .B(n[307]), .Z(n19369) );
  NAND U26845 ( .A(n21523), .B(n[307]), .Z(n25103) );
  XNOR U26846 ( .A(n25104), .B(n25101), .Z(n19370) );
  XOR U26847 ( .A(n25105), .B(n25106), .Z(n25101) );
  AND U26848 ( .A(n19377), .B(n25107), .Z(n25105) );
  XNOR U26849 ( .A(n19376), .B(n25106), .Z(n25107) );
  NAND U26850 ( .A(n25108), .B(n[306]), .Z(n19376) );
  NAND U26851 ( .A(n21523), .B(n[306]), .Z(n25108) );
  XNOR U26852 ( .A(n25109), .B(n25106), .Z(n19377) );
  XOR U26853 ( .A(n25110), .B(n25111), .Z(n25106) );
  AND U26854 ( .A(n19384), .B(n25112), .Z(n25110) );
  XNOR U26855 ( .A(n19383), .B(n25111), .Z(n25112) );
  NAND U26856 ( .A(n25113), .B(n[305]), .Z(n19383) );
  NAND U26857 ( .A(n21523), .B(n[305]), .Z(n25113) );
  XNOR U26858 ( .A(n25114), .B(n25111), .Z(n19384) );
  XOR U26859 ( .A(n25115), .B(n25116), .Z(n25111) );
  AND U26860 ( .A(n19391), .B(n25117), .Z(n25115) );
  XNOR U26861 ( .A(n19390), .B(n25116), .Z(n25117) );
  NAND U26862 ( .A(n25118), .B(n[304]), .Z(n19390) );
  NAND U26863 ( .A(n21523), .B(n[304]), .Z(n25118) );
  XNOR U26864 ( .A(n25119), .B(n25116), .Z(n19391) );
  XOR U26865 ( .A(n25120), .B(n25121), .Z(n25116) );
  AND U26866 ( .A(n19398), .B(n25122), .Z(n25120) );
  XNOR U26867 ( .A(n19397), .B(n25121), .Z(n25122) );
  NAND U26868 ( .A(n25123), .B(n[303]), .Z(n19397) );
  NAND U26869 ( .A(n21523), .B(n[303]), .Z(n25123) );
  XNOR U26870 ( .A(n25124), .B(n25121), .Z(n19398) );
  XOR U26871 ( .A(n25125), .B(n25126), .Z(n25121) );
  AND U26872 ( .A(n19405), .B(n25127), .Z(n25125) );
  XNOR U26873 ( .A(n19404), .B(n25126), .Z(n25127) );
  NAND U26874 ( .A(n25128), .B(n[302]), .Z(n19404) );
  NAND U26875 ( .A(n21523), .B(n[302]), .Z(n25128) );
  XNOR U26876 ( .A(n25129), .B(n25126), .Z(n19405) );
  XOR U26877 ( .A(n25130), .B(n25131), .Z(n25126) );
  AND U26878 ( .A(n19412), .B(n25132), .Z(n25130) );
  XNOR U26879 ( .A(n19411), .B(n25131), .Z(n25132) );
  NAND U26880 ( .A(n25133), .B(n[301]), .Z(n19411) );
  NAND U26881 ( .A(n21523), .B(n[301]), .Z(n25133) );
  XNOR U26882 ( .A(n25134), .B(n25131), .Z(n19412) );
  XOR U26883 ( .A(n25135), .B(n25136), .Z(n25131) );
  AND U26884 ( .A(n19419), .B(n25137), .Z(n25135) );
  XNOR U26885 ( .A(n19418), .B(n25136), .Z(n25137) );
  NAND U26886 ( .A(n25138), .B(n[300]), .Z(n19418) );
  NAND U26887 ( .A(n21523), .B(n[300]), .Z(n25138) );
  XNOR U26888 ( .A(n25139), .B(n25136), .Z(n19419) );
  XOR U26889 ( .A(n25140), .B(n25141), .Z(n25136) );
  AND U26890 ( .A(n19426), .B(n25142), .Z(n25140) );
  XNOR U26891 ( .A(n19425), .B(n25141), .Z(n25142) );
  NAND U26892 ( .A(n25143), .B(n[299]), .Z(n19425) );
  NAND U26893 ( .A(n21523), .B(n[299]), .Z(n25143) );
  XNOR U26894 ( .A(n25144), .B(n25141), .Z(n19426) );
  XOR U26895 ( .A(n25145), .B(n25146), .Z(n25141) );
  AND U26896 ( .A(n19433), .B(n25147), .Z(n25145) );
  XNOR U26897 ( .A(n19432), .B(n25146), .Z(n25147) );
  NAND U26898 ( .A(n25148), .B(n[298]), .Z(n19432) );
  NAND U26899 ( .A(n21523), .B(n[298]), .Z(n25148) );
  XNOR U26900 ( .A(n25149), .B(n25146), .Z(n19433) );
  XOR U26901 ( .A(n25150), .B(n25151), .Z(n25146) );
  AND U26902 ( .A(n19440), .B(n25152), .Z(n25150) );
  XNOR U26903 ( .A(n19439), .B(n25151), .Z(n25152) );
  NAND U26904 ( .A(n25153), .B(n[297]), .Z(n19439) );
  NAND U26905 ( .A(n21523), .B(n[297]), .Z(n25153) );
  XNOR U26906 ( .A(n25154), .B(n25151), .Z(n19440) );
  XOR U26907 ( .A(n25155), .B(n25156), .Z(n25151) );
  AND U26908 ( .A(n19447), .B(n25157), .Z(n25155) );
  XNOR U26909 ( .A(n19446), .B(n25156), .Z(n25157) );
  NAND U26910 ( .A(n25158), .B(n[296]), .Z(n19446) );
  NAND U26911 ( .A(n21523), .B(n[296]), .Z(n25158) );
  XNOR U26912 ( .A(n25159), .B(n25156), .Z(n19447) );
  XOR U26913 ( .A(n25160), .B(n25161), .Z(n25156) );
  AND U26914 ( .A(n19454), .B(n25162), .Z(n25160) );
  XNOR U26915 ( .A(n19453), .B(n25161), .Z(n25162) );
  NAND U26916 ( .A(n25163), .B(n[295]), .Z(n19453) );
  NAND U26917 ( .A(n21523), .B(n[295]), .Z(n25163) );
  XNOR U26918 ( .A(n25164), .B(n25161), .Z(n19454) );
  XOR U26919 ( .A(n25165), .B(n25166), .Z(n25161) );
  AND U26920 ( .A(n19461), .B(n25167), .Z(n25165) );
  XNOR U26921 ( .A(n19460), .B(n25166), .Z(n25167) );
  NAND U26922 ( .A(n25168), .B(n[294]), .Z(n19460) );
  NAND U26923 ( .A(n21523), .B(n[294]), .Z(n25168) );
  XNOR U26924 ( .A(n25169), .B(n25166), .Z(n19461) );
  XOR U26925 ( .A(n25170), .B(n25171), .Z(n25166) );
  AND U26926 ( .A(n19468), .B(n25172), .Z(n25170) );
  XNOR U26927 ( .A(n19467), .B(n25171), .Z(n25172) );
  NAND U26928 ( .A(n25173), .B(n[293]), .Z(n19467) );
  NAND U26929 ( .A(n21523), .B(n[293]), .Z(n25173) );
  XNOR U26930 ( .A(n25174), .B(n25171), .Z(n19468) );
  XOR U26931 ( .A(n25175), .B(n25176), .Z(n25171) );
  AND U26932 ( .A(n19475), .B(n25177), .Z(n25175) );
  XNOR U26933 ( .A(n19474), .B(n25176), .Z(n25177) );
  NAND U26934 ( .A(n25178), .B(n[292]), .Z(n19474) );
  NAND U26935 ( .A(n21523), .B(n[292]), .Z(n25178) );
  XNOR U26936 ( .A(n25179), .B(n25176), .Z(n19475) );
  XOR U26937 ( .A(n25180), .B(n25181), .Z(n25176) );
  AND U26938 ( .A(n19482), .B(n25182), .Z(n25180) );
  XNOR U26939 ( .A(n19481), .B(n25181), .Z(n25182) );
  NAND U26940 ( .A(n25183), .B(n[291]), .Z(n19481) );
  NAND U26941 ( .A(n21523), .B(n[291]), .Z(n25183) );
  XNOR U26942 ( .A(n25184), .B(n25181), .Z(n19482) );
  XOR U26943 ( .A(n25185), .B(n25186), .Z(n25181) );
  AND U26944 ( .A(n19489), .B(n25187), .Z(n25185) );
  XNOR U26945 ( .A(n19488), .B(n25186), .Z(n25187) );
  NAND U26946 ( .A(n25188), .B(n[290]), .Z(n19488) );
  NAND U26947 ( .A(n21523), .B(n[290]), .Z(n25188) );
  XNOR U26948 ( .A(n25189), .B(n25186), .Z(n19489) );
  XOR U26949 ( .A(n25190), .B(n25191), .Z(n25186) );
  AND U26950 ( .A(n19496), .B(n25192), .Z(n25190) );
  XNOR U26951 ( .A(n19495), .B(n25191), .Z(n25192) );
  NAND U26952 ( .A(n25193), .B(n[289]), .Z(n19495) );
  NAND U26953 ( .A(n21523), .B(n[289]), .Z(n25193) );
  XNOR U26954 ( .A(n25194), .B(n25191), .Z(n19496) );
  XOR U26955 ( .A(n25195), .B(n25196), .Z(n25191) );
  AND U26956 ( .A(n19503), .B(n25197), .Z(n25195) );
  XNOR U26957 ( .A(n19502), .B(n25196), .Z(n25197) );
  NAND U26958 ( .A(n25198), .B(n[288]), .Z(n19502) );
  NAND U26959 ( .A(n21523), .B(n[288]), .Z(n25198) );
  XNOR U26960 ( .A(n25199), .B(n25196), .Z(n19503) );
  XOR U26961 ( .A(n25200), .B(n25201), .Z(n25196) );
  AND U26962 ( .A(n19510), .B(n25202), .Z(n25200) );
  XNOR U26963 ( .A(n19509), .B(n25201), .Z(n25202) );
  NAND U26964 ( .A(n25203), .B(n[287]), .Z(n19509) );
  NAND U26965 ( .A(n21523), .B(n[287]), .Z(n25203) );
  XNOR U26966 ( .A(n25204), .B(n25201), .Z(n19510) );
  XOR U26967 ( .A(n25205), .B(n25206), .Z(n25201) );
  AND U26968 ( .A(n19517), .B(n25207), .Z(n25205) );
  XNOR U26969 ( .A(n19516), .B(n25206), .Z(n25207) );
  NAND U26970 ( .A(n25208), .B(n[286]), .Z(n19516) );
  NAND U26971 ( .A(n21523), .B(n[286]), .Z(n25208) );
  XNOR U26972 ( .A(n25209), .B(n25206), .Z(n19517) );
  XOR U26973 ( .A(n25210), .B(n25211), .Z(n25206) );
  AND U26974 ( .A(n19524), .B(n25212), .Z(n25210) );
  XNOR U26975 ( .A(n19523), .B(n25211), .Z(n25212) );
  NAND U26976 ( .A(n25213), .B(n[285]), .Z(n19523) );
  NAND U26977 ( .A(n21523), .B(n[285]), .Z(n25213) );
  XNOR U26978 ( .A(n25214), .B(n25211), .Z(n19524) );
  XOR U26979 ( .A(n25215), .B(n25216), .Z(n25211) );
  AND U26980 ( .A(n19531), .B(n25217), .Z(n25215) );
  XNOR U26981 ( .A(n19530), .B(n25216), .Z(n25217) );
  NAND U26982 ( .A(n25218), .B(n[284]), .Z(n19530) );
  NAND U26983 ( .A(n21523), .B(n[284]), .Z(n25218) );
  XNOR U26984 ( .A(n25219), .B(n25216), .Z(n19531) );
  XOR U26985 ( .A(n25220), .B(n25221), .Z(n25216) );
  AND U26986 ( .A(n19538), .B(n25222), .Z(n25220) );
  XNOR U26987 ( .A(n19537), .B(n25221), .Z(n25222) );
  NAND U26988 ( .A(n25223), .B(n[283]), .Z(n19537) );
  NAND U26989 ( .A(n21523), .B(n[283]), .Z(n25223) );
  XNOR U26990 ( .A(n25224), .B(n25221), .Z(n19538) );
  XOR U26991 ( .A(n25225), .B(n25226), .Z(n25221) );
  AND U26992 ( .A(n19545), .B(n25227), .Z(n25225) );
  XNOR U26993 ( .A(n19544), .B(n25226), .Z(n25227) );
  NAND U26994 ( .A(n25228), .B(n[282]), .Z(n19544) );
  NAND U26995 ( .A(n21523), .B(n[282]), .Z(n25228) );
  XNOR U26996 ( .A(n25229), .B(n25226), .Z(n19545) );
  XOR U26997 ( .A(n25230), .B(n25231), .Z(n25226) );
  AND U26998 ( .A(n19552), .B(n25232), .Z(n25230) );
  XNOR U26999 ( .A(n19551), .B(n25231), .Z(n25232) );
  NAND U27000 ( .A(n25233), .B(n[281]), .Z(n19551) );
  NAND U27001 ( .A(n21523), .B(n[281]), .Z(n25233) );
  XNOR U27002 ( .A(n25234), .B(n25231), .Z(n19552) );
  XOR U27003 ( .A(n25235), .B(n25236), .Z(n25231) );
  AND U27004 ( .A(n19559), .B(n25237), .Z(n25235) );
  XNOR U27005 ( .A(n19558), .B(n25236), .Z(n25237) );
  NAND U27006 ( .A(n25238), .B(n[280]), .Z(n19558) );
  NAND U27007 ( .A(n21523), .B(n[280]), .Z(n25238) );
  XNOR U27008 ( .A(n25239), .B(n25236), .Z(n19559) );
  XOR U27009 ( .A(n25240), .B(n25241), .Z(n25236) );
  AND U27010 ( .A(n19566), .B(n25242), .Z(n25240) );
  XNOR U27011 ( .A(n19565), .B(n25241), .Z(n25242) );
  NAND U27012 ( .A(n25243), .B(n[279]), .Z(n19565) );
  NAND U27013 ( .A(n21523), .B(n[279]), .Z(n25243) );
  XNOR U27014 ( .A(n25244), .B(n25241), .Z(n19566) );
  XOR U27015 ( .A(n25245), .B(n25246), .Z(n25241) );
  AND U27016 ( .A(n19573), .B(n25247), .Z(n25245) );
  XNOR U27017 ( .A(n19572), .B(n25246), .Z(n25247) );
  NAND U27018 ( .A(n25248), .B(n[278]), .Z(n19572) );
  NAND U27019 ( .A(n21523), .B(n[278]), .Z(n25248) );
  XNOR U27020 ( .A(n25249), .B(n25246), .Z(n19573) );
  XOR U27021 ( .A(n25250), .B(n25251), .Z(n25246) );
  AND U27022 ( .A(n19580), .B(n25252), .Z(n25250) );
  XNOR U27023 ( .A(n19579), .B(n25251), .Z(n25252) );
  NAND U27024 ( .A(n25253), .B(n[277]), .Z(n19579) );
  NAND U27025 ( .A(n21523), .B(n[277]), .Z(n25253) );
  XNOR U27026 ( .A(n25254), .B(n25251), .Z(n19580) );
  XOR U27027 ( .A(n25255), .B(n25256), .Z(n25251) );
  AND U27028 ( .A(n19587), .B(n25257), .Z(n25255) );
  XNOR U27029 ( .A(n19586), .B(n25256), .Z(n25257) );
  NAND U27030 ( .A(n25258), .B(n[276]), .Z(n19586) );
  NAND U27031 ( .A(n21523), .B(n[276]), .Z(n25258) );
  XNOR U27032 ( .A(n25259), .B(n25256), .Z(n19587) );
  XOR U27033 ( .A(n25260), .B(n25261), .Z(n25256) );
  AND U27034 ( .A(n19594), .B(n25262), .Z(n25260) );
  XNOR U27035 ( .A(n19593), .B(n25261), .Z(n25262) );
  NAND U27036 ( .A(n25263), .B(n[275]), .Z(n19593) );
  NAND U27037 ( .A(n21523), .B(n[275]), .Z(n25263) );
  XNOR U27038 ( .A(n25264), .B(n25261), .Z(n19594) );
  XOR U27039 ( .A(n25265), .B(n25266), .Z(n25261) );
  AND U27040 ( .A(n19601), .B(n25267), .Z(n25265) );
  XNOR U27041 ( .A(n19600), .B(n25266), .Z(n25267) );
  NAND U27042 ( .A(n25268), .B(n[274]), .Z(n19600) );
  NAND U27043 ( .A(n21523), .B(n[274]), .Z(n25268) );
  XNOR U27044 ( .A(n25269), .B(n25266), .Z(n19601) );
  XOR U27045 ( .A(n25270), .B(n25271), .Z(n25266) );
  AND U27046 ( .A(n19608), .B(n25272), .Z(n25270) );
  XNOR U27047 ( .A(n19607), .B(n25271), .Z(n25272) );
  NAND U27048 ( .A(n25273), .B(n[273]), .Z(n19607) );
  NAND U27049 ( .A(n21523), .B(n[273]), .Z(n25273) );
  XNOR U27050 ( .A(n25274), .B(n25271), .Z(n19608) );
  XOR U27051 ( .A(n25275), .B(n25276), .Z(n25271) );
  AND U27052 ( .A(n19615), .B(n25277), .Z(n25275) );
  XNOR U27053 ( .A(n19614), .B(n25276), .Z(n25277) );
  NAND U27054 ( .A(n25278), .B(n[272]), .Z(n19614) );
  NAND U27055 ( .A(n21523), .B(n[272]), .Z(n25278) );
  XNOR U27056 ( .A(n25279), .B(n25276), .Z(n19615) );
  XOR U27057 ( .A(n25280), .B(n25281), .Z(n25276) );
  AND U27058 ( .A(n19622), .B(n25282), .Z(n25280) );
  XNOR U27059 ( .A(n19621), .B(n25281), .Z(n25282) );
  NAND U27060 ( .A(n25283), .B(n[271]), .Z(n19621) );
  NAND U27061 ( .A(n21523), .B(n[271]), .Z(n25283) );
  XNOR U27062 ( .A(n25284), .B(n25281), .Z(n19622) );
  XOR U27063 ( .A(n25285), .B(n25286), .Z(n25281) );
  AND U27064 ( .A(n19629), .B(n25287), .Z(n25285) );
  XNOR U27065 ( .A(n19628), .B(n25286), .Z(n25287) );
  NAND U27066 ( .A(n25288), .B(n[270]), .Z(n19628) );
  NAND U27067 ( .A(n21523), .B(n[270]), .Z(n25288) );
  XNOR U27068 ( .A(n25289), .B(n25286), .Z(n19629) );
  XOR U27069 ( .A(n25290), .B(n25291), .Z(n25286) );
  AND U27070 ( .A(n19636), .B(n25292), .Z(n25290) );
  XNOR U27071 ( .A(n19635), .B(n25291), .Z(n25292) );
  NAND U27072 ( .A(n25293), .B(n[269]), .Z(n19635) );
  NAND U27073 ( .A(n21523), .B(n[269]), .Z(n25293) );
  XNOR U27074 ( .A(n25294), .B(n25291), .Z(n19636) );
  XOR U27075 ( .A(n25295), .B(n25296), .Z(n25291) );
  AND U27076 ( .A(n19643), .B(n25297), .Z(n25295) );
  XNOR U27077 ( .A(n19642), .B(n25296), .Z(n25297) );
  NAND U27078 ( .A(n25298), .B(n[268]), .Z(n19642) );
  NAND U27079 ( .A(n21523), .B(n[268]), .Z(n25298) );
  XNOR U27080 ( .A(n25299), .B(n25296), .Z(n19643) );
  XOR U27081 ( .A(n25300), .B(n25301), .Z(n25296) );
  AND U27082 ( .A(n19650), .B(n25302), .Z(n25300) );
  XNOR U27083 ( .A(n19649), .B(n25301), .Z(n25302) );
  NAND U27084 ( .A(n25303), .B(n[267]), .Z(n19649) );
  NAND U27085 ( .A(n21523), .B(n[267]), .Z(n25303) );
  XNOR U27086 ( .A(n25304), .B(n25301), .Z(n19650) );
  XOR U27087 ( .A(n25305), .B(n25306), .Z(n25301) );
  AND U27088 ( .A(n19657), .B(n25307), .Z(n25305) );
  XNOR U27089 ( .A(n19656), .B(n25306), .Z(n25307) );
  NAND U27090 ( .A(n25308), .B(n[266]), .Z(n19656) );
  NAND U27091 ( .A(n21523), .B(n[266]), .Z(n25308) );
  XNOR U27092 ( .A(n25309), .B(n25306), .Z(n19657) );
  XOR U27093 ( .A(n25310), .B(n25311), .Z(n25306) );
  AND U27094 ( .A(n19664), .B(n25312), .Z(n25310) );
  XNOR U27095 ( .A(n19663), .B(n25311), .Z(n25312) );
  NAND U27096 ( .A(n25313), .B(n[265]), .Z(n19663) );
  NAND U27097 ( .A(n21523), .B(n[265]), .Z(n25313) );
  XNOR U27098 ( .A(n25314), .B(n25311), .Z(n19664) );
  XOR U27099 ( .A(n25315), .B(n25316), .Z(n25311) );
  AND U27100 ( .A(n19671), .B(n25317), .Z(n25315) );
  XNOR U27101 ( .A(n19670), .B(n25316), .Z(n25317) );
  NAND U27102 ( .A(n25318), .B(n[264]), .Z(n19670) );
  NAND U27103 ( .A(n21523), .B(n[264]), .Z(n25318) );
  XNOR U27104 ( .A(n25319), .B(n25316), .Z(n19671) );
  XOR U27105 ( .A(n25320), .B(n25321), .Z(n25316) );
  AND U27106 ( .A(n19678), .B(n25322), .Z(n25320) );
  XNOR U27107 ( .A(n19677), .B(n25321), .Z(n25322) );
  NAND U27108 ( .A(n25323), .B(n[263]), .Z(n19677) );
  NAND U27109 ( .A(n21523), .B(n[263]), .Z(n25323) );
  XNOR U27110 ( .A(n25324), .B(n25321), .Z(n19678) );
  XOR U27111 ( .A(n25325), .B(n25326), .Z(n25321) );
  AND U27112 ( .A(n19685), .B(n25327), .Z(n25325) );
  XNOR U27113 ( .A(n19684), .B(n25326), .Z(n25327) );
  NAND U27114 ( .A(n25328), .B(n[262]), .Z(n19684) );
  NAND U27115 ( .A(n21523), .B(n[262]), .Z(n25328) );
  XNOR U27116 ( .A(n25329), .B(n25326), .Z(n19685) );
  XOR U27117 ( .A(n25330), .B(n25331), .Z(n25326) );
  AND U27118 ( .A(n19692), .B(n25332), .Z(n25330) );
  XNOR U27119 ( .A(n19691), .B(n25331), .Z(n25332) );
  NAND U27120 ( .A(n25333), .B(n[261]), .Z(n19691) );
  NAND U27121 ( .A(n21523), .B(n[261]), .Z(n25333) );
  XNOR U27122 ( .A(n25334), .B(n25331), .Z(n19692) );
  XOR U27123 ( .A(n25335), .B(n25336), .Z(n25331) );
  AND U27124 ( .A(n19699), .B(n25337), .Z(n25335) );
  XNOR U27125 ( .A(n19698), .B(n25336), .Z(n25337) );
  NAND U27126 ( .A(n25338), .B(n[260]), .Z(n19698) );
  NAND U27127 ( .A(n21523), .B(n[260]), .Z(n25338) );
  XNOR U27128 ( .A(n25339), .B(n25336), .Z(n19699) );
  XOR U27129 ( .A(n25340), .B(n25341), .Z(n25336) );
  AND U27130 ( .A(n19706), .B(n25342), .Z(n25340) );
  XNOR U27131 ( .A(n19705), .B(n25341), .Z(n25342) );
  NAND U27132 ( .A(n25343), .B(n[259]), .Z(n19705) );
  NAND U27133 ( .A(n21523), .B(n[259]), .Z(n25343) );
  XNOR U27134 ( .A(n25344), .B(n25341), .Z(n19706) );
  XOR U27135 ( .A(n25345), .B(n25346), .Z(n25341) );
  AND U27136 ( .A(n19713), .B(n25347), .Z(n25345) );
  XNOR U27137 ( .A(n19712), .B(n25346), .Z(n25347) );
  NAND U27138 ( .A(n25348), .B(n[258]), .Z(n19712) );
  NAND U27139 ( .A(n21523), .B(n[258]), .Z(n25348) );
  XNOR U27140 ( .A(n25349), .B(n25346), .Z(n19713) );
  XOR U27141 ( .A(n25350), .B(n25351), .Z(n25346) );
  AND U27142 ( .A(n19720), .B(n25352), .Z(n25350) );
  XNOR U27143 ( .A(n19719), .B(n25351), .Z(n25352) );
  NAND U27144 ( .A(n25353), .B(n[257]), .Z(n19719) );
  NAND U27145 ( .A(n21523), .B(n[257]), .Z(n25353) );
  XNOR U27146 ( .A(n25354), .B(n25351), .Z(n19720) );
  XOR U27147 ( .A(n25355), .B(n25356), .Z(n25351) );
  AND U27148 ( .A(n19727), .B(n25357), .Z(n25355) );
  XNOR U27149 ( .A(n19726), .B(n25356), .Z(n25357) );
  NAND U27150 ( .A(n25358), .B(n[256]), .Z(n19726) );
  NAND U27151 ( .A(n21523), .B(n[256]), .Z(n25358) );
  XNOR U27152 ( .A(n25359), .B(n25356), .Z(n19727) );
  XOR U27153 ( .A(n25360), .B(n25361), .Z(n25356) );
  AND U27154 ( .A(n19734), .B(n25362), .Z(n25360) );
  XNOR U27155 ( .A(n19733), .B(n25361), .Z(n25362) );
  NAND U27156 ( .A(n25363), .B(n[255]), .Z(n19733) );
  NAND U27157 ( .A(n21523), .B(n[255]), .Z(n25363) );
  XNOR U27158 ( .A(n25364), .B(n25361), .Z(n19734) );
  XOR U27159 ( .A(n25365), .B(n25366), .Z(n25361) );
  AND U27160 ( .A(n19741), .B(n25367), .Z(n25365) );
  XNOR U27161 ( .A(n19740), .B(n25366), .Z(n25367) );
  NAND U27162 ( .A(n25368), .B(n[254]), .Z(n19740) );
  NAND U27163 ( .A(n21523), .B(n[254]), .Z(n25368) );
  XNOR U27164 ( .A(n25369), .B(n25366), .Z(n19741) );
  XOR U27165 ( .A(n25370), .B(n25371), .Z(n25366) );
  AND U27166 ( .A(n19748), .B(n25372), .Z(n25370) );
  XNOR U27167 ( .A(n19747), .B(n25371), .Z(n25372) );
  NAND U27168 ( .A(n25373), .B(n[253]), .Z(n19747) );
  NAND U27169 ( .A(n21523), .B(n[253]), .Z(n25373) );
  XNOR U27170 ( .A(n25374), .B(n25371), .Z(n19748) );
  XOR U27171 ( .A(n25375), .B(n25376), .Z(n25371) );
  AND U27172 ( .A(n19755), .B(n25377), .Z(n25375) );
  XNOR U27173 ( .A(n19754), .B(n25376), .Z(n25377) );
  NAND U27174 ( .A(n25378), .B(n[252]), .Z(n19754) );
  NAND U27175 ( .A(n21523), .B(n[252]), .Z(n25378) );
  XNOR U27176 ( .A(n25379), .B(n25376), .Z(n19755) );
  XOR U27177 ( .A(n25380), .B(n25381), .Z(n25376) );
  AND U27178 ( .A(n19762), .B(n25382), .Z(n25380) );
  XNOR U27179 ( .A(n19761), .B(n25381), .Z(n25382) );
  NAND U27180 ( .A(n25383), .B(n[251]), .Z(n19761) );
  NAND U27181 ( .A(n21523), .B(n[251]), .Z(n25383) );
  XNOR U27182 ( .A(n25384), .B(n25381), .Z(n19762) );
  XOR U27183 ( .A(n25385), .B(n25386), .Z(n25381) );
  AND U27184 ( .A(n19769), .B(n25387), .Z(n25385) );
  XNOR U27185 ( .A(n19768), .B(n25386), .Z(n25387) );
  NAND U27186 ( .A(n25388), .B(n[250]), .Z(n19768) );
  NAND U27187 ( .A(n21523), .B(n[250]), .Z(n25388) );
  XNOR U27188 ( .A(n25389), .B(n25386), .Z(n19769) );
  XOR U27189 ( .A(n25390), .B(n25391), .Z(n25386) );
  AND U27190 ( .A(n19776), .B(n25392), .Z(n25390) );
  XNOR U27191 ( .A(n19775), .B(n25391), .Z(n25392) );
  NAND U27192 ( .A(n25393), .B(n[249]), .Z(n19775) );
  NAND U27193 ( .A(n21523), .B(n[249]), .Z(n25393) );
  XNOR U27194 ( .A(n25394), .B(n25391), .Z(n19776) );
  XOR U27195 ( .A(n25395), .B(n25396), .Z(n25391) );
  AND U27196 ( .A(n19783), .B(n25397), .Z(n25395) );
  XNOR U27197 ( .A(n19782), .B(n25396), .Z(n25397) );
  NAND U27198 ( .A(n25398), .B(n[248]), .Z(n19782) );
  NAND U27199 ( .A(n21523), .B(n[248]), .Z(n25398) );
  XNOR U27200 ( .A(n25399), .B(n25396), .Z(n19783) );
  XOR U27201 ( .A(n25400), .B(n25401), .Z(n25396) );
  AND U27202 ( .A(n19790), .B(n25402), .Z(n25400) );
  XNOR U27203 ( .A(n19789), .B(n25401), .Z(n25402) );
  NAND U27204 ( .A(n25403), .B(n[247]), .Z(n19789) );
  NAND U27205 ( .A(n21523), .B(n[247]), .Z(n25403) );
  XNOR U27206 ( .A(n25404), .B(n25401), .Z(n19790) );
  XOR U27207 ( .A(n25405), .B(n25406), .Z(n25401) );
  AND U27208 ( .A(n19797), .B(n25407), .Z(n25405) );
  XNOR U27209 ( .A(n19796), .B(n25406), .Z(n25407) );
  NAND U27210 ( .A(n25408), .B(n[246]), .Z(n19796) );
  NAND U27211 ( .A(n21523), .B(n[246]), .Z(n25408) );
  XNOR U27212 ( .A(n25409), .B(n25406), .Z(n19797) );
  XOR U27213 ( .A(n25410), .B(n25411), .Z(n25406) );
  AND U27214 ( .A(n19804), .B(n25412), .Z(n25410) );
  XNOR U27215 ( .A(n19803), .B(n25411), .Z(n25412) );
  NAND U27216 ( .A(n25413), .B(n[245]), .Z(n19803) );
  NAND U27217 ( .A(n21523), .B(n[245]), .Z(n25413) );
  XNOR U27218 ( .A(n25414), .B(n25411), .Z(n19804) );
  XOR U27219 ( .A(n25415), .B(n25416), .Z(n25411) );
  AND U27220 ( .A(n19811), .B(n25417), .Z(n25415) );
  XNOR U27221 ( .A(n19810), .B(n25416), .Z(n25417) );
  NAND U27222 ( .A(n25418), .B(n[244]), .Z(n19810) );
  NAND U27223 ( .A(n21523), .B(n[244]), .Z(n25418) );
  XNOR U27224 ( .A(n25419), .B(n25416), .Z(n19811) );
  XOR U27225 ( .A(n25420), .B(n25421), .Z(n25416) );
  AND U27226 ( .A(n19818), .B(n25422), .Z(n25420) );
  XNOR U27227 ( .A(n19817), .B(n25421), .Z(n25422) );
  NAND U27228 ( .A(n25423), .B(n[243]), .Z(n19817) );
  NAND U27229 ( .A(n21523), .B(n[243]), .Z(n25423) );
  XNOR U27230 ( .A(n25424), .B(n25421), .Z(n19818) );
  XOR U27231 ( .A(n25425), .B(n25426), .Z(n25421) );
  AND U27232 ( .A(n19825), .B(n25427), .Z(n25425) );
  XNOR U27233 ( .A(n19824), .B(n25426), .Z(n25427) );
  NAND U27234 ( .A(n25428), .B(n[242]), .Z(n19824) );
  NAND U27235 ( .A(n21523), .B(n[242]), .Z(n25428) );
  XNOR U27236 ( .A(n25429), .B(n25426), .Z(n19825) );
  XOR U27237 ( .A(n25430), .B(n25431), .Z(n25426) );
  AND U27238 ( .A(n19832), .B(n25432), .Z(n25430) );
  XNOR U27239 ( .A(n19831), .B(n25431), .Z(n25432) );
  NAND U27240 ( .A(n25433), .B(n[241]), .Z(n19831) );
  NAND U27241 ( .A(n21523), .B(n[241]), .Z(n25433) );
  XNOR U27242 ( .A(n25434), .B(n25431), .Z(n19832) );
  XOR U27243 ( .A(n25435), .B(n25436), .Z(n25431) );
  AND U27244 ( .A(n19839), .B(n25437), .Z(n25435) );
  XNOR U27245 ( .A(n19838), .B(n25436), .Z(n25437) );
  NAND U27246 ( .A(n25438), .B(n[240]), .Z(n19838) );
  NAND U27247 ( .A(n21523), .B(n[240]), .Z(n25438) );
  XNOR U27248 ( .A(n25439), .B(n25436), .Z(n19839) );
  XOR U27249 ( .A(n25440), .B(n25441), .Z(n25436) );
  AND U27250 ( .A(n19846), .B(n25442), .Z(n25440) );
  XNOR U27251 ( .A(n19845), .B(n25441), .Z(n25442) );
  NAND U27252 ( .A(n25443), .B(n[239]), .Z(n19845) );
  NAND U27253 ( .A(n21523), .B(n[239]), .Z(n25443) );
  XNOR U27254 ( .A(n25444), .B(n25441), .Z(n19846) );
  XOR U27255 ( .A(n25445), .B(n25446), .Z(n25441) );
  AND U27256 ( .A(n19853), .B(n25447), .Z(n25445) );
  XNOR U27257 ( .A(n19852), .B(n25446), .Z(n25447) );
  NAND U27258 ( .A(n25448), .B(n[238]), .Z(n19852) );
  NAND U27259 ( .A(n21523), .B(n[238]), .Z(n25448) );
  XNOR U27260 ( .A(n25449), .B(n25446), .Z(n19853) );
  XOR U27261 ( .A(n25450), .B(n25451), .Z(n25446) );
  AND U27262 ( .A(n19860), .B(n25452), .Z(n25450) );
  XNOR U27263 ( .A(n19859), .B(n25451), .Z(n25452) );
  NAND U27264 ( .A(n25453), .B(n[237]), .Z(n19859) );
  NAND U27265 ( .A(n21523), .B(n[237]), .Z(n25453) );
  XNOR U27266 ( .A(n25454), .B(n25451), .Z(n19860) );
  XOR U27267 ( .A(n25455), .B(n25456), .Z(n25451) );
  AND U27268 ( .A(n19867), .B(n25457), .Z(n25455) );
  XNOR U27269 ( .A(n19866), .B(n25456), .Z(n25457) );
  NAND U27270 ( .A(n25458), .B(n[236]), .Z(n19866) );
  NAND U27271 ( .A(n21523), .B(n[236]), .Z(n25458) );
  XNOR U27272 ( .A(n25459), .B(n25456), .Z(n19867) );
  XOR U27273 ( .A(n25460), .B(n25461), .Z(n25456) );
  AND U27274 ( .A(n19874), .B(n25462), .Z(n25460) );
  XNOR U27275 ( .A(n19873), .B(n25461), .Z(n25462) );
  NAND U27276 ( .A(n25463), .B(n[235]), .Z(n19873) );
  NAND U27277 ( .A(n21523), .B(n[235]), .Z(n25463) );
  XNOR U27278 ( .A(n25464), .B(n25461), .Z(n19874) );
  XOR U27279 ( .A(n25465), .B(n25466), .Z(n25461) );
  AND U27280 ( .A(n19881), .B(n25467), .Z(n25465) );
  XNOR U27281 ( .A(n19880), .B(n25466), .Z(n25467) );
  NAND U27282 ( .A(n25468), .B(n[234]), .Z(n19880) );
  NAND U27283 ( .A(n21523), .B(n[234]), .Z(n25468) );
  XNOR U27284 ( .A(n25469), .B(n25466), .Z(n19881) );
  XOR U27285 ( .A(n25470), .B(n25471), .Z(n25466) );
  AND U27286 ( .A(n19888), .B(n25472), .Z(n25470) );
  XNOR U27287 ( .A(n19887), .B(n25471), .Z(n25472) );
  NAND U27288 ( .A(n25473), .B(n[233]), .Z(n19887) );
  NAND U27289 ( .A(n21523), .B(n[233]), .Z(n25473) );
  XNOR U27290 ( .A(n25474), .B(n25471), .Z(n19888) );
  XOR U27291 ( .A(n25475), .B(n25476), .Z(n25471) );
  AND U27292 ( .A(n19895), .B(n25477), .Z(n25475) );
  XNOR U27293 ( .A(n19894), .B(n25476), .Z(n25477) );
  NAND U27294 ( .A(n25478), .B(n[232]), .Z(n19894) );
  NAND U27295 ( .A(n21523), .B(n[232]), .Z(n25478) );
  XNOR U27296 ( .A(n25479), .B(n25476), .Z(n19895) );
  XOR U27297 ( .A(n25480), .B(n25481), .Z(n25476) );
  AND U27298 ( .A(n19902), .B(n25482), .Z(n25480) );
  XNOR U27299 ( .A(n19901), .B(n25481), .Z(n25482) );
  NAND U27300 ( .A(n25483), .B(n[231]), .Z(n19901) );
  NAND U27301 ( .A(n21523), .B(n[231]), .Z(n25483) );
  XNOR U27302 ( .A(n25484), .B(n25481), .Z(n19902) );
  XOR U27303 ( .A(n25485), .B(n25486), .Z(n25481) );
  AND U27304 ( .A(n19909), .B(n25487), .Z(n25485) );
  XNOR U27305 ( .A(n19908), .B(n25486), .Z(n25487) );
  NAND U27306 ( .A(n25488), .B(n[230]), .Z(n19908) );
  NAND U27307 ( .A(n21523), .B(n[230]), .Z(n25488) );
  XNOR U27308 ( .A(n25489), .B(n25486), .Z(n19909) );
  XOR U27309 ( .A(n25490), .B(n25491), .Z(n25486) );
  AND U27310 ( .A(n19916), .B(n25492), .Z(n25490) );
  XNOR U27311 ( .A(n19915), .B(n25491), .Z(n25492) );
  NAND U27312 ( .A(n25493), .B(n[229]), .Z(n19915) );
  NAND U27313 ( .A(n21523), .B(n[229]), .Z(n25493) );
  XNOR U27314 ( .A(n25494), .B(n25491), .Z(n19916) );
  XOR U27315 ( .A(n25495), .B(n25496), .Z(n25491) );
  AND U27316 ( .A(n19923), .B(n25497), .Z(n25495) );
  XNOR U27317 ( .A(n19922), .B(n25496), .Z(n25497) );
  NAND U27318 ( .A(n25498), .B(n[228]), .Z(n19922) );
  NAND U27319 ( .A(n21523), .B(n[228]), .Z(n25498) );
  XNOR U27320 ( .A(n25499), .B(n25496), .Z(n19923) );
  XOR U27321 ( .A(n25500), .B(n25501), .Z(n25496) );
  AND U27322 ( .A(n19930), .B(n25502), .Z(n25500) );
  XNOR U27323 ( .A(n19929), .B(n25501), .Z(n25502) );
  NAND U27324 ( .A(n25503), .B(n[227]), .Z(n19929) );
  NAND U27325 ( .A(n21523), .B(n[227]), .Z(n25503) );
  XNOR U27326 ( .A(n25504), .B(n25501), .Z(n19930) );
  XOR U27327 ( .A(n25505), .B(n25506), .Z(n25501) );
  AND U27328 ( .A(n19937), .B(n25507), .Z(n25505) );
  XNOR U27329 ( .A(n19936), .B(n25506), .Z(n25507) );
  NAND U27330 ( .A(n25508), .B(n[226]), .Z(n19936) );
  NAND U27331 ( .A(n21523), .B(n[226]), .Z(n25508) );
  XNOR U27332 ( .A(n25509), .B(n25506), .Z(n19937) );
  XOR U27333 ( .A(n25510), .B(n25511), .Z(n25506) );
  AND U27334 ( .A(n19944), .B(n25512), .Z(n25510) );
  XNOR U27335 ( .A(n19943), .B(n25511), .Z(n25512) );
  NAND U27336 ( .A(n25513), .B(n[225]), .Z(n19943) );
  NAND U27337 ( .A(n21523), .B(n[225]), .Z(n25513) );
  XNOR U27338 ( .A(n25514), .B(n25511), .Z(n19944) );
  XOR U27339 ( .A(n25515), .B(n25516), .Z(n25511) );
  AND U27340 ( .A(n19951), .B(n25517), .Z(n25515) );
  XNOR U27341 ( .A(n19950), .B(n25516), .Z(n25517) );
  NAND U27342 ( .A(n25518), .B(n[224]), .Z(n19950) );
  NAND U27343 ( .A(n21523), .B(n[224]), .Z(n25518) );
  XNOR U27344 ( .A(n25519), .B(n25516), .Z(n19951) );
  XOR U27345 ( .A(n25520), .B(n25521), .Z(n25516) );
  AND U27346 ( .A(n19958), .B(n25522), .Z(n25520) );
  XNOR U27347 ( .A(n19957), .B(n25521), .Z(n25522) );
  NAND U27348 ( .A(n25523), .B(n[223]), .Z(n19957) );
  NAND U27349 ( .A(n21523), .B(n[223]), .Z(n25523) );
  XNOR U27350 ( .A(n25524), .B(n25521), .Z(n19958) );
  XOR U27351 ( .A(n25525), .B(n25526), .Z(n25521) );
  AND U27352 ( .A(n19965), .B(n25527), .Z(n25525) );
  XNOR U27353 ( .A(n19964), .B(n25526), .Z(n25527) );
  NAND U27354 ( .A(n25528), .B(n[222]), .Z(n19964) );
  NAND U27355 ( .A(n21523), .B(n[222]), .Z(n25528) );
  XNOR U27356 ( .A(n25529), .B(n25526), .Z(n19965) );
  XOR U27357 ( .A(n25530), .B(n25531), .Z(n25526) );
  AND U27358 ( .A(n19972), .B(n25532), .Z(n25530) );
  XNOR U27359 ( .A(n19971), .B(n25531), .Z(n25532) );
  NAND U27360 ( .A(n25533), .B(n[221]), .Z(n19971) );
  NAND U27361 ( .A(n21523), .B(n[221]), .Z(n25533) );
  XNOR U27362 ( .A(n25534), .B(n25531), .Z(n19972) );
  XOR U27363 ( .A(n25535), .B(n25536), .Z(n25531) );
  AND U27364 ( .A(n19979), .B(n25537), .Z(n25535) );
  XNOR U27365 ( .A(n19978), .B(n25536), .Z(n25537) );
  NAND U27366 ( .A(n25538), .B(n[220]), .Z(n19978) );
  NAND U27367 ( .A(n21523), .B(n[220]), .Z(n25538) );
  XNOR U27368 ( .A(n25539), .B(n25536), .Z(n19979) );
  XOR U27369 ( .A(n25540), .B(n25541), .Z(n25536) );
  AND U27370 ( .A(n19986), .B(n25542), .Z(n25540) );
  XNOR U27371 ( .A(n19985), .B(n25541), .Z(n25542) );
  NAND U27372 ( .A(n25543), .B(n[219]), .Z(n19985) );
  NAND U27373 ( .A(n21523), .B(n[219]), .Z(n25543) );
  XNOR U27374 ( .A(n25544), .B(n25541), .Z(n19986) );
  XOR U27375 ( .A(n25545), .B(n25546), .Z(n25541) );
  AND U27376 ( .A(n19993), .B(n25547), .Z(n25545) );
  XNOR U27377 ( .A(n19992), .B(n25546), .Z(n25547) );
  NAND U27378 ( .A(n25548), .B(n[218]), .Z(n19992) );
  NAND U27379 ( .A(n21523), .B(n[218]), .Z(n25548) );
  XNOR U27380 ( .A(n25549), .B(n25546), .Z(n19993) );
  XOR U27381 ( .A(n25550), .B(n25551), .Z(n25546) );
  AND U27382 ( .A(n20000), .B(n25552), .Z(n25550) );
  XNOR U27383 ( .A(n19999), .B(n25551), .Z(n25552) );
  NAND U27384 ( .A(n25553), .B(n[217]), .Z(n19999) );
  NAND U27385 ( .A(n21523), .B(n[217]), .Z(n25553) );
  XNOR U27386 ( .A(n25554), .B(n25551), .Z(n20000) );
  XOR U27387 ( .A(n25555), .B(n25556), .Z(n25551) );
  AND U27388 ( .A(n20007), .B(n25557), .Z(n25555) );
  XNOR U27389 ( .A(n20006), .B(n25556), .Z(n25557) );
  NAND U27390 ( .A(n25558), .B(n[216]), .Z(n20006) );
  NAND U27391 ( .A(n21523), .B(n[216]), .Z(n25558) );
  XNOR U27392 ( .A(n25559), .B(n25556), .Z(n20007) );
  XOR U27393 ( .A(n25560), .B(n25561), .Z(n25556) );
  AND U27394 ( .A(n20014), .B(n25562), .Z(n25560) );
  XNOR U27395 ( .A(n20013), .B(n25561), .Z(n25562) );
  NAND U27396 ( .A(n25563), .B(n[215]), .Z(n20013) );
  NAND U27397 ( .A(n21523), .B(n[215]), .Z(n25563) );
  XNOR U27398 ( .A(n25564), .B(n25561), .Z(n20014) );
  XOR U27399 ( .A(n25565), .B(n25566), .Z(n25561) );
  AND U27400 ( .A(n20021), .B(n25567), .Z(n25565) );
  XNOR U27401 ( .A(n20020), .B(n25566), .Z(n25567) );
  NAND U27402 ( .A(n25568), .B(n[214]), .Z(n20020) );
  NAND U27403 ( .A(n21523), .B(n[214]), .Z(n25568) );
  XNOR U27404 ( .A(n25569), .B(n25566), .Z(n20021) );
  XOR U27405 ( .A(n25570), .B(n25571), .Z(n25566) );
  AND U27406 ( .A(n20028), .B(n25572), .Z(n25570) );
  XNOR U27407 ( .A(n20027), .B(n25571), .Z(n25572) );
  NAND U27408 ( .A(n25573), .B(n[213]), .Z(n20027) );
  NAND U27409 ( .A(n21523), .B(n[213]), .Z(n25573) );
  XNOR U27410 ( .A(n25574), .B(n25571), .Z(n20028) );
  XOR U27411 ( .A(n25575), .B(n25576), .Z(n25571) );
  AND U27412 ( .A(n20035), .B(n25577), .Z(n25575) );
  XNOR U27413 ( .A(n20034), .B(n25576), .Z(n25577) );
  NAND U27414 ( .A(n25578), .B(n[212]), .Z(n20034) );
  NAND U27415 ( .A(n21523), .B(n[212]), .Z(n25578) );
  XNOR U27416 ( .A(n25579), .B(n25576), .Z(n20035) );
  XOR U27417 ( .A(n25580), .B(n25581), .Z(n25576) );
  AND U27418 ( .A(n20042), .B(n25582), .Z(n25580) );
  XNOR U27419 ( .A(n20041), .B(n25581), .Z(n25582) );
  NAND U27420 ( .A(n25583), .B(n[211]), .Z(n20041) );
  NAND U27421 ( .A(n21523), .B(n[211]), .Z(n25583) );
  XNOR U27422 ( .A(n25584), .B(n25581), .Z(n20042) );
  XOR U27423 ( .A(n25585), .B(n25586), .Z(n25581) );
  AND U27424 ( .A(n20049), .B(n25587), .Z(n25585) );
  XNOR U27425 ( .A(n20048), .B(n25586), .Z(n25587) );
  NAND U27426 ( .A(n25588), .B(n[210]), .Z(n20048) );
  NAND U27427 ( .A(n21523), .B(n[210]), .Z(n25588) );
  XNOR U27428 ( .A(n25589), .B(n25586), .Z(n20049) );
  XOR U27429 ( .A(n25590), .B(n25591), .Z(n25586) );
  AND U27430 ( .A(n20056), .B(n25592), .Z(n25590) );
  XNOR U27431 ( .A(n20055), .B(n25591), .Z(n25592) );
  NAND U27432 ( .A(n25593), .B(n[209]), .Z(n20055) );
  NAND U27433 ( .A(n21523), .B(n[209]), .Z(n25593) );
  XNOR U27434 ( .A(n25594), .B(n25591), .Z(n20056) );
  XOR U27435 ( .A(n25595), .B(n25596), .Z(n25591) );
  AND U27436 ( .A(n20063), .B(n25597), .Z(n25595) );
  XNOR U27437 ( .A(n20062), .B(n25596), .Z(n25597) );
  NAND U27438 ( .A(n25598), .B(n[208]), .Z(n20062) );
  NAND U27439 ( .A(n21523), .B(n[208]), .Z(n25598) );
  XNOR U27440 ( .A(n25599), .B(n25596), .Z(n20063) );
  XOR U27441 ( .A(n25600), .B(n25601), .Z(n25596) );
  AND U27442 ( .A(n20070), .B(n25602), .Z(n25600) );
  XNOR U27443 ( .A(n20069), .B(n25601), .Z(n25602) );
  NAND U27444 ( .A(n25603), .B(n[207]), .Z(n20069) );
  NAND U27445 ( .A(n21523), .B(n[207]), .Z(n25603) );
  XNOR U27446 ( .A(n25604), .B(n25601), .Z(n20070) );
  XOR U27447 ( .A(n25605), .B(n25606), .Z(n25601) );
  AND U27448 ( .A(n20077), .B(n25607), .Z(n25605) );
  XNOR U27449 ( .A(n20076), .B(n25606), .Z(n25607) );
  NAND U27450 ( .A(n25608), .B(n[206]), .Z(n20076) );
  NAND U27451 ( .A(n21523), .B(n[206]), .Z(n25608) );
  XNOR U27452 ( .A(n25609), .B(n25606), .Z(n20077) );
  XOR U27453 ( .A(n25610), .B(n25611), .Z(n25606) );
  AND U27454 ( .A(n20084), .B(n25612), .Z(n25610) );
  XNOR U27455 ( .A(n20083), .B(n25611), .Z(n25612) );
  NAND U27456 ( .A(n25613), .B(n[205]), .Z(n20083) );
  NAND U27457 ( .A(n21523), .B(n[205]), .Z(n25613) );
  XNOR U27458 ( .A(n25614), .B(n25611), .Z(n20084) );
  XOR U27459 ( .A(n25615), .B(n25616), .Z(n25611) );
  AND U27460 ( .A(n20091), .B(n25617), .Z(n25615) );
  XNOR U27461 ( .A(n20090), .B(n25616), .Z(n25617) );
  NAND U27462 ( .A(n25618), .B(n[204]), .Z(n20090) );
  NAND U27463 ( .A(n21523), .B(n[204]), .Z(n25618) );
  XNOR U27464 ( .A(n25619), .B(n25616), .Z(n20091) );
  XOR U27465 ( .A(n25620), .B(n25621), .Z(n25616) );
  AND U27466 ( .A(n20098), .B(n25622), .Z(n25620) );
  XNOR U27467 ( .A(n20097), .B(n25621), .Z(n25622) );
  NAND U27468 ( .A(n25623), .B(n[203]), .Z(n20097) );
  NAND U27469 ( .A(n21523), .B(n[203]), .Z(n25623) );
  XNOR U27470 ( .A(n25624), .B(n25621), .Z(n20098) );
  XOR U27471 ( .A(n25625), .B(n25626), .Z(n25621) );
  AND U27472 ( .A(n20105), .B(n25627), .Z(n25625) );
  XNOR U27473 ( .A(n20104), .B(n25626), .Z(n25627) );
  NAND U27474 ( .A(n25628), .B(n[202]), .Z(n20104) );
  NAND U27475 ( .A(n21523), .B(n[202]), .Z(n25628) );
  XNOR U27476 ( .A(n25629), .B(n25626), .Z(n20105) );
  XOR U27477 ( .A(n25630), .B(n25631), .Z(n25626) );
  AND U27478 ( .A(n20112), .B(n25632), .Z(n25630) );
  XNOR U27479 ( .A(n20111), .B(n25631), .Z(n25632) );
  NAND U27480 ( .A(n25633), .B(n[201]), .Z(n20111) );
  NAND U27481 ( .A(n21523), .B(n[201]), .Z(n25633) );
  XNOR U27482 ( .A(n25634), .B(n25631), .Z(n20112) );
  XOR U27483 ( .A(n25635), .B(n25636), .Z(n25631) );
  AND U27484 ( .A(n20119), .B(n25637), .Z(n25635) );
  XNOR U27485 ( .A(n20118), .B(n25636), .Z(n25637) );
  NAND U27486 ( .A(n25638), .B(n[200]), .Z(n20118) );
  NAND U27487 ( .A(n21523), .B(n[200]), .Z(n25638) );
  XNOR U27488 ( .A(n25639), .B(n25636), .Z(n20119) );
  XOR U27489 ( .A(n25640), .B(n25641), .Z(n25636) );
  AND U27490 ( .A(n20126), .B(n25642), .Z(n25640) );
  XNOR U27491 ( .A(n20125), .B(n25641), .Z(n25642) );
  NAND U27492 ( .A(n25643), .B(n[199]), .Z(n20125) );
  NAND U27493 ( .A(n21523), .B(n[199]), .Z(n25643) );
  XNOR U27494 ( .A(n25644), .B(n25641), .Z(n20126) );
  XOR U27495 ( .A(n25645), .B(n25646), .Z(n25641) );
  AND U27496 ( .A(n20133), .B(n25647), .Z(n25645) );
  XNOR U27497 ( .A(n20132), .B(n25646), .Z(n25647) );
  NAND U27498 ( .A(n25648), .B(n[198]), .Z(n20132) );
  NAND U27499 ( .A(n21523), .B(n[198]), .Z(n25648) );
  XNOR U27500 ( .A(n25649), .B(n25646), .Z(n20133) );
  XOR U27501 ( .A(n25650), .B(n25651), .Z(n25646) );
  AND U27502 ( .A(n20140), .B(n25652), .Z(n25650) );
  XNOR U27503 ( .A(n20139), .B(n25651), .Z(n25652) );
  NAND U27504 ( .A(n25653), .B(n[197]), .Z(n20139) );
  NAND U27505 ( .A(n21523), .B(n[197]), .Z(n25653) );
  XNOR U27506 ( .A(n25654), .B(n25651), .Z(n20140) );
  XOR U27507 ( .A(n25655), .B(n25656), .Z(n25651) );
  AND U27508 ( .A(n20147), .B(n25657), .Z(n25655) );
  XNOR U27509 ( .A(n20146), .B(n25656), .Z(n25657) );
  NAND U27510 ( .A(n25658), .B(n[196]), .Z(n20146) );
  NAND U27511 ( .A(n21523), .B(n[196]), .Z(n25658) );
  XNOR U27512 ( .A(n25659), .B(n25656), .Z(n20147) );
  XOR U27513 ( .A(n25660), .B(n25661), .Z(n25656) );
  AND U27514 ( .A(n20154), .B(n25662), .Z(n25660) );
  XNOR U27515 ( .A(n20153), .B(n25661), .Z(n25662) );
  NAND U27516 ( .A(n25663), .B(n[195]), .Z(n20153) );
  NAND U27517 ( .A(n21523), .B(n[195]), .Z(n25663) );
  XNOR U27518 ( .A(n25664), .B(n25661), .Z(n20154) );
  XOR U27519 ( .A(n25665), .B(n25666), .Z(n25661) );
  AND U27520 ( .A(n20161), .B(n25667), .Z(n25665) );
  XNOR U27521 ( .A(n20160), .B(n25666), .Z(n25667) );
  NAND U27522 ( .A(n25668), .B(n[194]), .Z(n20160) );
  NAND U27523 ( .A(n21523), .B(n[194]), .Z(n25668) );
  XNOR U27524 ( .A(n25669), .B(n25666), .Z(n20161) );
  XOR U27525 ( .A(n25670), .B(n25671), .Z(n25666) );
  AND U27526 ( .A(n20168), .B(n25672), .Z(n25670) );
  XNOR U27527 ( .A(n20167), .B(n25671), .Z(n25672) );
  NAND U27528 ( .A(n25673), .B(n[193]), .Z(n20167) );
  NAND U27529 ( .A(n21523), .B(n[193]), .Z(n25673) );
  XNOR U27530 ( .A(n25674), .B(n25671), .Z(n20168) );
  XOR U27531 ( .A(n25675), .B(n25676), .Z(n25671) );
  AND U27532 ( .A(n20175), .B(n25677), .Z(n25675) );
  XNOR U27533 ( .A(n20174), .B(n25676), .Z(n25677) );
  NAND U27534 ( .A(n25678), .B(n[192]), .Z(n20174) );
  NAND U27535 ( .A(n21523), .B(n[192]), .Z(n25678) );
  XNOR U27536 ( .A(n25679), .B(n25676), .Z(n20175) );
  XOR U27537 ( .A(n25680), .B(n25681), .Z(n25676) );
  AND U27538 ( .A(n20182), .B(n25682), .Z(n25680) );
  XNOR U27539 ( .A(n20181), .B(n25681), .Z(n25682) );
  NAND U27540 ( .A(n25683), .B(n[191]), .Z(n20181) );
  NAND U27541 ( .A(n21523), .B(n[191]), .Z(n25683) );
  XNOR U27542 ( .A(n25684), .B(n25681), .Z(n20182) );
  XOR U27543 ( .A(n25685), .B(n25686), .Z(n25681) );
  AND U27544 ( .A(n20189), .B(n25687), .Z(n25685) );
  XNOR U27545 ( .A(n20188), .B(n25686), .Z(n25687) );
  NAND U27546 ( .A(n25688), .B(n[190]), .Z(n20188) );
  NAND U27547 ( .A(n21523), .B(n[190]), .Z(n25688) );
  XNOR U27548 ( .A(n25689), .B(n25686), .Z(n20189) );
  XOR U27549 ( .A(n25690), .B(n25691), .Z(n25686) );
  AND U27550 ( .A(n20196), .B(n25692), .Z(n25690) );
  XNOR U27551 ( .A(n20195), .B(n25691), .Z(n25692) );
  NAND U27552 ( .A(n25693), .B(n[189]), .Z(n20195) );
  NAND U27553 ( .A(n21523), .B(n[189]), .Z(n25693) );
  XNOR U27554 ( .A(n25694), .B(n25691), .Z(n20196) );
  XOR U27555 ( .A(n25695), .B(n25696), .Z(n25691) );
  AND U27556 ( .A(n20203), .B(n25697), .Z(n25695) );
  XNOR U27557 ( .A(n20202), .B(n25696), .Z(n25697) );
  NAND U27558 ( .A(n25698), .B(n[188]), .Z(n20202) );
  NAND U27559 ( .A(n21523), .B(n[188]), .Z(n25698) );
  XNOR U27560 ( .A(n25699), .B(n25696), .Z(n20203) );
  XOR U27561 ( .A(n25700), .B(n25701), .Z(n25696) );
  AND U27562 ( .A(n20210), .B(n25702), .Z(n25700) );
  XNOR U27563 ( .A(n20209), .B(n25701), .Z(n25702) );
  NAND U27564 ( .A(n25703), .B(n[187]), .Z(n20209) );
  NAND U27565 ( .A(n21523), .B(n[187]), .Z(n25703) );
  XNOR U27566 ( .A(n25704), .B(n25701), .Z(n20210) );
  XOR U27567 ( .A(n25705), .B(n25706), .Z(n25701) );
  AND U27568 ( .A(n20217), .B(n25707), .Z(n25705) );
  XNOR U27569 ( .A(n20216), .B(n25706), .Z(n25707) );
  NAND U27570 ( .A(n25708), .B(n[186]), .Z(n20216) );
  NAND U27571 ( .A(n21523), .B(n[186]), .Z(n25708) );
  XNOR U27572 ( .A(n25709), .B(n25706), .Z(n20217) );
  XOR U27573 ( .A(n25710), .B(n25711), .Z(n25706) );
  AND U27574 ( .A(n20224), .B(n25712), .Z(n25710) );
  XNOR U27575 ( .A(n20223), .B(n25711), .Z(n25712) );
  NAND U27576 ( .A(n25713), .B(n[185]), .Z(n20223) );
  NAND U27577 ( .A(n21523), .B(n[185]), .Z(n25713) );
  XNOR U27578 ( .A(n25714), .B(n25711), .Z(n20224) );
  XOR U27579 ( .A(n25715), .B(n25716), .Z(n25711) );
  AND U27580 ( .A(n20231), .B(n25717), .Z(n25715) );
  XNOR U27581 ( .A(n20230), .B(n25716), .Z(n25717) );
  NAND U27582 ( .A(n25718), .B(n[184]), .Z(n20230) );
  NAND U27583 ( .A(n21523), .B(n[184]), .Z(n25718) );
  XNOR U27584 ( .A(n25719), .B(n25716), .Z(n20231) );
  XOR U27585 ( .A(n25720), .B(n25721), .Z(n25716) );
  AND U27586 ( .A(n20238), .B(n25722), .Z(n25720) );
  XNOR U27587 ( .A(n20237), .B(n25721), .Z(n25722) );
  NAND U27588 ( .A(n25723), .B(n[183]), .Z(n20237) );
  NAND U27589 ( .A(n21523), .B(n[183]), .Z(n25723) );
  XNOR U27590 ( .A(n25724), .B(n25721), .Z(n20238) );
  XOR U27591 ( .A(n25725), .B(n25726), .Z(n25721) );
  AND U27592 ( .A(n20245), .B(n25727), .Z(n25725) );
  XNOR U27593 ( .A(n20244), .B(n25726), .Z(n25727) );
  NAND U27594 ( .A(n25728), .B(n[182]), .Z(n20244) );
  NAND U27595 ( .A(n21523), .B(n[182]), .Z(n25728) );
  XNOR U27596 ( .A(n25729), .B(n25726), .Z(n20245) );
  XOR U27597 ( .A(n25730), .B(n25731), .Z(n25726) );
  AND U27598 ( .A(n20252), .B(n25732), .Z(n25730) );
  XNOR U27599 ( .A(n20251), .B(n25731), .Z(n25732) );
  NAND U27600 ( .A(n25733), .B(n[181]), .Z(n20251) );
  NAND U27601 ( .A(n21523), .B(n[181]), .Z(n25733) );
  XNOR U27602 ( .A(n25734), .B(n25731), .Z(n20252) );
  XOR U27603 ( .A(n25735), .B(n25736), .Z(n25731) );
  AND U27604 ( .A(n20259), .B(n25737), .Z(n25735) );
  XNOR U27605 ( .A(n20258), .B(n25736), .Z(n25737) );
  NAND U27606 ( .A(n25738), .B(n[180]), .Z(n20258) );
  NAND U27607 ( .A(n21523), .B(n[180]), .Z(n25738) );
  XNOR U27608 ( .A(n25739), .B(n25736), .Z(n20259) );
  XOR U27609 ( .A(n25740), .B(n25741), .Z(n25736) );
  AND U27610 ( .A(n20266), .B(n25742), .Z(n25740) );
  XNOR U27611 ( .A(n20265), .B(n25741), .Z(n25742) );
  NAND U27612 ( .A(n25743), .B(n[179]), .Z(n20265) );
  NAND U27613 ( .A(n21523), .B(n[179]), .Z(n25743) );
  XNOR U27614 ( .A(n25744), .B(n25741), .Z(n20266) );
  XOR U27615 ( .A(n25745), .B(n25746), .Z(n25741) );
  AND U27616 ( .A(n20273), .B(n25747), .Z(n25745) );
  XNOR U27617 ( .A(n20272), .B(n25746), .Z(n25747) );
  NAND U27618 ( .A(n25748), .B(n[178]), .Z(n20272) );
  NAND U27619 ( .A(n21523), .B(n[178]), .Z(n25748) );
  XNOR U27620 ( .A(n25749), .B(n25746), .Z(n20273) );
  XOR U27621 ( .A(n25750), .B(n25751), .Z(n25746) );
  AND U27622 ( .A(n20280), .B(n25752), .Z(n25750) );
  XNOR U27623 ( .A(n20279), .B(n25751), .Z(n25752) );
  NAND U27624 ( .A(n25753), .B(n[177]), .Z(n20279) );
  NAND U27625 ( .A(n21523), .B(n[177]), .Z(n25753) );
  XNOR U27626 ( .A(n25754), .B(n25751), .Z(n20280) );
  XOR U27627 ( .A(n25755), .B(n25756), .Z(n25751) );
  AND U27628 ( .A(n20287), .B(n25757), .Z(n25755) );
  XNOR U27629 ( .A(n20286), .B(n25756), .Z(n25757) );
  NAND U27630 ( .A(n25758), .B(n[176]), .Z(n20286) );
  NAND U27631 ( .A(n21523), .B(n[176]), .Z(n25758) );
  XNOR U27632 ( .A(n25759), .B(n25756), .Z(n20287) );
  XOR U27633 ( .A(n25760), .B(n25761), .Z(n25756) );
  AND U27634 ( .A(n20294), .B(n25762), .Z(n25760) );
  XNOR U27635 ( .A(n20293), .B(n25761), .Z(n25762) );
  NAND U27636 ( .A(n25763), .B(n[175]), .Z(n20293) );
  NAND U27637 ( .A(n21523), .B(n[175]), .Z(n25763) );
  XNOR U27638 ( .A(n25764), .B(n25761), .Z(n20294) );
  XOR U27639 ( .A(n25765), .B(n25766), .Z(n25761) );
  AND U27640 ( .A(n20301), .B(n25767), .Z(n25765) );
  XNOR U27641 ( .A(n20300), .B(n25766), .Z(n25767) );
  NAND U27642 ( .A(n25768), .B(n[174]), .Z(n20300) );
  NAND U27643 ( .A(n21523), .B(n[174]), .Z(n25768) );
  XNOR U27644 ( .A(n25769), .B(n25766), .Z(n20301) );
  XOR U27645 ( .A(n25770), .B(n25771), .Z(n25766) );
  AND U27646 ( .A(n20308), .B(n25772), .Z(n25770) );
  XNOR U27647 ( .A(n20307), .B(n25771), .Z(n25772) );
  NAND U27648 ( .A(n25773), .B(n[173]), .Z(n20307) );
  NAND U27649 ( .A(n21523), .B(n[173]), .Z(n25773) );
  XNOR U27650 ( .A(n25774), .B(n25771), .Z(n20308) );
  XOR U27651 ( .A(n25775), .B(n25776), .Z(n25771) );
  AND U27652 ( .A(n20315), .B(n25777), .Z(n25775) );
  XNOR U27653 ( .A(n20314), .B(n25776), .Z(n25777) );
  NAND U27654 ( .A(n25778), .B(n[172]), .Z(n20314) );
  NAND U27655 ( .A(n21523), .B(n[172]), .Z(n25778) );
  XNOR U27656 ( .A(n25779), .B(n25776), .Z(n20315) );
  XOR U27657 ( .A(n25780), .B(n25781), .Z(n25776) );
  AND U27658 ( .A(n20322), .B(n25782), .Z(n25780) );
  XNOR U27659 ( .A(n20321), .B(n25781), .Z(n25782) );
  NAND U27660 ( .A(n25783), .B(n[171]), .Z(n20321) );
  NAND U27661 ( .A(n21523), .B(n[171]), .Z(n25783) );
  XNOR U27662 ( .A(n25784), .B(n25781), .Z(n20322) );
  XOR U27663 ( .A(n25785), .B(n25786), .Z(n25781) );
  AND U27664 ( .A(n20329), .B(n25787), .Z(n25785) );
  XNOR U27665 ( .A(n20328), .B(n25786), .Z(n25787) );
  NAND U27666 ( .A(n25788), .B(n[170]), .Z(n20328) );
  NAND U27667 ( .A(n21523), .B(n[170]), .Z(n25788) );
  XNOR U27668 ( .A(n25789), .B(n25786), .Z(n20329) );
  XOR U27669 ( .A(n25790), .B(n25791), .Z(n25786) );
  AND U27670 ( .A(n20336), .B(n25792), .Z(n25790) );
  XNOR U27671 ( .A(n20335), .B(n25791), .Z(n25792) );
  NAND U27672 ( .A(n25793), .B(n[169]), .Z(n20335) );
  NAND U27673 ( .A(n21523), .B(n[169]), .Z(n25793) );
  XNOR U27674 ( .A(n25794), .B(n25791), .Z(n20336) );
  XOR U27675 ( .A(n25795), .B(n25796), .Z(n25791) );
  AND U27676 ( .A(n20343), .B(n25797), .Z(n25795) );
  XNOR U27677 ( .A(n20342), .B(n25796), .Z(n25797) );
  NAND U27678 ( .A(n25798), .B(n[168]), .Z(n20342) );
  NAND U27679 ( .A(n21523), .B(n[168]), .Z(n25798) );
  XNOR U27680 ( .A(n25799), .B(n25796), .Z(n20343) );
  XOR U27681 ( .A(n25800), .B(n25801), .Z(n25796) );
  AND U27682 ( .A(n20350), .B(n25802), .Z(n25800) );
  XNOR U27683 ( .A(n20349), .B(n25801), .Z(n25802) );
  NAND U27684 ( .A(n25803), .B(n[167]), .Z(n20349) );
  NAND U27685 ( .A(n21523), .B(n[167]), .Z(n25803) );
  XNOR U27686 ( .A(n25804), .B(n25801), .Z(n20350) );
  XOR U27687 ( .A(n25805), .B(n25806), .Z(n25801) );
  AND U27688 ( .A(n20357), .B(n25807), .Z(n25805) );
  XNOR U27689 ( .A(n20356), .B(n25806), .Z(n25807) );
  NAND U27690 ( .A(n25808), .B(n[166]), .Z(n20356) );
  NAND U27691 ( .A(n21523), .B(n[166]), .Z(n25808) );
  XNOR U27692 ( .A(n25809), .B(n25806), .Z(n20357) );
  XOR U27693 ( .A(n25810), .B(n25811), .Z(n25806) );
  AND U27694 ( .A(n20364), .B(n25812), .Z(n25810) );
  XNOR U27695 ( .A(n20363), .B(n25811), .Z(n25812) );
  NAND U27696 ( .A(n25813), .B(n[165]), .Z(n20363) );
  NAND U27697 ( .A(n21523), .B(n[165]), .Z(n25813) );
  XNOR U27698 ( .A(n25814), .B(n25811), .Z(n20364) );
  XOR U27699 ( .A(n25815), .B(n25816), .Z(n25811) );
  AND U27700 ( .A(n20371), .B(n25817), .Z(n25815) );
  XNOR U27701 ( .A(n20370), .B(n25816), .Z(n25817) );
  NAND U27702 ( .A(n25818), .B(n[164]), .Z(n20370) );
  NAND U27703 ( .A(n21523), .B(n[164]), .Z(n25818) );
  XNOR U27704 ( .A(n25819), .B(n25816), .Z(n20371) );
  XOR U27705 ( .A(n25820), .B(n25821), .Z(n25816) );
  AND U27706 ( .A(n20378), .B(n25822), .Z(n25820) );
  XNOR U27707 ( .A(n20377), .B(n25821), .Z(n25822) );
  NAND U27708 ( .A(n25823), .B(n[163]), .Z(n20377) );
  NAND U27709 ( .A(n21523), .B(n[163]), .Z(n25823) );
  XNOR U27710 ( .A(n25824), .B(n25821), .Z(n20378) );
  XOR U27711 ( .A(n25825), .B(n25826), .Z(n25821) );
  AND U27712 ( .A(n20385), .B(n25827), .Z(n25825) );
  XNOR U27713 ( .A(n20384), .B(n25826), .Z(n25827) );
  NAND U27714 ( .A(n25828), .B(n[162]), .Z(n20384) );
  NAND U27715 ( .A(n21523), .B(n[162]), .Z(n25828) );
  XNOR U27716 ( .A(n25829), .B(n25826), .Z(n20385) );
  XOR U27717 ( .A(n25830), .B(n25831), .Z(n25826) );
  AND U27718 ( .A(n20392), .B(n25832), .Z(n25830) );
  XNOR U27719 ( .A(n20391), .B(n25831), .Z(n25832) );
  NAND U27720 ( .A(n25833), .B(n[161]), .Z(n20391) );
  NAND U27721 ( .A(n21523), .B(n[161]), .Z(n25833) );
  XNOR U27722 ( .A(n25834), .B(n25831), .Z(n20392) );
  XOR U27723 ( .A(n25835), .B(n25836), .Z(n25831) );
  AND U27724 ( .A(n20399), .B(n25837), .Z(n25835) );
  XNOR U27725 ( .A(n20398), .B(n25836), .Z(n25837) );
  NAND U27726 ( .A(n25838), .B(n[160]), .Z(n20398) );
  NAND U27727 ( .A(n21523), .B(n[160]), .Z(n25838) );
  XNOR U27728 ( .A(n25839), .B(n25836), .Z(n20399) );
  XOR U27729 ( .A(n25840), .B(n25841), .Z(n25836) );
  AND U27730 ( .A(n20406), .B(n25842), .Z(n25840) );
  XNOR U27731 ( .A(n20405), .B(n25841), .Z(n25842) );
  NAND U27732 ( .A(n25843), .B(n[159]), .Z(n20405) );
  NAND U27733 ( .A(n21523), .B(n[159]), .Z(n25843) );
  XNOR U27734 ( .A(n25844), .B(n25841), .Z(n20406) );
  XOR U27735 ( .A(n25845), .B(n25846), .Z(n25841) );
  AND U27736 ( .A(n20413), .B(n25847), .Z(n25845) );
  XNOR U27737 ( .A(n20412), .B(n25846), .Z(n25847) );
  NAND U27738 ( .A(n25848), .B(n[158]), .Z(n20412) );
  NAND U27739 ( .A(n21523), .B(n[158]), .Z(n25848) );
  XNOR U27740 ( .A(n25849), .B(n25846), .Z(n20413) );
  XOR U27741 ( .A(n25850), .B(n25851), .Z(n25846) );
  AND U27742 ( .A(n20420), .B(n25852), .Z(n25850) );
  XNOR U27743 ( .A(n20419), .B(n25851), .Z(n25852) );
  NAND U27744 ( .A(n25853), .B(n[157]), .Z(n20419) );
  NAND U27745 ( .A(n21523), .B(n[157]), .Z(n25853) );
  XNOR U27746 ( .A(n25854), .B(n25851), .Z(n20420) );
  XOR U27747 ( .A(n25855), .B(n25856), .Z(n25851) );
  AND U27748 ( .A(n20427), .B(n25857), .Z(n25855) );
  XNOR U27749 ( .A(n20426), .B(n25856), .Z(n25857) );
  NAND U27750 ( .A(n25858), .B(n[156]), .Z(n20426) );
  NAND U27751 ( .A(n21523), .B(n[156]), .Z(n25858) );
  XNOR U27752 ( .A(n25859), .B(n25856), .Z(n20427) );
  XOR U27753 ( .A(n25860), .B(n25861), .Z(n25856) );
  AND U27754 ( .A(n20434), .B(n25862), .Z(n25860) );
  XNOR U27755 ( .A(n20433), .B(n25861), .Z(n25862) );
  NAND U27756 ( .A(n25863), .B(n[155]), .Z(n20433) );
  NAND U27757 ( .A(n21523), .B(n[155]), .Z(n25863) );
  XNOR U27758 ( .A(n25864), .B(n25861), .Z(n20434) );
  XOR U27759 ( .A(n25865), .B(n25866), .Z(n25861) );
  AND U27760 ( .A(n20441), .B(n25867), .Z(n25865) );
  XNOR U27761 ( .A(n20440), .B(n25866), .Z(n25867) );
  NAND U27762 ( .A(n25868), .B(n[154]), .Z(n20440) );
  NAND U27763 ( .A(n21523), .B(n[154]), .Z(n25868) );
  XNOR U27764 ( .A(n25869), .B(n25866), .Z(n20441) );
  XOR U27765 ( .A(n25870), .B(n25871), .Z(n25866) );
  AND U27766 ( .A(n20448), .B(n25872), .Z(n25870) );
  XNOR U27767 ( .A(n20447), .B(n25871), .Z(n25872) );
  NAND U27768 ( .A(n25873), .B(n[153]), .Z(n20447) );
  NAND U27769 ( .A(n21523), .B(n[153]), .Z(n25873) );
  XNOR U27770 ( .A(n25874), .B(n25871), .Z(n20448) );
  XOR U27771 ( .A(n25875), .B(n25876), .Z(n25871) );
  AND U27772 ( .A(n20455), .B(n25877), .Z(n25875) );
  XNOR U27773 ( .A(n20454), .B(n25876), .Z(n25877) );
  NAND U27774 ( .A(n25878), .B(n[152]), .Z(n20454) );
  NAND U27775 ( .A(n21523), .B(n[152]), .Z(n25878) );
  XNOR U27776 ( .A(n25879), .B(n25876), .Z(n20455) );
  XOR U27777 ( .A(n25880), .B(n25881), .Z(n25876) );
  AND U27778 ( .A(n20462), .B(n25882), .Z(n25880) );
  XNOR U27779 ( .A(n20461), .B(n25881), .Z(n25882) );
  NAND U27780 ( .A(n25883), .B(n[151]), .Z(n20461) );
  NAND U27781 ( .A(n21523), .B(n[151]), .Z(n25883) );
  XNOR U27782 ( .A(n25884), .B(n25881), .Z(n20462) );
  XOR U27783 ( .A(n25885), .B(n25886), .Z(n25881) );
  AND U27784 ( .A(n20469), .B(n25887), .Z(n25885) );
  XNOR U27785 ( .A(n20468), .B(n25886), .Z(n25887) );
  NAND U27786 ( .A(n25888), .B(n[150]), .Z(n20468) );
  NAND U27787 ( .A(n21523), .B(n[150]), .Z(n25888) );
  XNOR U27788 ( .A(n25889), .B(n25886), .Z(n20469) );
  XOR U27789 ( .A(n25890), .B(n25891), .Z(n25886) );
  AND U27790 ( .A(n20476), .B(n25892), .Z(n25890) );
  XNOR U27791 ( .A(n20475), .B(n25891), .Z(n25892) );
  NAND U27792 ( .A(n25893), .B(n[149]), .Z(n20475) );
  NAND U27793 ( .A(n21523), .B(n[149]), .Z(n25893) );
  XNOR U27794 ( .A(n25894), .B(n25891), .Z(n20476) );
  XOR U27795 ( .A(n25895), .B(n25896), .Z(n25891) );
  AND U27796 ( .A(n20483), .B(n25897), .Z(n25895) );
  XNOR U27797 ( .A(n20482), .B(n25896), .Z(n25897) );
  NAND U27798 ( .A(n25898), .B(n[148]), .Z(n20482) );
  NAND U27799 ( .A(n21523), .B(n[148]), .Z(n25898) );
  XNOR U27800 ( .A(n25899), .B(n25896), .Z(n20483) );
  XOR U27801 ( .A(n25900), .B(n25901), .Z(n25896) );
  AND U27802 ( .A(n20490), .B(n25902), .Z(n25900) );
  XNOR U27803 ( .A(n20489), .B(n25901), .Z(n25902) );
  NAND U27804 ( .A(n25903), .B(n[147]), .Z(n20489) );
  NAND U27805 ( .A(n21523), .B(n[147]), .Z(n25903) );
  XNOR U27806 ( .A(n25904), .B(n25901), .Z(n20490) );
  XOR U27807 ( .A(n25905), .B(n25906), .Z(n25901) );
  AND U27808 ( .A(n20497), .B(n25907), .Z(n25905) );
  XNOR U27809 ( .A(n20496), .B(n25906), .Z(n25907) );
  NAND U27810 ( .A(n25908), .B(n[146]), .Z(n20496) );
  NAND U27811 ( .A(n21523), .B(n[146]), .Z(n25908) );
  XNOR U27812 ( .A(n25909), .B(n25906), .Z(n20497) );
  XOR U27813 ( .A(n25910), .B(n25911), .Z(n25906) );
  AND U27814 ( .A(n20504), .B(n25912), .Z(n25910) );
  XNOR U27815 ( .A(n20503), .B(n25911), .Z(n25912) );
  NAND U27816 ( .A(n25913), .B(n[145]), .Z(n20503) );
  NAND U27817 ( .A(n21523), .B(n[145]), .Z(n25913) );
  XNOR U27818 ( .A(n25914), .B(n25911), .Z(n20504) );
  XOR U27819 ( .A(n25915), .B(n25916), .Z(n25911) );
  AND U27820 ( .A(n20511), .B(n25917), .Z(n25915) );
  XNOR U27821 ( .A(n20510), .B(n25916), .Z(n25917) );
  NAND U27822 ( .A(n25918), .B(n[144]), .Z(n20510) );
  NAND U27823 ( .A(n21523), .B(n[144]), .Z(n25918) );
  XNOR U27824 ( .A(n25919), .B(n25916), .Z(n20511) );
  XOR U27825 ( .A(n25920), .B(n25921), .Z(n25916) );
  AND U27826 ( .A(n20518), .B(n25922), .Z(n25920) );
  XNOR U27827 ( .A(n20517), .B(n25921), .Z(n25922) );
  NAND U27828 ( .A(n25923), .B(n[143]), .Z(n20517) );
  NAND U27829 ( .A(n21523), .B(n[143]), .Z(n25923) );
  XNOR U27830 ( .A(n25924), .B(n25921), .Z(n20518) );
  XOR U27831 ( .A(n25925), .B(n25926), .Z(n25921) );
  AND U27832 ( .A(n20525), .B(n25927), .Z(n25925) );
  XNOR U27833 ( .A(n20524), .B(n25926), .Z(n25927) );
  NAND U27834 ( .A(n25928), .B(n[142]), .Z(n20524) );
  NAND U27835 ( .A(n21523), .B(n[142]), .Z(n25928) );
  XNOR U27836 ( .A(n25929), .B(n25926), .Z(n20525) );
  XOR U27837 ( .A(n25930), .B(n25931), .Z(n25926) );
  AND U27838 ( .A(n20532), .B(n25932), .Z(n25930) );
  XNOR U27839 ( .A(n20531), .B(n25931), .Z(n25932) );
  NAND U27840 ( .A(n25933), .B(n[141]), .Z(n20531) );
  NAND U27841 ( .A(n21523), .B(n[141]), .Z(n25933) );
  XNOR U27842 ( .A(n25934), .B(n25931), .Z(n20532) );
  XOR U27843 ( .A(n25935), .B(n25936), .Z(n25931) );
  AND U27844 ( .A(n20539), .B(n25937), .Z(n25935) );
  XNOR U27845 ( .A(n20538), .B(n25936), .Z(n25937) );
  NAND U27846 ( .A(n25938), .B(n[140]), .Z(n20538) );
  NAND U27847 ( .A(n21523), .B(n[140]), .Z(n25938) );
  XNOR U27848 ( .A(n25939), .B(n25936), .Z(n20539) );
  XOR U27849 ( .A(n25940), .B(n25941), .Z(n25936) );
  AND U27850 ( .A(n20546), .B(n25942), .Z(n25940) );
  XNOR U27851 ( .A(n20545), .B(n25941), .Z(n25942) );
  NAND U27852 ( .A(n25943), .B(n[139]), .Z(n20545) );
  NAND U27853 ( .A(n21523), .B(n[139]), .Z(n25943) );
  XNOR U27854 ( .A(n25944), .B(n25941), .Z(n20546) );
  XOR U27855 ( .A(n25945), .B(n25946), .Z(n25941) );
  AND U27856 ( .A(n20553), .B(n25947), .Z(n25945) );
  XNOR U27857 ( .A(n20552), .B(n25946), .Z(n25947) );
  NAND U27858 ( .A(n25948), .B(n[138]), .Z(n20552) );
  NAND U27859 ( .A(n21523), .B(n[138]), .Z(n25948) );
  XNOR U27860 ( .A(n25949), .B(n25946), .Z(n20553) );
  XOR U27861 ( .A(n25950), .B(n25951), .Z(n25946) );
  AND U27862 ( .A(n20560), .B(n25952), .Z(n25950) );
  XNOR U27863 ( .A(n20559), .B(n25951), .Z(n25952) );
  NAND U27864 ( .A(n25953), .B(n[137]), .Z(n20559) );
  NAND U27865 ( .A(n21523), .B(n[137]), .Z(n25953) );
  XNOR U27866 ( .A(n25954), .B(n25951), .Z(n20560) );
  XOR U27867 ( .A(n25955), .B(n25956), .Z(n25951) );
  AND U27868 ( .A(n20567), .B(n25957), .Z(n25955) );
  XNOR U27869 ( .A(n20566), .B(n25956), .Z(n25957) );
  NAND U27870 ( .A(n25958), .B(n[136]), .Z(n20566) );
  NAND U27871 ( .A(n21523), .B(n[136]), .Z(n25958) );
  XNOR U27872 ( .A(n25959), .B(n25956), .Z(n20567) );
  XOR U27873 ( .A(n25960), .B(n25961), .Z(n25956) );
  AND U27874 ( .A(n20574), .B(n25962), .Z(n25960) );
  XNOR U27875 ( .A(n20573), .B(n25961), .Z(n25962) );
  NAND U27876 ( .A(n25963), .B(n[135]), .Z(n20573) );
  NAND U27877 ( .A(n21523), .B(n[135]), .Z(n25963) );
  XNOR U27878 ( .A(n25964), .B(n25961), .Z(n20574) );
  XOR U27879 ( .A(n25965), .B(n25966), .Z(n25961) );
  AND U27880 ( .A(n20581), .B(n25967), .Z(n25965) );
  XNOR U27881 ( .A(n20580), .B(n25966), .Z(n25967) );
  NAND U27882 ( .A(n25968), .B(n[134]), .Z(n20580) );
  NAND U27883 ( .A(n21523), .B(n[134]), .Z(n25968) );
  XNOR U27884 ( .A(n25969), .B(n25966), .Z(n20581) );
  XOR U27885 ( .A(n25970), .B(n25971), .Z(n25966) );
  AND U27886 ( .A(n20588), .B(n25972), .Z(n25970) );
  XNOR U27887 ( .A(n20587), .B(n25971), .Z(n25972) );
  NAND U27888 ( .A(n25973), .B(n[133]), .Z(n20587) );
  NAND U27889 ( .A(n21523), .B(n[133]), .Z(n25973) );
  XNOR U27890 ( .A(n25974), .B(n25971), .Z(n20588) );
  XOR U27891 ( .A(n25975), .B(n25976), .Z(n25971) );
  AND U27892 ( .A(n20595), .B(n25977), .Z(n25975) );
  XNOR U27893 ( .A(n20594), .B(n25976), .Z(n25977) );
  NAND U27894 ( .A(n25978), .B(n[132]), .Z(n20594) );
  NAND U27895 ( .A(n21523), .B(n[132]), .Z(n25978) );
  XNOR U27896 ( .A(n25979), .B(n25976), .Z(n20595) );
  XOR U27897 ( .A(n25980), .B(n25981), .Z(n25976) );
  AND U27898 ( .A(n20602), .B(n25982), .Z(n25980) );
  XNOR U27899 ( .A(n20601), .B(n25981), .Z(n25982) );
  NAND U27900 ( .A(n25983), .B(n[131]), .Z(n20601) );
  NAND U27901 ( .A(n21523), .B(n[131]), .Z(n25983) );
  XNOR U27902 ( .A(n25984), .B(n25981), .Z(n20602) );
  XOR U27903 ( .A(n25985), .B(n25986), .Z(n25981) );
  AND U27904 ( .A(n20609), .B(n25987), .Z(n25985) );
  XNOR U27905 ( .A(n20608), .B(n25986), .Z(n25987) );
  NAND U27906 ( .A(n25988), .B(n[130]), .Z(n20608) );
  NAND U27907 ( .A(n21523), .B(n[130]), .Z(n25988) );
  XNOR U27908 ( .A(n25989), .B(n25986), .Z(n20609) );
  XOR U27909 ( .A(n25990), .B(n25991), .Z(n25986) );
  AND U27910 ( .A(n20616), .B(n25992), .Z(n25990) );
  XNOR U27911 ( .A(n20615), .B(n25991), .Z(n25992) );
  NAND U27912 ( .A(n25993), .B(n[129]), .Z(n20615) );
  NAND U27913 ( .A(n21523), .B(n[129]), .Z(n25993) );
  XNOR U27914 ( .A(n25994), .B(n25991), .Z(n20616) );
  XOR U27915 ( .A(n25995), .B(n25996), .Z(n25991) );
  AND U27916 ( .A(n20623), .B(n25997), .Z(n25995) );
  XNOR U27917 ( .A(n20622), .B(n25996), .Z(n25997) );
  NAND U27918 ( .A(n25998), .B(n[128]), .Z(n20622) );
  NAND U27919 ( .A(n21523), .B(n[128]), .Z(n25998) );
  XNOR U27920 ( .A(n25999), .B(n25996), .Z(n20623) );
  XOR U27921 ( .A(n26000), .B(n26001), .Z(n25996) );
  AND U27922 ( .A(n20630), .B(n26002), .Z(n26000) );
  XNOR U27923 ( .A(n20629), .B(n26001), .Z(n26002) );
  NAND U27924 ( .A(n26003), .B(n[127]), .Z(n20629) );
  NAND U27925 ( .A(n21523), .B(n[127]), .Z(n26003) );
  XNOR U27926 ( .A(n26004), .B(n26001), .Z(n20630) );
  XOR U27927 ( .A(n26005), .B(n26006), .Z(n26001) );
  AND U27928 ( .A(n20637), .B(n26007), .Z(n26005) );
  XNOR U27929 ( .A(n20636), .B(n26006), .Z(n26007) );
  NAND U27930 ( .A(n26008), .B(n[126]), .Z(n20636) );
  NAND U27931 ( .A(n21523), .B(n[126]), .Z(n26008) );
  XNOR U27932 ( .A(n26009), .B(n26006), .Z(n20637) );
  XOR U27933 ( .A(n26010), .B(n26011), .Z(n26006) );
  AND U27934 ( .A(n20644), .B(n26012), .Z(n26010) );
  XNOR U27935 ( .A(n20643), .B(n26011), .Z(n26012) );
  NAND U27936 ( .A(n26013), .B(n[125]), .Z(n20643) );
  NAND U27937 ( .A(n21523), .B(n[125]), .Z(n26013) );
  XNOR U27938 ( .A(n26014), .B(n26011), .Z(n20644) );
  XOR U27939 ( .A(n26015), .B(n26016), .Z(n26011) );
  AND U27940 ( .A(n20651), .B(n26017), .Z(n26015) );
  XNOR U27941 ( .A(n20650), .B(n26016), .Z(n26017) );
  NAND U27942 ( .A(n26018), .B(n[124]), .Z(n20650) );
  NAND U27943 ( .A(n21523), .B(n[124]), .Z(n26018) );
  XNOR U27944 ( .A(n26019), .B(n26016), .Z(n20651) );
  XOR U27945 ( .A(n26020), .B(n26021), .Z(n26016) );
  AND U27946 ( .A(n20658), .B(n26022), .Z(n26020) );
  XNOR U27947 ( .A(n20657), .B(n26021), .Z(n26022) );
  NAND U27948 ( .A(n26023), .B(n[123]), .Z(n20657) );
  NAND U27949 ( .A(n21523), .B(n[123]), .Z(n26023) );
  XNOR U27950 ( .A(n26024), .B(n26021), .Z(n20658) );
  XOR U27951 ( .A(n26025), .B(n26026), .Z(n26021) );
  AND U27952 ( .A(n20665), .B(n26027), .Z(n26025) );
  XNOR U27953 ( .A(n20664), .B(n26026), .Z(n26027) );
  NAND U27954 ( .A(n26028), .B(n[122]), .Z(n20664) );
  NAND U27955 ( .A(n21523), .B(n[122]), .Z(n26028) );
  XNOR U27956 ( .A(n26029), .B(n26026), .Z(n20665) );
  XOR U27957 ( .A(n26030), .B(n26031), .Z(n26026) );
  AND U27958 ( .A(n20672), .B(n26032), .Z(n26030) );
  XNOR U27959 ( .A(n20671), .B(n26031), .Z(n26032) );
  NAND U27960 ( .A(n26033), .B(n[121]), .Z(n20671) );
  NAND U27961 ( .A(n21523), .B(n[121]), .Z(n26033) );
  XNOR U27962 ( .A(n26034), .B(n26031), .Z(n20672) );
  XOR U27963 ( .A(n26035), .B(n26036), .Z(n26031) );
  AND U27964 ( .A(n20679), .B(n26037), .Z(n26035) );
  XNOR U27965 ( .A(n20678), .B(n26036), .Z(n26037) );
  NAND U27966 ( .A(n26038), .B(n[120]), .Z(n20678) );
  NAND U27967 ( .A(n21523), .B(n[120]), .Z(n26038) );
  XNOR U27968 ( .A(n26039), .B(n26036), .Z(n20679) );
  XOR U27969 ( .A(n26040), .B(n26041), .Z(n26036) );
  AND U27970 ( .A(n20686), .B(n26042), .Z(n26040) );
  XNOR U27971 ( .A(n20685), .B(n26041), .Z(n26042) );
  NAND U27972 ( .A(n26043), .B(n[119]), .Z(n20685) );
  NAND U27973 ( .A(n21523), .B(n[119]), .Z(n26043) );
  XNOR U27974 ( .A(n26044), .B(n26041), .Z(n20686) );
  XOR U27975 ( .A(n26045), .B(n26046), .Z(n26041) );
  AND U27976 ( .A(n20693), .B(n26047), .Z(n26045) );
  XNOR U27977 ( .A(n20692), .B(n26046), .Z(n26047) );
  NAND U27978 ( .A(n26048), .B(n[118]), .Z(n20692) );
  NAND U27979 ( .A(n21523), .B(n[118]), .Z(n26048) );
  XNOR U27980 ( .A(n26049), .B(n26046), .Z(n20693) );
  XOR U27981 ( .A(n26050), .B(n26051), .Z(n26046) );
  AND U27982 ( .A(n20700), .B(n26052), .Z(n26050) );
  XNOR U27983 ( .A(n20699), .B(n26051), .Z(n26052) );
  NAND U27984 ( .A(n26053), .B(n[117]), .Z(n20699) );
  NAND U27985 ( .A(n21523), .B(n[117]), .Z(n26053) );
  XNOR U27986 ( .A(n26054), .B(n26051), .Z(n20700) );
  XOR U27987 ( .A(n26055), .B(n26056), .Z(n26051) );
  AND U27988 ( .A(n20707), .B(n26057), .Z(n26055) );
  XNOR U27989 ( .A(n20706), .B(n26056), .Z(n26057) );
  NAND U27990 ( .A(n26058), .B(n[116]), .Z(n20706) );
  NAND U27991 ( .A(n21523), .B(n[116]), .Z(n26058) );
  XNOR U27992 ( .A(n26059), .B(n26056), .Z(n20707) );
  XOR U27993 ( .A(n26060), .B(n26061), .Z(n26056) );
  AND U27994 ( .A(n20714), .B(n26062), .Z(n26060) );
  XNOR U27995 ( .A(n20713), .B(n26061), .Z(n26062) );
  NAND U27996 ( .A(n26063), .B(n[115]), .Z(n20713) );
  NAND U27997 ( .A(n21523), .B(n[115]), .Z(n26063) );
  XNOR U27998 ( .A(n26064), .B(n26061), .Z(n20714) );
  XOR U27999 ( .A(n26065), .B(n26066), .Z(n26061) );
  AND U28000 ( .A(n20721), .B(n26067), .Z(n26065) );
  XNOR U28001 ( .A(n20720), .B(n26066), .Z(n26067) );
  NAND U28002 ( .A(n26068), .B(n[114]), .Z(n20720) );
  NAND U28003 ( .A(n21523), .B(n[114]), .Z(n26068) );
  XNOR U28004 ( .A(n26069), .B(n26066), .Z(n20721) );
  XOR U28005 ( .A(n26070), .B(n26071), .Z(n26066) );
  AND U28006 ( .A(n20728), .B(n26072), .Z(n26070) );
  XNOR U28007 ( .A(n20727), .B(n26071), .Z(n26072) );
  NAND U28008 ( .A(n26073), .B(n[113]), .Z(n20727) );
  NAND U28009 ( .A(n21523), .B(n[113]), .Z(n26073) );
  XNOR U28010 ( .A(n26074), .B(n26071), .Z(n20728) );
  XOR U28011 ( .A(n26075), .B(n26076), .Z(n26071) );
  AND U28012 ( .A(n20735), .B(n26077), .Z(n26075) );
  XNOR U28013 ( .A(n20734), .B(n26076), .Z(n26077) );
  NAND U28014 ( .A(n26078), .B(n[112]), .Z(n20734) );
  NAND U28015 ( .A(n21523), .B(n[112]), .Z(n26078) );
  XNOR U28016 ( .A(n26079), .B(n26076), .Z(n20735) );
  XOR U28017 ( .A(n26080), .B(n26081), .Z(n26076) );
  AND U28018 ( .A(n20742), .B(n26082), .Z(n26080) );
  XNOR U28019 ( .A(n20741), .B(n26081), .Z(n26082) );
  NAND U28020 ( .A(n26083), .B(n[111]), .Z(n20741) );
  NAND U28021 ( .A(n21523), .B(n[111]), .Z(n26083) );
  XNOR U28022 ( .A(n26084), .B(n26081), .Z(n20742) );
  XOR U28023 ( .A(n26085), .B(n26086), .Z(n26081) );
  AND U28024 ( .A(n20749), .B(n26087), .Z(n26085) );
  XNOR U28025 ( .A(n20748), .B(n26086), .Z(n26087) );
  NAND U28026 ( .A(n26088), .B(n[110]), .Z(n20748) );
  NAND U28027 ( .A(n21523), .B(n[110]), .Z(n26088) );
  XNOR U28028 ( .A(n26089), .B(n26086), .Z(n20749) );
  XOR U28029 ( .A(n26090), .B(n26091), .Z(n26086) );
  AND U28030 ( .A(n20756), .B(n26092), .Z(n26090) );
  XNOR U28031 ( .A(n20755), .B(n26091), .Z(n26092) );
  NAND U28032 ( .A(n26093), .B(n[109]), .Z(n20755) );
  NAND U28033 ( .A(n21523), .B(n[109]), .Z(n26093) );
  XNOR U28034 ( .A(n26094), .B(n26091), .Z(n20756) );
  XOR U28035 ( .A(n26095), .B(n26096), .Z(n26091) );
  AND U28036 ( .A(n20763), .B(n26097), .Z(n26095) );
  XNOR U28037 ( .A(n20762), .B(n26096), .Z(n26097) );
  NAND U28038 ( .A(n26098), .B(n[108]), .Z(n20762) );
  NAND U28039 ( .A(n21523), .B(n[108]), .Z(n26098) );
  XNOR U28040 ( .A(n26099), .B(n26096), .Z(n20763) );
  XOR U28041 ( .A(n26100), .B(n26101), .Z(n26096) );
  AND U28042 ( .A(n20770), .B(n26102), .Z(n26100) );
  XNOR U28043 ( .A(n20769), .B(n26101), .Z(n26102) );
  NAND U28044 ( .A(n26103), .B(n[107]), .Z(n20769) );
  NAND U28045 ( .A(n21523), .B(n[107]), .Z(n26103) );
  XNOR U28046 ( .A(n26104), .B(n26101), .Z(n20770) );
  XOR U28047 ( .A(n26105), .B(n26106), .Z(n26101) );
  AND U28048 ( .A(n20777), .B(n26107), .Z(n26105) );
  XNOR U28049 ( .A(n20776), .B(n26106), .Z(n26107) );
  NAND U28050 ( .A(n26108), .B(n[106]), .Z(n20776) );
  NAND U28051 ( .A(n21523), .B(n[106]), .Z(n26108) );
  XNOR U28052 ( .A(n26109), .B(n26106), .Z(n20777) );
  XOR U28053 ( .A(n26110), .B(n26111), .Z(n26106) );
  AND U28054 ( .A(n20784), .B(n26112), .Z(n26110) );
  XNOR U28055 ( .A(n20783), .B(n26111), .Z(n26112) );
  NAND U28056 ( .A(n26113), .B(n[105]), .Z(n20783) );
  NAND U28057 ( .A(n21523), .B(n[105]), .Z(n26113) );
  XNOR U28058 ( .A(n26114), .B(n26111), .Z(n20784) );
  XOR U28059 ( .A(n26115), .B(n26116), .Z(n26111) );
  AND U28060 ( .A(n20791), .B(n26117), .Z(n26115) );
  XNOR U28061 ( .A(n20790), .B(n26116), .Z(n26117) );
  NAND U28062 ( .A(n26118), .B(n[104]), .Z(n20790) );
  NAND U28063 ( .A(n21523), .B(n[104]), .Z(n26118) );
  XNOR U28064 ( .A(n26119), .B(n26116), .Z(n20791) );
  XOR U28065 ( .A(n26120), .B(n26121), .Z(n26116) );
  AND U28066 ( .A(n20798), .B(n26122), .Z(n26120) );
  XNOR U28067 ( .A(n20797), .B(n26121), .Z(n26122) );
  NAND U28068 ( .A(n26123), .B(n[103]), .Z(n20797) );
  NAND U28069 ( .A(n21523), .B(n[103]), .Z(n26123) );
  XNOR U28070 ( .A(n26124), .B(n26121), .Z(n20798) );
  XOR U28071 ( .A(n26125), .B(n26126), .Z(n26121) );
  AND U28072 ( .A(n20805), .B(n26127), .Z(n26125) );
  XNOR U28073 ( .A(n20804), .B(n26126), .Z(n26127) );
  NAND U28074 ( .A(n26128), .B(n[102]), .Z(n20804) );
  NAND U28075 ( .A(n21523), .B(n[102]), .Z(n26128) );
  XNOR U28076 ( .A(n26129), .B(n26126), .Z(n20805) );
  XOR U28077 ( .A(n26130), .B(n26131), .Z(n26126) );
  AND U28078 ( .A(n20812), .B(n26132), .Z(n26130) );
  XNOR U28079 ( .A(n20811), .B(n26131), .Z(n26132) );
  NAND U28080 ( .A(n26133), .B(n[101]), .Z(n20811) );
  NAND U28081 ( .A(n21523), .B(n[101]), .Z(n26133) );
  XNOR U28082 ( .A(n26134), .B(n26131), .Z(n20812) );
  XOR U28083 ( .A(n26135), .B(n26136), .Z(n26131) );
  AND U28084 ( .A(n20819), .B(n26137), .Z(n26135) );
  XNOR U28085 ( .A(n20818), .B(n26136), .Z(n26137) );
  NAND U28086 ( .A(n26138), .B(n[100]), .Z(n20818) );
  NAND U28087 ( .A(n21523), .B(n[100]), .Z(n26138) );
  XNOR U28088 ( .A(n26139), .B(n26136), .Z(n20819) );
  XOR U28089 ( .A(n26140), .B(n26141), .Z(n26136) );
  AND U28090 ( .A(n20826), .B(n26142), .Z(n26140) );
  XNOR U28091 ( .A(n20825), .B(n26141), .Z(n26142) );
  NAND U28092 ( .A(n26143), .B(n[99]), .Z(n20825) );
  NAND U28093 ( .A(n21523), .B(n[99]), .Z(n26143) );
  XNOR U28094 ( .A(n26144), .B(n26141), .Z(n20826) );
  XOR U28095 ( .A(n26145), .B(n26146), .Z(n26141) );
  AND U28096 ( .A(n20833), .B(n26147), .Z(n26145) );
  XNOR U28097 ( .A(n20832), .B(n26146), .Z(n26147) );
  NAND U28098 ( .A(n26148), .B(n[98]), .Z(n20832) );
  NAND U28099 ( .A(n21523), .B(n[98]), .Z(n26148) );
  XNOR U28100 ( .A(n26149), .B(n26146), .Z(n20833) );
  XOR U28101 ( .A(n26150), .B(n26151), .Z(n26146) );
  AND U28102 ( .A(n20840), .B(n26152), .Z(n26150) );
  XNOR U28103 ( .A(n20839), .B(n26151), .Z(n26152) );
  NAND U28104 ( .A(n26153), .B(n[97]), .Z(n20839) );
  NAND U28105 ( .A(n21523), .B(n[97]), .Z(n26153) );
  XNOR U28106 ( .A(n26154), .B(n26151), .Z(n20840) );
  XOR U28107 ( .A(n26155), .B(n26156), .Z(n26151) );
  AND U28108 ( .A(n20847), .B(n26157), .Z(n26155) );
  XNOR U28109 ( .A(n20846), .B(n26156), .Z(n26157) );
  NAND U28110 ( .A(n26158), .B(n[96]), .Z(n20846) );
  NAND U28111 ( .A(n21523), .B(n[96]), .Z(n26158) );
  XNOR U28112 ( .A(n26159), .B(n26156), .Z(n20847) );
  XOR U28113 ( .A(n26160), .B(n26161), .Z(n26156) );
  AND U28114 ( .A(n20854), .B(n26162), .Z(n26160) );
  XNOR U28115 ( .A(n20853), .B(n26161), .Z(n26162) );
  NAND U28116 ( .A(n26163), .B(n[95]), .Z(n20853) );
  NAND U28117 ( .A(n21523), .B(n[95]), .Z(n26163) );
  XNOR U28118 ( .A(n26164), .B(n26161), .Z(n20854) );
  XOR U28119 ( .A(n26165), .B(n26166), .Z(n26161) );
  AND U28120 ( .A(n20861), .B(n26167), .Z(n26165) );
  XNOR U28121 ( .A(n20860), .B(n26166), .Z(n26167) );
  NAND U28122 ( .A(n26168), .B(n[94]), .Z(n20860) );
  NAND U28123 ( .A(n21523), .B(n[94]), .Z(n26168) );
  XNOR U28124 ( .A(n26169), .B(n26166), .Z(n20861) );
  XOR U28125 ( .A(n26170), .B(n26171), .Z(n26166) );
  AND U28126 ( .A(n20868), .B(n26172), .Z(n26170) );
  XNOR U28127 ( .A(n20867), .B(n26171), .Z(n26172) );
  NAND U28128 ( .A(n26173), .B(n[93]), .Z(n20867) );
  NAND U28129 ( .A(n21523), .B(n[93]), .Z(n26173) );
  XNOR U28130 ( .A(n26174), .B(n26171), .Z(n20868) );
  XOR U28131 ( .A(n26175), .B(n26176), .Z(n26171) );
  AND U28132 ( .A(n20875), .B(n26177), .Z(n26175) );
  XNOR U28133 ( .A(n20874), .B(n26176), .Z(n26177) );
  NAND U28134 ( .A(n26178), .B(n[92]), .Z(n20874) );
  NAND U28135 ( .A(n21523), .B(n[92]), .Z(n26178) );
  XNOR U28136 ( .A(n26179), .B(n26176), .Z(n20875) );
  XOR U28137 ( .A(n26180), .B(n26181), .Z(n26176) );
  AND U28138 ( .A(n20882), .B(n26182), .Z(n26180) );
  XNOR U28139 ( .A(n20881), .B(n26181), .Z(n26182) );
  NAND U28140 ( .A(n26183), .B(n[91]), .Z(n20881) );
  NAND U28141 ( .A(n21523), .B(n[91]), .Z(n26183) );
  XNOR U28142 ( .A(n26184), .B(n26181), .Z(n20882) );
  XOR U28143 ( .A(n26185), .B(n26186), .Z(n26181) );
  AND U28144 ( .A(n20889), .B(n26187), .Z(n26185) );
  XNOR U28145 ( .A(n20888), .B(n26186), .Z(n26187) );
  NAND U28146 ( .A(n26188), .B(n[90]), .Z(n20888) );
  NAND U28147 ( .A(n21523), .B(n[90]), .Z(n26188) );
  XNOR U28148 ( .A(n26189), .B(n26186), .Z(n20889) );
  XOR U28149 ( .A(n26190), .B(n26191), .Z(n26186) );
  AND U28150 ( .A(n20896), .B(n26192), .Z(n26190) );
  XNOR U28151 ( .A(n20895), .B(n26191), .Z(n26192) );
  NAND U28152 ( .A(n26193), .B(n[89]), .Z(n20895) );
  NAND U28153 ( .A(n21523), .B(n[89]), .Z(n26193) );
  XNOR U28154 ( .A(n26194), .B(n26191), .Z(n20896) );
  XOR U28155 ( .A(n26195), .B(n26196), .Z(n26191) );
  AND U28156 ( .A(n20903), .B(n26197), .Z(n26195) );
  XNOR U28157 ( .A(n20902), .B(n26196), .Z(n26197) );
  NAND U28158 ( .A(n26198), .B(n[88]), .Z(n20902) );
  NAND U28159 ( .A(n21523), .B(n[88]), .Z(n26198) );
  XNOR U28160 ( .A(n26199), .B(n26196), .Z(n20903) );
  XOR U28161 ( .A(n26200), .B(n26201), .Z(n26196) );
  AND U28162 ( .A(n20910), .B(n26202), .Z(n26200) );
  XNOR U28163 ( .A(n20909), .B(n26201), .Z(n26202) );
  NAND U28164 ( .A(n26203), .B(n[87]), .Z(n20909) );
  NAND U28165 ( .A(n21523), .B(n[87]), .Z(n26203) );
  XNOR U28166 ( .A(n26204), .B(n26201), .Z(n20910) );
  XOR U28167 ( .A(n26205), .B(n26206), .Z(n26201) );
  AND U28168 ( .A(n20917), .B(n26207), .Z(n26205) );
  XNOR U28169 ( .A(n20916), .B(n26206), .Z(n26207) );
  NAND U28170 ( .A(n26208), .B(n[86]), .Z(n20916) );
  NAND U28171 ( .A(n21523), .B(n[86]), .Z(n26208) );
  XNOR U28172 ( .A(n26209), .B(n26206), .Z(n20917) );
  XOR U28173 ( .A(n26210), .B(n26211), .Z(n26206) );
  AND U28174 ( .A(n20924), .B(n26212), .Z(n26210) );
  XNOR U28175 ( .A(n20923), .B(n26211), .Z(n26212) );
  NAND U28176 ( .A(n26213), .B(n[85]), .Z(n20923) );
  NAND U28177 ( .A(n21523), .B(n[85]), .Z(n26213) );
  XNOR U28178 ( .A(n26214), .B(n26211), .Z(n20924) );
  XOR U28179 ( .A(n26215), .B(n26216), .Z(n26211) );
  AND U28180 ( .A(n20931), .B(n26217), .Z(n26215) );
  XNOR U28181 ( .A(n20930), .B(n26216), .Z(n26217) );
  NAND U28182 ( .A(n26218), .B(n[84]), .Z(n20930) );
  NAND U28183 ( .A(n21523), .B(n[84]), .Z(n26218) );
  XNOR U28184 ( .A(n26219), .B(n26216), .Z(n20931) );
  XOR U28185 ( .A(n26220), .B(n26221), .Z(n26216) );
  AND U28186 ( .A(n20938), .B(n26222), .Z(n26220) );
  XNOR U28187 ( .A(n20937), .B(n26221), .Z(n26222) );
  NAND U28188 ( .A(n26223), .B(n[83]), .Z(n20937) );
  NAND U28189 ( .A(n21523), .B(n[83]), .Z(n26223) );
  XNOR U28190 ( .A(n26224), .B(n26221), .Z(n20938) );
  XOR U28191 ( .A(n26225), .B(n26226), .Z(n26221) );
  AND U28192 ( .A(n20945), .B(n26227), .Z(n26225) );
  XNOR U28193 ( .A(n20944), .B(n26226), .Z(n26227) );
  NAND U28194 ( .A(n26228), .B(n[82]), .Z(n20944) );
  NAND U28195 ( .A(n21523), .B(n[82]), .Z(n26228) );
  XNOR U28196 ( .A(n26229), .B(n26226), .Z(n20945) );
  XOR U28197 ( .A(n26230), .B(n26231), .Z(n26226) );
  AND U28198 ( .A(n20952), .B(n26232), .Z(n26230) );
  XNOR U28199 ( .A(n20951), .B(n26231), .Z(n26232) );
  NAND U28200 ( .A(n26233), .B(n[81]), .Z(n20951) );
  NAND U28201 ( .A(n21523), .B(n[81]), .Z(n26233) );
  XNOR U28202 ( .A(n26234), .B(n26231), .Z(n20952) );
  XOR U28203 ( .A(n26235), .B(n26236), .Z(n26231) );
  AND U28204 ( .A(n20959), .B(n26237), .Z(n26235) );
  XNOR U28205 ( .A(n20958), .B(n26236), .Z(n26237) );
  NAND U28206 ( .A(n26238), .B(n[80]), .Z(n20958) );
  NAND U28207 ( .A(n21523), .B(n[80]), .Z(n26238) );
  XNOR U28208 ( .A(n26239), .B(n26236), .Z(n20959) );
  XOR U28209 ( .A(n26240), .B(n26241), .Z(n26236) );
  AND U28210 ( .A(n20966), .B(n26242), .Z(n26240) );
  XNOR U28211 ( .A(n20965), .B(n26241), .Z(n26242) );
  NAND U28212 ( .A(n26243), .B(n[79]), .Z(n20965) );
  NAND U28213 ( .A(n21523), .B(n[79]), .Z(n26243) );
  XNOR U28214 ( .A(n26244), .B(n26241), .Z(n20966) );
  XOR U28215 ( .A(n26245), .B(n26246), .Z(n26241) );
  AND U28216 ( .A(n20973), .B(n26247), .Z(n26245) );
  XNOR U28217 ( .A(n20972), .B(n26246), .Z(n26247) );
  NAND U28218 ( .A(n26248), .B(n[78]), .Z(n20972) );
  NAND U28219 ( .A(n21523), .B(n[78]), .Z(n26248) );
  XNOR U28220 ( .A(n26249), .B(n26246), .Z(n20973) );
  XOR U28221 ( .A(n26250), .B(n26251), .Z(n26246) );
  AND U28222 ( .A(n20980), .B(n26252), .Z(n26250) );
  XNOR U28223 ( .A(n20979), .B(n26251), .Z(n26252) );
  NAND U28224 ( .A(n26253), .B(n[77]), .Z(n20979) );
  NAND U28225 ( .A(n21523), .B(n[77]), .Z(n26253) );
  XNOR U28226 ( .A(n26254), .B(n26251), .Z(n20980) );
  XOR U28227 ( .A(n26255), .B(n26256), .Z(n26251) );
  AND U28228 ( .A(n20987), .B(n26257), .Z(n26255) );
  XNOR U28229 ( .A(n20986), .B(n26256), .Z(n26257) );
  NAND U28230 ( .A(n26258), .B(n[76]), .Z(n20986) );
  NAND U28231 ( .A(n21523), .B(n[76]), .Z(n26258) );
  XNOR U28232 ( .A(n26259), .B(n26256), .Z(n20987) );
  XOR U28233 ( .A(n26260), .B(n26261), .Z(n26256) );
  AND U28234 ( .A(n20994), .B(n26262), .Z(n26260) );
  XNOR U28235 ( .A(n20993), .B(n26261), .Z(n26262) );
  NAND U28236 ( .A(n26263), .B(n[75]), .Z(n20993) );
  NAND U28237 ( .A(n21523), .B(n[75]), .Z(n26263) );
  XNOR U28238 ( .A(n26264), .B(n26261), .Z(n20994) );
  XOR U28239 ( .A(n26265), .B(n26266), .Z(n26261) );
  AND U28240 ( .A(n21001), .B(n26267), .Z(n26265) );
  XNOR U28241 ( .A(n21000), .B(n26266), .Z(n26267) );
  NAND U28242 ( .A(n26268), .B(n[74]), .Z(n21000) );
  NAND U28243 ( .A(n21523), .B(n[74]), .Z(n26268) );
  XNOR U28244 ( .A(n26269), .B(n26266), .Z(n21001) );
  XOR U28245 ( .A(n26270), .B(n26271), .Z(n26266) );
  AND U28246 ( .A(n21008), .B(n26272), .Z(n26270) );
  XNOR U28247 ( .A(n21007), .B(n26271), .Z(n26272) );
  NAND U28248 ( .A(n26273), .B(n[73]), .Z(n21007) );
  NAND U28249 ( .A(n21523), .B(n[73]), .Z(n26273) );
  XNOR U28250 ( .A(n26274), .B(n26271), .Z(n21008) );
  XOR U28251 ( .A(n26275), .B(n26276), .Z(n26271) );
  AND U28252 ( .A(n21015), .B(n26277), .Z(n26275) );
  XNOR U28253 ( .A(n21014), .B(n26276), .Z(n26277) );
  NAND U28254 ( .A(n26278), .B(n[72]), .Z(n21014) );
  NAND U28255 ( .A(n21523), .B(n[72]), .Z(n26278) );
  XNOR U28256 ( .A(n26279), .B(n26276), .Z(n21015) );
  XOR U28257 ( .A(n26280), .B(n26281), .Z(n26276) );
  AND U28258 ( .A(n21022), .B(n26282), .Z(n26280) );
  XNOR U28259 ( .A(n21021), .B(n26281), .Z(n26282) );
  NAND U28260 ( .A(n26283), .B(n[71]), .Z(n21021) );
  NAND U28261 ( .A(n21523), .B(n[71]), .Z(n26283) );
  XNOR U28262 ( .A(n26284), .B(n26281), .Z(n21022) );
  XOR U28263 ( .A(n26285), .B(n26286), .Z(n26281) );
  AND U28264 ( .A(n21029), .B(n26287), .Z(n26285) );
  XNOR U28265 ( .A(n21028), .B(n26286), .Z(n26287) );
  NAND U28266 ( .A(n26288), .B(n[70]), .Z(n21028) );
  NAND U28267 ( .A(n21523), .B(n[70]), .Z(n26288) );
  XNOR U28268 ( .A(n26289), .B(n26286), .Z(n21029) );
  XOR U28269 ( .A(n26290), .B(n26291), .Z(n26286) );
  AND U28270 ( .A(n21036), .B(n26292), .Z(n26290) );
  XNOR U28271 ( .A(n21035), .B(n26291), .Z(n26292) );
  NAND U28272 ( .A(n26293), .B(n[69]), .Z(n21035) );
  NAND U28273 ( .A(n21523), .B(n[69]), .Z(n26293) );
  XNOR U28274 ( .A(n26294), .B(n26291), .Z(n21036) );
  XOR U28275 ( .A(n26295), .B(n26296), .Z(n26291) );
  AND U28276 ( .A(n21043), .B(n26297), .Z(n26295) );
  XNOR U28277 ( .A(n21042), .B(n26296), .Z(n26297) );
  NAND U28278 ( .A(n26298), .B(n[68]), .Z(n21042) );
  NAND U28279 ( .A(n21523), .B(n[68]), .Z(n26298) );
  XNOR U28280 ( .A(n26299), .B(n26296), .Z(n21043) );
  XOR U28281 ( .A(n26300), .B(n26301), .Z(n26296) );
  AND U28282 ( .A(n21050), .B(n26302), .Z(n26300) );
  XNOR U28283 ( .A(n21049), .B(n26301), .Z(n26302) );
  NAND U28284 ( .A(n26303), .B(n[67]), .Z(n21049) );
  NAND U28285 ( .A(n21523), .B(n[67]), .Z(n26303) );
  XNOR U28286 ( .A(n26304), .B(n26301), .Z(n21050) );
  XOR U28287 ( .A(n26305), .B(n26306), .Z(n26301) );
  AND U28288 ( .A(n21057), .B(n26307), .Z(n26305) );
  XNOR U28289 ( .A(n21056), .B(n26306), .Z(n26307) );
  NAND U28290 ( .A(n26308), .B(n[66]), .Z(n21056) );
  NAND U28291 ( .A(n21523), .B(n[66]), .Z(n26308) );
  XNOR U28292 ( .A(n26309), .B(n26306), .Z(n21057) );
  XOR U28293 ( .A(n26310), .B(n26311), .Z(n26306) );
  AND U28294 ( .A(n21064), .B(n26312), .Z(n26310) );
  XNOR U28295 ( .A(n21063), .B(n26311), .Z(n26312) );
  NAND U28296 ( .A(n26313), .B(n[65]), .Z(n21063) );
  NAND U28297 ( .A(n21523), .B(n[65]), .Z(n26313) );
  XNOR U28298 ( .A(n26314), .B(n26311), .Z(n21064) );
  XOR U28299 ( .A(n26315), .B(n26316), .Z(n26311) );
  AND U28300 ( .A(n21071), .B(n26317), .Z(n26315) );
  XNOR U28301 ( .A(n21070), .B(n26316), .Z(n26317) );
  NAND U28302 ( .A(n26318), .B(n[64]), .Z(n21070) );
  NAND U28303 ( .A(n21523), .B(n[64]), .Z(n26318) );
  XNOR U28304 ( .A(n26319), .B(n26316), .Z(n21071) );
  XOR U28305 ( .A(n26320), .B(n26321), .Z(n26316) );
  AND U28306 ( .A(n21078), .B(n26322), .Z(n26320) );
  XNOR U28307 ( .A(n21077), .B(n26321), .Z(n26322) );
  NAND U28308 ( .A(n26323), .B(n[63]), .Z(n21077) );
  NAND U28309 ( .A(n21523), .B(n[63]), .Z(n26323) );
  XNOR U28310 ( .A(n26324), .B(n26321), .Z(n21078) );
  XOR U28311 ( .A(n26325), .B(n26326), .Z(n26321) );
  AND U28312 ( .A(n21085), .B(n26327), .Z(n26325) );
  XNOR U28313 ( .A(n21084), .B(n26326), .Z(n26327) );
  NAND U28314 ( .A(n26328), .B(n[62]), .Z(n21084) );
  NAND U28315 ( .A(n21523), .B(n[62]), .Z(n26328) );
  XNOR U28316 ( .A(n26329), .B(n26326), .Z(n21085) );
  XOR U28317 ( .A(n26330), .B(n26331), .Z(n26326) );
  AND U28318 ( .A(n21092), .B(n26332), .Z(n26330) );
  XNOR U28319 ( .A(n21091), .B(n26331), .Z(n26332) );
  NAND U28320 ( .A(n26333), .B(n[61]), .Z(n21091) );
  NAND U28321 ( .A(n21523), .B(n[61]), .Z(n26333) );
  XNOR U28322 ( .A(n26334), .B(n26331), .Z(n21092) );
  XOR U28323 ( .A(n26335), .B(n26336), .Z(n26331) );
  AND U28324 ( .A(n21099), .B(n26337), .Z(n26335) );
  XNOR U28325 ( .A(n21098), .B(n26336), .Z(n26337) );
  NAND U28326 ( .A(n26338), .B(n[60]), .Z(n21098) );
  NAND U28327 ( .A(n21523), .B(n[60]), .Z(n26338) );
  XNOR U28328 ( .A(n26339), .B(n26336), .Z(n21099) );
  XOR U28329 ( .A(n26340), .B(n26341), .Z(n26336) );
  AND U28330 ( .A(n21106), .B(n26342), .Z(n26340) );
  XNOR U28331 ( .A(n21105), .B(n26341), .Z(n26342) );
  NAND U28332 ( .A(n26343), .B(n[59]), .Z(n21105) );
  NAND U28333 ( .A(n21523), .B(n[59]), .Z(n26343) );
  XNOR U28334 ( .A(n26344), .B(n26341), .Z(n21106) );
  XOR U28335 ( .A(n26345), .B(n26346), .Z(n26341) );
  AND U28336 ( .A(n21113), .B(n26347), .Z(n26345) );
  XNOR U28337 ( .A(n21112), .B(n26346), .Z(n26347) );
  NAND U28338 ( .A(n26348), .B(n[58]), .Z(n21112) );
  NAND U28339 ( .A(n21523), .B(n[58]), .Z(n26348) );
  XNOR U28340 ( .A(n26349), .B(n26346), .Z(n21113) );
  XOR U28341 ( .A(n26350), .B(n26351), .Z(n26346) );
  AND U28342 ( .A(n21120), .B(n26352), .Z(n26350) );
  XNOR U28343 ( .A(n21119), .B(n26351), .Z(n26352) );
  NAND U28344 ( .A(n26353), .B(n[57]), .Z(n21119) );
  NAND U28345 ( .A(n21523), .B(n[57]), .Z(n26353) );
  XNOR U28346 ( .A(n26354), .B(n26351), .Z(n21120) );
  XOR U28347 ( .A(n26355), .B(n26356), .Z(n26351) );
  AND U28348 ( .A(n21127), .B(n26357), .Z(n26355) );
  XNOR U28349 ( .A(n21126), .B(n26356), .Z(n26357) );
  NAND U28350 ( .A(n26358), .B(n[56]), .Z(n21126) );
  NAND U28351 ( .A(n21523), .B(n[56]), .Z(n26358) );
  XNOR U28352 ( .A(n26359), .B(n26356), .Z(n21127) );
  XOR U28353 ( .A(n26360), .B(n26361), .Z(n26356) );
  AND U28354 ( .A(n21134), .B(n26362), .Z(n26360) );
  XNOR U28355 ( .A(n21133), .B(n26361), .Z(n26362) );
  NAND U28356 ( .A(n26363), .B(n[55]), .Z(n21133) );
  NAND U28357 ( .A(n21523), .B(n[55]), .Z(n26363) );
  XNOR U28358 ( .A(n26364), .B(n26361), .Z(n21134) );
  XOR U28359 ( .A(n26365), .B(n26366), .Z(n26361) );
  AND U28360 ( .A(n21141), .B(n26367), .Z(n26365) );
  XNOR U28361 ( .A(n21140), .B(n26366), .Z(n26367) );
  NAND U28362 ( .A(n26368), .B(n[54]), .Z(n21140) );
  NAND U28363 ( .A(n21523), .B(n[54]), .Z(n26368) );
  XNOR U28364 ( .A(n26369), .B(n26366), .Z(n21141) );
  XOR U28365 ( .A(n26370), .B(n26371), .Z(n26366) );
  AND U28366 ( .A(n21148), .B(n26372), .Z(n26370) );
  XNOR U28367 ( .A(n21147), .B(n26371), .Z(n26372) );
  NAND U28368 ( .A(n26373), .B(n[53]), .Z(n21147) );
  NAND U28369 ( .A(n21523), .B(n[53]), .Z(n26373) );
  XNOR U28370 ( .A(n26374), .B(n26371), .Z(n21148) );
  XOR U28371 ( .A(n26375), .B(n26376), .Z(n26371) );
  AND U28372 ( .A(n21155), .B(n26377), .Z(n26375) );
  XNOR U28373 ( .A(n21154), .B(n26376), .Z(n26377) );
  NAND U28374 ( .A(n26378), .B(n[52]), .Z(n21154) );
  NAND U28375 ( .A(n21523), .B(n[52]), .Z(n26378) );
  XNOR U28376 ( .A(n26379), .B(n26376), .Z(n21155) );
  XOR U28377 ( .A(n26380), .B(n26381), .Z(n26376) );
  AND U28378 ( .A(n21162), .B(n26382), .Z(n26380) );
  XNOR U28379 ( .A(n21161), .B(n26381), .Z(n26382) );
  NAND U28380 ( .A(n26383), .B(n[51]), .Z(n21161) );
  NAND U28381 ( .A(n21523), .B(n[51]), .Z(n26383) );
  XNOR U28382 ( .A(n26384), .B(n26381), .Z(n21162) );
  XOR U28383 ( .A(n26385), .B(n26386), .Z(n26381) );
  AND U28384 ( .A(n21169), .B(n26387), .Z(n26385) );
  XNOR U28385 ( .A(n21168), .B(n26386), .Z(n26387) );
  NAND U28386 ( .A(n26388), .B(n[50]), .Z(n21168) );
  NAND U28387 ( .A(n21523), .B(n[50]), .Z(n26388) );
  XNOR U28388 ( .A(n26389), .B(n26386), .Z(n21169) );
  XOR U28389 ( .A(n26390), .B(n26391), .Z(n26386) );
  AND U28390 ( .A(n21176), .B(n26392), .Z(n26390) );
  XNOR U28391 ( .A(n21175), .B(n26391), .Z(n26392) );
  NAND U28392 ( .A(n26393), .B(n[49]), .Z(n21175) );
  NAND U28393 ( .A(n21523), .B(n[49]), .Z(n26393) );
  XNOR U28394 ( .A(n26394), .B(n26391), .Z(n21176) );
  XOR U28395 ( .A(n26395), .B(n26396), .Z(n26391) );
  AND U28396 ( .A(n21183), .B(n26397), .Z(n26395) );
  XNOR U28397 ( .A(n21182), .B(n26396), .Z(n26397) );
  NAND U28398 ( .A(n26398), .B(n[48]), .Z(n21182) );
  NAND U28399 ( .A(n21523), .B(n[48]), .Z(n26398) );
  XNOR U28400 ( .A(n26399), .B(n26396), .Z(n21183) );
  XOR U28401 ( .A(n26400), .B(n26401), .Z(n26396) );
  AND U28402 ( .A(n21190), .B(n26402), .Z(n26400) );
  XNOR U28403 ( .A(n21189), .B(n26401), .Z(n26402) );
  NAND U28404 ( .A(n26403), .B(n[47]), .Z(n21189) );
  NAND U28405 ( .A(n21523), .B(n[47]), .Z(n26403) );
  XNOR U28406 ( .A(n26404), .B(n26401), .Z(n21190) );
  XOR U28407 ( .A(n26405), .B(n26406), .Z(n26401) );
  AND U28408 ( .A(n21197), .B(n26407), .Z(n26405) );
  XNOR U28409 ( .A(n21196), .B(n26406), .Z(n26407) );
  NAND U28410 ( .A(n26408), .B(n[46]), .Z(n21196) );
  NAND U28411 ( .A(n21523), .B(n[46]), .Z(n26408) );
  XNOR U28412 ( .A(n26409), .B(n26406), .Z(n21197) );
  XOR U28413 ( .A(n26410), .B(n26411), .Z(n26406) );
  AND U28414 ( .A(n21204), .B(n26412), .Z(n26410) );
  XNOR U28415 ( .A(n21203), .B(n26411), .Z(n26412) );
  NAND U28416 ( .A(n26413), .B(n[45]), .Z(n21203) );
  NAND U28417 ( .A(n21523), .B(n[45]), .Z(n26413) );
  XNOR U28418 ( .A(n26414), .B(n26411), .Z(n21204) );
  XOR U28419 ( .A(n26415), .B(n26416), .Z(n26411) );
  AND U28420 ( .A(n21211), .B(n26417), .Z(n26415) );
  XNOR U28421 ( .A(n21210), .B(n26416), .Z(n26417) );
  NAND U28422 ( .A(n26418), .B(n[44]), .Z(n21210) );
  NAND U28423 ( .A(n21523), .B(n[44]), .Z(n26418) );
  XNOR U28424 ( .A(n26419), .B(n26416), .Z(n21211) );
  XOR U28425 ( .A(n26420), .B(n26421), .Z(n26416) );
  AND U28426 ( .A(n21218), .B(n26422), .Z(n26420) );
  XNOR U28427 ( .A(n21217), .B(n26421), .Z(n26422) );
  NAND U28428 ( .A(n26423), .B(n[43]), .Z(n21217) );
  NAND U28429 ( .A(n21523), .B(n[43]), .Z(n26423) );
  XNOR U28430 ( .A(n26424), .B(n26421), .Z(n21218) );
  XOR U28431 ( .A(n26425), .B(n26426), .Z(n26421) );
  AND U28432 ( .A(n21225), .B(n26427), .Z(n26425) );
  XNOR U28433 ( .A(n21224), .B(n26426), .Z(n26427) );
  NAND U28434 ( .A(n26428), .B(n[42]), .Z(n21224) );
  NAND U28435 ( .A(n21523), .B(n[42]), .Z(n26428) );
  XNOR U28436 ( .A(n26429), .B(n26426), .Z(n21225) );
  XOR U28437 ( .A(n26430), .B(n26431), .Z(n26426) );
  AND U28438 ( .A(n21232), .B(n26432), .Z(n26430) );
  XNOR U28439 ( .A(n21231), .B(n26431), .Z(n26432) );
  NAND U28440 ( .A(n26433), .B(n[41]), .Z(n21231) );
  NAND U28441 ( .A(n21523), .B(n[41]), .Z(n26433) );
  XNOR U28442 ( .A(n26434), .B(n26431), .Z(n21232) );
  XOR U28443 ( .A(n26435), .B(n26436), .Z(n26431) );
  AND U28444 ( .A(n21239), .B(n26437), .Z(n26435) );
  XNOR U28445 ( .A(n21238), .B(n26436), .Z(n26437) );
  NAND U28446 ( .A(n26438), .B(n[40]), .Z(n21238) );
  NAND U28447 ( .A(n21523), .B(n[40]), .Z(n26438) );
  XNOR U28448 ( .A(n26439), .B(n26436), .Z(n21239) );
  XOR U28449 ( .A(n26440), .B(n26441), .Z(n26436) );
  AND U28450 ( .A(n21246), .B(n26442), .Z(n26440) );
  XNOR U28451 ( .A(n21245), .B(n26441), .Z(n26442) );
  NAND U28452 ( .A(n26443), .B(n[39]), .Z(n21245) );
  NAND U28453 ( .A(n21523), .B(n[39]), .Z(n26443) );
  XNOR U28454 ( .A(n26444), .B(n26441), .Z(n21246) );
  XOR U28455 ( .A(n26445), .B(n26446), .Z(n26441) );
  AND U28456 ( .A(n21253), .B(n26447), .Z(n26445) );
  XNOR U28457 ( .A(n21252), .B(n26446), .Z(n26447) );
  NAND U28458 ( .A(n26448), .B(n[38]), .Z(n21252) );
  NAND U28459 ( .A(n21523), .B(n[38]), .Z(n26448) );
  XNOR U28460 ( .A(n26449), .B(n26446), .Z(n21253) );
  XOR U28461 ( .A(n26450), .B(n26451), .Z(n26446) );
  AND U28462 ( .A(n21260), .B(n26452), .Z(n26450) );
  XNOR U28463 ( .A(n21259), .B(n26451), .Z(n26452) );
  NAND U28464 ( .A(n26453), .B(n[37]), .Z(n21259) );
  NAND U28465 ( .A(n21523), .B(n[37]), .Z(n26453) );
  XNOR U28466 ( .A(n26454), .B(n26451), .Z(n21260) );
  XOR U28467 ( .A(n26455), .B(n26456), .Z(n26451) );
  AND U28468 ( .A(n21267), .B(n26457), .Z(n26455) );
  XNOR U28469 ( .A(n21266), .B(n26456), .Z(n26457) );
  NAND U28470 ( .A(n26458), .B(n[36]), .Z(n21266) );
  NAND U28471 ( .A(n21523), .B(n[36]), .Z(n26458) );
  XNOR U28472 ( .A(n26459), .B(n26456), .Z(n21267) );
  XOR U28473 ( .A(n26460), .B(n26461), .Z(n26456) );
  AND U28474 ( .A(n21274), .B(n26462), .Z(n26460) );
  XNOR U28475 ( .A(n21273), .B(n26461), .Z(n26462) );
  NAND U28476 ( .A(n26463), .B(n[35]), .Z(n21273) );
  NAND U28477 ( .A(n21523), .B(n[35]), .Z(n26463) );
  XNOR U28478 ( .A(n26464), .B(n26461), .Z(n21274) );
  XOR U28479 ( .A(n26465), .B(n26466), .Z(n26461) );
  AND U28480 ( .A(n21281), .B(n26467), .Z(n26465) );
  XNOR U28481 ( .A(n21280), .B(n26466), .Z(n26467) );
  NAND U28482 ( .A(n26468), .B(n[34]), .Z(n21280) );
  NAND U28483 ( .A(n21523), .B(n[34]), .Z(n26468) );
  XNOR U28484 ( .A(n26469), .B(n26466), .Z(n21281) );
  XOR U28485 ( .A(n26470), .B(n26471), .Z(n26466) );
  AND U28486 ( .A(n21288), .B(n26472), .Z(n26470) );
  XNOR U28487 ( .A(n21287), .B(n26471), .Z(n26472) );
  NAND U28488 ( .A(n26473), .B(n[33]), .Z(n21287) );
  NAND U28489 ( .A(n21523), .B(n[33]), .Z(n26473) );
  XNOR U28490 ( .A(n26474), .B(n26471), .Z(n21288) );
  XOR U28491 ( .A(n26475), .B(n26476), .Z(n26471) );
  AND U28492 ( .A(n21295), .B(n26477), .Z(n26475) );
  XNOR U28493 ( .A(n21294), .B(n26476), .Z(n26477) );
  NAND U28494 ( .A(n26478), .B(n[32]), .Z(n21294) );
  NAND U28495 ( .A(n21523), .B(n[32]), .Z(n26478) );
  XNOR U28496 ( .A(n26479), .B(n26476), .Z(n21295) );
  XOR U28497 ( .A(n26480), .B(n26481), .Z(n26476) );
  AND U28498 ( .A(n21302), .B(n26482), .Z(n26480) );
  XNOR U28499 ( .A(n21301), .B(n26481), .Z(n26482) );
  NAND U28500 ( .A(n26483), .B(n[31]), .Z(n21301) );
  NAND U28501 ( .A(n21523), .B(n[31]), .Z(n26483) );
  XNOR U28502 ( .A(n26484), .B(n26481), .Z(n21302) );
  XOR U28503 ( .A(n26485), .B(n26486), .Z(n26481) );
  AND U28504 ( .A(n21309), .B(n26487), .Z(n26485) );
  XNOR U28505 ( .A(n21308), .B(n26486), .Z(n26487) );
  NAND U28506 ( .A(n26488), .B(n[30]), .Z(n21308) );
  NAND U28507 ( .A(n21523), .B(n[30]), .Z(n26488) );
  XNOR U28508 ( .A(n26489), .B(n26486), .Z(n21309) );
  XOR U28509 ( .A(n26490), .B(n26491), .Z(n26486) );
  AND U28510 ( .A(n21316), .B(n26492), .Z(n26490) );
  XNOR U28511 ( .A(n21315), .B(n26491), .Z(n26492) );
  NAND U28512 ( .A(n26493), .B(n[29]), .Z(n21315) );
  NAND U28513 ( .A(n21523), .B(n[29]), .Z(n26493) );
  XNOR U28514 ( .A(n26494), .B(n26491), .Z(n21316) );
  XOR U28515 ( .A(n26495), .B(n26496), .Z(n26491) );
  AND U28516 ( .A(n21323), .B(n26497), .Z(n26495) );
  XNOR U28517 ( .A(n21322), .B(n26496), .Z(n26497) );
  NAND U28518 ( .A(n26498), .B(n[28]), .Z(n21322) );
  NAND U28519 ( .A(n21523), .B(n[28]), .Z(n26498) );
  XNOR U28520 ( .A(n26499), .B(n26496), .Z(n21323) );
  XOR U28521 ( .A(n26500), .B(n26501), .Z(n26496) );
  AND U28522 ( .A(n21330), .B(n26502), .Z(n26500) );
  XNOR U28523 ( .A(n21329), .B(n26501), .Z(n26502) );
  NAND U28524 ( .A(n26503), .B(n[27]), .Z(n21329) );
  NAND U28525 ( .A(n21523), .B(n[27]), .Z(n26503) );
  XNOR U28526 ( .A(n26504), .B(n26501), .Z(n21330) );
  XOR U28527 ( .A(n26505), .B(n26506), .Z(n26501) );
  AND U28528 ( .A(n21337), .B(n26507), .Z(n26505) );
  XNOR U28529 ( .A(n21336), .B(n26506), .Z(n26507) );
  NAND U28530 ( .A(n26508), .B(n[26]), .Z(n21336) );
  NAND U28531 ( .A(n21523), .B(n[26]), .Z(n26508) );
  XNOR U28532 ( .A(n26509), .B(n26506), .Z(n21337) );
  XOR U28533 ( .A(n26510), .B(n26511), .Z(n26506) );
  AND U28534 ( .A(n21344), .B(n26512), .Z(n26510) );
  XNOR U28535 ( .A(n21343), .B(n26511), .Z(n26512) );
  NAND U28536 ( .A(n26513), .B(n[25]), .Z(n21343) );
  NAND U28537 ( .A(n21523), .B(n[25]), .Z(n26513) );
  XNOR U28538 ( .A(n26514), .B(n26511), .Z(n21344) );
  XOR U28539 ( .A(n26515), .B(n26516), .Z(n26511) );
  AND U28540 ( .A(n21351), .B(n26517), .Z(n26515) );
  XNOR U28541 ( .A(n21350), .B(n26516), .Z(n26517) );
  NAND U28542 ( .A(n26518), .B(n[24]), .Z(n21350) );
  NAND U28543 ( .A(n21523), .B(n[24]), .Z(n26518) );
  XNOR U28544 ( .A(n26519), .B(n26516), .Z(n21351) );
  XOR U28545 ( .A(n26520), .B(n26521), .Z(n26516) );
  AND U28546 ( .A(n21358), .B(n26522), .Z(n26520) );
  XNOR U28547 ( .A(n21357), .B(n26521), .Z(n26522) );
  NAND U28548 ( .A(n26523), .B(n[23]), .Z(n21357) );
  NAND U28549 ( .A(n21523), .B(n[23]), .Z(n26523) );
  XNOR U28550 ( .A(n26524), .B(n26521), .Z(n21358) );
  XOR U28551 ( .A(n26525), .B(n26526), .Z(n26521) );
  AND U28552 ( .A(n21365), .B(n26527), .Z(n26525) );
  XNOR U28553 ( .A(n21364), .B(n26526), .Z(n26527) );
  NAND U28554 ( .A(n26528), .B(n[22]), .Z(n21364) );
  NAND U28555 ( .A(n21523), .B(n[22]), .Z(n26528) );
  XNOR U28556 ( .A(n26529), .B(n26526), .Z(n21365) );
  XOR U28557 ( .A(n26530), .B(n26531), .Z(n26526) );
  AND U28558 ( .A(n21372), .B(n26532), .Z(n26530) );
  XNOR U28559 ( .A(n21371), .B(n26531), .Z(n26532) );
  NAND U28560 ( .A(n26533), .B(n[21]), .Z(n21371) );
  NAND U28561 ( .A(n21523), .B(n[21]), .Z(n26533) );
  XNOR U28562 ( .A(n26534), .B(n26531), .Z(n21372) );
  XOR U28563 ( .A(n26535), .B(n26536), .Z(n26531) );
  AND U28564 ( .A(n21379), .B(n26537), .Z(n26535) );
  XNOR U28565 ( .A(n21378), .B(n26536), .Z(n26537) );
  NAND U28566 ( .A(n26538), .B(n[20]), .Z(n21378) );
  NAND U28567 ( .A(n21523), .B(n[20]), .Z(n26538) );
  XNOR U28568 ( .A(n26539), .B(n26536), .Z(n21379) );
  XOR U28569 ( .A(n26540), .B(n26541), .Z(n26536) );
  AND U28570 ( .A(n21386), .B(n26542), .Z(n26540) );
  XNOR U28571 ( .A(n21385), .B(n26541), .Z(n26542) );
  NAND U28572 ( .A(n26543), .B(n[19]), .Z(n21385) );
  NAND U28573 ( .A(n21523), .B(n[19]), .Z(n26543) );
  XNOR U28574 ( .A(n26544), .B(n26541), .Z(n21386) );
  XOR U28575 ( .A(n26545), .B(n26546), .Z(n26541) );
  AND U28576 ( .A(n21393), .B(n26547), .Z(n26545) );
  XNOR U28577 ( .A(n21392), .B(n26546), .Z(n26547) );
  NAND U28578 ( .A(n26548), .B(n[18]), .Z(n21392) );
  NAND U28579 ( .A(n21523), .B(n[18]), .Z(n26548) );
  XNOR U28580 ( .A(n26549), .B(n26546), .Z(n21393) );
  XOR U28581 ( .A(n26550), .B(n26551), .Z(n26546) );
  AND U28582 ( .A(n21400), .B(n26552), .Z(n26550) );
  XNOR U28583 ( .A(n21399), .B(n26551), .Z(n26552) );
  NAND U28584 ( .A(n26553), .B(n[17]), .Z(n21399) );
  NAND U28585 ( .A(n21523), .B(n[17]), .Z(n26553) );
  XNOR U28586 ( .A(n26554), .B(n26551), .Z(n21400) );
  XOR U28587 ( .A(n26555), .B(n26556), .Z(n26551) );
  AND U28588 ( .A(n21407), .B(n26557), .Z(n26555) );
  XNOR U28589 ( .A(n21406), .B(n26556), .Z(n26557) );
  NAND U28590 ( .A(n26558), .B(n[16]), .Z(n21406) );
  NAND U28591 ( .A(n21523), .B(n[16]), .Z(n26558) );
  XNOR U28592 ( .A(n26559), .B(n26556), .Z(n21407) );
  XOR U28593 ( .A(n26560), .B(n26561), .Z(n26556) );
  AND U28594 ( .A(n21414), .B(n26562), .Z(n26560) );
  XNOR U28595 ( .A(n21413), .B(n26561), .Z(n26562) );
  NAND U28596 ( .A(n26563), .B(n[15]), .Z(n21413) );
  NAND U28597 ( .A(n21523), .B(n[15]), .Z(n26563) );
  XNOR U28598 ( .A(n26564), .B(n26561), .Z(n21414) );
  XOR U28599 ( .A(n26565), .B(n26566), .Z(n26561) );
  AND U28600 ( .A(n21421), .B(n26567), .Z(n26565) );
  XNOR U28601 ( .A(n21420), .B(n26566), .Z(n26567) );
  NAND U28602 ( .A(n26568), .B(n[14]), .Z(n21420) );
  NAND U28603 ( .A(n21523), .B(n[14]), .Z(n26568) );
  XNOR U28604 ( .A(n26569), .B(n26566), .Z(n21421) );
  XOR U28605 ( .A(n26570), .B(n26571), .Z(n26566) );
  AND U28606 ( .A(n21428), .B(n26572), .Z(n26570) );
  XNOR U28607 ( .A(n21427), .B(n26571), .Z(n26572) );
  NAND U28608 ( .A(n26573), .B(n[13]), .Z(n21427) );
  NAND U28609 ( .A(n21523), .B(n[13]), .Z(n26573) );
  XNOR U28610 ( .A(n26574), .B(n26571), .Z(n21428) );
  XOR U28611 ( .A(n26575), .B(n26576), .Z(n26571) );
  AND U28612 ( .A(n21435), .B(n26577), .Z(n26575) );
  XNOR U28613 ( .A(n21434), .B(n26576), .Z(n26577) );
  NAND U28614 ( .A(n26578), .B(n[12]), .Z(n21434) );
  NAND U28615 ( .A(n21523), .B(n[12]), .Z(n26578) );
  XNOR U28616 ( .A(n26579), .B(n26576), .Z(n21435) );
  XOR U28617 ( .A(n26580), .B(n26581), .Z(n26576) );
  AND U28618 ( .A(n21442), .B(n26582), .Z(n26580) );
  XNOR U28619 ( .A(n21441), .B(n26581), .Z(n26582) );
  NAND U28620 ( .A(n26583), .B(n[11]), .Z(n21441) );
  NAND U28621 ( .A(n21523), .B(n[11]), .Z(n26583) );
  XNOR U28622 ( .A(n26584), .B(n26581), .Z(n21442) );
  XOR U28623 ( .A(n26585), .B(n26586), .Z(n26581) );
  AND U28624 ( .A(n21449), .B(n26587), .Z(n26585) );
  XNOR U28625 ( .A(n21448), .B(n26586), .Z(n26587) );
  NAND U28626 ( .A(n26588), .B(n[10]), .Z(n21448) );
  NAND U28627 ( .A(n21523), .B(n[10]), .Z(n26588) );
  XNOR U28628 ( .A(n26589), .B(n26586), .Z(n21449) );
  XOR U28629 ( .A(n26590), .B(n26591), .Z(n26586) );
  AND U28630 ( .A(n21456), .B(n26592), .Z(n26590) );
  XNOR U28631 ( .A(n21455), .B(n26591), .Z(n26592) );
  NAND U28632 ( .A(n26593), .B(n[9]), .Z(n21455) );
  NAND U28633 ( .A(n21523), .B(n[9]), .Z(n26593) );
  XNOR U28634 ( .A(n26594), .B(n26591), .Z(n21456) );
  XOR U28635 ( .A(n26595), .B(n26596), .Z(n26591) );
  AND U28636 ( .A(n21463), .B(n26597), .Z(n26595) );
  XNOR U28637 ( .A(n21462), .B(n26596), .Z(n26597) );
  NAND U28638 ( .A(n26598), .B(n[8]), .Z(n21462) );
  NAND U28639 ( .A(n21523), .B(n[8]), .Z(n26598) );
  XNOR U28640 ( .A(n26599), .B(n26596), .Z(n21463) );
  XOR U28641 ( .A(n26600), .B(n26601), .Z(n26596) );
  AND U28642 ( .A(n21470), .B(n26602), .Z(n26600) );
  XNOR U28643 ( .A(n21469), .B(n26601), .Z(n26602) );
  NAND U28644 ( .A(n26603), .B(n[7]), .Z(n21469) );
  NAND U28645 ( .A(n21523), .B(n[7]), .Z(n26603) );
  XNOR U28646 ( .A(n26604), .B(n26601), .Z(n21470) );
  XOR U28647 ( .A(n26605), .B(n26606), .Z(n26601) );
  AND U28648 ( .A(n21477), .B(n26607), .Z(n26605) );
  XNOR U28649 ( .A(n21476), .B(n26606), .Z(n26607) );
  NAND U28650 ( .A(n26608), .B(n[6]), .Z(n21476) );
  NAND U28651 ( .A(n21523), .B(n[6]), .Z(n26608) );
  XNOR U28652 ( .A(n26609), .B(n26606), .Z(n21477) );
  XOR U28653 ( .A(n26610), .B(n26611), .Z(n26606) );
  AND U28654 ( .A(n21484), .B(n26612), .Z(n26610) );
  XNOR U28655 ( .A(n21483), .B(n26611), .Z(n26612) );
  NAND U28656 ( .A(n26613), .B(n[5]), .Z(n21483) );
  NAND U28657 ( .A(n21523), .B(n[5]), .Z(n26613) );
  XNOR U28658 ( .A(n26614), .B(n26611), .Z(n21484) );
  XOR U28659 ( .A(n26615), .B(n26616), .Z(n26611) );
  AND U28660 ( .A(n21491), .B(n26617), .Z(n26615) );
  XNOR U28661 ( .A(n21490), .B(n26616), .Z(n26617) );
  NAND U28662 ( .A(n26618), .B(n[4]), .Z(n21490) );
  NAND U28663 ( .A(n21523), .B(n[4]), .Z(n26618) );
  XNOR U28664 ( .A(n26619), .B(n26616), .Z(n21491) );
  XOR U28665 ( .A(n26620), .B(n26621), .Z(n26616) );
  AND U28666 ( .A(n21498), .B(n26622), .Z(n26620) );
  XNOR U28667 ( .A(n21497), .B(n26621), .Z(n26622) );
  NAND U28668 ( .A(n26623), .B(n[3]), .Z(n21497) );
  NAND U28669 ( .A(n21523), .B(n[3]), .Z(n26623) );
  XNOR U28670 ( .A(n26624), .B(n26621), .Z(n21498) );
  XOR U28671 ( .A(n26625), .B(n26626), .Z(n26621) );
  AND U28672 ( .A(n21505), .B(n26627), .Z(n26625) );
  XNOR U28673 ( .A(n21504), .B(n26626), .Z(n26627) );
  NAND U28674 ( .A(n26628), .B(n[2]), .Z(n21504) );
  NAND U28675 ( .A(n21523), .B(n[2]), .Z(n26628) );
  XOR U28676 ( .A(n26629), .B(n26626), .Z(n21505) );
  XNOR U28677 ( .A(n26630), .B(n26631), .Z(n26626) );
  NANDN U28678 ( .A(n21511), .B(n26632), .Z(n26631) );
  XNOR U28679 ( .A(n26630), .B(n21510), .Z(n26632) );
  NAND U28680 ( .A(n26633), .B(n[1]), .Z(n21510) );
  NAND U28681 ( .A(n21523), .B(n[1]), .Z(n26633) );
  XOR U28682 ( .A(n26630), .B(n26634), .Z(n21511) );
  NOR U28683 ( .A(n21514), .B(n21512), .Z(n26630) );
  NAND U28684 ( .A(n26635), .B(n[0]), .Z(n21512) );
  NAND U28685 ( .A(n21523), .B(n[0]), .Z(n26635) );
  NAND U28686 ( .A(n26636), .B(n26637), .Z(n21523) );
  NAND U28687 ( .A(n26638), .B(n26637), .Z(n26636) );
  XOR U28688 ( .A(n26637), .B(n21516), .Z(n26638) );
  XNOR U28689 ( .A(n26639), .B(n26640), .Z(n21516) );
  XOR U28690 ( .A(\modmult_1/zin[0][1024] ), .B(n26641), .Z(n26640) );
  NANDN U28691 ( .A(n26639), .B(n21518), .Z(n26641) );
  AND U28692 ( .A(n26642), .B(n26643), .Z(n26637) );
  NAND U28693 ( .A(n26644), .B(n26643), .Z(n26642) );
  XNOR U28694 ( .A(n26643), .B(n21518), .Z(n26644) );
  XOR U28695 ( .A(\modmult_1/zin[0][1023] ), .B(n26645), .Z(n21518) );
  IV U28696 ( .A(n26639), .Z(n26645) );
  XOR U28697 ( .A(n26646), .B(n26647), .Z(n26639) );
  ANDN U28698 ( .B(n26648), .A(n26649), .Z(n26646) );
  XOR U28699 ( .A(n26647), .B(n26650), .Z(n26648) );
  XOR U28700 ( .A(n26651), .B(n26652), .Z(n26643) );
  AND U28701 ( .A(n26653), .B(n26654), .Z(n26651) );
  XOR U28702 ( .A(n[1023]), .B(n26652), .Z(n26654) );
  XNOR U28703 ( .A(n26652), .B(n21524), .Z(n26653) );
  XOR U28704 ( .A(n26655), .B(n26656), .Z(n26652) );
  AND U28705 ( .A(n26657), .B(n26658), .Z(n26655) );
  XOR U28706 ( .A(n[1022]), .B(n26656), .Z(n26658) );
  XNOR U28707 ( .A(n26656), .B(n21529), .Z(n26657) );
  XOR U28708 ( .A(n26659), .B(n26660), .Z(n26656) );
  AND U28709 ( .A(n26661), .B(n26662), .Z(n26659) );
  XOR U28710 ( .A(n[1021]), .B(n26660), .Z(n26662) );
  XNOR U28711 ( .A(n26660), .B(n21534), .Z(n26661) );
  XOR U28712 ( .A(n26663), .B(n26664), .Z(n26660) );
  AND U28713 ( .A(n26665), .B(n26666), .Z(n26663) );
  XOR U28714 ( .A(n[1020]), .B(n26664), .Z(n26666) );
  XNOR U28715 ( .A(n26664), .B(n21539), .Z(n26665) );
  XOR U28716 ( .A(n26667), .B(n26668), .Z(n26664) );
  AND U28717 ( .A(n26669), .B(n26670), .Z(n26667) );
  XOR U28718 ( .A(n[1019]), .B(n26668), .Z(n26670) );
  XNOR U28719 ( .A(n26668), .B(n21544), .Z(n26669) );
  XOR U28720 ( .A(n26671), .B(n26672), .Z(n26668) );
  AND U28721 ( .A(n26673), .B(n26674), .Z(n26671) );
  XOR U28722 ( .A(n[1018]), .B(n26672), .Z(n26674) );
  XNOR U28723 ( .A(n26672), .B(n21549), .Z(n26673) );
  XOR U28724 ( .A(n26675), .B(n26676), .Z(n26672) );
  AND U28725 ( .A(n26677), .B(n26678), .Z(n26675) );
  XOR U28726 ( .A(n[1017]), .B(n26676), .Z(n26678) );
  XNOR U28727 ( .A(n26676), .B(n21554), .Z(n26677) );
  XOR U28728 ( .A(n26679), .B(n26680), .Z(n26676) );
  AND U28729 ( .A(n26681), .B(n26682), .Z(n26679) );
  XOR U28730 ( .A(n[1016]), .B(n26680), .Z(n26682) );
  XNOR U28731 ( .A(n26680), .B(n21559), .Z(n26681) );
  XOR U28732 ( .A(n26683), .B(n26684), .Z(n26680) );
  AND U28733 ( .A(n26685), .B(n26686), .Z(n26683) );
  XOR U28734 ( .A(n[1015]), .B(n26684), .Z(n26686) );
  XNOR U28735 ( .A(n26684), .B(n21564), .Z(n26685) );
  XOR U28736 ( .A(n26687), .B(n26688), .Z(n26684) );
  AND U28737 ( .A(n26689), .B(n26690), .Z(n26687) );
  XOR U28738 ( .A(n[1014]), .B(n26688), .Z(n26690) );
  XNOR U28739 ( .A(n26688), .B(n21569), .Z(n26689) );
  XOR U28740 ( .A(n26691), .B(n26692), .Z(n26688) );
  AND U28741 ( .A(n26693), .B(n26694), .Z(n26691) );
  XOR U28742 ( .A(n[1013]), .B(n26692), .Z(n26694) );
  XNOR U28743 ( .A(n26692), .B(n21574), .Z(n26693) );
  XOR U28744 ( .A(n26695), .B(n26696), .Z(n26692) );
  AND U28745 ( .A(n26697), .B(n26698), .Z(n26695) );
  XOR U28746 ( .A(n[1012]), .B(n26696), .Z(n26698) );
  XNOR U28747 ( .A(n26696), .B(n21579), .Z(n26697) );
  XOR U28748 ( .A(n26699), .B(n26700), .Z(n26696) );
  AND U28749 ( .A(n26701), .B(n26702), .Z(n26699) );
  XOR U28750 ( .A(n[1011]), .B(n26700), .Z(n26702) );
  XNOR U28751 ( .A(n26700), .B(n21584), .Z(n26701) );
  XOR U28752 ( .A(n26703), .B(n26704), .Z(n26700) );
  AND U28753 ( .A(n26705), .B(n26706), .Z(n26703) );
  XOR U28754 ( .A(n[1010]), .B(n26704), .Z(n26706) );
  XNOR U28755 ( .A(n26704), .B(n21589), .Z(n26705) );
  XOR U28756 ( .A(n26707), .B(n26708), .Z(n26704) );
  AND U28757 ( .A(n26709), .B(n26710), .Z(n26707) );
  XOR U28758 ( .A(n[1009]), .B(n26708), .Z(n26710) );
  XNOR U28759 ( .A(n26708), .B(n21594), .Z(n26709) );
  XOR U28760 ( .A(n26711), .B(n26712), .Z(n26708) );
  AND U28761 ( .A(n26713), .B(n26714), .Z(n26711) );
  XOR U28762 ( .A(n[1008]), .B(n26712), .Z(n26714) );
  XNOR U28763 ( .A(n26712), .B(n21599), .Z(n26713) );
  XOR U28764 ( .A(n26715), .B(n26716), .Z(n26712) );
  AND U28765 ( .A(n26717), .B(n26718), .Z(n26715) );
  XOR U28766 ( .A(n[1007]), .B(n26716), .Z(n26718) );
  XNOR U28767 ( .A(n26716), .B(n21604), .Z(n26717) );
  XOR U28768 ( .A(n26719), .B(n26720), .Z(n26716) );
  AND U28769 ( .A(n26721), .B(n26722), .Z(n26719) );
  XOR U28770 ( .A(n[1006]), .B(n26720), .Z(n26722) );
  XNOR U28771 ( .A(n26720), .B(n21609), .Z(n26721) );
  XOR U28772 ( .A(n26723), .B(n26724), .Z(n26720) );
  AND U28773 ( .A(n26725), .B(n26726), .Z(n26723) );
  XOR U28774 ( .A(n[1005]), .B(n26724), .Z(n26726) );
  XNOR U28775 ( .A(n26724), .B(n21614), .Z(n26725) );
  XOR U28776 ( .A(n26727), .B(n26728), .Z(n26724) );
  AND U28777 ( .A(n26729), .B(n26730), .Z(n26727) );
  XOR U28778 ( .A(n[1004]), .B(n26728), .Z(n26730) );
  XNOR U28779 ( .A(n26728), .B(n21619), .Z(n26729) );
  XOR U28780 ( .A(n26731), .B(n26732), .Z(n26728) );
  AND U28781 ( .A(n26733), .B(n26734), .Z(n26731) );
  XOR U28782 ( .A(n[1003]), .B(n26732), .Z(n26734) );
  XNOR U28783 ( .A(n26732), .B(n21624), .Z(n26733) );
  XOR U28784 ( .A(n26735), .B(n26736), .Z(n26732) );
  AND U28785 ( .A(n26737), .B(n26738), .Z(n26735) );
  XOR U28786 ( .A(n[1002]), .B(n26736), .Z(n26738) );
  XNOR U28787 ( .A(n26736), .B(n21629), .Z(n26737) );
  XOR U28788 ( .A(n26739), .B(n26740), .Z(n26736) );
  AND U28789 ( .A(n26741), .B(n26742), .Z(n26739) );
  XOR U28790 ( .A(n[1001]), .B(n26740), .Z(n26742) );
  XNOR U28791 ( .A(n26740), .B(n21634), .Z(n26741) );
  XOR U28792 ( .A(n26743), .B(n26744), .Z(n26740) );
  AND U28793 ( .A(n26745), .B(n26746), .Z(n26743) );
  XOR U28794 ( .A(n[1000]), .B(n26744), .Z(n26746) );
  XNOR U28795 ( .A(n26744), .B(n21639), .Z(n26745) );
  XOR U28796 ( .A(n26747), .B(n26748), .Z(n26744) );
  AND U28797 ( .A(n26749), .B(n26750), .Z(n26747) );
  XOR U28798 ( .A(n[999]), .B(n26748), .Z(n26750) );
  XNOR U28799 ( .A(n26748), .B(n21644), .Z(n26749) );
  XOR U28800 ( .A(n26751), .B(n26752), .Z(n26748) );
  AND U28801 ( .A(n26753), .B(n26754), .Z(n26751) );
  XOR U28802 ( .A(n[998]), .B(n26752), .Z(n26754) );
  XNOR U28803 ( .A(n26752), .B(n21649), .Z(n26753) );
  XOR U28804 ( .A(n26755), .B(n26756), .Z(n26752) );
  AND U28805 ( .A(n26757), .B(n26758), .Z(n26755) );
  XOR U28806 ( .A(n[997]), .B(n26756), .Z(n26758) );
  XNOR U28807 ( .A(n26756), .B(n21654), .Z(n26757) );
  XOR U28808 ( .A(n26759), .B(n26760), .Z(n26756) );
  AND U28809 ( .A(n26761), .B(n26762), .Z(n26759) );
  XOR U28810 ( .A(n[996]), .B(n26760), .Z(n26762) );
  XNOR U28811 ( .A(n26760), .B(n21659), .Z(n26761) );
  XOR U28812 ( .A(n26763), .B(n26764), .Z(n26760) );
  AND U28813 ( .A(n26765), .B(n26766), .Z(n26763) );
  XOR U28814 ( .A(n[995]), .B(n26764), .Z(n26766) );
  XNOR U28815 ( .A(n26764), .B(n21664), .Z(n26765) );
  XOR U28816 ( .A(n26767), .B(n26768), .Z(n26764) );
  AND U28817 ( .A(n26769), .B(n26770), .Z(n26767) );
  XOR U28818 ( .A(n[994]), .B(n26768), .Z(n26770) );
  XNOR U28819 ( .A(n26768), .B(n21669), .Z(n26769) );
  XOR U28820 ( .A(n26771), .B(n26772), .Z(n26768) );
  AND U28821 ( .A(n26773), .B(n26774), .Z(n26771) );
  XOR U28822 ( .A(n[993]), .B(n26772), .Z(n26774) );
  XNOR U28823 ( .A(n26772), .B(n21674), .Z(n26773) );
  XOR U28824 ( .A(n26775), .B(n26776), .Z(n26772) );
  AND U28825 ( .A(n26777), .B(n26778), .Z(n26775) );
  XOR U28826 ( .A(n[992]), .B(n26776), .Z(n26778) );
  XNOR U28827 ( .A(n26776), .B(n21679), .Z(n26777) );
  XOR U28828 ( .A(n26779), .B(n26780), .Z(n26776) );
  AND U28829 ( .A(n26781), .B(n26782), .Z(n26779) );
  XOR U28830 ( .A(n[991]), .B(n26780), .Z(n26782) );
  XNOR U28831 ( .A(n26780), .B(n21684), .Z(n26781) );
  XOR U28832 ( .A(n26783), .B(n26784), .Z(n26780) );
  AND U28833 ( .A(n26785), .B(n26786), .Z(n26783) );
  XOR U28834 ( .A(n[990]), .B(n26784), .Z(n26786) );
  XNOR U28835 ( .A(n26784), .B(n21689), .Z(n26785) );
  XOR U28836 ( .A(n26787), .B(n26788), .Z(n26784) );
  AND U28837 ( .A(n26789), .B(n26790), .Z(n26787) );
  XOR U28838 ( .A(n[989]), .B(n26788), .Z(n26790) );
  XNOR U28839 ( .A(n26788), .B(n21694), .Z(n26789) );
  XOR U28840 ( .A(n26791), .B(n26792), .Z(n26788) );
  AND U28841 ( .A(n26793), .B(n26794), .Z(n26791) );
  XOR U28842 ( .A(n[988]), .B(n26792), .Z(n26794) );
  XNOR U28843 ( .A(n26792), .B(n21699), .Z(n26793) );
  XOR U28844 ( .A(n26795), .B(n26796), .Z(n26792) );
  AND U28845 ( .A(n26797), .B(n26798), .Z(n26795) );
  XOR U28846 ( .A(n[987]), .B(n26796), .Z(n26798) );
  XNOR U28847 ( .A(n26796), .B(n21704), .Z(n26797) );
  XOR U28848 ( .A(n26799), .B(n26800), .Z(n26796) );
  AND U28849 ( .A(n26801), .B(n26802), .Z(n26799) );
  XOR U28850 ( .A(n[986]), .B(n26800), .Z(n26802) );
  XNOR U28851 ( .A(n26800), .B(n21709), .Z(n26801) );
  XOR U28852 ( .A(n26803), .B(n26804), .Z(n26800) );
  AND U28853 ( .A(n26805), .B(n26806), .Z(n26803) );
  XOR U28854 ( .A(n[985]), .B(n26804), .Z(n26806) );
  XNOR U28855 ( .A(n26804), .B(n21714), .Z(n26805) );
  XOR U28856 ( .A(n26807), .B(n26808), .Z(n26804) );
  AND U28857 ( .A(n26809), .B(n26810), .Z(n26807) );
  XOR U28858 ( .A(n[984]), .B(n26808), .Z(n26810) );
  XNOR U28859 ( .A(n26808), .B(n21719), .Z(n26809) );
  XOR U28860 ( .A(n26811), .B(n26812), .Z(n26808) );
  AND U28861 ( .A(n26813), .B(n26814), .Z(n26811) );
  XOR U28862 ( .A(n[983]), .B(n26812), .Z(n26814) );
  XNOR U28863 ( .A(n26812), .B(n21724), .Z(n26813) );
  XOR U28864 ( .A(n26815), .B(n26816), .Z(n26812) );
  AND U28865 ( .A(n26817), .B(n26818), .Z(n26815) );
  XOR U28866 ( .A(n[982]), .B(n26816), .Z(n26818) );
  XNOR U28867 ( .A(n26816), .B(n21729), .Z(n26817) );
  XOR U28868 ( .A(n26819), .B(n26820), .Z(n26816) );
  AND U28869 ( .A(n26821), .B(n26822), .Z(n26819) );
  XOR U28870 ( .A(n[981]), .B(n26820), .Z(n26822) );
  XNOR U28871 ( .A(n26820), .B(n21734), .Z(n26821) );
  XOR U28872 ( .A(n26823), .B(n26824), .Z(n26820) );
  AND U28873 ( .A(n26825), .B(n26826), .Z(n26823) );
  XOR U28874 ( .A(n[980]), .B(n26824), .Z(n26826) );
  XNOR U28875 ( .A(n26824), .B(n21739), .Z(n26825) );
  XOR U28876 ( .A(n26827), .B(n26828), .Z(n26824) );
  AND U28877 ( .A(n26829), .B(n26830), .Z(n26827) );
  XOR U28878 ( .A(n[979]), .B(n26828), .Z(n26830) );
  XNOR U28879 ( .A(n26828), .B(n21744), .Z(n26829) );
  XOR U28880 ( .A(n26831), .B(n26832), .Z(n26828) );
  AND U28881 ( .A(n26833), .B(n26834), .Z(n26831) );
  XOR U28882 ( .A(n[978]), .B(n26832), .Z(n26834) );
  XNOR U28883 ( .A(n26832), .B(n21749), .Z(n26833) );
  XOR U28884 ( .A(n26835), .B(n26836), .Z(n26832) );
  AND U28885 ( .A(n26837), .B(n26838), .Z(n26835) );
  XOR U28886 ( .A(n[977]), .B(n26836), .Z(n26838) );
  XNOR U28887 ( .A(n26836), .B(n21754), .Z(n26837) );
  XOR U28888 ( .A(n26839), .B(n26840), .Z(n26836) );
  AND U28889 ( .A(n26841), .B(n26842), .Z(n26839) );
  XOR U28890 ( .A(n[976]), .B(n26840), .Z(n26842) );
  XNOR U28891 ( .A(n26840), .B(n21759), .Z(n26841) );
  XOR U28892 ( .A(n26843), .B(n26844), .Z(n26840) );
  AND U28893 ( .A(n26845), .B(n26846), .Z(n26843) );
  XOR U28894 ( .A(n[975]), .B(n26844), .Z(n26846) );
  XNOR U28895 ( .A(n26844), .B(n21764), .Z(n26845) );
  XOR U28896 ( .A(n26847), .B(n26848), .Z(n26844) );
  AND U28897 ( .A(n26849), .B(n26850), .Z(n26847) );
  XOR U28898 ( .A(n[974]), .B(n26848), .Z(n26850) );
  XNOR U28899 ( .A(n26848), .B(n21769), .Z(n26849) );
  XOR U28900 ( .A(n26851), .B(n26852), .Z(n26848) );
  AND U28901 ( .A(n26853), .B(n26854), .Z(n26851) );
  XOR U28902 ( .A(n[973]), .B(n26852), .Z(n26854) );
  XNOR U28903 ( .A(n26852), .B(n21774), .Z(n26853) );
  XOR U28904 ( .A(n26855), .B(n26856), .Z(n26852) );
  AND U28905 ( .A(n26857), .B(n26858), .Z(n26855) );
  XOR U28906 ( .A(n[972]), .B(n26856), .Z(n26858) );
  XNOR U28907 ( .A(n26856), .B(n21779), .Z(n26857) );
  XOR U28908 ( .A(n26859), .B(n26860), .Z(n26856) );
  AND U28909 ( .A(n26861), .B(n26862), .Z(n26859) );
  XOR U28910 ( .A(n[971]), .B(n26860), .Z(n26862) );
  XNOR U28911 ( .A(n26860), .B(n21784), .Z(n26861) );
  XOR U28912 ( .A(n26863), .B(n26864), .Z(n26860) );
  AND U28913 ( .A(n26865), .B(n26866), .Z(n26863) );
  XOR U28914 ( .A(n[970]), .B(n26864), .Z(n26866) );
  XNOR U28915 ( .A(n26864), .B(n21789), .Z(n26865) );
  XOR U28916 ( .A(n26867), .B(n26868), .Z(n26864) );
  AND U28917 ( .A(n26869), .B(n26870), .Z(n26867) );
  XOR U28918 ( .A(n[969]), .B(n26868), .Z(n26870) );
  XNOR U28919 ( .A(n26868), .B(n21794), .Z(n26869) );
  XOR U28920 ( .A(n26871), .B(n26872), .Z(n26868) );
  AND U28921 ( .A(n26873), .B(n26874), .Z(n26871) );
  XOR U28922 ( .A(n[968]), .B(n26872), .Z(n26874) );
  XNOR U28923 ( .A(n26872), .B(n21799), .Z(n26873) );
  XOR U28924 ( .A(n26875), .B(n26876), .Z(n26872) );
  AND U28925 ( .A(n26877), .B(n26878), .Z(n26875) );
  XOR U28926 ( .A(n[967]), .B(n26876), .Z(n26878) );
  XNOR U28927 ( .A(n26876), .B(n21804), .Z(n26877) );
  XOR U28928 ( .A(n26879), .B(n26880), .Z(n26876) );
  AND U28929 ( .A(n26881), .B(n26882), .Z(n26879) );
  XOR U28930 ( .A(n[966]), .B(n26880), .Z(n26882) );
  XNOR U28931 ( .A(n26880), .B(n21809), .Z(n26881) );
  XOR U28932 ( .A(n26883), .B(n26884), .Z(n26880) );
  AND U28933 ( .A(n26885), .B(n26886), .Z(n26883) );
  XOR U28934 ( .A(n[965]), .B(n26884), .Z(n26886) );
  XNOR U28935 ( .A(n26884), .B(n21814), .Z(n26885) );
  XOR U28936 ( .A(n26887), .B(n26888), .Z(n26884) );
  AND U28937 ( .A(n26889), .B(n26890), .Z(n26887) );
  XOR U28938 ( .A(n[964]), .B(n26888), .Z(n26890) );
  XNOR U28939 ( .A(n26888), .B(n21819), .Z(n26889) );
  XOR U28940 ( .A(n26891), .B(n26892), .Z(n26888) );
  AND U28941 ( .A(n26893), .B(n26894), .Z(n26891) );
  XOR U28942 ( .A(n[963]), .B(n26892), .Z(n26894) );
  XNOR U28943 ( .A(n26892), .B(n21824), .Z(n26893) );
  XOR U28944 ( .A(n26895), .B(n26896), .Z(n26892) );
  AND U28945 ( .A(n26897), .B(n26898), .Z(n26895) );
  XOR U28946 ( .A(n[962]), .B(n26896), .Z(n26898) );
  XNOR U28947 ( .A(n26896), .B(n21829), .Z(n26897) );
  XOR U28948 ( .A(n26899), .B(n26900), .Z(n26896) );
  AND U28949 ( .A(n26901), .B(n26902), .Z(n26899) );
  XOR U28950 ( .A(n[961]), .B(n26900), .Z(n26902) );
  XNOR U28951 ( .A(n26900), .B(n21834), .Z(n26901) );
  XOR U28952 ( .A(n26903), .B(n26904), .Z(n26900) );
  AND U28953 ( .A(n26905), .B(n26906), .Z(n26903) );
  XOR U28954 ( .A(n[960]), .B(n26904), .Z(n26906) );
  XNOR U28955 ( .A(n26904), .B(n21839), .Z(n26905) );
  XOR U28956 ( .A(n26907), .B(n26908), .Z(n26904) );
  AND U28957 ( .A(n26909), .B(n26910), .Z(n26907) );
  XOR U28958 ( .A(n[959]), .B(n26908), .Z(n26910) );
  XNOR U28959 ( .A(n26908), .B(n21844), .Z(n26909) );
  XOR U28960 ( .A(n26911), .B(n26912), .Z(n26908) );
  AND U28961 ( .A(n26913), .B(n26914), .Z(n26911) );
  XOR U28962 ( .A(n[958]), .B(n26912), .Z(n26914) );
  XNOR U28963 ( .A(n26912), .B(n21849), .Z(n26913) );
  XOR U28964 ( .A(n26915), .B(n26916), .Z(n26912) );
  AND U28965 ( .A(n26917), .B(n26918), .Z(n26915) );
  XOR U28966 ( .A(n[957]), .B(n26916), .Z(n26918) );
  XNOR U28967 ( .A(n26916), .B(n21854), .Z(n26917) );
  XOR U28968 ( .A(n26919), .B(n26920), .Z(n26916) );
  AND U28969 ( .A(n26921), .B(n26922), .Z(n26919) );
  XOR U28970 ( .A(n[956]), .B(n26920), .Z(n26922) );
  XNOR U28971 ( .A(n26920), .B(n21859), .Z(n26921) );
  XOR U28972 ( .A(n26923), .B(n26924), .Z(n26920) );
  AND U28973 ( .A(n26925), .B(n26926), .Z(n26923) );
  XOR U28974 ( .A(n[955]), .B(n26924), .Z(n26926) );
  XNOR U28975 ( .A(n26924), .B(n21864), .Z(n26925) );
  XOR U28976 ( .A(n26927), .B(n26928), .Z(n26924) );
  AND U28977 ( .A(n26929), .B(n26930), .Z(n26927) );
  XOR U28978 ( .A(n[954]), .B(n26928), .Z(n26930) );
  XNOR U28979 ( .A(n26928), .B(n21869), .Z(n26929) );
  XOR U28980 ( .A(n26931), .B(n26932), .Z(n26928) );
  AND U28981 ( .A(n26933), .B(n26934), .Z(n26931) );
  XOR U28982 ( .A(n[953]), .B(n26932), .Z(n26934) );
  XNOR U28983 ( .A(n26932), .B(n21874), .Z(n26933) );
  XOR U28984 ( .A(n26935), .B(n26936), .Z(n26932) );
  AND U28985 ( .A(n26937), .B(n26938), .Z(n26935) );
  XOR U28986 ( .A(n[952]), .B(n26936), .Z(n26938) );
  XNOR U28987 ( .A(n26936), .B(n21879), .Z(n26937) );
  XOR U28988 ( .A(n26939), .B(n26940), .Z(n26936) );
  AND U28989 ( .A(n26941), .B(n26942), .Z(n26939) );
  XOR U28990 ( .A(n[951]), .B(n26940), .Z(n26942) );
  XNOR U28991 ( .A(n26940), .B(n21884), .Z(n26941) );
  XOR U28992 ( .A(n26943), .B(n26944), .Z(n26940) );
  AND U28993 ( .A(n26945), .B(n26946), .Z(n26943) );
  XOR U28994 ( .A(n[950]), .B(n26944), .Z(n26946) );
  XNOR U28995 ( .A(n26944), .B(n21889), .Z(n26945) );
  XOR U28996 ( .A(n26947), .B(n26948), .Z(n26944) );
  AND U28997 ( .A(n26949), .B(n26950), .Z(n26947) );
  XOR U28998 ( .A(n[949]), .B(n26948), .Z(n26950) );
  XNOR U28999 ( .A(n26948), .B(n21894), .Z(n26949) );
  XOR U29000 ( .A(n26951), .B(n26952), .Z(n26948) );
  AND U29001 ( .A(n26953), .B(n26954), .Z(n26951) );
  XOR U29002 ( .A(n[948]), .B(n26952), .Z(n26954) );
  XNOR U29003 ( .A(n26952), .B(n21899), .Z(n26953) );
  XOR U29004 ( .A(n26955), .B(n26956), .Z(n26952) );
  AND U29005 ( .A(n26957), .B(n26958), .Z(n26955) );
  XOR U29006 ( .A(n[947]), .B(n26956), .Z(n26958) );
  XNOR U29007 ( .A(n26956), .B(n21904), .Z(n26957) );
  XOR U29008 ( .A(n26959), .B(n26960), .Z(n26956) );
  AND U29009 ( .A(n26961), .B(n26962), .Z(n26959) );
  XOR U29010 ( .A(n[946]), .B(n26960), .Z(n26962) );
  XNOR U29011 ( .A(n26960), .B(n21909), .Z(n26961) );
  XOR U29012 ( .A(n26963), .B(n26964), .Z(n26960) );
  AND U29013 ( .A(n26965), .B(n26966), .Z(n26963) );
  XOR U29014 ( .A(n[945]), .B(n26964), .Z(n26966) );
  XNOR U29015 ( .A(n26964), .B(n21914), .Z(n26965) );
  XOR U29016 ( .A(n26967), .B(n26968), .Z(n26964) );
  AND U29017 ( .A(n26969), .B(n26970), .Z(n26967) );
  XOR U29018 ( .A(n[944]), .B(n26968), .Z(n26970) );
  XNOR U29019 ( .A(n26968), .B(n21919), .Z(n26969) );
  XOR U29020 ( .A(n26971), .B(n26972), .Z(n26968) );
  AND U29021 ( .A(n26973), .B(n26974), .Z(n26971) );
  XOR U29022 ( .A(n[943]), .B(n26972), .Z(n26974) );
  XNOR U29023 ( .A(n26972), .B(n21924), .Z(n26973) );
  XOR U29024 ( .A(n26975), .B(n26976), .Z(n26972) );
  AND U29025 ( .A(n26977), .B(n26978), .Z(n26975) );
  XOR U29026 ( .A(n[942]), .B(n26976), .Z(n26978) );
  XNOR U29027 ( .A(n26976), .B(n21929), .Z(n26977) );
  XOR U29028 ( .A(n26979), .B(n26980), .Z(n26976) );
  AND U29029 ( .A(n26981), .B(n26982), .Z(n26979) );
  XOR U29030 ( .A(n[941]), .B(n26980), .Z(n26982) );
  XNOR U29031 ( .A(n26980), .B(n21934), .Z(n26981) );
  XOR U29032 ( .A(n26983), .B(n26984), .Z(n26980) );
  AND U29033 ( .A(n26985), .B(n26986), .Z(n26983) );
  XOR U29034 ( .A(n[940]), .B(n26984), .Z(n26986) );
  XNOR U29035 ( .A(n26984), .B(n21939), .Z(n26985) );
  XOR U29036 ( .A(n26987), .B(n26988), .Z(n26984) );
  AND U29037 ( .A(n26989), .B(n26990), .Z(n26987) );
  XOR U29038 ( .A(n[939]), .B(n26988), .Z(n26990) );
  XNOR U29039 ( .A(n26988), .B(n21944), .Z(n26989) );
  XOR U29040 ( .A(n26991), .B(n26992), .Z(n26988) );
  AND U29041 ( .A(n26993), .B(n26994), .Z(n26991) );
  XOR U29042 ( .A(n[938]), .B(n26992), .Z(n26994) );
  XNOR U29043 ( .A(n26992), .B(n21949), .Z(n26993) );
  XOR U29044 ( .A(n26995), .B(n26996), .Z(n26992) );
  AND U29045 ( .A(n26997), .B(n26998), .Z(n26995) );
  XOR U29046 ( .A(n[937]), .B(n26996), .Z(n26998) );
  XNOR U29047 ( .A(n26996), .B(n21954), .Z(n26997) );
  XOR U29048 ( .A(n26999), .B(n27000), .Z(n26996) );
  AND U29049 ( .A(n27001), .B(n27002), .Z(n26999) );
  XOR U29050 ( .A(n[936]), .B(n27000), .Z(n27002) );
  XNOR U29051 ( .A(n27000), .B(n21959), .Z(n27001) );
  XOR U29052 ( .A(n27003), .B(n27004), .Z(n27000) );
  AND U29053 ( .A(n27005), .B(n27006), .Z(n27003) );
  XOR U29054 ( .A(n[935]), .B(n27004), .Z(n27006) );
  XNOR U29055 ( .A(n27004), .B(n21964), .Z(n27005) );
  XOR U29056 ( .A(n27007), .B(n27008), .Z(n27004) );
  AND U29057 ( .A(n27009), .B(n27010), .Z(n27007) );
  XOR U29058 ( .A(n[934]), .B(n27008), .Z(n27010) );
  XNOR U29059 ( .A(n27008), .B(n21969), .Z(n27009) );
  XOR U29060 ( .A(n27011), .B(n27012), .Z(n27008) );
  AND U29061 ( .A(n27013), .B(n27014), .Z(n27011) );
  XOR U29062 ( .A(n[933]), .B(n27012), .Z(n27014) );
  XNOR U29063 ( .A(n27012), .B(n21974), .Z(n27013) );
  XOR U29064 ( .A(n27015), .B(n27016), .Z(n27012) );
  AND U29065 ( .A(n27017), .B(n27018), .Z(n27015) );
  XOR U29066 ( .A(n[932]), .B(n27016), .Z(n27018) );
  XNOR U29067 ( .A(n27016), .B(n21979), .Z(n27017) );
  XOR U29068 ( .A(n27019), .B(n27020), .Z(n27016) );
  AND U29069 ( .A(n27021), .B(n27022), .Z(n27019) );
  XOR U29070 ( .A(n[931]), .B(n27020), .Z(n27022) );
  XNOR U29071 ( .A(n27020), .B(n21984), .Z(n27021) );
  XOR U29072 ( .A(n27023), .B(n27024), .Z(n27020) );
  AND U29073 ( .A(n27025), .B(n27026), .Z(n27023) );
  XOR U29074 ( .A(n[930]), .B(n27024), .Z(n27026) );
  XNOR U29075 ( .A(n27024), .B(n21989), .Z(n27025) );
  XOR U29076 ( .A(n27027), .B(n27028), .Z(n27024) );
  AND U29077 ( .A(n27029), .B(n27030), .Z(n27027) );
  XOR U29078 ( .A(n[929]), .B(n27028), .Z(n27030) );
  XNOR U29079 ( .A(n27028), .B(n21994), .Z(n27029) );
  XOR U29080 ( .A(n27031), .B(n27032), .Z(n27028) );
  AND U29081 ( .A(n27033), .B(n27034), .Z(n27031) );
  XOR U29082 ( .A(n[928]), .B(n27032), .Z(n27034) );
  XNOR U29083 ( .A(n27032), .B(n21999), .Z(n27033) );
  XOR U29084 ( .A(n27035), .B(n27036), .Z(n27032) );
  AND U29085 ( .A(n27037), .B(n27038), .Z(n27035) );
  XOR U29086 ( .A(n[927]), .B(n27036), .Z(n27038) );
  XNOR U29087 ( .A(n27036), .B(n22004), .Z(n27037) );
  XOR U29088 ( .A(n27039), .B(n27040), .Z(n27036) );
  AND U29089 ( .A(n27041), .B(n27042), .Z(n27039) );
  XOR U29090 ( .A(n[926]), .B(n27040), .Z(n27042) );
  XNOR U29091 ( .A(n27040), .B(n22009), .Z(n27041) );
  XOR U29092 ( .A(n27043), .B(n27044), .Z(n27040) );
  AND U29093 ( .A(n27045), .B(n27046), .Z(n27043) );
  XOR U29094 ( .A(n[925]), .B(n27044), .Z(n27046) );
  XNOR U29095 ( .A(n27044), .B(n22014), .Z(n27045) );
  XOR U29096 ( .A(n27047), .B(n27048), .Z(n27044) );
  AND U29097 ( .A(n27049), .B(n27050), .Z(n27047) );
  XOR U29098 ( .A(n[924]), .B(n27048), .Z(n27050) );
  XNOR U29099 ( .A(n27048), .B(n22019), .Z(n27049) );
  XOR U29100 ( .A(n27051), .B(n27052), .Z(n27048) );
  AND U29101 ( .A(n27053), .B(n27054), .Z(n27051) );
  XOR U29102 ( .A(n[923]), .B(n27052), .Z(n27054) );
  XNOR U29103 ( .A(n27052), .B(n22024), .Z(n27053) );
  XOR U29104 ( .A(n27055), .B(n27056), .Z(n27052) );
  AND U29105 ( .A(n27057), .B(n27058), .Z(n27055) );
  XOR U29106 ( .A(n[922]), .B(n27056), .Z(n27058) );
  XNOR U29107 ( .A(n27056), .B(n22029), .Z(n27057) );
  XOR U29108 ( .A(n27059), .B(n27060), .Z(n27056) );
  AND U29109 ( .A(n27061), .B(n27062), .Z(n27059) );
  XOR U29110 ( .A(n[921]), .B(n27060), .Z(n27062) );
  XNOR U29111 ( .A(n27060), .B(n22034), .Z(n27061) );
  XOR U29112 ( .A(n27063), .B(n27064), .Z(n27060) );
  AND U29113 ( .A(n27065), .B(n27066), .Z(n27063) );
  XOR U29114 ( .A(n[920]), .B(n27064), .Z(n27066) );
  XNOR U29115 ( .A(n27064), .B(n22039), .Z(n27065) );
  XOR U29116 ( .A(n27067), .B(n27068), .Z(n27064) );
  AND U29117 ( .A(n27069), .B(n27070), .Z(n27067) );
  XOR U29118 ( .A(n[919]), .B(n27068), .Z(n27070) );
  XNOR U29119 ( .A(n27068), .B(n22044), .Z(n27069) );
  XOR U29120 ( .A(n27071), .B(n27072), .Z(n27068) );
  AND U29121 ( .A(n27073), .B(n27074), .Z(n27071) );
  XOR U29122 ( .A(n[918]), .B(n27072), .Z(n27074) );
  XNOR U29123 ( .A(n27072), .B(n22049), .Z(n27073) );
  XOR U29124 ( .A(n27075), .B(n27076), .Z(n27072) );
  AND U29125 ( .A(n27077), .B(n27078), .Z(n27075) );
  XOR U29126 ( .A(n[917]), .B(n27076), .Z(n27078) );
  XNOR U29127 ( .A(n27076), .B(n22054), .Z(n27077) );
  XOR U29128 ( .A(n27079), .B(n27080), .Z(n27076) );
  AND U29129 ( .A(n27081), .B(n27082), .Z(n27079) );
  XOR U29130 ( .A(n[916]), .B(n27080), .Z(n27082) );
  XNOR U29131 ( .A(n27080), .B(n22059), .Z(n27081) );
  XOR U29132 ( .A(n27083), .B(n27084), .Z(n27080) );
  AND U29133 ( .A(n27085), .B(n27086), .Z(n27083) );
  XOR U29134 ( .A(n[915]), .B(n27084), .Z(n27086) );
  XNOR U29135 ( .A(n27084), .B(n22064), .Z(n27085) );
  XOR U29136 ( .A(n27087), .B(n27088), .Z(n27084) );
  AND U29137 ( .A(n27089), .B(n27090), .Z(n27087) );
  XOR U29138 ( .A(n[914]), .B(n27088), .Z(n27090) );
  XNOR U29139 ( .A(n27088), .B(n22069), .Z(n27089) );
  XOR U29140 ( .A(n27091), .B(n27092), .Z(n27088) );
  AND U29141 ( .A(n27093), .B(n27094), .Z(n27091) );
  XOR U29142 ( .A(n[913]), .B(n27092), .Z(n27094) );
  XNOR U29143 ( .A(n27092), .B(n22074), .Z(n27093) );
  XOR U29144 ( .A(n27095), .B(n27096), .Z(n27092) );
  AND U29145 ( .A(n27097), .B(n27098), .Z(n27095) );
  XOR U29146 ( .A(n[912]), .B(n27096), .Z(n27098) );
  XNOR U29147 ( .A(n27096), .B(n22079), .Z(n27097) );
  XOR U29148 ( .A(n27099), .B(n27100), .Z(n27096) );
  AND U29149 ( .A(n27101), .B(n27102), .Z(n27099) );
  XOR U29150 ( .A(n[911]), .B(n27100), .Z(n27102) );
  XNOR U29151 ( .A(n27100), .B(n22084), .Z(n27101) );
  XOR U29152 ( .A(n27103), .B(n27104), .Z(n27100) );
  AND U29153 ( .A(n27105), .B(n27106), .Z(n27103) );
  XOR U29154 ( .A(n[910]), .B(n27104), .Z(n27106) );
  XNOR U29155 ( .A(n27104), .B(n22089), .Z(n27105) );
  XOR U29156 ( .A(n27107), .B(n27108), .Z(n27104) );
  AND U29157 ( .A(n27109), .B(n27110), .Z(n27107) );
  XOR U29158 ( .A(n[909]), .B(n27108), .Z(n27110) );
  XNOR U29159 ( .A(n27108), .B(n22094), .Z(n27109) );
  XOR U29160 ( .A(n27111), .B(n27112), .Z(n27108) );
  AND U29161 ( .A(n27113), .B(n27114), .Z(n27111) );
  XOR U29162 ( .A(n[908]), .B(n27112), .Z(n27114) );
  XNOR U29163 ( .A(n27112), .B(n22099), .Z(n27113) );
  XOR U29164 ( .A(n27115), .B(n27116), .Z(n27112) );
  AND U29165 ( .A(n27117), .B(n27118), .Z(n27115) );
  XOR U29166 ( .A(n[907]), .B(n27116), .Z(n27118) );
  XNOR U29167 ( .A(n27116), .B(n22104), .Z(n27117) );
  XOR U29168 ( .A(n27119), .B(n27120), .Z(n27116) );
  AND U29169 ( .A(n27121), .B(n27122), .Z(n27119) );
  XOR U29170 ( .A(n[906]), .B(n27120), .Z(n27122) );
  XNOR U29171 ( .A(n27120), .B(n22109), .Z(n27121) );
  XOR U29172 ( .A(n27123), .B(n27124), .Z(n27120) );
  AND U29173 ( .A(n27125), .B(n27126), .Z(n27123) );
  XOR U29174 ( .A(n[905]), .B(n27124), .Z(n27126) );
  XNOR U29175 ( .A(n27124), .B(n22114), .Z(n27125) );
  XOR U29176 ( .A(n27127), .B(n27128), .Z(n27124) );
  AND U29177 ( .A(n27129), .B(n27130), .Z(n27127) );
  XOR U29178 ( .A(n[904]), .B(n27128), .Z(n27130) );
  XNOR U29179 ( .A(n27128), .B(n22119), .Z(n27129) );
  XOR U29180 ( .A(n27131), .B(n27132), .Z(n27128) );
  AND U29181 ( .A(n27133), .B(n27134), .Z(n27131) );
  XOR U29182 ( .A(n[903]), .B(n27132), .Z(n27134) );
  XNOR U29183 ( .A(n27132), .B(n22124), .Z(n27133) );
  XOR U29184 ( .A(n27135), .B(n27136), .Z(n27132) );
  AND U29185 ( .A(n27137), .B(n27138), .Z(n27135) );
  XOR U29186 ( .A(n[902]), .B(n27136), .Z(n27138) );
  XNOR U29187 ( .A(n27136), .B(n22129), .Z(n27137) );
  XOR U29188 ( .A(n27139), .B(n27140), .Z(n27136) );
  AND U29189 ( .A(n27141), .B(n27142), .Z(n27139) );
  XOR U29190 ( .A(n[901]), .B(n27140), .Z(n27142) );
  XNOR U29191 ( .A(n27140), .B(n22134), .Z(n27141) );
  XOR U29192 ( .A(n27143), .B(n27144), .Z(n27140) );
  AND U29193 ( .A(n27145), .B(n27146), .Z(n27143) );
  XOR U29194 ( .A(n[900]), .B(n27144), .Z(n27146) );
  XNOR U29195 ( .A(n27144), .B(n22139), .Z(n27145) );
  XOR U29196 ( .A(n27147), .B(n27148), .Z(n27144) );
  AND U29197 ( .A(n27149), .B(n27150), .Z(n27147) );
  XOR U29198 ( .A(n[899]), .B(n27148), .Z(n27150) );
  XNOR U29199 ( .A(n27148), .B(n22144), .Z(n27149) );
  XOR U29200 ( .A(n27151), .B(n27152), .Z(n27148) );
  AND U29201 ( .A(n27153), .B(n27154), .Z(n27151) );
  XOR U29202 ( .A(n[898]), .B(n27152), .Z(n27154) );
  XNOR U29203 ( .A(n27152), .B(n22149), .Z(n27153) );
  XOR U29204 ( .A(n27155), .B(n27156), .Z(n27152) );
  AND U29205 ( .A(n27157), .B(n27158), .Z(n27155) );
  XOR U29206 ( .A(n[897]), .B(n27156), .Z(n27158) );
  XNOR U29207 ( .A(n27156), .B(n22154), .Z(n27157) );
  XOR U29208 ( .A(n27159), .B(n27160), .Z(n27156) );
  AND U29209 ( .A(n27161), .B(n27162), .Z(n27159) );
  XOR U29210 ( .A(n[896]), .B(n27160), .Z(n27162) );
  XNOR U29211 ( .A(n27160), .B(n22159), .Z(n27161) );
  XOR U29212 ( .A(n27163), .B(n27164), .Z(n27160) );
  AND U29213 ( .A(n27165), .B(n27166), .Z(n27163) );
  XOR U29214 ( .A(n[895]), .B(n27164), .Z(n27166) );
  XNOR U29215 ( .A(n27164), .B(n22164), .Z(n27165) );
  XOR U29216 ( .A(n27167), .B(n27168), .Z(n27164) );
  AND U29217 ( .A(n27169), .B(n27170), .Z(n27167) );
  XOR U29218 ( .A(n[894]), .B(n27168), .Z(n27170) );
  XNOR U29219 ( .A(n27168), .B(n22169), .Z(n27169) );
  XOR U29220 ( .A(n27171), .B(n27172), .Z(n27168) );
  AND U29221 ( .A(n27173), .B(n27174), .Z(n27171) );
  XOR U29222 ( .A(n[893]), .B(n27172), .Z(n27174) );
  XNOR U29223 ( .A(n27172), .B(n22174), .Z(n27173) );
  XOR U29224 ( .A(n27175), .B(n27176), .Z(n27172) );
  AND U29225 ( .A(n27177), .B(n27178), .Z(n27175) );
  XOR U29226 ( .A(n[892]), .B(n27176), .Z(n27178) );
  XNOR U29227 ( .A(n27176), .B(n22179), .Z(n27177) );
  XOR U29228 ( .A(n27179), .B(n27180), .Z(n27176) );
  AND U29229 ( .A(n27181), .B(n27182), .Z(n27179) );
  XOR U29230 ( .A(n[891]), .B(n27180), .Z(n27182) );
  XNOR U29231 ( .A(n27180), .B(n22184), .Z(n27181) );
  XOR U29232 ( .A(n27183), .B(n27184), .Z(n27180) );
  AND U29233 ( .A(n27185), .B(n27186), .Z(n27183) );
  XOR U29234 ( .A(n[890]), .B(n27184), .Z(n27186) );
  XNOR U29235 ( .A(n27184), .B(n22189), .Z(n27185) );
  XOR U29236 ( .A(n27187), .B(n27188), .Z(n27184) );
  AND U29237 ( .A(n27189), .B(n27190), .Z(n27187) );
  XOR U29238 ( .A(n[889]), .B(n27188), .Z(n27190) );
  XNOR U29239 ( .A(n27188), .B(n22194), .Z(n27189) );
  XOR U29240 ( .A(n27191), .B(n27192), .Z(n27188) );
  AND U29241 ( .A(n27193), .B(n27194), .Z(n27191) );
  XOR U29242 ( .A(n[888]), .B(n27192), .Z(n27194) );
  XNOR U29243 ( .A(n27192), .B(n22199), .Z(n27193) );
  XOR U29244 ( .A(n27195), .B(n27196), .Z(n27192) );
  AND U29245 ( .A(n27197), .B(n27198), .Z(n27195) );
  XOR U29246 ( .A(n[887]), .B(n27196), .Z(n27198) );
  XNOR U29247 ( .A(n27196), .B(n22204), .Z(n27197) );
  XOR U29248 ( .A(n27199), .B(n27200), .Z(n27196) );
  AND U29249 ( .A(n27201), .B(n27202), .Z(n27199) );
  XOR U29250 ( .A(n[886]), .B(n27200), .Z(n27202) );
  XNOR U29251 ( .A(n27200), .B(n22209), .Z(n27201) );
  XOR U29252 ( .A(n27203), .B(n27204), .Z(n27200) );
  AND U29253 ( .A(n27205), .B(n27206), .Z(n27203) );
  XOR U29254 ( .A(n[885]), .B(n27204), .Z(n27206) );
  XNOR U29255 ( .A(n27204), .B(n22214), .Z(n27205) );
  XOR U29256 ( .A(n27207), .B(n27208), .Z(n27204) );
  AND U29257 ( .A(n27209), .B(n27210), .Z(n27207) );
  XOR U29258 ( .A(n[884]), .B(n27208), .Z(n27210) );
  XNOR U29259 ( .A(n27208), .B(n22219), .Z(n27209) );
  XOR U29260 ( .A(n27211), .B(n27212), .Z(n27208) );
  AND U29261 ( .A(n27213), .B(n27214), .Z(n27211) );
  XOR U29262 ( .A(n[883]), .B(n27212), .Z(n27214) );
  XNOR U29263 ( .A(n27212), .B(n22224), .Z(n27213) );
  XOR U29264 ( .A(n27215), .B(n27216), .Z(n27212) );
  AND U29265 ( .A(n27217), .B(n27218), .Z(n27215) );
  XOR U29266 ( .A(n[882]), .B(n27216), .Z(n27218) );
  XNOR U29267 ( .A(n27216), .B(n22229), .Z(n27217) );
  XOR U29268 ( .A(n27219), .B(n27220), .Z(n27216) );
  AND U29269 ( .A(n27221), .B(n27222), .Z(n27219) );
  XOR U29270 ( .A(n[881]), .B(n27220), .Z(n27222) );
  XNOR U29271 ( .A(n27220), .B(n22234), .Z(n27221) );
  XOR U29272 ( .A(n27223), .B(n27224), .Z(n27220) );
  AND U29273 ( .A(n27225), .B(n27226), .Z(n27223) );
  XOR U29274 ( .A(n[880]), .B(n27224), .Z(n27226) );
  XNOR U29275 ( .A(n27224), .B(n22239), .Z(n27225) );
  XOR U29276 ( .A(n27227), .B(n27228), .Z(n27224) );
  AND U29277 ( .A(n27229), .B(n27230), .Z(n27227) );
  XOR U29278 ( .A(n[879]), .B(n27228), .Z(n27230) );
  XNOR U29279 ( .A(n27228), .B(n22244), .Z(n27229) );
  XOR U29280 ( .A(n27231), .B(n27232), .Z(n27228) );
  AND U29281 ( .A(n27233), .B(n27234), .Z(n27231) );
  XOR U29282 ( .A(n[878]), .B(n27232), .Z(n27234) );
  XNOR U29283 ( .A(n27232), .B(n22249), .Z(n27233) );
  XOR U29284 ( .A(n27235), .B(n27236), .Z(n27232) );
  AND U29285 ( .A(n27237), .B(n27238), .Z(n27235) );
  XOR U29286 ( .A(n[877]), .B(n27236), .Z(n27238) );
  XNOR U29287 ( .A(n27236), .B(n22254), .Z(n27237) );
  XOR U29288 ( .A(n27239), .B(n27240), .Z(n27236) );
  AND U29289 ( .A(n27241), .B(n27242), .Z(n27239) );
  XOR U29290 ( .A(n[876]), .B(n27240), .Z(n27242) );
  XNOR U29291 ( .A(n27240), .B(n22259), .Z(n27241) );
  XOR U29292 ( .A(n27243), .B(n27244), .Z(n27240) );
  AND U29293 ( .A(n27245), .B(n27246), .Z(n27243) );
  XOR U29294 ( .A(n[875]), .B(n27244), .Z(n27246) );
  XNOR U29295 ( .A(n27244), .B(n22264), .Z(n27245) );
  XOR U29296 ( .A(n27247), .B(n27248), .Z(n27244) );
  AND U29297 ( .A(n27249), .B(n27250), .Z(n27247) );
  XOR U29298 ( .A(n[874]), .B(n27248), .Z(n27250) );
  XNOR U29299 ( .A(n27248), .B(n22269), .Z(n27249) );
  XOR U29300 ( .A(n27251), .B(n27252), .Z(n27248) );
  AND U29301 ( .A(n27253), .B(n27254), .Z(n27251) );
  XOR U29302 ( .A(n[873]), .B(n27252), .Z(n27254) );
  XNOR U29303 ( .A(n27252), .B(n22274), .Z(n27253) );
  XOR U29304 ( .A(n27255), .B(n27256), .Z(n27252) );
  AND U29305 ( .A(n27257), .B(n27258), .Z(n27255) );
  XOR U29306 ( .A(n[872]), .B(n27256), .Z(n27258) );
  XNOR U29307 ( .A(n27256), .B(n22279), .Z(n27257) );
  XOR U29308 ( .A(n27259), .B(n27260), .Z(n27256) );
  AND U29309 ( .A(n27261), .B(n27262), .Z(n27259) );
  XOR U29310 ( .A(n[871]), .B(n27260), .Z(n27262) );
  XNOR U29311 ( .A(n27260), .B(n22284), .Z(n27261) );
  XOR U29312 ( .A(n27263), .B(n27264), .Z(n27260) );
  AND U29313 ( .A(n27265), .B(n27266), .Z(n27263) );
  XOR U29314 ( .A(n[870]), .B(n27264), .Z(n27266) );
  XNOR U29315 ( .A(n27264), .B(n22289), .Z(n27265) );
  XOR U29316 ( .A(n27267), .B(n27268), .Z(n27264) );
  AND U29317 ( .A(n27269), .B(n27270), .Z(n27267) );
  XOR U29318 ( .A(n[869]), .B(n27268), .Z(n27270) );
  XNOR U29319 ( .A(n27268), .B(n22294), .Z(n27269) );
  XOR U29320 ( .A(n27271), .B(n27272), .Z(n27268) );
  AND U29321 ( .A(n27273), .B(n27274), .Z(n27271) );
  XOR U29322 ( .A(n[868]), .B(n27272), .Z(n27274) );
  XNOR U29323 ( .A(n27272), .B(n22299), .Z(n27273) );
  XOR U29324 ( .A(n27275), .B(n27276), .Z(n27272) );
  AND U29325 ( .A(n27277), .B(n27278), .Z(n27275) );
  XOR U29326 ( .A(n[867]), .B(n27276), .Z(n27278) );
  XNOR U29327 ( .A(n27276), .B(n22304), .Z(n27277) );
  XOR U29328 ( .A(n27279), .B(n27280), .Z(n27276) );
  AND U29329 ( .A(n27281), .B(n27282), .Z(n27279) );
  XOR U29330 ( .A(n[866]), .B(n27280), .Z(n27282) );
  XNOR U29331 ( .A(n27280), .B(n22309), .Z(n27281) );
  XOR U29332 ( .A(n27283), .B(n27284), .Z(n27280) );
  AND U29333 ( .A(n27285), .B(n27286), .Z(n27283) );
  XOR U29334 ( .A(n[865]), .B(n27284), .Z(n27286) );
  XNOR U29335 ( .A(n27284), .B(n22314), .Z(n27285) );
  XOR U29336 ( .A(n27287), .B(n27288), .Z(n27284) );
  AND U29337 ( .A(n27289), .B(n27290), .Z(n27287) );
  XOR U29338 ( .A(n[864]), .B(n27288), .Z(n27290) );
  XNOR U29339 ( .A(n27288), .B(n22319), .Z(n27289) );
  XOR U29340 ( .A(n27291), .B(n27292), .Z(n27288) );
  AND U29341 ( .A(n27293), .B(n27294), .Z(n27291) );
  XOR U29342 ( .A(n[863]), .B(n27292), .Z(n27294) );
  XNOR U29343 ( .A(n27292), .B(n22324), .Z(n27293) );
  XOR U29344 ( .A(n27295), .B(n27296), .Z(n27292) );
  AND U29345 ( .A(n27297), .B(n27298), .Z(n27295) );
  XOR U29346 ( .A(n[862]), .B(n27296), .Z(n27298) );
  XNOR U29347 ( .A(n27296), .B(n22329), .Z(n27297) );
  XOR U29348 ( .A(n27299), .B(n27300), .Z(n27296) );
  AND U29349 ( .A(n27301), .B(n27302), .Z(n27299) );
  XOR U29350 ( .A(n[861]), .B(n27300), .Z(n27302) );
  XNOR U29351 ( .A(n27300), .B(n22334), .Z(n27301) );
  XOR U29352 ( .A(n27303), .B(n27304), .Z(n27300) );
  AND U29353 ( .A(n27305), .B(n27306), .Z(n27303) );
  XOR U29354 ( .A(n[860]), .B(n27304), .Z(n27306) );
  XNOR U29355 ( .A(n27304), .B(n22339), .Z(n27305) );
  XOR U29356 ( .A(n27307), .B(n27308), .Z(n27304) );
  AND U29357 ( .A(n27309), .B(n27310), .Z(n27307) );
  XOR U29358 ( .A(n[859]), .B(n27308), .Z(n27310) );
  XNOR U29359 ( .A(n27308), .B(n22344), .Z(n27309) );
  XOR U29360 ( .A(n27311), .B(n27312), .Z(n27308) );
  AND U29361 ( .A(n27313), .B(n27314), .Z(n27311) );
  XOR U29362 ( .A(n[858]), .B(n27312), .Z(n27314) );
  XNOR U29363 ( .A(n27312), .B(n22349), .Z(n27313) );
  XOR U29364 ( .A(n27315), .B(n27316), .Z(n27312) );
  AND U29365 ( .A(n27317), .B(n27318), .Z(n27315) );
  XOR U29366 ( .A(n[857]), .B(n27316), .Z(n27318) );
  XNOR U29367 ( .A(n27316), .B(n22354), .Z(n27317) );
  XOR U29368 ( .A(n27319), .B(n27320), .Z(n27316) );
  AND U29369 ( .A(n27321), .B(n27322), .Z(n27319) );
  XOR U29370 ( .A(n[856]), .B(n27320), .Z(n27322) );
  XNOR U29371 ( .A(n27320), .B(n22359), .Z(n27321) );
  XOR U29372 ( .A(n27323), .B(n27324), .Z(n27320) );
  AND U29373 ( .A(n27325), .B(n27326), .Z(n27323) );
  XOR U29374 ( .A(n[855]), .B(n27324), .Z(n27326) );
  XNOR U29375 ( .A(n27324), .B(n22364), .Z(n27325) );
  XOR U29376 ( .A(n27327), .B(n27328), .Z(n27324) );
  AND U29377 ( .A(n27329), .B(n27330), .Z(n27327) );
  XOR U29378 ( .A(n[854]), .B(n27328), .Z(n27330) );
  XNOR U29379 ( .A(n27328), .B(n22369), .Z(n27329) );
  XOR U29380 ( .A(n27331), .B(n27332), .Z(n27328) );
  AND U29381 ( .A(n27333), .B(n27334), .Z(n27331) );
  XOR U29382 ( .A(n[853]), .B(n27332), .Z(n27334) );
  XNOR U29383 ( .A(n27332), .B(n22374), .Z(n27333) );
  XOR U29384 ( .A(n27335), .B(n27336), .Z(n27332) );
  AND U29385 ( .A(n27337), .B(n27338), .Z(n27335) );
  XOR U29386 ( .A(n[852]), .B(n27336), .Z(n27338) );
  XNOR U29387 ( .A(n27336), .B(n22379), .Z(n27337) );
  XOR U29388 ( .A(n27339), .B(n27340), .Z(n27336) );
  AND U29389 ( .A(n27341), .B(n27342), .Z(n27339) );
  XOR U29390 ( .A(n[851]), .B(n27340), .Z(n27342) );
  XNOR U29391 ( .A(n27340), .B(n22384), .Z(n27341) );
  XOR U29392 ( .A(n27343), .B(n27344), .Z(n27340) );
  AND U29393 ( .A(n27345), .B(n27346), .Z(n27343) );
  XOR U29394 ( .A(n[850]), .B(n27344), .Z(n27346) );
  XNOR U29395 ( .A(n27344), .B(n22389), .Z(n27345) );
  XOR U29396 ( .A(n27347), .B(n27348), .Z(n27344) );
  AND U29397 ( .A(n27349), .B(n27350), .Z(n27347) );
  XOR U29398 ( .A(n[849]), .B(n27348), .Z(n27350) );
  XNOR U29399 ( .A(n27348), .B(n22394), .Z(n27349) );
  XOR U29400 ( .A(n27351), .B(n27352), .Z(n27348) );
  AND U29401 ( .A(n27353), .B(n27354), .Z(n27351) );
  XOR U29402 ( .A(n[848]), .B(n27352), .Z(n27354) );
  XNOR U29403 ( .A(n27352), .B(n22399), .Z(n27353) );
  XOR U29404 ( .A(n27355), .B(n27356), .Z(n27352) );
  AND U29405 ( .A(n27357), .B(n27358), .Z(n27355) );
  XOR U29406 ( .A(n[847]), .B(n27356), .Z(n27358) );
  XNOR U29407 ( .A(n27356), .B(n22404), .Z(n27357) );
  XOR U29408 ( .A(n27359), .B(n27360), .Z(n27356) );
  AND U29409 ( .A(n27361), .B(n27362), .Z(n27359) );
  XOR U29410 ( .A(n[846]), .B(n27360), .Z(n27362) );
  XNOR U29411 ( .A(n27360), .B(n22409), .Z(n27361) );
  XOR U29412 ( .A(n27363), .B(n27364), .Z(n27360) );
  AND U29413 ( .A(n27365), .B(n27366), .Z(n27363) );
  XOR U29414 ( .A(n[845]), .B(n27364), .Z(n27366) );
  XNOR U29415 ( .A(n27364), .B(n22414), .Z(n27365) );
  XOR U29416 ( .A(n27367), .B(n27368), .Z(n27364) );
  AND U29417 ( .A(n27369), .B(n27370), .Z(n27367) );
  XOR U29418 ( .A(n[844]), .B(n27368), .Z(n27370) );
  XNOR U29419 ( .A(n27368), .B(n22419), .Z(n27369) );
  XOR U29420 ( .A(n27371), .B(n27372), .Z(n27368) );
  AND U29421 ( .A(n27373), .B(n27374), .Z(n27371) );
  XOR U29422 ( .A(n[843]), .B(n27372), .Z(n27374) );
  XNOR U29423 ( .A(n27372), .B(n22424), .Z(n27373) );
  XOR U29424 ( .A(n27375), .B(n27376), .Z(n27372) );
  AND U29425 ( .A(n27377), .B(n27378), .Z(n27375) );
  XOR U29426 ( .A(n[842]), .B(n27376), .Z(n27378) );
  XNOR U29427 ( .A(n27376), .B(n22429), .Z(n27377) );
  XOR U29428 ( .A(n27379), .B(n27380), .Z(n27376) );
  AND U29429 ( .A(n27381), .B(n27382), .Z(n27379) );
  XOR U29430 ( .A(n[841]), .B(n27380), .Z(n27382) );
  XNOR U29431 ( .A(n27380), .B(n22434), .Z(n27381) );
  XOR U29432 ( .A(n27383), .B(n27384), .Z(n27380) );
  AND U29433 ( .A(n27385), .B(n27386), .Z(n27383) );
  XOR U29434 ( .A(n[840]), .B(n27384), .Z(n27386) );
  XNOR U29435 ( .A(n27384), .B(n22439), .Z(n27385) );
  XOR U29436 ( .A(n27387), .B(n27388), .Z(n27384) );
  AND U29437 ( .A(n27389), .B(n27390), .Z(n27387) );
  XOR U29438 ( .A(n[839]), .B(n27388), .Z(n27390) );
  XNOR U29439 ( .A(n27388), .B(n22444), .Z(n27389) );
  XOR U29440 ( .A(n27391), .B(n27392), .Z(n27388) );
  AND U29441 ( .A(n27393), .B(n27394), .Z(n27391) );
  XOR U29442 ( .A(n[838]), .B(n27392), .Z(n27394) );
  XNOR U29443 ( .A(n27392), .B(n22449), .Z(n27393) );
  XOR U29444 ( .A(n27395), .B(n27396), .Z(n27392) );
  AND U29445 ( .A(n27397), .B(n27398), .Z(n27395) );
  XOR U29446 ( .A(n[837]), .B(n27396), .Z(n27398) );
  XNOR U29447 ( .A(n27396), .B(n22454), .Z(n27397) );
  XOR U29448 ( .A(n27399), .B(n27400), .Z(n27396) );
  AND U29449 ( .A(n27401), .B(n27402), .Z(n27399) );
  XOR U29450 ( .A(n[836]), .B(n27400), .Z(n27402) );
  XNOR U29451 ( .A(n27400), .B(n22459), .Z(n27401) );
  XOR U29452 ( .A(n27403), .B(n27404), .Z(n27400) );
  AND U29453 ( .A(n27405), .B(n27406), .Z(n27403) );
  XOR U29454 ( .A(n[835]), .B(n27404), .Z(n27406) );
  XNOR U29455 ( .A(n27404), .B(n22464), .Z(n27405) );
  XOR U29456 ( .A(n27407), .B(n27408), .Z(n27404) );
  AND U29457 ( .A(n27409), .B(n27410), .Z(n27407) );
  XOR U29458 ( .A(n[834]), .B(n27408), .Z(n27410) );
  XNOR U29459 ( .A(n27408), .B(n22469), .Z(n27409) );
  XOR U29460 ( .A(n27411), .B(n27412), .Z(n27408) );
  AND U29461 ( .A(n27413), .B(n27414), .Z(n27411) );
  XOR U29462 ( .A(n[833]), .B(n27412), .Z(n27414) );
  XNOR U29463 ( .A(n27412), .B(n22474), .Z(n27413) );
  XOR U29464 ( .A(n27415), .B(n27416), .Z(n27412) );
  AND U29465 ( .A(n27417), .B(n27418), .Z(n27415) );
  XOR U29466 ( .A(n[832]), .B(n27416), .Z(n27418) );
  XNOR U29467 ( .A(n27416), .B(n22479), .Z(n27417) );
  XOR U29468 ( .A(n27419), .B(n27420), .Z(n27416) );
  AND U29469 ( .A(n27421), .B(n27422), .Z(n27419) );
  XOR U29470 ( .A(n[831]), .B(n27420), .Z(n27422) );
  XNOR U29471 ( .A(n27420), .B(n22484), .Z(n27421) );
  XOR U29472 ( .A(n27423), .B(n27424), .Z(n27420) );
  AND U29473 ( .A(n27425), .B(n27426), .Z(n27423) );
  XOR U29474 ( .A(n[830]), .B(n27424), .Z(n27426) );
  XNOR U29475 ( .A(n27424), .B(n22489), .Z(n27425) );
  XOR U29476 ( .A(n27427), .B(n27428), .Z(n27424) );
  AND U29477 ( .A(n27429), .B(n27430), .Z(n27427) );
  XOR U29478 ( .A(n[829]), .B(n27428), .Z(n27430) );
  XNOR U29479 ( .A(n27428), .B(n22494), .Z(n27429) );
  XOR U29480 ( .A(n27431), .B(n27432), .Z(n27428) );
  AND U29481 ( .A(n27433), .B(n27434), .Z(n27431) );
  XOR U29482 ( .A(n[828]), .B(n27432), .Z(n27434) );
  XNOR U29483 ( .A(n27432), .B(n22499), .Z(n27433) );
  XOR U29484 ( .A(n27435), .B(n27436), .Z(n27432) );
  AND U29485 ( .A(n27437), .B(n27438), .Z(n27435) );
  XOR U29486 ( .A(n[827]), .B(n27436), .Z(n27438) );
  XNOR U29487 ( .A(n27436), .B(n22504), .Z(n27437) );
  XOR U29488 ( .A(n27439), .B(n27440), .Z(n27436) );
  AND U29489 ( .A(n27441), .B(n27442), .Z(n27439) );
  XOR U29490 ( .A(n[826]), .B(n27440), .Z(n27442) );
  XNOR U29491 ( .A(n27440), .B(n22509), .Z(n27441) );
  XOR U29492 ( .A(n27443), .B(n27444), .Z(n27440) );
  AND U29493 ( .A(n27445), .B(n27446), .Z(n27443) );
  XOR U29494 ( .A(n[825]), .B(n27444), .Z(n27446) );
  XNOR U29495 ( .A(n27444), .B(n22514), .Z(n27445) );
  XOR U29496 ( .A(n27447), .B(n27448), .Z(n27444) );
  AND U29497 ( .A(n27449), .B(n27450), .Z(n27447) );
  XOR U29498 ( .A(n[824]), .B(n27448), .Z(n27450) );
  XNOR U29499 ( .A(n27448), .B(n22519), .Z(n27449) );
  XOR U29500 ( .A(n27451), .B(n27452), .Z(n27448) );
  AND U29501 ( .A(n27453), .B(n27454), .Z(n27451) );
  XOR U29502 ( .A(n[823]), .B(n27452), .Z(n27454) );
  XNOR U29503 ( .A(n27452), .B(n22524), .Z(n27453) );
  XOR U29504 ( .A(n27455), .B(n27456), .Z(n27452) );
  AND U29505 ( .A(n27457), .B(n27458), .Z(n27455) );
  XOR U29506 ( .A(n[822]), .B(n27456), .Z(n27458) );
  XNOR U29507 ( .A(n27456), .B(n22529), .Z(n27457) );
  XOR U29508 ( .A(n27459), .B(n27460), .Z(n27456) );
  AND U29509 ( .A(n27461), .B(n27462), .Z(n27459) );
  XOR U29510 ( .A(n[821]), .B(n27460), .Z(n27462) );
  XNOR U29511 ( .A(n27460), .B(n22534), .Z(n27461) );
  XOR U29512 ( .A(n27463), .B(n27464), .Z(n27460) );
  AND U29513 ( .A(n27465), .B(n27466), .Z(n27463) );
  XOR U29514 ( .A(n[820]), .B(n27464), .Z(n27466) );
  XNOR U29515 ( .A(n27464), .B(n22539), .Z(n27465) );
  XOR U29516 ( .A(n27467), .B(n27468), .Z(n27464) );
  AND U29517 ( .A(n27469), .B(n27470), .Z(n27467) );
  XOR U29518 ( .A(n[819]), .B(n27468), .Z(n27470) );
  XNOR U29519 ( .A(n27468), .B(n22544), .Z(n27469) );
  XOR U29520 ( .A(n27471), .B(n27472), .Z(n27468) );
  AND U29521 ( .A(n27473), .B(n27474), .Z(n27471) );
  XOR U29522 ( .A(n[818]), .B(n27472), .Z(n27474) );
  XNOR U29523 ( .A(n27472), .B(n22549), .Z(n27473) );
  XOR U29524 ( .A(n27475), .B(n27476), .Z(n27472) );
  AND U29525 ( .A(n27477), .B(n27478), .Z(n27475) );
  XOR U29526 ( .A(n[817]), .B(n27476), .Z(n27478) );
  XNOR U29527 ( .A(n27476), .B(n22554), .Z(n27477) );
  XOR U29528 ( .A(n27479), .B(n27480), .Z(n27476) );
  AND U29529 ( .A(n27481), .B(n27482), .Z(n27479) );
  XOR U29530 ( .A(n[816]), .B(n27480), .Z(n27482) );
  XNOR U29531 ( .A(n27480), .B(n22559), .Z(n27481) );
  XOR U29532 ( .A(n27483), .B(n27484), .Z(n27480) );
  AND U29533 ( .A(n27485), .B(n27486), .Z(n27483) );
  XOR U29534 ( .A(n[815]), .B(n27484), .Z(n27486) );
  XNOR U29535 ( .A(n27484), .B(n22564), .Z(n27485) );
  XOR U29536 ( .A(n27487), .B(n27488), .Z(n27484) );
  AND U29537 ( .A(n27489), .B(n27490), .Z(n27487) );
  XOR U29538 ( .A(n[814]), .B(n27488), .Z(n27490) );
  XNOR U29539 ( .A(n27488), .B(n22569), .Z(n27489) );
  XOR U29540 ( .A(n27491), .B(n27492), .Z(n27488) );
  AND U29541 ( .A(n27493), .B(n27494), .Z(n27491) );
  XOR U29542 ( .A(n[813]), .B(n27492), .Z(n27494) );
  XNOR U29543 ( .A(n27492), .B(n22574), .Z(n27493) );
  XOR U29544 ( .A(n27495), .B(n27496), .Z(n27492) );
  AND U29545 ( .A(n27497), .B(n27498), .Z(n27495) );
  XOR U29546 ( .A(n[812]), .B(n27496), .Z(n27498) );
  XNOR U29547 ( .A(n27496), .B(n22579), .Z(n27497) );
  XOR U29548 ( .A(n27499), .B(n27500), .Z(n27496) );
  AND U29549 ( .A(n27501), .B(n27502), .Z(n27499) );
  XOR U29550 ( .A(n[811]), .B(n27500), .Z(n27502) );
  XNOR U29551 ( .A(n27500), .B(n22584), .Z(n27501) );
  XOR U29552 ( .A(n27503), .B(n27504), .Z(n27500) );
  AND U29553 ( .A(n27505), .B(n27506), .Z(n27503) );
  XOR U29554 ( .A(n[810]), .B(n27504), .Z(n27506) );
  XNOR U29555 ( .A(n27504), .B(n22589), .Z(n27505) );
  XOR U29556 ( .A(n27507), .B(n27508), .Z(n27504) );
  AND U29557 ( .A(n27509), .B(n27510), .Z(n27507) );
  XOR U29558 ( .A(n[809]), .B(n27508), .Z(n27510) );
  XNOR U29559 ( .A(n27508), .B(n22594), .Z(n27509) );
  XOR U29560 ( .A(n27511), .B(n27512), .Z(n27508) );
  AND U29561 ( .A(n27513), .B(n27514), .Z(n27511) );
  XOR U29562 ( .A(n[808]), .B(n27512), .Z(n27514) );
  XNOR U29563 ( .A(n27512), .B(n22599), .Z(n27513) );
  XOR U29564 ( .A(n27515), .B(n27516), .Z(n27512) );
  AND U29565 ( .A(n27517), .B(n27518), .Z(n27515) );
  XOR U29566 ( .A(n[807]), .B(n27516), .Z(n27518) );
  XNOR U29567 ( .A(n27516), .B(n22604), .Z(n27517) );
  XOR U29568 ( .A(n27519), .B(n27520), .Z(n27516) );
  AND U29569 ( .A(n27521), .B(n27522), .Z(n27519) );
  XOR U29570 ( .A(n[806]), .B(n27520), .Z(n27522) );
  XNOR U29571 ( .A(n27520), .B(n22609), .Z(n27521) );
  XOR U29572 ( .A(n27523), .B(n27524), .Z(n27520) );
  AND U29573 ( .A(n27525), .B(n27526), .Z(n27523) );
  XOR U29574 ( .A(n[805]), .B(n27524), .Z(n27526) );
  XNOR U29575 ( .A(n27524), .B(n22614), .Z(n27525) );
  XOR U29576 ( .A(n27527), .B(n27528), .Z(n27524) );
  AND U29577 ( .A(n27529), .B(n27530), .Z(n27527) );
  XOR U29578 ( .A(n[804]), .B(n27528), .Z(n27530) );
  XNOR U29579 ( .A(n27528), .B(n22619), .Z(n27529) );
  XOR U29580 ( .A(n27531), .B(n27532), .Z(n27528) );
  AND U29581 ( .A(n27533), .B(n27534), .Z(n27531) );
  XOR U29582 ( .A(n[803]), .B(n27532), .Z(n27534) );
  XNOR U29583 ( .A(n27532), .B(n22624), .Z(n27533) );
  XOR U29584 ( .A(n27535), .B(n27536), .Z(n27532) );
  AND U29585 ( .A(n27537), .B(n27538), .Z(n27535) );
  XOR U29586 ( .A(n[802]), .B(n27536), .Z(n27538) );
  XNOR U29587 ( .A(n27536), .B(n22629), .Z(n27537) );
  XOR U29588 ( .A(n27539), .B(n27540), .Z(n27536) );
  AND U29589 ( .A(n27541), .B(n27542), .Z(n27539) );
  XOR U29590 ( .A(n[801]), .B(n27540), .Z(n27542) );
  XNOR U29591 ( .A(n27540), .B(n22634), .Z(n27541) );
  XOR U29592 ( .A(n27543), .B(n27544), .Z(n27540) );
  AND U29593 ( .A(n27545), .B(n27546), .Z(n27543) );
  XOR U29594 ( .A(n[800]), .B(n27544), .Z(n27546) );
  XNOR U29595 ( .A(n27544), .B(n22639), .Z(n27545) );
  XOR U29596 ( .A(n27547), .B(n27548), .Z(n27544) );
  AND U29597 ( .A(n27549), .B(n27550), .Z(n27547) );
  XOR U29598 ( .A(n[799]), .B(n27548), .Z(n27550) );
  XNOR U29599 ( .A(n27548), .B(n22644), .Z(n27549) );
  XOR U29600 ( .A(n27551), .B(n27552), .Z(n27548) );
  AND U29601 ( .A(n27553), .B(n27554), .Z(n27551) );
  XOR U29602 ( .A(n[798]), .B(n27552), .Z(n27554) );
  XNOR U29603 ( .A(n27552), .B(n22649), .Z(n27553) );
  XOR U29604 ( .A(n27555), .B(n27556), .Z(n27552) );
  AND U29605 ( .A(n27557), .B(n27558), .Z(n27555) );
  XOR U29606 ( .A(n[797]), .B(n27556), .Z(n27558) );
  XNOR U29607 ( .A(n27556), .B(n22654), .Z(n27557) );
  XOR U29608 ( .A(n27559), .B(n27560), .Z(n27556) );
  AND U29609 ( .A(n27561), .B(n27562), .Z(n27559) );
  XOR U29610 ( .A(n[796]), .B(n27560), .Z(n27562) );
  XNOR U29611 ( .A(n27560), .B(n22659), .Z(n27561) );
  XOR U29612 ( .A(n27563), .B(n27564), .Z(n27560) );
  AND U29613 ( .A(n27565), .B(n27566), .Z(n27563) );
  XOR U29614 ( .A(n[795]), .B(n27564), .Z(n27566) );
  XNOR U29615 ( .A(n27564), .B(n22664), .Z(n27565) );
  XOR U29616 ( .A(n27567), .B(n27568), .Z(n27564) );
  AND U29617 ( .A(n27569), .B(n27570), .Z(n27567) );
  XOR U29618 ( .A(n[794]), .B(n27568), .Z(n27570) );
  XNOR U29619 ( .A(n27568), .B(n22669), .Z(n27569) );
  XOR U29620 ( .A(n27571), .B(n27572), .Z(n27568) );
  AND U29621 ( .A(n27573), .B(n27574), .Z(n27571) );
  XOR U29622 ( .A(n[793]), .B(n27572), .Z(n27574) );
  XNOR U29623 ( .A(n27572), .B(n22674), .Z(n27573) );
  XOR U29624 ( .A(n27575), .B(n27576), .Z(n27572) );
  AND U29625 ( .A(n27577), .B(n27578), .Z(n27575) );
  XOR U29626 ( .A(n[792]), .B(n27576), .Z(n27578) );
  XNOR U29627 ( .A(n27576), .B(n22679), .Z(n27577) );
  XOR U29628 ( .A(n27579), .B(n27580), .Z(n27576) );
  AND U29629 ( .A(n27581), .B(n27582), .Z(n27579) );
  XOR U29630 ( .A(n[791]), .B(n27580), .Z(n27582) );
  XNOR U29631 ( .A(n27580), .B(n22684), .Z(n27581) );
  XOR U29632 ( .A(n27583), .B(n27584), .Z(n27580) );
  AND U29633 ( .A(n27585), .B(n27586), .Z(n27583) );
  XOR U29634 ( .A(n[790]), .B(n27584), .Z(n27586) );
  XNOR U29635 ( .A(n27584), .B(n22689), .Z(n27585) );
  XOR U29636 ( .A(n27587), .B(n27588), .Z(n27584) );
  AND U29637 ( .A(n27589), .B(n27590), .Z(n27587) );
  XOR U29638 ( .A(n[789]), .B(n27588), .Z(n27590) );
  XNOR U29639 ( .A(n27588), .B(n22694), .Z(n27589) );
  XOR U29640 ( .A(n27591), .B(n27592), .Z(n27588) );
  AND U29641 ( .A(n27593), .B(n27594), .Z(n27591) );
  XOR U29642 ( .A(n[788]), .B(n27592), .Z(n27594) );
  XNOR U29643 ( .A(n27592), .B(n22699), .Z(n27593) );
  XOR U29644 ( .A(n27595), .B(n27596), .Z(n27592) );
  AND U29645 ( .A(n27597), .B(n27598), .Z(n27595) );
  XOR U29646 ( .A(n[787]), .B(n27596), .Z(n27598) );
  XNOR U29647 ( .A(n27596), .B(n22704), .Z(n27597) );
  XOR U29648 ( .A(n27599), .B(n27600), .Z(n27596) );
  AND U29649 ( .A(n27601), .B(n27602), .Z(n27599) );
  XOR U29650 ( .A(n[786]), .B(n27600), .Z(n27602) );
  XNOR U29651 ( .A(n27600), .B(n22709), .Z(n27601) );
  XOR U29652 ( .A(n27603), .B(n27604), .Z(n27600) );
  AND U29653 ( .A(n27605), .B(n27606), .Z(n27603) );
  XOR U29654 ( .A(n[785]), .B(n27604), .Z(n27606) );
  XNOR U29655 ( .A(n27604), .B(n22714), .Z(n27605) );
  XOR U29656 ( .A(n27607), .B(n27608), .Z(n27604) );
  AND U29657 ( .A(n27609), .B(n27610), .Z(n27607) );
  XOR U29658 ( .A(n[784]), .B(n27608), .Z(n27610) );
  XNOR U29659 ( .A(n27608), .B(n22719), .Z(n27609) );
  XOR U29660 ( .A(n27611), .B(n27612), .Z(n27608) );
  AND U29661 ( .A(n27613), .B(n27614), .Z(n27611) );
  XOR U29662 ( .A(n[783]), .B(n27612), .Z(n27614) );
  XNOR U29663 ( .A(n27612), .B(n22724), .Z(n27613) );
  XOR U29664 ( .A(n27615), .B(n27616), .Z(n27612) );
  AND U29665 ( .A(n27617), .B(n27618), .Z(n27615) );
  XOR U29666 ( .A(n[782]), .B(n27616), .Z(n27618) );
  XNOR U29667 ( .A(n27616), .B(n22729), .Z(n27617) );
  XOR U29668 ( .A(n27619), .B(n27620), .Z(n27616) );
  AND U29669 ( .A(n27621), .B(n27622), .Z(n27619) );
  XOR U29670 ( .A(n[781]), .B(n27620), .Z(n27622) );
  XNOR U29671 ( .A(n27620), .B(n22734), .Z(n27621) );
  XOR U29672 ( .A(n27623), .B(n27624), .Z(n27620) );
  AND U29673 ( .A(n27625), .B(n27626), .Z(n27623) );
  XOR U29674 ( .A(n[780]), .B(n27624), .Z(n27626) );
  XNOR U29675 ( .A(n27624), .B(n22739), .Z(n27625) );
  XOR U29676 ( .A(n27627), .B(n27628), .Z(n27624) );
  AND U29677 ( .A(n27629), .B(n27630), .Z(n27627) );
  XOR U29678 ( .A(n[779]), .B(n27628), .Z(n27630) );
  XNOR U29679 ( .A(n27628), .B(n22744), .Z(n27629) );
  XOR U29680 ( .A(n27631), .B(n27632), .Z(n27628) );
  AND U29681 ( .A(n27633), .B(n27634), .Z(n27631) );
  XOR U29682 ( .A(n[778]), .B(n27632), .Z(n27634) );
  XNOR U29683 ( .A(n27632), .B(n22749), .Z(n27633) );
  XOR U29684 ( .A(n27635), .B(n27636), .Z(n27632) );
  AND U29685 ( .A(n27637), .B(n27638), .Z(n27635) );
  XOR U29686 ( .A(n[777]), .B(n27636), .Z(n27638) );
  XNOR U29687 ( .A(n27636), .B(n22754), .Z(n27637) );
  XOR U29688 ( .A(n27639), .B(n27640), .Z(n27636) );
  AND U29689 ( .A(n27641), .B(n27642), .Z(n27639) );
  XOR U29690 ( .A(n[776]), .B(n27640), .Z(n27642) );
  XNOR U29691 ( .A(n27640), .B(n22759), .Z(n27641) );
  XOR U29692 ( .A(n27643), .B(n27644), .Z(n27640) );
  AND U29693 ( .A(n27645), .B(n27646), .Z(n27643) );
  XOR U29694 ( .A(n[775]), .B(n27644), .Z(n27646) );
  XNOR U29695 ( .A(n27644), .B(n22764), .Z(n27645) );
  XOR U29696 ( .A(n27647), .B(n27648), .Z(n27644) );
  AND U29697 ( .A(n27649), .B(n27650), .Z(n27647) );
  XOR U29698 ( .A(n[774]), .B(n27648), .Z(n27650) );
  XNOR U29699 ( .A(n27648), .B(n22769), .Z(n27649) );
  XOR U29700 ( .A(n27651), .B(n27652), .Z(n27648) );
  AND U29701 ( .A(n27653), .B(n27654), .Z(n27651) );
  XOR U29702 ( .A(n[773]), .B(n27652), .Z(n27654) );
  XNOR U29703 ( .A(n27652), .B(n22774), .Z(n27653) );
  XOR U29704 ( .A(n27655), .B(n27656), .Z(n27652) );
  AND U29705 ( .A(n27657), .B(n27658), .Z(n27655) );
  XOR U29706 ( .A(n[772]), .B(n27656), .Z(n27658) );
  XNOR U29707 ( .A(n27656), .B(n22779), .Z(n27657) );
  XOR U29708 ( .A(n27659), .B(n27660), .Z(n27656) );
  AND U29709 ( .A(n27661), .B(n27662), .Z(n27659) );
  XOR U29710 ( .A(n[771]), .B(n27660), .Z(n27662) );
  XNOR U29711 ( .A(n27660), .B(n22784), .Z(n27661) );
  XOR U29712 ( .A(n27663), .B(n27664), .Z(n27660) );
  AND U29713 ( .A(n27665), .B(n27666), .Z(n27663) );
  XOR U29714 ( .A(n[770]), .B(n27664), .Z(n27666) );
  XNOR U29715 ( .A(n27664), .B(n22789), .Z(n27665) );
  XOR U29716 ( .A(n27667), .B(n27668), .Z(n27664) );
  AND U29717 ( .A(n27669), .B(n27670), .Z(n27667) );
  XOR U29718 ( .A(n[769]), .B(n27668), .Z(n27670) );
  XNOR U29719 ( .A(n27668), .B(n22794), .Z(n27669) );
  XOR U29720 ( .A(n27671), .B(n27672), .Z(n27668) );
  AND U29721 ( .A(n27673), .B(n27674), .Z(n27671) );
  XOR U29722 ( .A(n[768]), .B(n27672), .Z(n27674) );
  XNOR U29723 ( .A(n27672), .B(n22799), .Z(n27673) );
  XOR U29724 ( .A(n27675), .B(n27676), .Z(n27672) );
  AND U29725 ( .A(n27677), .B(n27678), .Z(n27675) );
  XOR U29726 ( .A(n[767]), .B(n27676), .Z(n27678) );
  XNOR U29727 ( .A(n27676), .B(n22804), .Z(n27677) );
  XOR U29728 ( .A(n27679), .B(n27680), .Z(n27676) );
  AND U29729 ( .A(n27681), .B(n27682), .Z(n27679) );
  XOR U29730 ( .A(n[766]), .B(n27680), .Z(n27682) );
  XNOR U29731 ( .A(n27680), .B(n22809), .Z(n27681) );
  XOR U29732 ( .A(n27683), .B(n27684), .Z(n27680) );
  AND U29733 ( .A(n27685), .B(n27686), .Z(n27683) );
  XOR U29734 ( .A(n[765]), .B(n27684), .Z(n27686) );
  XNOR U29735 ( .A(n27684), .B(n22814), .Z(n27685) );
  XOR U29736 ( .A(n27687), .B(n27688), .Z(n27684) );
  AND U29737 ( .A(n27689), .B(n27690), .Z(n27687) );
  XOR U29738 ( .A(n[764]), .B(n27688), .Z(n27690) );
  XNOR U29739 ( .A(n27688), .B(n22819), .Z(n27689) );
  XOR U29740 ( .A(n27691), .B(n27692), .Z(n27688) );
  AND U29741 ( .A(n27693), .B(n27694), .Z(n27691) );
  XOR U29742 ( .A(n[763]), .B(n27692), .Z(n27694) );
  XNOR U29743 ( .A(n27692), .B(n22824), .Z(n27693) );
  XOR U29744 ( .A(n27695), .B(n27696), .Z(n27692) );
  AND U29745 ( .A(n27697), .B(n27698), .Z(n27695) );
  XOR U29746 ( .A(n[762]), .B(n27696), .Z(n27698) );
  XNOR U29747 ( .A(n27696), .B(n22829), .Z(n27697) );
  XOR U29748 ( .A(n27699), .B(n27700), .Z(n27696) );
  AND U29749 ( .A(n27701), .B(n27702), .Z(n27699) );
  XOR U29750 ( .A(n[761]), .B(n27700), .Z(n27702) );
  XNOR U29751 ( .A(n27700), .B(n22834), .Z(n27701) );
  XOR U29752 ( .A(n27703), .B(n27704), .Z(n27700) );
  AND U29753 ( .A(n27705), .B(n27706), .Z(n27703) );
  XOR U29754 ( .A(n[760]), .B(n27704), .Z(n27706) );
  XNOR U29755 ( .A(n27704), .B(n22839), .Z(n27705) );
  XOR U29756 ( .A(n27707), .B(n27708), .Z(n27704) );
  AND U29757 ( .A(n27709), .B(n27710), .Z(n27707) );
  XOR U29758 ( .A(n[759]), .B(n27708), .Z(n27710) );
  XNOR U29759 ( .A(n27708), .B(n22844), .Z(n27709) );
  XOR U29760 ( .A(n27711), .B(n27712), .Z(n27708) );
  AND U29761 ( .A(n27713), .B(n27714), .Z(n27711) );
  XOR U29762 ( .A(n[758]), .B(n27712), .Z(n27714) );
  XNOR U29763 ( .A(n27712), .B(n22849), .Z(n27713) );
  XOR U29764 ( .A(n27715), .B(n27716), .Z(n27712) );
  AND U29765 ( .A(n27717), .B(n27718), .Z(n27715) );
  XOR U29766 ( .A(n[757]), .B(n27716), .Z(n27718) );
  XNOR U29767 ( .A(n27716), .B(n22854), .Z(n27717) );
  XOR U29768 ( .A(n27719), .B(n27720), .Z(n27716) );
  AND U29769 ( .A(n27721), .B(n27722), .Z(n27719) );
  XOR U29770 ( .A(n[756]), .B(n27720), .Z(n27722) );
  XNOR U29771 ( .A(n27720), .B(n22859), .Z(n27721) );
  XOR U29772 ( .A(n27723), .B(n27724), .Z(n27720) );
  AND U29773 ( .A(n27725), .B(n27726), .Z(n27723) );
  XOR U29774 ( .A(n[755]), .B(n27724), .Z(n27726) );
  XNOR U29775 ( .A(n27724), .B(n22864), .Z(n27725) );
  XOR U29776 ( .A(n27727), .B(n27728), .Z(n27724) );
  AND U29777 ( .A(n27729), .B(n27730), .Z(n27727) );
  XOR U29778 ( .A(n[754]), .B(n27728), .Z(n27730) );
  XNOR U29779 ( .A(n27728), .B(n22869), .Z(n27729) );
  XOR U29780 ( .A(n27731), .B(n27732), .Z(n27728) );
  AND U29781 ( .A(n27733), .B(n27734), .Z(n27731) );
  XOR U29782 ( .A(n[753]), .B(n27732), .Z(n27734) );
  XNOR U29783 ( .A(n27732), .B(n22874), .Z(n27733) );
  XOR U29784 ( .A(n27735), .B(n27736), .Z(n27732) );
  AND U29785 ( .A(n27737), .B(n27738), .Z(n27735) );
  XOR U29786 ( .A(n[752]), .B(n27736), .Z(n27738) );
  XNOR U29787 ( .A(n27736), .B(n22879), .Z(n27737) );
  XOR U29788 ( .A(n27739), .B(n27740), .Z(n27736) );
  AND U29789 ( .A(n27741), .B(n27742), .Z(n27739) );
  XOR U29790 ( .A(n[751]), .B(n27740), .Z(n27742) );
  XNOR U29791 ( .A(n27740), .B(n22884), .Z(n27741) );
  XOR U29792 ( .A(n27743), .B(n27744), .Z(n27740) );
  AND U29793 ( .A(n27745), .B(n27746), .Z(n27743) );
  XOR U29794 ( .A(n[750]), .B(n27744), .Z(n27746) );
  XNOR U29795 ( .A(n27744), .B(n22889), .Z(n27745) );
  XOR U29796 ( .A(n27747), .B(n27748), .Z(n27744) );
  AND U29797 ( .A(n27749), .B(n27750), .Z(n27747) );
  XOR U29798 ( .A(n[749]), .B(n27748), .Z(n27750) );
  XNOR U29799 ( .A(n27748), .B(n22894), .Z(n27749) );
  XOR U29800 ( .A(n27751), .B(n27752), .Z(n27748) );
  AND U29801 ( .A(n27753), .B(n27754), .Z(n27751) );
  XOR U29802 ( .A(n[748]), .B(n27752), .Z(n27754) );
  XNOR U29803 ( .A(n27752), .B(n22899), .Z(n27753) );
  XOR U29804 ( .A(n27755), .B(n27756), .Z(n27752) );
  AND U29805 ( .A(n27757), .B(n27758), .Z(n27755) );
  XOR U29806 ( .A(n[747]), .B(n27756), .Z(n27758) );
  XNOR U29807 ( .A(n27756), .B(n22904), .Z(n27757) );
  XOR U29808 ( .A(n27759), .B(n27760), .Z(n27756) );
  AND U29809 ( .A(n27761), .B(n27762), .Z(n27759) );
  XOR U29810 ( .A(n[746]), .B(n27760), .Z(n27762) );
  XNOR U29811 ( .A(n27760), .B(n22909), .Z(n27761) );
  XOR U29812 ( .A(n27763), .B(n27764), .Z(n27760) );
  AND U29813 ( .A(n27765), .B(n27766), .Z(n27763) );
  XOR U29814 ( .A(n[745]), .B(n27764), .Z(n27766) );
  XNOR U29815 ( .A(n27764), .B(n22914), .Z(n27765) );
  XOR U29816 ( .A(n27767), .B(n27768), .Z(n27764) );
  AND U29817 ( .A(n27769), .B(n27770), .Z(n27767) );
  XOR U29818 ( .A(n[744]), .B(n27768), .Z(n27770) );
  XNOR U29819 ( .A(n27768), .B(n22919), .Z(n27769) );
  XOR U29820 ( .A(n27771), .B(n27772), .Z(n27768) );
  AND U29821 ( .A(n27773), .B(n27774), .Z(n27771) );
  XOR U29822 ( .A(n[743]), .B(n27772), .Z(n27774) );
  XNOR U29823 ( .A(n27772), .B(n22924), .Z(n27773) );
  XOR U29824 ( .A(n27775), .B(n27776), .Z(n27772) );
  AND U29825 ( .A(n27777), .B(n27778), .Z(n27775) );
  XOR U29826 ( .A(n[742]), .B(n27776), .Z(n27778) );
  XNOR U29827 ( .A(n27776), .B(n22929), .Z(n27777) );
  XOR U29828 ( .A(n27779), .B(n27780), .Z(n27776) );
  AND U29829 ( .A(n27781), .B(n27782), .Z(n27779) );
  XOR U29830 ( .A(n[741]), .B(n27780), .Z(n27782) );
  XNOR U29831 ( .A(n27780), .B(n22934), .Z(n27781) );
  XOR U29832 ( .A(n27783), .B(n27784), .Z(n27780) );
  AND U29833 ( .A(n27785), .B(n27786), .Z(n27783) );
  XOR U29834 ( .A(n[740]), .B(n27784), .Z(n27786) );
  XNOR U29835 ( .A(n27784), .B(n22939), .Z(n27785) );
  XOR U29836 ( .A(n27787), .B(n27788), .Z(n27784) );
  AND U29837 ( .A(n27789), .B(n27790), .Z(n27787) );
  XOR U29838 ( .A(n[739]), .B(n27788), .Z(n27790) );
  XNOR U29839 ( .A(n27788), .B(n22944), .Z(n27789) );
  XOR U29840 ( .A(n27791), .B(n27792), .Z(n27788) );
  AND U29841 ( .A(n27793), .B(n27794), .Z(n27791) );
  XOR U29842 ( .A(n[738]), .B(n27792), .Z(n27794) );
  XNOR U29843 ( .A(n27792), .B(n22949), .Z(n27793) );
  XOR U29844 ( .A(n27795), .B(n27796), .Z(n27792) );
  AND U29845 ( .A(n27797), .B(n27798), .Z(n27795) );
  XOR U29846 ( .A(n[737]), .B(n27796), .Z(n27798) );
  XNOR U29847 ( .A(n27796), .B(n22954), .Z(n27797) );
  XOR U29848 ( .A(n27799), .B(n27800), .Z(n27796) );
  AND U29849 ( .A(n27801), .B(n27802), .Z(n27799) );
  XOR U29850 ( .A(n[736]), .B(n27800), .Z(n27802) );
  XNOR U29851 ( .A(n27800), .B(n22959), .Z(n27801) );
  XOR U29852 ( .A(n27803), .B(n27804), .Z(n27800) );
  AND U29853 ( .A(n27805), .B(n27806), .Z(n27803) );
  XOR U29854 ( .A(n[735]), .B(n27804), .Z(n27806) );
  XNOR U29855 ( .A(n27804), .B(n22964), .Z(n27805) );
  XOR U29856 ( .A(n27807), .B(n27808), .Z(n27804) );
  AND U29857 ( .A(n27809), .B(n27810), .Z(n27807) );
  XOR U29858 ( .A(n[734]), .B(n27808), .Z(n27810) );
  XNOR U29859 ( .A(n27808), .B(n22969), .Z(n27809) );
  XOR U29860 ( .A(n27811), .B(n27812), .Z(n27808) );
  AND U29861 ( .A(n27813), .B(n27814), .Z(n27811) );
  XOR U29862 ( .A(n[733]), .B(n27812), .Z(n27814) );
  XNOR U29863 ( .A(n27812), .B(n22974), .Z(n27813) );
  XOR U29864 ( .A(n27815), .B(n27816), .Z(n27812) );
  AND U29865 ( .A(n27817), .B(n27818), .Z(n27815) );
  XOR U29866 ( .A(n[732]), .B(n27816), .Z(n27818) );
  XNOR U29867 ( .A(n27816), .B(n22979), .Z(n27817) );
  XOR U29868 ( .A(n27819), .B(n27820), .Z(n27816) );
  AND U29869 ( .A(n27821), .B(n27822), .Z(n27819) );
  XOR U29870 ( .A(n[731]), .B(n27820), .Z(n27822) );
  XNOR U29871 ( .A(n27820), .B(n22984), .Z(n27821) );
  XOR U29872 ( .A(n27823), .B(n27824), .Z(n27820) );
  AND U29873 ( .A(n27825), .B(n27826), .Z(n27823) );
  XOR U29874 ( .A(n[730]), .B(n27824), .Z(n27826) );
  XNOR U29875 ( .A(n27824), .B(n22989), .Z(n27825) );
  XOR U29876 ( .A(n27827), .B(n27828), .Z(n27824) );
  AND U29877 ( .A(n27829), .B(n27830), .Z(n27827) );
  XOR U29878 ( .A(n[729]), .B(n27828), .Z(n27830) );
  XNOR U29879 ( .A(n27828), .B(n22994), .Z(n27829) );
  XOR U29880 ( .A(n27831), .B(n27832), .Z(n27828) );
  AND U29881 ( .A(n27833), .B(n27834), .Z(n27831) );
  XOR U29882 ( .A(n[728]), .B(n27832), .Z(n27834) );
  XNOR U29883 ( .A(n27832), .B(n22999), .Z(n27833) );
  XOR U29884 ( .A(n27835), .B(n27836), .Z(n27832) );
  AND U29885 ( .A(n27837), .B(n27838), .Z(n27835) );
  XOR U29886 ( .A(n[727]), .B(n27836), .Z(n27838) );
  XNOR U29887 ( .A(n27836), .B(n23004), .Z(n27837) );
  XOR U29888 ( .A(n27839), .B(n27840), .Z(n27836) );
  AND U29889 ( .A(n27841), .B(n27842), .Z(n27839) );
  XOR U29890 ( .A(n[726]), .B(n27840), .Z(n27842) );
  XNOR U29891 ( .A(n27840), .B(n23009), .Z(n27841) );
  XOR U29892 ( .A(n27843), .B(n27844), .Z(n27840) );
  AND U29893 ( .A(n27845), .B(n27846), .Z(n27843) );
  XOR U29894 ( .A(n[725]), .B(n27844), .Z(n27846) );
  XNOR U29895 ( .A(n27844), .B(n23014), .Z(n27845) );
  XOR U29896 ( .A(n27847), .B(n27848), .Z(n27844) );
  AND U29897 ( .A(n27849), .B(n27850), .Z(n27847) );
  XOR U29898 ( .A(n[724]), .B(n27848), .Z(n27850) );
  XNOR U29899 ( .A(n27848), .B(n23019), .Z(n27849) );
  XOR U29900 ( .A(n27851), .B(n27852), .Z(n27848) );
  AND U29901 ( .A(n27853), .B(n27854), .Z(n27851) );
  XOR U29902 ( .A(n[723]), .B(n27852), .Z(n27854) );
  XNOR U29903 ( .A(n27852), .B(n23024), .Z(n27853) );
  XOR U29904 ( .A(n27855), .B(n27856), .Z(n27852) );
  AND U29905 ( .A(n27857), .B(n27858), .Z(n27855) );
  XOR U29906 ( .A(n[722]), .B(n27856), .Z(n27858) );
  XNOR U29907 ( .A(n27856), .B(n23029), .Z(n27857) );
  XOR U29908 ( .A(n27859), .B(n27860), .Z(n27856) );
  AND U29909 ( .A(n27861), .B(n27862), .Z(n27859) );
  XOR U29910 ( .A(n[721]), .B(n27860), .Z(n27862) );
  XNOR U29911 ( .A(n27860), .B(n23034), .Z(n27861) );
  XOR U29912 ( .A(n27863), .B(n27864), .Z(n27860) );
  AND U29913 ( .A(n27865), .B(n27866), .Z(n27863) );
  XOR U29914 ( .A(n[720]), .B(n27864), .Z(n27866) );
  XNOR U29915 ( .A(n27864), .B(n23039), .Z(n27865) );
  XOR U29916 ( .A(n27867), .B(n27868), .Z(n27864) );
  AND U29917 ( .A(n27869), .B(n27870), .Z(n27867) );
  XOR U29918 ( .A(n[719]), .B(n27868), .Z(n27870) );
  XNOR U29919 ( .A(n27868), .B(n23044), .Z(n27869) );
  XOR U29920 ( .A(n27871), .B(n27872), .Z(n27868) );
  AND U29921 ( .A(n27873), .B(n27874), .Z(n27871) );
  XOR U29922 ( .A(n[718]), .B(n27872), .Z(n27874) );
  XNOR U29923 ( .A(n27872), .B(n23049), .Z(n27873) );
  XOR U29924 ( .A(n27875), .B(n27876), .Z(n27872) );
  AND U29925 ( .A(n27877), .B(n27878), .Z(n27875) );
  XOR U29926 ( .A(n[717]), .B(n27876), .Z(n27878) );
  XNOR U29927 ( .A(n27876), .B(n23054), .Z(n27877) );
  XOR U29928 ( .A(n27879), .B(n27880), .Z(n27876) );
  AND U29929 ( .A(n27881), .B(n27882), .Z(n27879) );
  XOR U29930 ( .A(n[716]), .B(n27880), .Z(n27882) );
  XNOR U29931 ( .A(n27880), .B(n23059), .Z(n27881) );
  XOR U29932 ( .A(n27883), .B(n27884), .Z(n27880) );
  AND U29933 ( .A(n27885), .B(n27886), .Z(n27883) );
  XOR U29934 ( .A(n[715]), .B(n27884), .Z(n27886) );
  XNOR U29935 ( .A(n27884), .B(n23064), .Z(n27885) );
  XOR U29936 ( .A(n27887), .B(n27888), .Z(n27884) );
  AND U29937 ( .A(n27889), .B(n27890), .Z(n27887) );
  XOR U29938 ( .A(n[714]), .B(n27888), .Z(n27890) );
  XNOR U29939 ( .A(n27888), .B(n23069), .Z(n27889) );
  XOR U29940 ( .A(n27891), .B(n27892), .Z(n27888) );
  AND U29941 ( .A(n27893), .B(n27894), .Z(n27891) );
  XOR U29942 ( .A(n[713]), .B(n27892), .Z(n27894) );
  XNOR U29943 ( .A(n27892), .B(n23074), .Z(n27893) );
  XOR U29944 ( .A(n27895), .B(n27896), .Z(n27892) );
  AND U29945 ( .A(n27897), .B(n27898), .Z(n27895) );
  XOR U29946 ( .A(n[712]), .B(n27896), .Z(n27898) );
  XNOR U29947 ( .A(n27896), .B(n23079), .Z(n27897) );
  XOR U29948 ( .A(n27899), .B(n27900), .Z(n27896) );
  AND U29949 ( .A(n27901), .B(n27902), .Z(n27899) );
  XOR U29950 ( .A(n[711]), .B(n27900), .Z(n27902) );
  XNOR U29951 ( .A(n27900), .B(n23084), .Z(n27901) );
  XOR U29952 ( .A(n27903), .B(n27904), .Z(n27900) );
  AND U29953 ( .A(n27905), .B(n27906), .Z(n27903) );
  XOR U29954 ( .A(n[710]), .B(n27904), .Z(n27906) );
  XNOR U29955 ( .A(n27904), .B(n23089), .Z(n27905) );
  XOR U29956 ( .A(n27907), .B(n27908), .Z(n27904) );
  AND U29957 ( .A(n27909), .B(n27910), .Z(n27907) );
  XOR U29958 ( .A(n[709]), .B(n27908), .Z(n27910) );
  XNOR U29959 ( .A(n27908), .B(n23094), .Z(n27909) );
  XOR U29960 ( .A(n27911), .B(n27912), .Z(n27908) );
  AND U29961 ( .A(n27913), .B(n27914), .Z(n27911) );
  XOR U29962 ( .A(n[708]), .B(n27912), .Z(n27914) );
  XNOR U29963 ( .A(n27912), .B(n23099), .Z(n27913) );
  XOR U29964 ( .A(n27915), .B(n27916), .Z(n27912) );
  AND U29965 ( .A(n27917), .B(n27918), .Z(n27915) );
  XOR U29966 ( .A(n[707]), .B(n27916), .Z(n27918) );
  XNOR U29967 ( .A(n27916), .B(n23104), .Z(n27917) );
  XOR U29968 ( .A(n27919), .B(n27920), .Z(n27916) );
  AND U29969 ( .A(n27921), .B(n27922), .Z(n27919) );
  XOR U29970 ( .A(n[706]), .B(n27920), .Z(n27922) );
  XNOR U29971 ( .A(n27920), .B(n23109), .Z(n27921) );
  XOR U29972 ( .A(n27923), .B(n27924), .Z(n27920) );
  AND U29973 ( .A(n27925), .B(n27926), .Z(n27923) );
  XOR U29974 ( .A(n[705]), .B(n27924), .Z(n27926) );
  XNOR U29975 ( .A(n27924), .B(n23114), .Z(n27925) );
  XOR U29976 ( .A(n27927), .B(n27928), .Z(n27924) );
  AND U29977 ( .A(n27929), .B(n27930), .Z(n27927) );
  XOR U29978 ( .A(n[704]), .B(n27928), .Z(n27930) );
  XNOR U29979 ( .A(n27928), .B(n23119), .Z(n27929) );
  XOR U29980 ( .A(n27931), .B(n27932), .Z(n27928) );
  AND U29981 ( .A(n27933), .B(n27934), .Z(n27931) );
  XOR U29982 ( .A(n[703]), .B(n27932), .Z(n27934) );
  XNOR U29983 ( .A(n27932), .B(n23124), .Z(n27933) );
  XOR U29984 ( .A(n27935), .B(n27936), .Z(n27932) );
  AND U29985 ( .A(n27937), .B(n27938), .Z(n27935) );
  XOR U29986 ( .A(n[702]), .B(n27936), .Z(n27938) );
  XNOR U29987 ( .A(n27936), .B(n23129), .Z(n27937) );
  XOR U29988 ( .A(n27939), .B(n27940), .Z(n27936) );
  AND U29989 ( .A(n27941), .B(n27942), .Z(n27939) );
  XOR U29990 ( .A(n[701]), .B(n27940), .Z(n27942) );
  XNOR U29991 ( .A(n27940), .B(n23134), .Z(n27941) );
  XOR U29992 ( .A(n27943), .B(n27944), .Z(n27940) );
  AND U29993 ( .A(n27945), .B(n27946), .Z(n27943) );
  XOR U29994 ( .A(n[700]), .B(n27944), .Z(n27946) );
  XNOR U29995 ( .A(n27944), .B(n23139), .Z(n27945) );
  XOR U29996 ( .A(n27947), .B(n27948), .Z(n27944) );
  AND U29997 ( .A(n27949), .B(n27950), .Z(n27947) );
  XOR U29998 ( .A(n[699]), .B(n27948), .Z(n27950) );
  XNOR U29999 ( .A(n27948), .B(n23144), .Z(n27949) );
  XOR U30000 ( .A(n27951), .B(n27952), .Z(n27948) );
  AND U30001 ( .A(n27953), .B(n27954), .Z(n27951) );
  XOR U30002 ( .A(n[698]), .B(n27952), .Z(n27954) );
  XNOR U30003 ( .A(n27952), .B(n23149), .Z(n27953) );
  XOR U30004 ( .A(n27955), .B(n27956), .Z(n27952) );
  AND U30005 ( .A(n27957), .B(n27958), .Z(n27955) );
  XOR U30006 ( .A(n[697]), .B(n27956), .Z(n27958) );
  XNOR U30007 ( .A(n27956), .B(n23154), .Z(n27957) );
  XOR U30008 ( .A(n27959), .B(n27960), .Z(n27956) );
  AND U30009 ( .A(n27961), .B(n27962), .Z(n27959) );
  XOR U30010 ( .A(n[696]), .B(n27960), .Z(n27962) );
  XNOR U30011 ( .A(n27960), .B(n23159), .Z(n27961) );
  XOR U30012 ( .A(n27963), .B(n27964), .Z(n27960) );
  AND U30013 ( .A(n27965), .B(n27966), .Z(n27963) );
  XOR U30014 ( .A(n[695]), .B(n27964), .Z(n27966) );
  XNOR U30015 ( .A(n27964), .B(n23164), .Z(n27965) );
  XOR U30016 ( .A(n27967), .B(n27968), .Z(n27964) );
  AND U30017 ( .A(n27969), .B(n27970), .Z(n27967) );
  XOR U30018 ( .A(n[694]), .B(n27968), .Z(n27970) );
  XNOR U30019 ( .A(n27968), .B(n23169), .Z(n27969) );
  XOR U30020 ( .A(n27971), .B(n27972), .Z(n27968) );
  AND U30021 ( .A(n27973), .B(n27974), .Z(n27971) );
  XOR U30022 ( .A(n[693]), .B(n27972), .Z(n27974) );
  XNOR U30023 ( .A(n27972), .B(n23174), .Z(n27973) );
  XOR U30024 ( .A(n27975), .B(n27976), .Z(n27972) );
  AND U30025 ( .A(n27977), .B(n27978), .Z(n27975) );
  XOR U30026 ( .A(n[692]), .B(n27976), .Z(n27978) );
  XNOR U30027 ( .A(n27976), .B(n23179), .Z(n27977) );
  XOR U30028 ( .A(n27979), .B(n27980), .Z(n27976) );
  AND U30029 ( .A(n27981), .B(n27982), .Z(n27979) );
  XOR U30030 ( .A(n[691]), .B(n27980), .Z(n27982) );
  XNOR U30031 ( .A(n27980), .B(n23184), .Z(n27981) );
  XOR U30032 ( .A(n27983), .B(n27984), .Z(n27980) );
  AND U30033 ( .A(n27985), .B(n27986), .Z(n27983) );
  XOR U30034 ( .A(n[690]), .B(n27984), .Z(n27986) );
  XNOR U30035 ( .A(n27984), .B(n23189), .Z(n27985) );
  XOR U30036 ( .A(n27987), .B(n27988), .Z(n27984) );
  AND U30037 ( .A(n27989), .B(n27990), .Z(n27987) );
  XOR U30038 ( .A(n[689]), .B(n27988), .Z(n27990) );
  XNOR U30039 ( .A(n27988), .B(n23194), .Z(n27989) );
  XOR U30040 ( .A(n27991), .B(n27992), .Z(n27988) );
  AND U30041 ( .A(n27993), .B(n27994), .Z(n27991) );
  XOR U30042 ( .A(n[688]), .B(n27992), .Z(n27994) );
  XNOR U30043 ( .A(n27992), .B(n23199), .Z(n27993) );
  XOR U30044 ( .A(n27995), .B(n27996), .Z(n27992) );
  AND U30045 ( .A(n27997), .B(n27998), .Z(n27995) );
  XOR U30046 ( .A(n[687]), .B(n27996), .Z(n27998) );
  XNOR U30047 ( .A(n27996), .B(n23204), .Z(n27997) );
  XOR U30048 ( .A(n27999), .B(n28000), .Z(n27996) );
  AND U30049 ( .A(n28001), .B(n28002), .Z(n27999) );
  XOR U30050 ( .A(n[686]), .B(n28000), .Z(n28002) );
  XNOR U30051 ( .A(n28000), .B(n23209), .Z(n28001) );
  XOR U30052 ( .A(n28003), .B(n28004), .Z(n28000) );
  AND U30053 ( .A(n28005), .B(n28006), .Z(n28003) );
  XOR U30054 ( .A(n[685]), .B(n28004), .Z(n28006) );
  XNOR U30055 ( .A(n28004), .B(n23214), .Z(n28005) );
  XOR U30056 ( .A(n28007), .B(n28008), .Z(n28004) );
  AND U30057 ( .A(n28009), .B(n28010), .Z(n28007) );
  XOR U30058 ( .A(n[684]), .B(n28008), .Z(n28010) );
  XNOR U30059 ( .A(n28008), .B(n23219), .Z(n28009) );
  XOR U30060 ( .A(n28011), .B(n28012), .Z(n28008) );
  AND U30061 ( .A(n28013), .B(n28014), .Z(n28011) );
  XOR U30062 ( .A(n[683]), .B(n28012), .Z(n28014) );
  XNOR U30063 ( .A(n28012), .B(n23224), .Z(n28013) );
  XOR U30064 ( .A(n28015), .B(n28016), .Z(n28012) );
  AND U30065 ( .A(n28017), .B(n28018), .Z(n28015) );
  XOR U30066 ( .A(n[682]), .B(n28016), .Z(n28018) );
  XNOR U30067 ( .A(n28016), .B(n23229), .Z(n28017) );
  XOR U30068 ( .A(n28019), .B(n28020), .Z(n28016) );
  AND U30069 ( .A(n28021), .B(n28022), .Z(n28019) );
  XOR U30070 ( .A(n[681]), .B(n28020), .Z(n28022) );
  XNOR U30071 ( .A(n28020), .B(n23234), .Z(n28021) );
  XOR U30072 ( .A(n28023), .B(n28024), .Z(n28020) );
  AND U30073 ( .A(n28025), .B(n28026), .Z(n28023) );
  XOR U30074 ( .A(n[680]), .B(n28024), .Z(n28026) );
  XNOR U30075 ( .A(n28024), .B(n23239), .Z(n28025) );
  XOR U30076 ( .A(n28027), .B(n28028), .Z(n28024) );
  AND U30077 ( .A(n28029), .B(n28030), .Z(n28027) );
  XOR U30078 ( .A(n[679]), .B(n28028), .Z(n28030) );
  XNOR U30079 ( .A(n28028), .B(n23244), .Z(n28029) );
  XOR U30080 ( .A(n28031), .B(n28032), .Z(n28028) );
  AND U30081 ( .A(n28033), .B(n28034), .Z(n28031) );
  XOR U30082 ( .A(n[678]), .B(n28032), .Z(n28034) );
  XNOR U30083 ( .A(n28032), .B(n23249), .Z(n28033) );
  XOR U30084 ( .A(n28035), .B(n28036), .Z(n28032) );
  AND U30085 ( .A(n28037), .B(n28038), .Z(n28035) );
  XOR U30086 ( .A(n[677]), .B(n28036), .Z(n28038) );
  XNOR U30087 ( .A(n28036), .B(n23254), .Z(n28037) );
  XOR U30088 ( .A(n28039), .B(n28040), .Z(n28036) );
  AND U30089 ( .A(n28041), .B(n28042), .Z(n28039) );
  XOR U30090 ( .A(n[676]), .B(n28040), .Z(n28042) );
  XNOR U30091 ( .A(n28040), .B(n23259), .Z(n28041) );
  XOR U30092 ( .A(n28043), .B(n28044), .Z(n28040) );
  AND U30093 ( .A(n28045), .B(n28046), .Z(n28043) );
  XOR U30094 ( .A(n[675]), .B(n28044), .Z(n28046) );
  XNOR U30095 ( .A(n28044), .B(n23264), .Z(n28045) );
  XOR U30096 ( .A(n28047), .B(n28048), .Z(n28044) );
  AND U30097 ( .A(n28049), .B(n28050), .Z(n28047) );
  XOR U30098 ( .A(n[674]), .B(n28048), .Z(n28050) );
  XNOR U30099 ( .A(n28048), .B(n23269), .Z(n28049) );
  XOR U30100 ( .A(n28051), .B(n28052), .Z(n28048) );
  AND U30101 ( .A(n28053), .B(n28054), .Z(n28051) );
  XOR U30102 ( .A(n[673]), .B(n28052), .Z(n28054) );
  XNOR U30103 ( .A(n28052), .B(n23274), .Z(n28053) );
  XOR U30104 ( .A(n28055), .B(n28056), .Z(n28052) );
  AND U30105 ( .A(n28057), .B(n28058), .Z(n28055) );
  XOR U30106 ( .A(n[672]), .B(n28056), .Z(n28058) );
  XNOR U30107 ( .A(n28056), .B(n23279), .Z(n28057) );
  XOR U30108 ( .A(n28059), .B(n28060), .Z(n28056) );
  AND U30109 ( .A(n28061), .B(n28062), .Z(n28059) );
  XOR U30110 ( .A(n[671]), .B(n28060), .Z(n28062) );
  XNOR U30111 ( .A(n28060), .B(n23284), .Z(n28061) );
  XOR U30112 ( .A(n28063), .B(n28064), .Z(n28060) );
  AND U30113 ( .A(n28065), .B(n28066), .Z(n28063) );
  XOR U30114 ( .A(n[670]), .B(n28064), .Z(n28066) );
  XNOR U30115 ( .A(n28064), .B(n23289), .Z(n28065) );
  XOR U30116 ( .A(n28067), .B(n28068), .Z(n28064) );
  AND U30117 ( .A(n28069), .B(n28070), .Z(n28067) );
  XOR U30118 ( .A(n[669]), .B(n28068), .Z(n28070) );
  XNOR U30119 ( .A(n28068), .B(n23294), .Z(n28069) );
  XOR U30120 ( .A(n28071), .B(n28072), .Z(n28068) );
  AND U30121 ( .A(n28073), .B(n28074), .Z(n28071) );
  XOR U30122 ( .A(n[668]), .B(n28072), .Z(n28074) );
  XNOR U30123 ( .A(n28072), .B(n23299), .Z(n28073) );
  XOR U30124 ( .A(n28075), .B(n28076), .Z(n28072) );
  AND U30125 ( .A(n28077), .B(n28078), .Z(n28075) );
  XOR U30126 ( .A(n[667]), .B(n28076), .Z(n28078) );
  XNOR U30127 ( .A(n28076), .B(n23304), .Z(n28077) );
  XOR U30128 ( .A(n28079), .B(n28080), .Z(n28076) );
  AND U30129 ( .A(n28081), .B(n28082), .Z(n28079) );
  XOR U30130 ( .A(n[666]), .B(n28080), .Z(n28082) );
  XNOR U30131 ( .A(n28080), .B(n23309), .Z(n28081) );
  XOR U30132 ( .A(n28083), .B(n28084), .Z(n28080) );
  AND U30133 ( .A(n28085), .B(n28086), .Z(n28083) );
  XOR U30134 ( .A(n[665]), .B(n28084), .Z(n28086) );
  XNOR U30135 ( .A(n28084), .B(n23314), .Z(n28085) );
  XOR U30136 ( .A(n28087), .B(n28088), .Z(n28084) );
  AND U30137 ( .A(n28089), .B(n28090), .Z(n28087) );
  XOR U30138 ( .A(n[664]), .B(n28088), .Z(n28090) );
  XNOR U30139 ( .A(n28088), .B(n23319), .Z(n28089) );
  XOR U30140 ( .A(n28091), .B(n28092), .Z(n28088) );
  AND U30141 ( .A(n28093), .B(n28094), .Z(n28091) );
  XOR U30142 ( .A(n[663]), .B(n28092), .Z(n28094) );
  XNOR U30143 ( .A(n28092), .B(n23324), .Z(n28093) );
  XOR U30144 ( .A(n28095), .B(n28096), .Z(n28092) );
  AND U30145 ( .A(n28097), .B(n28098), .Z(n28095) );
  XOR U30146 ( .A(n[662]), .B(n28096), .Z(n28098) );
  XNOR U30147 ( .A(n28096), .B(n23329), .Z(n28097) );
  XOR U30148 ( .A(n28099), .B(n28100), .Z(n28096) );
  AND U30149 ( .A(n28101), .B(n28102), .Z(n28099) );
  XOR U30150 ( .A(n[661]), .B(n28100), .Z(n28102) );
  XNOR U30151 ( .A(n28100), .B(n23334), .Z(n28101) );
  XOR U30152 ( .A(n28103), .B(n28104), .Z(n28100) );
  AND U30153 ( .A(n28105), .B(n28106), .Z(n28103) );
  XOR U30154 ( .A(n[660]), .B(n28104), .Z(n28106) );
  XNOR U30155 ( .A(n28104), .B(n23339), .Z(n28105) );
  XOR U30156 ( .A(n28107), .B(n28108), .Z(n28104) );
  AND U30157 ( .A(n28109), .B(n28110), .Z(n28107) );
  XOR U30158 ( .A(n[659]), .B(n28108), .Z(n28110) );
  XNOR U30159 ( .A(n28108), .B(n23344), .Z(n28109) );
  XOR U30160 ( .A(n28111), .B(n28112), .Z(n28108) );
  AND U30161 ( .A(n28113), .B(n28114), .Z(n28111) );
  XOR U30162 ( .A(n[658]), .B(n28112), .Z(n28114) );
  XNOR U30163 ( .A(n28112), .B(n23349), .Z(n28113) );
  XOR U30164 ( .A(n28115), .B(n28116), .Z(n28112) );
  AND U30165 ( .A(n28117), .B(n28118), .Z(n28115) );
  XOR U30166 ( .A(n[657]), .B(n28116), .Z(n28118) );
  XNOR U30167 ( .A(n28116), .B(n23354), .Z(n28117) );
  XOR U30168 ( .A(n28119), .B(n28120), .Z(n28116) );
  AND U30169 ( .A(n28121), .B(n28122), .Z(n28119) );
  XOR U30170 ( .A(n[656]), .B(n28120), .Z(n28122) );
  XNOR U30171 ( .A(n28120), .B(n23359), .Z(n28121) );
  XOR U30172 ( .A(n28123), .B(n28124), .Z(n28120) );
  AND U30173 ( .A(n28125), .B(n28126), .Z(n28123) );
  XOR U30174 ( .A(n[655]), .B(n28124), .Z(n28126) );
  XNOR U30175 ( .A(n28124), .B(n23364), .Z(n28125) );
  XOR U30176 ( .A(n28127), .B(n28128), .Z(n28124) );
  AND U30177 ( .A(n28129), .B(n28130), .Z(n28127) );
  XOR U30178 ( .A(n[654]), .B(n28128), .Z(n28130) );
  XNOR U30179 ( .A(n28128), .B(n23369), .Z(n28129) );
  XOR U30180 ( .A(n28131), .B(n28132), .Z(n28128) );
  AND U30181 ( .A(n28133), .B(n28134), .Z(n28131) );
  XOR U30182 ( .A(n[653]), .B(n28132), .Z(n28134) );
  XNOR U30183 ( .A(n28132), .B(n23374), .Z(n28133) );
  XOR U30184 ( .A(n28135), .B(n28136), .Z(n28132) );
  AND U30185 ( .A(n28137), .B(n28138), .Z(n28135) );
  XOR U30186 ( .A(n[652]), .B(n28136), .Z(n28138) );
  XNOR U30187 ( .A(n28136), .B(n23379), .Z(n28137) );
  XOR U30188 ( .A(n28139), .B(n28140), .Z(n28136) );
  AND U30189 ( .A(n28141), .B(n28142), .Z(n28139) );
  XOR U30190 ( .A(n[651]), .B(n28140), .Z(n28142) );
  XNOR U30191 ( .A(n28140), .B(n23384), .Z(n28141) );
  XOR U30192 ( .A(n28143), .B(n28144), .Z(n28140) );
  AND U30193 ( .A(n28145), .B(n28146), .Z(n28143) );
  XOR U30194 ( .A(n[650]), .B(n28144), .Z(n28146) );
  XNOR U30195 ( .A(n28144), .B(n23389), .Z(n28145) );
  XOR U30196 ( .A(n28147), .B(n28148), .Z(n28144) );
  AND U30197 ( .A(n28149), .B(n28150), .Z(n28147) );
  XOR U30198 ( .A(n[649]), .B(n28148), .Z(n28150) );
  XNOR U30199 ( .A(n28148), .B(n23394), .Z(n28149) );
  XOR U30200 ( .A(n28151), .B(n28152), .Z(n28148) );
  AND U30201 ( .A(n28153), .B(n28154), .Z(n28151) );
  XOR U30202 ( .A(n[648]), .B(n28152), .Z(n28154) );
  XNOR U30203 ( .A(n28152), .B(n23399), .Z(n28153) );
  XOR U30204 ( .A(n28155), .B(n28156), .Z(n28152) );
  AND U30205 ( .A(n28157), .B(n28158), .Z(n28155) );
  XOR U30206 ( .A(n[647]), .B(n28156), .Z(n28158) );
  XNOR U30207 ( .A(n28156), .B(n23404), .Z(n28157) );
  XOR U30208 ( .A(n28159), .B(n28160), .Z(n28156) );
  AND U30209 ( .A(n28161), .B(n28162), .Z(n28159) );
  XOR U30210 ( .A(n[646]), .B(n28160), .Z(n28162) );
  XNOR U30211 ( .A(n28160), .B(n23409), .Z(n28161) );
  XOR U30212 ( .A(n28163), .B(n28164), .Z(n28160) );
  AND U30213 ( .A(n28165), .B(n28166), .Z(n28163) );
  XOR U30214 ( .A(n[645]), .B(n28164), .Z(n28166) );
  XNOR U30215 ( .A(n28164), .B(n23414), .Z(n28165) );
  XOR U30216 ( .A(n28167), .B(n28168), .Z(n28164) );
  AND U30217 ( .A(n28169), .B(n28170), .Z(n28167) );
  XOR U30218 ( .A(n[644]), .B(n28168), .Z(n28170) );
  XNOR U30219 ( .A(n28168), .B(n23419), .Z(n28169) );
  XOR U30220 ( .A(n28171), .B(n28172), .Z(n28168) );
  AND U30221 ( .A(n28173), .B(n28174), .Z(n28171) );
  XOR U30222 ( .A(n[643]), .B(n28172), .Z(n28174) );
  XNOR U30223 ( .A(n28172), .B(n23424), .Z(n28173) );
  XOR U30224 ( .A(n28175), .B(n28176), .Z(n28172) );
  AND U30225 ( .A(n28177), .B(n28178), .Z(n28175) );
  XOR U30226 ( .A(n[642]), .B(n28176), .Z(n28178) );
  XNOR U30227 ( .A(n28176), .B(n23429), .Z(n28177) );
  XOR U30228 ( .A(n28179), .B(n28180), .Z(n28176) );
  AND U30229 ( .A(n28181), .B(n28182), .Z(n28179) );
  XOR U30230 ( .A(n[641]), .B(n28180), .Z(n28182) );
  XNOR U30231 ( .A(n28180), .B(n23434), .Z(n28181) );
  XOR U30232 ( .A(n28183), .B(n28184), .Z(n28180) );
  AND U30233 ( .A(n28185), .B(n28186), .Z(n28183) );
  XOR U30234 ( .A(n[640]), .B(n28184), .Z(n28186) );
  XNOR U30235 ( .A(n28184), .B(n23439), .Z(n28185) );
  XOR U30236 ( .A(n28187), .B(n28188), .Z(n28184) );
  AND U30237 ( .A(n28189), .B(n28190), .Z(n28187) );
  XOR U30238 ( .A(n[639]), .B(n28188), .Z(n28190) );
  XNOR U30239 ( .A(n28188), .B(n23444), .Z(n28189) );
  XOR U30240 ( .A(n28191), .B(n28192), .Z(n28188) );
  AND U30241 ( .A(n28193), .B(n28194), .Z(n28191) );
  XOR U30242 ( .A(n[638]), .B(n28192), .Z(n28194) );
  XNOR U30243 ( .A(n28192), .B(n23449), .Z(n28193) );
  XOR U30244 ( .A(n28195), .B(n28196), .Z(n28192) );
  AND U30245 ( .A(n28197), .B(n28198), .Z(n28195) );
  XOR U30246 ( .A(n[637]), .B(n28196), .Z(n28198) );
  XNOR U30247 ( .A(n28196), .B(n23454), .Z(n28197) );
  XOR U30248 ( .A(n28199), .B(n28200), .Z(n28196) );
  AND U30249 ( .A(n28201), .B(n28202), .Z(n28199) );
  XOR U30250 ( .A(n[636]), .B(n28200), .Z(n28202) );
  XNOR U30251 ( .A(n28200), .B(n23459), .Z(n28201) );
  XOR U30252 ( .A(n28203), .B(n28204), .Z(n28200) );
  AND U30253 ( .A(n28205), .B(n28206), .Z(n28203) );
  XOR U30254 ( .A(n[635]), .B(n28204), .Z(n28206) );
  XNOR U30255 ( .A(n28204), .B(n23464), .Z(n28205) );
  XOR U30256 ( .A(n28207), .B(n28208), .Z(n28204) );
  AND U30257 ( .A(n28209), .B(n28210), .Z(n28207) );
  XOR U30258 ( .A(n[634]), .B(n28208), .Z(n28210) );
  XNOR U30259 ( .A(n28208), .B(n23469), .Z(n28209) );
  XOR U30260 ( .A(n28211), .B(n28212), .Z(n28208) );
  AND U30261 ( .A(n28213), .B(n28214), .Z(n28211) );
  XOR U30262 ( .A(n[633]), .B(n28212), .Z(n28214) );
  XNOR U30263 ( .A(n28212), .B(n23474), .Z(n28213) );
  XOR U30264 ( .A(n28215), .B(n28216), .Z(n28212) );
  AND U30265 ( .A(n28217), .B(n28218), .Z(n28215) );
  XOR U30266 ( .A(n[632]), .B(n28216), .Z(n28218) );
  XNOR U30267 ( .A(n28216), .B(n23479), .Z(n28217) );
  XOR U30268 ( .A(n28219), .B(n28220), .Z(n28216) );
  AND U30269 ( .A(n28221), .B(n28222), .Z(n28219) );
  XOR U30270 ( .A(n[631]), .B(n28220), .Z(n28222) );
  XNOR U30271 ( .A(n28220), .B(n23484), .Z(n28221) );
  XOR U30272 ( .A(n28223), .B(n28224), .Z(n28220) );
  AND U30273 ( .A(n28225), .B(n28226), .Z(n28223) );
  XOR U30274 ( .A(n[630]), .B(n28224), .Z(n28226) );
  XNOR U30275 ( .A(n28224), .B(n23489), .Z(n28225) );
  XOR U30276 ( .A(n28227), .B(n28228), .Z(n28224) );
  AND U30277 ( .A(n28229), .B(n28230), .Z(n28227) );
  XOR U30278 ( .A(n[629]), .B(n28228), .Z(n28230) );
  XNOR U30279 ( .A(n28228), .B(n23494), .Z(n28229) );
  XOR U30280 ( .A(n28231), .B(n28232), .Z(n28228) );
  AND U30281 ( .A(n28233), .B(n28234), .Z(n28231) );
  XOR U30282 ( .A(n[628]), .B(n28232), .Z(n28234) );
  XNOR U30283 ( .A(n28232), .B(n23499), .Z(n28233) );
  XOR U30284 ( .A(n28235), .B(n28236), .Z(n28232) );
  AND U30285 ( .A(n28237), .B(n28238), .Z(n28235) );
  XOR U30286 ( .A(n[627]), .B(n28236), .Z(n28238) );
  XNOR U30287 ( .A(n28236), .B(n23504), .Z(n28237) );
  XOR U30288 ( .A(n28239), .B(n28240), .Z(n28236) );
  AND U30289 ( .A(n28241), .B(n28242), .Z(n28239) );
  XOR U30290 ( .A(n[626]), .B(n28240), .Z(n28242) );
  XNOR U30291 ( .A(n28240), .B(n23509), .Z(n28241) );
  XOR U30292 ( .A(n28243), .B(n28244), .Z(n28240) );
  AND U30293 ( .A(n28245), .B(n28246), .Z(n28243) );
  XOR U30294 ( .A(n[625]), .B(n28244), .Z(n28246) );
  XNOR U30295 ( .A(n28244), .B(n23514), .Z(n28245) );
  XOR U30296 ( .A(n28247), .B(n28248), .Z(n28244) );
  AND U30297 ( .A(n28249), .B(n28250), .Z(n28247) );
  XOR U30298 ( .A(n[624]), .B(n28248), .Z(n28250) );
  XNOR U30299 ( .A(n28248), .B(n23519), .Z(n28249) );
  XOR U30300 ( .A(n28251), .B(n28252), .Z(n28248) );
  AND U30301 ( .A(n28253), .B(n28254), .Z(n28251) );
  XOR U30302 ( .A(n[623]), .B(n28252), .Z(n28254) );
  XNOR U30303 ( .A(n28252), .B(n23524), .Z(n28253) );
  XOR U30304 ( .A(n28255), .B(n28256), .Z(n28252) );
  AND U30305 ( .A(n28257), .B(n28258), .Z(n28255) );
  XOR U30306 ( .A(n[622]), .B(n28256), .Z(n28258) );
  XNOR U30307 ( .A(n28256), .B(n23529), .Z(n28257) );
  XOR U30308 ( .A(n28259), .B(n28260), .Z(n28256) );
  AND U30309 ( .A(n28261), .B(n28262), .Z(n28259) );
  XOR U30310 ( .A(n[621]), .B(n28260), .Z(n28262) );
  XNOR U30311 ( .A(n28260), .B(n23534), .Z(n28261) );
  XOR U30312 ( .A(n28263), .B(n28264), .Z(n28260) );
  AND U30313 ( .A(n28265), .B(n28266), .Z(n28263) );
  XOR U30314 ( .A(n[620]), .B(n28264), .Z(n28266) );
  XNOR U30315 ( .A(n28264), .B(n23539), .Z(n28265) );
  XOR U30316 ( .A(n28267), .B(n28268), .Z(n28264) );
  AND U30317 ( .A(n28269), .B(n28270), .Z(n28267) );
  XOR U30318 ( .A(n[619]), .B(n28268), .Z(n28270) );
  XNOR U30319 ( .A(n28268), .B(n23544), .Z(n28269) );
  XOR U30320 ( .A(n28271), .B(n28272), .Z(n28268) );
  AND U30321 ( .A(n28273), .B(n28274), .Z(n28271) );
  XOR U30322 ( .A(n[618]), .B(n28272), .Z(n28274) );
  XNOR U30323 ( .A(n28272), .B(n23549), .Z(n28273) );
  XOR U30324 ( .A(n28275), .B(n28276), .Z(n28272) );
  AND U30325 ( .A(n28277), .B(n28278), .Z(n28275) );
  XOR U30326 ( .A(n[617]), .B(n28276), .Z(n28278) );
  XNOR U30327 ( .A(n28276), .B(n23554), .Z(n28277) );
  XOR U30328 ( .A(n28279), .B(n28280), .Z(n28276) );
  AND U30329 ( .A(n28281), .B(n28282), .Z(n28279) );
  XOR U30330 ( .A(n[616]), .B(n28280), .Z(n28282) );
  XNOR U30331 ( .A(n28280), .B(n23559), .Z(n28281) );
  XOR U30332 ( .A(n28283), .B(n28284), .Z(n28280) );
  AND U30333 ( .A(n28285), .B(n28286), .Z(n28283) );
  XOR U30334 ( .A(n[615]), .B(n28284), .Z(n28286) );
  XNOR U30335 ( .A(n28284), .B(n23564), .Z(n28285) );
  XOR U30336 ( .A(n28287), .B(n28288), .Z(n28284) );
  AND U30337 ( .A(n28289), .B(n28290), .Z(n28287) );
  XOR U30338 ( .A(n[614]), .B(n28288), .Z(n28290) );
  XNOR U30339 ( .A(n28288), .B(n23569), .Z(n28289) );
  XOR U30340 ( .A(n28291), .B(n28292), .Z(n28288) );
  AND U30341 ( .A(n28293), .B(n28294), .Z(n28291) );
  XOR U30342 ( .A(n[613]), .B(n28292), .Z(n28294) );
  XNOR U30343 ( .A(n28292), .B(n23574), .Z(n28293) );
  XOR U30344 ( .A(n28295), .B(n28296), .Z(n28292) );
  AND U30345 ( .A(n28297), .B(n28298), .Z(n28295) );
  XOR U30346 ( .A(n[612]), .B(n28296), .Z(n28298) );
  XNOR U30347 ( .A(n28296), .B(n23579), .Z(n28297) );
  XOR U30348 ( .A(n28299), .B(n28300), .Z(n28296) );
  AND U30349 ( .A(n28301), .B(n28302), .Z(n28299) );
  XOR U30350 ( .A(n[611]), .B(n28300), .Z(n28302) );
  XNOR U30351 ( .A(n28300), .B(n23584), .Z(n28301) );
  XOR U30352 ( .A(n28303), .B(n28304), .Z(n28300) );
  AND U30353 ( .A(n28305), .B(n28306), .Z(n28303) );
  XOR U30354 ( .A(n[610]), .B(n28304), .Z(n28306) );
  XNOR U30355 ( .A(n28304), .B(n23589), .Z(n28305) );
  XOR U30356 ( .A(n28307), .B(n28308), .Z(n28304) );
  AND U30357 ( .A(n28309), .B(n28310), .Z(n28307) );
  XOR U30358 ( .A(n[609]), .B(n28308), .Z(n28310) );
  XNOR U30359 ( .A(n28308), .B(n23594), .Z(n28309) );
  XOR U30360 ( .A(n28311), .B(n28312), .Z(n28308) );
  AND U30361 ( .A(n28313), .B(n28314), .Z(n28311) );
  XOR U30362 ( .A(n[608]), .B(n28312), .Z(n28314) );
  XNOR U30363 ( .A(n28312), .B(n23599), .Z(n28313) );
  XOR U30364 ( .A(n28315), .B(n28316), .Z(n28312) );
  AND U30365 ( .A(n28317), .B(n28318), .Z(n28315) );
  XOR U30366 ( .A(n[607]), .B(n28316), .Z(n28318) );
  XNOR U30367 ( .A(n28316), .B(n23604), .Z(n28317) );
  XOR U30368 ( .A(n28319), .B(n28320), .Z(n28316) );
  AND U30369 ( .A(n28321), .B(n28322), .Z(n28319) );
  XOR U30370 ( .A(n[606]), .B(n28320), .Z(n28322) );
  XNOR U30371 ( .A(n28320), .B(n23609), .Z(n28321) );
  XOR U30372 ( .A(n28323), .B(n28324), .Z(n28320) );
  AND U30373 ( .A(n28325), .B(n28326), .Z(n28323) );
  XOR U30374 ( .A(n[605]), .B(n28324), .Z(n28326) );
  XNOR U30375 ( .A(n28324), .B(n23614), .Z(n28325) );
  XOR U30376 ( .A(n28327), .B(n28328), .Z(n28324) );
  AND U30377 ( .A(n28329), .B(n28330), .Z(n28327) );
  XOR U30378 ( .A(n[604]), .B(n28328), .Z(n28330) );
  XNOR U30379 ( .A(n28328), .B(n23619), .Z(n28329) );
  XOR U30380 ( .A(n28331), .B(n28332), .Z(n28328) );
  AND U30381 ( .A(n28333), .B(n28334), .Z(n28331) );
  XOR U30382 ( .A(n[603]), .B(n28332), .Z(n28334) );
  XNOR U30383 ( .A(n28332), .B(n23624), .Z(n28333) );
  XOR U30384 ( .A(n28335), .B(n28336), .Z(n28332) );
  AND U30385 ( .A(n28337), .B(n28338), .Z(n28335) );
  XOR U30386 ( .A(n[602]), .B(n28336), .Z(n28338) );
  XNOR U30387 ( .A(n28336), .B(n23629), .Z(n28337) );
  XOR U30388 ( .A(n28339), .B(n28340), .Z(n28336) );
  AND U30389 ( .A(n28341), .B(n28342), .Z(n28339) );
  XOR U30390 ( .A(n[601]), .B(n28340), .Z(n28342) );
  XNOR U30391 ( .A(n28340), .B(n23634), .Z(n28341) );
  XOR U30392 ( .A(n28343), .B(n28344), .Z(n28340) );
  AND U30393 ( .A(n28345), .B(n28346), .Z(n28343) );
  XOR U30394 ( .A(n[600]), .B(n28344), .Z(n28346) );
  XNOR U30395 ( .A(n28344), .B(n23639), .Z(n28345) );
  XOR U30396 ( .A(n28347), .B(n28348), .Z(n28344) );
  AND U30397 ( .A(n28349), .B(n28350), .Z(n28347) );
  XOR U30398 ( .A(n[599]), .B(n28348), .Z(n28350) );
  XNOR U30399 ( .A(n28348), .B(n23644), .Z(n28349) );
  XOR U30400 ( .A(n28351), .B(n28352), .Z(n28348) );
  AND U30401 ( .A(n28353), .B(n28354), .Z(n28351) );
  XOR U30402 ( .A(n[598]), .B(n28352), .Z(n28354) );
  XNOR U30403 ( .A(n28352), .B(n23649), .Z(n28353) );
  XOR U30404 ( .A(n28355), .B(n28356), .Z(n28352) );
  AND U30405 ( .A(n28357), .B(n28358), .Z(n28355) );
  XOR U30406 ( .A(n[597]), .B(n28356), .Z(n28358) );
  XNOR U30407 ( .A(n28356), .B(n23654), .Z(n28357) );
  XOR U30408 ( .A(n28359), .B(n28360), .Z(n28356) );
  AND U30409 ( .A(n28361), .B(n28362), .Z(n28359) );
  XOR U30410 ( .A(n[596]), .B(n28360), .Z(n28362) );
  XNOR U30411 ( .A(n28360), .B(n23659), .Z(n28361) );
  XOR U30412 ( .A(n28363), .B(n28364), .Z(n28360) );
  AND U30413 ( .A(n28365), .B(n28366), .Z(n28363) );
  XOR U30414 ( .A(n[595]), .B(n28364), .Z(n28366) );
  XNOR U30415 ( .A(n28364), .B(n23664), .Z(n28365) );
  XOR U30416 ( .A(n28367), .B(n28368), .Z(n28364) );
  AND U30417 ( .A(n28369), .B(n28370), .Z(n28367) );
  XOR U30418 ( .A(n[594]), .B(n28368), .Z(n28370) );
  XNOR U30419 ( .A(n28368), .B(n23669), .Z(n28369) );
  XOR U30420 ( .A(n28371), .B(n28372), .Z(n28368) );
  AND U30421 ( .A(n28373), .B(n28374), .Z(n28371) );
  XOR U30422 ( .A(n[593]), .B(n28372), .Z(n28374) );
  XNOR U30423 ( .A(n28372), .B(n23674), .Z(n28373) );
  XOR U30424 ( .A(n28375), .B(n28376), .Z(n28372) );
  AND U30425 ( .A(n28377), .B(n28378), .Z(n28375) );
  XOR U30426 ( .A(n[592]), .B(n28376), .Z(n28378) );
  XNOR U30427 ( .A(n28376), .B(n23679), .Z(n28377) );
  XOR U30428 ( .A(n28379), .B(n28380), .Z(n28376) );
  AND U30429 ( .A(n28381), .B(n28382), .Z(n28379) );
  XOR U30430 ( .A(n[591]), .B(n28380), .Z(n28382) );
  XNOR U30431 ( .A(n28380), .B(n23684), .Z(n28381) );
  XOR U30432 ( .A(n28383), .B(n28384), .Z(n28380) );
  AND U30433 ( .A(n28385), .B(n28386), .Z(n28383) );
  XOR U30434 ( .A(n[590]), .B(n28384), .Z(n28386) );
  XNOR U30435 ( .A(n28384), .B(n23689), .Z(n28385) );
  XOR U30436 ( .A(n28387), .B(n28388), .Z(n28384) );
  AND U30437 ( .A(n28389), .B(n28390), .Z(n28387) );
  XOR U30438 ( .A(n[589]), .B(n28388), .Z(n28390) );
  XNOR U30439 ( .A(n28388), .B(n23694), .Z(n28389) );
  XOR U30440 ( .A(n28391), .B(n28392), .Z(n28388) );
  AND U30441 ( .A(n28393), .B(n28394), .Z(n28391) );
  XOR U30442 ( .A(n[588]), .B(n28392), .Z(n28394) );
  XNOR U30443 ( .A(n28392), .B(n23699), .Z(n28393) );
  XOR U30444 ( .A(n28395), .B(n28396), .Z(n28392) );
  AND U30445 ( .A(n28397), .B(n28398), .Z(n28395) );
  XOR U30446 ( .A(n[587]), .B(n28396), .Z(n28398) );
  XNOR U30447 ( .A(n28396), .B(n23704), .Z(n28397) );
  XOR U30448 ( .A(n28399), .B(n28400), .Z(n28396) );
  AND U30449 ( .A(n28401), .B(n28402), .Z(n28399) );
  XOR U30450 ( .A(n[586]), .B(n28400), .Z(n28402) );
  XNOR U30451 ( .A(n28400), .B(n23709), .Z(n28401) );
  XOR U30452 ( .A(n28403), .B(n28404), .Z(n28400) );
  AND U30453 ( .A(n28405), .B(n28406), .Z(n28403) );
  XOR U30454 ( .A(n[585]), .B(n28404), .Z(n28406) );
  XNOR U30455 ( .A(n28404), .B(n23714), .Z(n28405) );
  XOR U30456 ( .A(n28407), .B(n28408), .Z(n28404) );
  AND U30457 ( .A(n28409), .B(n28410), .Z(n28407) );
  XOR U30458 ( .A(n[584]), .B(n28408), .Z(n28410) );
  XNOR U30459 ( .A(n28408), .B(n23719), .Z(n28409) );
  XOR U30460 ( .A(n28411), .B(n28412), .Z(n28408) );
  AND U30461 ( .A(n28413), .B(n28414), .Z(n28411) );
  XOR U30462 ( .A(n[583]), .B(n28412), .Z(n28414) );
  XNOR U30463 ( .A(n28412), .B(n23724), .Z(n28413) );
  XOR U30464 ( .A(n28415), .B(n28416), .Z(n28412) );
  AND U30465 ( .A(n28417), .B(n28418), .Z(n28415) );
  XOR U30466 ( .A(n[582]), .B(n28416), .Z(n28418) );
  XNOR U30467 ( .A(n28416), .B(n23729), .Z(n28417) );
  XOR U30468 ( .A(n28419), .B(n28420), .Z(n28416) );
  AND U30469 ( .A(n28421), .B(n28422), .Z(n28419) );
  XOR U30470 ( .A(n[581]), .B(n28420), .Z(n28422) );
  XNOR U30471 ( .A(n28420), .B(n23734), .Z(n28421) );
  XOR U30472 ( .A(n28423), .B(n28424), .Z(n28420) );
  AND U30473 ( .A(n28425), .B(n28426), .Z(n28423) );
  XOR U30474 ( .A(n[580]), .B(n28424), .Z(n28426) );
  XNOR U30475 ( .A(n28424), .B(n23739), .Z(n28425) );
  XOR U30476 ( .A(n28427), .B(n28428), .Z(n28424) );
  AND U30477 ( .A(n28429), .B(n28430), .Z(n28427) );
  XOR U30478 ( .A(n[579]), .B(n28428), .Z(n28430) );
  XNOR U30479 ( .A(n28428), .B(n23744), .Z(n28429) );
  XOR U30480 ( .A(n28431), .B(n28432), .Z(n28428) );
  AND U30481 ( .A(n28433), .B(n28434), .Z(n28431) );
  XOR U30482 ( .A(n[578]), .B(n28432), .Z(n28434) );
  XNOR U30483 ( .A(n28432), .B(n23749), .Z(n28433) );
  XOR U30484 ( .A(n28435), .B(n28436), .Z(n28432) );
  AND U30485 ( .A(n28437), .B(n28438), .Z(n28435) );
  XOR U30486 ( .A(n[577]), .B(n28436), .Z(n28438) );
  XNOR U30487 ( .A(n28436), .B(n23754), .Z(n28437) );
  XOR U30488 ( .A(n28439), .B(n28440), .Z(n28436) );
  AND U30489 ( .A(n28441), .B(n28442), .Z(n28439) );
  XOR U30490 ( .A(n[576]), .B(n28440), .Z(n28442) );
  XNOR U30491 ( .A(n28440), .B(n23759), .Z(n28441) );
  XOR U30492 ( .A(n28443), .B(n28444), .Z(n28440) );
  AND U30493 ( .A(n28445), .B(n28446), .Z(n28443) );
  XOR U30494 ( .A(n[575]), .B(n28444), .Z(n28446) );
  XNOR U30495 ( .A(n28444), .B(n23764), .Z(n28445) );
  XOR U30496 ( .A(n28447), .B(n28448), .Z(n28444) );
  AND U30497 ( .A(n28449), .B(n28450), .Z(n28447) );
  XOR U30498 ( .A(n[574]), .B(n28448), .Z(n28450) );
  XNOR U30499 ( .A(n28448), .B(n23769), .Z(n28449) );
  XOR U30500 ( .A(n28451), .B(n28452), .Z(n28448) );
  AND U30501 ( .A(n28453), .B(n28454), .Z(n28451) );
  XOR U30502 ( .A(n[573]), .B(n28452), .Z(n28454) );
  XNOR U30503 ( .A(n28452), .B(n23774), .Z(n28453) );
  XOR U30504 ( .A(n28455), .B(n28456), .Z(n28452) );
  AND U30505 ( .A(n28457), .B(n28458), .Z(n28455) );
  XOR U30506 ( .A(n[572]), .B(n28456), .Z(n28458) );
  XNOR U30507 ( .A(n28456), .B(n23779), .Z(n28457) );
  XOR U30508 ( .A(n28459), .B(n28460), .Z(n28456) );
  AND U30509 ( .A(n28461), .B(n28462), .Z(n28459) );
  XOR U30510 ( .A(n[571]), .B(n28460), .Z(n28462) );
  XNOR U30511 ( .A(n28460), .B(n23784), .Z(n28461) );
  XOR U30512 ( .A(n28463), .B(n28464), .Z(n28460) );
  AND U30513 ( .A(n28465), .B(n28466), .Z(n28463) );
  XOR U30514 ( .A(n[570]), .B(n28464), .Z(n28466) );
  XNOR U30515 ( .A(n28464), .B(n23789), .Z(n28465) );
  XOR U30516 ( .A(n28467), .B(n28468), .Z(n28464) );
  AND U30517 ( .A(n28469), .B(n28470), .Z(n28467) );
  XOR U30518 ( .A(n[569]), .B(n28468), .Z(n28470) );
  XNOR U30519 ( .A(n28468), .B(n23794), .Z(n28469) );
  XOR U30520 ( .A(n28471), .B(n28472), .Z(n28468) );
  AND U30521 ( .A(n28473), .B(n28474), .Z(n28471) );
  XOR U30522 ( .A(n[568]), .B(n28472), .Z(n28474) );
  XNOR U30523 ( .A(n28472), .B(n23799), .Z(n28473) );
  XOR U30524 ( .A(n28475), .B(n28476), .Z(n28472) );
  AND U30525 ( .A(n28477), .B(n28478), .Z(n28475) );
  XOR U30526 ( .A(n[567]), .B(n28476), .Z(n28478) );
  XNOR U30527 ( .A(n28476), .B(n23804), .Z(n28477) );
  XOR U30528 ( .A(n28479), .B(n28480), .Z(n28476) );
  AND U30529 ( .A(n28481), .B(n28482), .Z(n28479) );
  XOR U30530 ( .A(n[566]), .B(n28480), .Z(n28482) );
  XNOR U30531 ( .A(n28480), .B(n23809), .Z(n28481) );
  XOR U30532 ( .A(n28483), .B(n28484), .Z(n28480) );
  AND U30533 ( .A(n28485), .B(n28486), .Z(n28483) );
  XOR U30534 ( .A(n[565]), .B(n28484), .Z(n28486) );
  XNOR U30535 ( .A(n28484), .B(n23814), .Z(n28485) );
  XOR U30536 ( .A(n28487), .B(n28488), .Z(n28484) );
  AND U30537 ( .A(n28489), .B(n28490), .Z(n28487) );
  XOR U30538 ( .A(n[564]), .B(n28488), .Z(n28490) );
  XNOR U30539 ( .A(n28488), .B(n23819), .Z(n28489) );
  XOR U30540 ( .A(n28491), .B(n28492), .Z(n28488) );
  AND U30541 ( .A(n28493), .B(n28494), .Z(n28491) );
  XOR U30542 ( .A(n[563]), .B(n28492), .Z(n28494) );
  XNOR U30543 ( .A(n28492), .B(n23824), .Z(n28493) );
  XOR U30544 ( .A(n28495), .B(n28496), .Z(n28492) );
  AND U30545 ( .A(n28497), .B(n28498), .Z(n28495) );
  XOR U30546 ( .A(n[562]), .B(n28496), .Z(n28498) );
  XNOR U30547 ( .A(n28496), .B(n23829), .Z(n28497) );
  XOR U30548 ( .A(n28499), .B(n28500), .Z(n28496) );
  AND U30549 ( .A(n28501), .B(n28502), .Z(n28499) );
  XOR U30550 ( .A(n[561]), .B(n28500), .Z(n28502) );
  XNOR U30551 ( .A(n28500), .B(n23834), .Z(n28501) );
  XOR U30552 ( .A(n28503), .B(n28504), .Z(n28500) );
  AND U30553 ( .A(n28505), .B(n28506), .Z(n28503) );
  XOR U30554 ( .A(n[560]), .B(n28504), .Z(n28506) );
  XNOR U30555 ( .A(n28504), .B(n23839), .Z(n28505) );
  XOR U30556 ( .A(n28507), .B(n28508), .Z(n28504) );
  AND U30557 ( .A(n28509), .B(n28510), .Z(n28507) );
  XOR U30558 ( .A(n[559]), .B(n28508), .Z(n28510) );
  XNOR U30559 ( .A(n28508), .B(n23844), .Z(n28509) );
  XOR U30560 ( .A(n28511), .B(n28512), .Z(n28508) );
  AND U30561 ( .A(n28513), .B(n28514), .Z(n28511) );
  XOR U30562 ( .A(n[558]), .B(n28512), .Z(n28514) );
  XNOR U30563 ( .A(n28512), .B(n23849), .Z(n28513) );
  XOR U30564 ( .A(n28515), .B(n28516), .Z(n28512) );
  AND U30565 ( .A(n28517), .B(n28518), .Z(n28515) );
  XOR U30566 ( .A(n[557]), .B(n28516), .Z(n28518) );
  XNOR U30567 ( .A(n28516), .B(n23854), .Z(n28517) );
  XOR U30568 ( .A(n28519), .B(n28520), .Z(n28516) );
  AND U30569 ( .A(n28521), .B(n28522), .Z(n28519) );
  XOR U30570 ( .A(n[556]), .B(n28520), .Z(n28522) );
  XNOR U30571 ( .A(n28520), .B(n23859), .Z(n28521) );
  XOR U30572 ( .A(n28523), .B(n28524), .Z(n28520) );
  AND U30573 ( .A(n28525), .B(n28526), .Z(n28523) );
  XOR U30574 ( .A(n[555]), .B(n28524), .Z(n28526) );
  XNOR U30575 ( .A(n28524), .B(n23864), .Z(n28525) );
  XOR U30576 ( .A(n28527), .B(n28528), .Z(n28524) );
  AND U30577 ( .A(n28529), .B(n28530), .Z(n28527) );
  XOR U30578 ( .A(n[554]), .B(n28528), .Z(n28530) );
  XNOR U30579 ( .A(n28528), .B(n23869), .Z(n28529) );
  XOR U30580 ( .A(n28531), .B(n28532), .Z(n28528) );
  AND U30581 ( .A(n28533), .B(n28534), .Z(n28531) );
  XOR U30582 ( .A(n[553]), .B(n28532), .Z(n28534) );
  XNOR U30583 ( .A(n28532), .B(n23874), .Z(n28533) );
  XOR U30584 ( .A(n28535), .B(n28536), .Z(n28532) );
  AND U30585 ( .A(n28537), .B(n28538), .Z(n28535) );
  XOR U30586 ( .A(n[552]), .B(n28536), .Z(n28538) );
  XNOR U30587 ( .A(n28536), .B(n23879), .Z(n28537) );
  XOR U30588 ( .A(n28539), .B(n28540), .Z(n28536) );
  AND U30589 ( .A(n28541), .B(n28542), .Z(n28539) );
  XOR U30590 ( .A(n[551]), .B(n28540), .Z(n28542) );
  XNOR U30591 ( .A(n28540), .B(n23884), .Z(n28541) );
  XOR U30592 ( .A(n28543), .B(n28544), .Z(n28540) );
  AND U30593 ( .A(n28545), .B(n28546), .Z(n28543) );
  XOR U30594 ( .A(n[550]), .B(n28544), .Z(n28546) );
  XNOR U30595 ( .A(n28544), .B(n23889), .Z(n28545) );
  XOR U30596 ( .A(n28547), .B(n28548), .Z(n28544) );
  AND U30597 ( .A(n28549), .B(n28550), .Z(n28547) );
  XOR U30598 ( .A(n[549]), .B(n28548), .Z(n28550) );
  XNOR U30599 ( .A(n28548), .B(n23894), .Z(n28549) );
  XOR U30600 ( .A(n28551), .B(n28552), .Z(n28548) );
  AND U30601 ( .A(n28553), .B(n28554), .Z(n28551) );
  XOR U30602 ( .A(n[548]), .B(n28552), .Z(n28554) );
  XNOR U30603 ( .A(n28552), .B(n23899), .Z(n28553) );
  XOR U30604 ( .A(n28555), .B(n28556), .Z(n28552) );
  AND U30605 ( .A(n28557), .B(n28558), .Z(n28555) );
  XOR U30606 ( .A(n[547]), .B(n28556), .Z(n28558) );
  XNOR U30607 ( .A(n28556), .B(n23904), .Z(n28557) );
  XOR U30608 ( .A(n28559), .B(n28560), .Z(n28556) );
  AND U30609 ( .A(n28561), .B(n28562), .Z(n28559) );
  XOR U30610 ( .A(n[546]), .B(n28560), .Z(n28562) );
  XNOR U30611 ( .A(n28560), .B(n23909), .Z(n28561) );
  XOR U30612 ( .A(n28563), .B(n28564), .Z(n28560) );
  AND U30613 ( .A(n28565), .B(n28566), .Z(n28563) );
  XOR U30614 ( .A(n[545]), .B(n28564), .Z(n28566) );
  XNOR U30615 ( .A(n28564), .B(n23914), .Z(n28565) );
  XOR U30616 ( .A(n28567), .B(n28568), .Z(n28564) );
  AND U30617 ( .A(n28569), .B(n28570), .Z(n28567) );
  XOR U30618 ( .A(n[544]), .B(n28568), .Z(n28570) );
  XNOR U30619 ( .A(n28568), .B(n23919), .Z(n28569) );
  XOR U30620 ( .A(n28571), .B(n28572), .Z(n28568) );
  AND U30621 ( .A(n28573), .B(n28574), .Z(n28571) );
  XOR U30622 ( .A(n[543]), .B(n28572), .Z(n28574) );
  XNOR U30623 ( .A(n28572), .B(n23924), .Z(n28573) );
  XOR U30624 ( .A(n28575), .B(n28576), .Z(n28572) );
  AND U30625 ( .A(n28577), .B(n28578), .Z(n28575) );
  XOR U30626 ( .A(n[542]), .B(n28576), .Z(n28578) );
  XNOR U30627 ( .A(n28576), .B(n23929), .Z(n28577) );
  XOR U30628 ( .A(n28579), .B(n28580), .Z(n28576) );
  AND U30629 ( .A(n28581), .B(n28582), .Z(n28579) );
  XOR U30630 ( .A(n[541]), .B(n28580), .Z(n28582) );
  XNOR U30631 ( .A(n28580), .B(n23934), .Z(n28581) );
  XOR U30632 ( .A(n28583), .B(n28584), .Z(n28580) );
  AND U30633 ( .A(n28585), .B(n28586), .Z(n28583) );
  XOR U30634 ( .A(n[540]), .B(n28584), .Z(n28586) );
  XNOR U30635 ( .A(n28584), .B(n23939), .Z(n28585) );
  XOR U30636 ( .A(n28587), .B(n28588), .Z(n28584) );
  AND U30637 ( .A(n28589), .B(n28590), .Z(n28587) );
  XOR U30638 ( .A(n[539]), .B(n28588), .Z(n28590) );
  XNOR U30639 ( .A(n28588), .B(n23944), .Z(n28589) );
  XOR U30640 ( .A(n28591), .B(n28592), .Z(n28588) );
  AND U30641 ( .A(n28593), .B(n28594), .Z(n28591) );
  XOR U30642 ( .A(n[538]), .B(n28592), .Z(n28594) );
  XNOR U30643 ( .A(n28592), .B(n23949), .Z(n28593) );
  XOR U30644 ( .A(n28595), .B(n28596), .Z(n28592) );
  AND U30645 ( .A(n28597), .B(n28598), .Z(n28595) );
  XOR U30646 ( .A(n[537]), .B(n28596), .Z(n28598) );
  XNOR U30647 ( .A(n28596), .B(n23954), .Z(n28597) );
  XOR U30648 ( .A(n28599), .B(n28600), .Z(n28596) );
  AND U30649 ( .A(n28601), .B(n28602), .Z(n28599) );
  XOR U30650 ( .A(n[536]), .B(n28600), .Z(n28602) );
  XNOR U30651 ( .A(n28600), .B(n23959), .Z(n28601) );
  XOR U30652 ( .A(n28603), .B(n28604), .Z(n28600) );
  AND U30653 ( .A(n28605), .B(n28606), .Z(n28603) );
  XOR U30654 ( .A(n[535]), .B(n28604), .Z(n28606) );
  XNOR U30655 ( .A(n28604), .B(n23964), .Z(n28605) );
  XOR U30656 ( .A(n28607), .B(n28608), .Z(n28604) );
  AND U30657 ( .A(n28609), .B(n28610), .Z(n28607) );
  XOR U30658 ( .A(n[534]), .B(n28608), .Z(n28610) );
  XNOR U30659 ( .A(n28608), .B(n23969), .Z(n28609) );
  XOR U30660 ( .A(n28611), .B(n28612), .Z(n28608) );
  AND U30661 ( .A(n28613), .B(n28614), .Z(n28611) );
  XOR U30662 ( .A(n[533]), .B(n28612), .Z(n28614) );
  XNOR U30663 ( .A(n28612), .B(n23974), .Z(n28613) );
  XOR U30664 ( .A(n28615), .B(n28616), .Z(n28612) );
  AND U30665 ( .A(n28617), .B(n28618), .Z(n28615) );
  XOR U30666 ( .A(n[532]), .B(n28616), .Z(n28618) );
  XNOR U30667 ( .A(n28616), .B(n23979), .Z(n28617) );
  XOR U30668 ( .A(n28619), .B(n28620), .Z(n28616) );
  AND U30669 ( .A(n28621), .B(n28622), .Z(n28619) );
  XOR U30670 ( .A(n[531]), .B(n28620), .Z(n28622) );
  XNOR U30671 ( .A(n28620), .B(n23984), .Z(n28621) );
  XOR U30672 ( .A(n28623), .B(n28624), .Z(n28620) );
  AND U30673 ( .A(n28625), .B(n28626), .Z(n28623) );
  XOR U30674 ( .A(n[530]), .B(n28624), .Z(n28626) );
  XNOR U30675 ( .A(n28624), .B(n23989), .Z(n28625) );
  XOR U30676 ( .A(n28627), .B(n28628), .Z(n28624) );
  AND U30677 ( .A(n28629), .B(n28630), .Z(n28627) );
  XOR U30678 ( .A(n[529]), .B(n28628), .Z(n28630) );
  XNOR U30679 ( .A(n28628), .B(n23994), .Z(n28629) );
  XOR U30680 ( .A(n28631), .B(n28632), .Z(n28628) );
  AND U30681 ( .A(n28633), .B(n28634), .Z(n28631) );
  XOR U30682 ( .A(n[528]), .B(n28632), .Z(n28634) );
  XNOR U30683 ( .A(n28632), .B(n23999), .Z(n28633) );
  XOR U30684 ( .A(n28635), .B(n28636), .Z(n28632) );
  AND U30685 ( .A(n28637), .B(n28638), .Z(n28635) );
  XOR U30686 ( .A(n[527]), .B(n28636), .Z(n28638) );
  XNOR U30687 ( .A(n28636), .B(n24004), .Z(n28637) );
  XOR U30688 ( .A(n28639), .B(n28640), .Z(n28636) );
  AND U30689 ( .A(n28641), .B(n28642), .Z(n28639) );
  XOR U30690 ( .A(n[526]), .B(n28640), .Z(n28642) );
  XNOR U30691 ( .A(n28640), .B(n24009), .Z(n28641) );
  XOR U30692 ( .A(n28643), .B(n28644), .Z(n28640) );
  AND U30693 ( .A(n28645), .B(n28646), .Z(n28643) );
  XOR U30694 ( .A(n[525]), .B(n28644), .Z(n28646) );
  XNOR U30695 ( .A(n28644), .B(n24014), .Z(n28645) );
  XOR U30696 ( .A(n28647), .B(n28648), .Z(n28644) );
  AND U30697 ( .A(n28649), .B(n28650), .Z(n28647) );
  XOR U30698 ( .A(n[524]), .B(n28648), .Z(n28650) );
  XNOR U30699 ( .A(n28648), .B(n24019), .Z(n28649) );
  XOR U30700 ( .A(n28651), .B(n28652), .Z(n28648) );
  AND U30701 ( .A(n28653), .B(n28654), .Z(n28651) );
  XOR U30702 ( .A(n[523]), .B(n28652), .Z(n28654) );
  XNOR U30703 ( .A(n28652), .B(n24024), .Z(n28653) );
  XOR U30704 ( .A(n28655), .B(n28656), .Z(n28652) );
  AND U30705 ( .A(n28657), .B(n28658), .Z(n28655) );
  XOR U30706 ( .A(n[522]), .B(n28656), .Z(n28658) );
  XNOR U30707 ( .A(n28656), .B(n24029), .Z(n28657) );
  XOR U30708 ( .A(n28659), .B(n28660), .Z(n28656) );
  AND U30709 ( .A(n28661), .B(n28662), .Z(n28659) );
  XOR U30710 ( .A(n[521]), .B(n28660), .Z(n28662) );
  XNOR U30711 ( .A(n28660), .B(n24034), .Z(n28661) );
  XOR U30712 ( .A(n28663), .B(n28664), .Z(n28660) );
  AND U30713 ( .A(n28665), .B(n28666), .Z(n28663) );
  XOR U30714 ( .A(n[520]), .B(n28664), .Z(n28666) );
  XNOR U30715 ( .A(n28664), .B(n24039), .Z(n28665) );
  XOR U30716 ( .A(n28667), .B(n28668), .Z(n28664) );
  AND U30717 ( .A(n28669), .B(n28670), .Z(n28667) );
  XOR U30718 ( .A(n[519]), .B(n28668), .Z(n28670) );
  XNOR U30719 ( .A(n28668), .B(n24044), .Z(n28669) );
  XOR U30720 ( .A(n28671), .B(n28672), .Z(n28668) );
  AND U30721 ( .A(n28673), .B(n28674), .Z(n28671) );
  XOR U30722 ( .A(n[518]), .B(n28672), .Z(n28674) );
  XNOR U30723 ( .A(n28672), .B(n24049), .Z(n28673) );
  XOR U30724 ( .A(n28675), .B(n28676), .Z(n28672) );
  AND U30725 ( .A(n28677), .B(n28678), .Z(n28675) );
  XOR U30726 ( .A(n[517]), .B(n28676), .Z(n28678) );
  XNOR U30727 ( .A(n28676), .B(n24054), .Z(n28677) );
  XOR U30728 ( .A(n28679), .B(n28680), .Z(n28676) );
  AND U30729 ( .A(n28681), .B(n28682), .Z(n28679) );
  XOR U30730 ( .A(n[516]), .B(n28680), .Z(n28682) );
  XNOR U30731 ( .A(n28680), .B(n24059), .Z(n28681) );
  XOR U30732 ( .A(n28683), .B(n28684), .Z(n28680) );
  AND U30733 ( .A(n28685), .B(n28686), .Z(n28683) );
  XOR U30734 ( .A(n[515]), .B(n28684), .Z(n28686) );
  XNOR U30735 ( .A(n28684), .B(n24064), .Z(n28685) );
  XOR U30736 ( .A(n28687), .B(n28688), .Z(n28684) );
  AND U30737 ( .A(n28689), .B(n28690), .Z(n28687) );
  XOR U30738 ( .A(n[514]), .B(n28688), .Z(n28690) );
  XNOR U30739 ( .A(n28688), .B(n24069), .Z(n28689) );
  XOR U30740 ( .A(n28691), .B(n28692), .Z(n28688) );
  AND U30741 ( .A(n28693), .B(n28694), .Z(n28691) );
  XOR U30742 ( .A(n[513]), .B(n28692), .Z(n28694) );
  XNOR U30743 ( .A(n28692), .B(n24074), .Z(n28693) );
  XOR U30744 ( .A(n28695), .B(n28696), .Z(n28692) );
  AND U30745 ( .A(n28697), .B(n28698), .Z(n28695) );
  XOR U30746 ( .A(n[512]), .B(n28696), .Z(n28698) );
  XNOR U30747 ( .A(n28696), .B(n24079), .Z(n28697) );
  XOR U30748 ( .A(n28699), .B(n28700), .Z(n28696) );
  AND U30749 ( .A(n28701), .B(n28702), .Z(n28699) );
  XOR U30750 ( .A(n[511]), .B(n28700), .Z(n28702) );
  XNOR U30751 ( .A(n28700), .B(n24084), .Z(n28701) );
  XOR U30752 ( .A(n28703), .B(n28704), .Z(n28700) );
  AND U30753 ( .A(n28705), .B(n28706), .Z(n28703) );
  XOR U30754 ( .A(n[510]), .B(n28704), .Z(n28706) );
  XNOR U30755 ( .A(n28704), .B(n24089), .Z(n28705) );
  XOR U30756 ( .A(n28707), .B(n28708), .Z(n28704) );
  AND U30757 ( .A(n28709), .B(n28710), .Z(n28707) );
  XOR U30758 ( .A(n[509]), .B(n28708), .Z(n28710) );
  XNOR U30759 ( .A(n28708), .B(n24094), .Z(n28709) );
  XOR U30760 ( .A(n28711), .B(n28712), .Z(n28708) );
  AND U30761 ( .A(n28713), .B(n28714), .Z(n28711) );
  XOR U30762 ( .A(n[508]), .B(n28712), .Z(n28714) );
  XNOR U30763 ( .A(n28712), .B(n24099), .Z(n28713) );
  XOR U30764 ( .A(n28715), .B(n28716), .Z(n28712) );
  AND U30765 ( .A(n28717), .B(n28718), .Z(n28715) );
  XOR U30766 ( .A(n[507]), .B(n28716), .Z(n28718) );
  XNOR U30767 ( .A(n28716), .B(n24104), .Z(n28717) );
  XOR U30768 ( .A(n28719), .B(n28720), .Z(n28716) );
  AND U30769 ( .A(n28721), .B(n28722), .Z(n28719) );
  XOR U30770 ( .A(n[506]), .B(n28720), .Z(n28722) );
  XNOR U30771 ( .A(n28720), .B(n24109), .Z(n28721) );
  XOR U30772 ( .A(n28723), .B(n28724), .Z(n28720) );
  AND U30773 ( .A(n28725), .B(n28726), .Z(n28723) );
  XOR U30774 ( .A(n[505]), .B(n28724), .Z(n28726) );
  XNOR U30775 ( .A(n28724), .B(n24114), .Z(n28725) );
  XOR U30776 ( .A(n28727), .B(n28728), .Z(n28724) );
  AND U30777 ( .A(n28729), .B(n28730), .Z(n28727) );
  XOR U30778 ( .A(n[504]), .B(n28728), .Z(n28730) );
  XNOR U30779 ( .A(n28728), .B(n24119), .Z(n28729) );
  XOR U30780 ( .A(n28731), .B(n28732), .Z(n28728) );
  AND U30781 ( .A(n28733), .B(n28734), .Z(n28731) );
  XOR U30782 ( .A(n[503]), .B(n28732), .Z(n28734) );
  XNOR U30783 ( .A(n28732), .B(n24124), .Z(n28733) );
  XOR U30784 ( .A(n28735), .B(n28736), .Z(n28732) );
  AND U30785 ( .A(n28737), .B(n28738), .Z(n28735) );
  XOR U30786 ( .A(n[502]), .B(n28736), .Z(n28738) );
  XNOR U30787 ( .A(n28736), .B(n24129), .Z(n28737) );
  XOR U30788 ( .A(n28739), .B(n28740), .Z(n28736) );
  AND U30789 ( .A(n28741), .B(n28742), .Z(n28739) );
  XOR U30790 ( .A(n[501]), .B(n28740), .Z(n28742) );
  XNOR U30791 ( .A(n28740), .B(n24134), .Z(n28741) );
  XOR U30792 ( .A(n28743), .B(n28744), .Z(n28740) );
  AND U30793 ( .A(n28745), .B(n28746), .Z(n28743) );
  XOR U30794 ( .A(n[500]), .B(n28744), .Z(n28746) );
  XNOR U30795 ( .A(n28744), .B(n24139), .Z(n28745) );
  XOR U30796 ( .A(n28747), .B(n28748), .Z(n28744) );
  AND U30797 ( .A(n28749), .B(n28750), .Z(n28747) );
  XOR U30798 ( .A(n[499]), .B(n28748), .Z(n28750) );
  XNOR U30799 ( .A(n28748), .B(n24144), .Z(n28749) );
  XOR U30800 ( .A(n28751), .B(n28752), .Z(n28748) );
  AND U30801 ( .A(n28753), .B(n28754), .Z(n28751) );
  XOR U30802 ( .A(n[498]), .B(n28752), .Z(n28754) );
  XNOR U30803 ( .A(n28752), .B(n24149), .Z(n28753) );
  XOR U30804 ( .A(n28755), .B(n28756), .Z(n28752) );
  AND U30805 ( .A(n28757), .B(n28758), .Z(n28755) );
  XOR U30806 ( .A(n[497]), .B(n28756), .Z(n28758) );
  XNOR U30807 ( .A(n28756), .B(n24154), .Z(n28757) );
  XOR U30808 ( .A(n28759), .B(n28760), .Z(n28756) );
  AND U30809 ( .A(n28761), .B(n28762), .Z(n28759) );
  XOR U30810 ( .A(n[496]), .B(n28760), .Z(n28762) );
  XNOR U30811 ( .A(n28760), .B(n24159), .Z(n28761) );
  XOR U30812 ( .A(n28763), .B(n28764), .Z(n28760) );
  AND U30813 ( .A(n28765), .B(n28766), .Z(n28763) );
  XOR U30814 ( .A(n[495]), .B(n28764), .Z(n28766) );
  XNOR U30815 ( .A(n28764), .B(n24164), .Z(n28765) );
  XOR U30816 ( .A(n28767), .B(n28768), .Z(n28764) );
  AND U30817 ( .A(n28769), .B(n28770), .Z(n28767) );
  XOR U30818 ( .A(n[494]), .B(n28768), .Z(n28770) );
  XNOR U30819 ( .A(n28768), .B(n24169), .Z(n28769) );
  XOR U30820 ( .A(n28771), .B(n28772), .Z(n28768) );
  AND U30821 ( .A(n28773), .B(n28774), .Z(n28771) );
  XOR U30822 ( .A(n[493]), .B(n28772), .Z(n28774) );
  XNOR U30823 ( .A(n28772), .B(n24174), .Z(n28773) );
  XOR U30824 ( .A(n28775), .B(n28776), .Z(n28772) );
  AND U30825 ( .A(n28777), .B(n28778), .Z(n28775) );
  XOR U30826 ( .A(n[492]), .B(n28776), .Z(n28778) );
  XNOR U30827 ( .A(n28776), .B(n24179), .Z(n28777) );
  XOR U30828 ( .A(n28779), .B(n28780), .Z(n28776) );
  AND U30829 ( .A(n28781), .B(n28782), .Z(n28779) );
  XOR U30830 ( .A(n[491]), .B(n28780), .Z(n28782) );
  XNOR U30831 ( .A(n28780), .B(n24184), .Z(n28781) );
  XOR U30832 ( .A(n28783), .B(n28784), .Z(n28780) );
  AND U30833 ( .A(n28785), .B(n28786), .Z(n28783) );
  XOR U30834 ( .A(n[490]), .B(n28784), .Z(n28786) );
  XNOR U30835 ( .A(n28784), .B(n24189), .Z(n28785) );
  XOR U30836 ( .A(n28787), .B(n28788), .Z(n28784) );
  AND U30837 ( .A(n28789), .B(n28790), .Z(n28787) );
  XOR U30838 ( .A(n[489]), .B(n28788), .Z(n28790) );
  XNOR U30839 ( .A(n28788), .B(n24194), .Z(n28789) );
  XOR U30840 ( .A(n28791), .B(n28792), .Z(n28788) );
  AND U30841 ( .A(n28793), .B(n28794), .Z(n28791) );
  XOR U30842 ( .A(n[488]), .B(n28792), .Z(n28794) );
  XNOR U30843 ( .A(n28792), .B(n24199), .Z(n28793) );
  XOR U30844 ( .A(n28795), .B(n28796), .Z(n28792) );
  AND U30845 ( .A(n28797), .B(n28798), .Z(n28795) );
  XOR U30846 ( .A(n[487]), .B(n28796), .Z(n28798) );
  XNOR U30847 ( .A(n28796), .B(n24204), .Z(n28797) );
  XOR U30848 ( .A(n28799), .B(n28800), .Z(n28796) );
  AND U30849 ( .A(n28801), .B(n28802), .Z(n28799) );
  XOR U30850 ( .A(n[486]), .B(n28800), .Z(n28802) );
  XNOR U30851 ( .A(n28800), .B(n24209), .Z(n28801) );
  XOR U30852 ( .A(n28803), .B(n28804), .Z(n28800) );
  AND U30853 ( .A(n28805), .B(n28806), .Z(n28803) );
  XOR U30854 ( .A(n[485]), .B(n28804), .Z(n28806) );
  XNOR U30855 ( .A(n28804), .B(n24214), .Z(n28805) );
  XOR U30856 ( .A(n28807), .B(n28808), .Z(n28804) );
  AND U30857 ( .A(n28809), .B(n28810), .Z(n28807) );
  XOR U30858 ( .A(n[484]), .B(n28808), .Z(n28810) );
  XNOR U30859 ( .A(n28808), .B(n24219), .Z(n28809) );
  XOR U30860 ( .A(n28811), .B(n28812), .Z(n28808) );
  AND U30861 ( .A(n28813), .B(n28814), .Z(n28811) );
  XOR U30862 ( .A(n[483]), .B(n28812), .Z(n28814) );
  XNOR U30863 ( .A(n28812), .B(n24224), .Z(n28813) );
  XOR U30864 ( .A(n28815), .B(n28816), .Z(n28812) );
  AND U30865 ( .A(n28817), .B(n28818), .Z(n28815) );
  XOR U30866 ( .A(n[482]), .B(n28816), .Z(n28818) );
  XNOR U30867 ( .A(n28816), .B(n24229), .Z(n28817) );
  XOR U30868 ( .A(n28819), .B(n28820), .Z(n28816) );
  AND U30869 ( .A(n28821), .B(n28822), .Z(n28819) );
  XOR U30870 ( .A(n[481]), .B(n28820), .Z(n28822) );
  XNOR U30871 ( .A(n28820), .B(n24234), .Z(n28821) );
  XOR U30872 ( .A(n28823), .B(n28824), .Z(n28820) );
  AND U30873 ( .A(n28825), .B(n28826), .Z(n28823) );
  XOR U30874 ( .A(n[480]), .B(n28824), .Z(n28826) );
  XNOR U30875 ( .A(n28824), .B(n24239), .Z(n28825) );
  XOR U30876 ( .A(n28827), .B(n28828), .Z(n28824) );
  AND U30877 ( .A(n28829), .B(n28830), .Z(n28827) );
  XOR U30878 ( .A(n[479]), .B(n28828), .Z(n28830) );
  XNOR U30879 ( .A(n28828), .B(n24244), .Z(n28829) );
  XOR U30880 ( .A(n28831), .B(n28832), .Z(n28828) );
  AND U30881 ( .A(n28833), .B(n28834), .Z(n28831) );
  XOR U30882 ( .A(n[478]), .B(n28832), .Z(n28834) );
  XNOR U30883 ( .A(n28832), .B(n24249), .Z(n28833) );
  XOR U30884 ( .A(n28835), .B(n28836), .Z(n28832) );
  AND U30885 ( .A(n28837), .B(n28838), .Z(n28835) );
  XOR U30886 ( .A(n[477]), .B(n28836), .Z(n28838) );
  XNOR U30887 ( .A(n28836), .B(n24254), .Z(n28837) );
  XOR U30888 ( .A(n28839), .B(n28840), .Z(n28836) );
  AND U30889 ( .A(n28841), .B(n28842), .Z(n28839) );
  XOR U30890 ( .A(n[476]), .B(n28840), .Z(n28842) );
  XNOR U30891 ( .A(n28840), .B(n24259), .Z(n28841) );
  XOR U30892 ( .A(n28843), .B(n28844), .Z(n28840) );
  AND U30893 ( .A(n28845), .B(n28846), .Z(n28843) );
  XOR U30894 ( .A(n[475]), .B(n28844), .Z(n28846) );
  XNOR U30895 ( .A(n28844), .B(n24264), .Z(n28845) );
  XOR U30896 ( .A(n28847), .B(n28848), .Z(n28844) );
  AND U30897 ( .A(n28849), .B(n28850), .Z(n28847) );
  XOR U30898 ( .A(n[474]), .B(n28848), .Z(n28850) );
  XNOR U30899 ( .A(n28848), .B(n24269), .Z(n28849) );
  XOR U30900 ( .A(n28851), .B(n28852), .Z(n28848) );
  AND U30901 ( .A(n28853), .B(n28854), .Z(n28851) );
  XOR U30902 ( .A(n[473]), .B(n28852), .Z(n28854) );
  XNOR U30903 ( .A(n28852), .B(n24274), .Z(n28853) );
  XOR U30904 ( .A(n28855), .B(n28856), .Z(n28852) );
  AND U30905 ( .A(n28857), .B(n28858), .Z(n28855) );
  XOR U30906 ( .A(n[472]), .B(n28856), .Z(n28858) );
  XNOR U30907 ( .A(n28856), .B(n24279), .Z(n28857) );
  XOR U30908 ( .A(n28859), .B(n28860), .Z(n28856) );
  AND U30909 ( .A(n28861), .B(n28862), .Z(n28859) );
  XOR U30910 ( .A(n[471]), .B(n28860), .Z(n28862) );
  XNOR U30911 ( .A(n28860), .B(n24284), .Z(n28861) );
  XOR U30912 ( .A(n28863), .B(n28864), .Z(n28860) );
  AND U30913 ( .A(n28865), .B(n28866), .Z(n28863) );
  XOR U30914 ( .A(n[470]), .B(n28864), .Z(n28866) );
  XNOR U30915 ( .A(n28864), .B(n24289), .Z(n28865) );
  XOR U30916 ( .A(n28867), .B(n28868), .Z(n28864) );
  AND U30917 ( .A(n28869), .B(n28870), .Z(n28867) );
  XOR U30918 ( .A(n[469]), .B(n28868), .Z(n28870) );
  XNOR U30919 ( .A(n28868), .B(n24294), .Z(n28869) );
  XOR U30920 ( .A(n28871), .B(n28872), .Z(n28868) );
  AND U30921 ( .A(n28873), .B(n28874), .Z(n28871) );
  XOR U30922 ( .A(n[468]), .B(n28872), .Z(n28874) );
  XNOR U30923 ( .A(n28872), .B(n24299), .Z(n28873) );
  XOR U30924 ( .A(n28875), .B(n28876), .Z(n28872) );
  AND U30925 ( .A(n28877), .B(n28878), .Z(n28875) );
  XOR U30926 ( .A(n[467]), .B(n28876), .Z(n28878) );
  XNOR U30927 ( .A(n28876), .B(n24304), .Z(n28877) );
  XOR U30928 ( .A(n28879), .B(n28880), .Z(n28876) );
  AND U30929 ( .A(n28881), .B(n28882), .Z(n28879) );
  XOR U30930 ( .A(n[466]), .B(n28880), .Z(n28882) );
  XNOR U30931 ( .A(n28880), .B(n24309), .Z(n28881) );
  XOR U30932 ( .A(n28883), .B(n28884), .Z(n28880) );
  AND U30933 ( .A(n28885), .B(n28886), .Z(n28883) );
  XOR U30934 ( .A(n[465]), .B(n28884), .Z(n28886) );
  XNOR U30935 ( .A(n28884), .B(n24314), .Z(n28885) );
  XOR U30936 ( .A(n28887), .B(n28888), .Z(n28884) );
  AND U30937 ( .A(n28889), .B(n28890), .Z(n28887) );
  XOR U30938 ( .A(n[464]), .B(n28888), .Z(n28890) );
  XNOR U30939 ( .A(n28888), .B(n24319), .Z(n28889) );
  XOR U30940 ( .A(n28891), .B(n28892), .Z(n28888) );
  AND U30941 ( .A(n28893), .B(n28894), .Z(n28891) );
  XOR U30942 ( .A(n[463]), .B(n28892), .Z(n28894) );
  XNOR U30943 ( .A(n28892), .B(n24324), .Z(n28893) );
  XOR U30944 ( .A(n28895), .B(n28896), .Z(n28892) );
  AND U30945 ( .A(n28897), .B(n28898), .Z(n28895) );
  XOR U30946 ( .A(n[462]), .B(n28896), .Z(n28898) );
  XNOR U30947 ( .A(n28896), .B(n24329), .Z(n28897) );
  XOR U30948 ( .A(n28899), .B(n28900), .Z(n28896) );
  AND U30949 ( .A(n28901), .B(n28902), .Z(n28899) );
  XOR U30950 ( .A(n[461]), .B(n28900), .Z(n28902) );
  XNOR U30951 ( .A(n28900), .B(n24334), .Z(n28901) );
  XOR U30952 ( .A(n28903), .B(n28904), .Z(n28900) );
  AND U30953 ( .A(n28905), .B(n28906), .Z(n28903) );
  XOR U30954 ( .A(n[460]), .B(n28904), .Z(n28906) );
  XNOR U30955 ( .A(n28904), .B(n24339), .Z(n28905) );
  XOR U30956 ( .A(n28907), .B(n28908), .Z(n28904) );
  AND U30957 ( .A(n28909), .B(n28910), .Z(n28907) );
  XOR U30958 ( .A(n[459]), .B(n28908), .Z(n28910) );
  XNOR U30959 ( .A(n28908), .B(n24344), .Z(n28909) );
  XOR U30960 ( .A(n28911), .B(n28912), .Z(n28908) );
  AND U30961 ( .A(n28913), .B(n28914), .Z(n28911) );
  XOR U30962 ( .A(n[458]), .B(n28912), .Z(n28914) );
  XNOR U30963 ( .A(n28912), .B(n24349), .Z(n28913) );
  XOR U30964 ( .A(n28915), .B(n28916), .Z(n28912) );
  AND U30965 ( .A(n28917), .B(n28918), .Z(n28915) );
  XOR U30966 ( .A(n[457]), .B(n28916), .Z(n28918) );
  XNOR U30967 ( .A(n28916), .B(n24354), .Z(n28917) );
  XOR U30968 ( .A(n28919), .B(n28920), .Z(n28916) );
  AND U30969 ( .A(n28921), .B(n28922), .Z(n28919) );
  XOR U30970 ( .A(n[456]), .B(n28920), .Z(n28922) );
  XNOR U30971 ( .A(n28920), .B(n24359), .Z(n28921) );
  XOR U30972 ( .A(n28923), .B(n28924), .Z(n28920) );
  AND U30973 ( .A(n28925), .B(n28926), .Z(n28923) );
  XOR U30974 ( .A(n[455]), .B(n28924), .Z(n28926) );
  XNOR U30975 ( .A(n28924), .B(n24364), .Z(n28925) );
  XOR U30976 ( .A(n28927), .B(n28928), .Z(n28924) );
  AND U30977 ( .A(n28929), .B(n28930), .Z(n28927) );
  XOR U30978 ( .A(n[454]), .B(n28928), .Z(n28930) );
  XNOR U30979 ( .A(n28928), .B(n24369), .Z(n28929) );
  XOR U30980 ( .A(n28931), .B(n28932), .Z(n28928) );
  AND U30981 ( .A(n28933), .B(n28934), .Z(n28931) );
  XOR U30982 ( .A(n[453]), .B(n28932), .Z(n28934) );
  XNOR U30983 ( .A(n28932), .B(n24374), .Z(n28933) );
  XOR U30984 ( .A(n28935), .B(n28936), .Z(n28932) );
  AND U30985 ( .A(n28937), .B(n28938), .Z(n28935) );
  XOR U30986 ( .A(n[452]), .B(n28936), .Z(n28938) );
  XNOR U30987 ( .A(n28936), .B(n24379), .Z(n28937) );
  XOR U30988 ( .A(n28939), .B(n28940), .Z(n28936) );
  AND U30989 ( .A(n28941), .B(n28942), .Z(n28939) );
  XOR U30990 ( .A(n[451]), .B(n28940), .Z(n28942) );
  XNOR U30991 ( .A(n28940), .B(n24384), .Z(n28941) );
  XOR U30992 ( .A(n28943), .B(n28944), .Z(n28940) );
  AND U30993 ( .A(n28945), .B(n28946), .Z(n28943) );
  XOR U30994 ( .A(n[450]), .B(n28944), .Z(n28946) );
  XNOR U30995 ( .A(n28944), .B(n24389), .Z(n28945) );
  XOR U30996 ( .A(n28947), .B(n28948), .Z(n28944) );
  AND U30997 ( .A(n28949), .B(n28950), .Z(n28947) );
  XOR U30998 ( .A(n[449]), .B(n28948), .Z(n28950) );
  XNOR U30999 ( .A(n28948), .B(n24394), .Z(n28949) );
  XOR U31000 ( .A(n28951), .B(n28952), .Z(n28948) );
  AND U31001 ( .A(n28953), .B(n28954), .Z(n28951) );
  XOR U31002 ( .A(n[448]), .B(n28952), .Z(n28954) );
  XNOR U31003 ( .A(n28952), .B(n24399), .Z(n28953) );
  XOR U31004 ( .A(n28955), .B(n28956), .Z(n28952) );
  AND U31005 ( .A(n28957), .B(n28958), .Z(n28955) );
  XOR U31006 ( .A(n[447]), .B(n28956), .Z(n28958) );
  XNOR U31007 ( .A(n28956), .B(n24404), .Z(n28957) );
  XOR U31008 ( .A(n28959), .B(n28960), .Z(n28956) );
  AND U31009 ( .A(n28961), .B(n28962), .Z(n28959) );
  XOR U31010 ( .A(n[446]), .B(n28960), .Z(n28962) );
  XNOR U31011 ( .A(n28960), .B(n24409), .Z(n28961) );
  XOR U31012 ( .A(n28963), .B(n28964), .Z(n28960) );
  AND U31013 ( .A(n28965), .B(n28966), .Z(n28963) );
  XOR U31014 ( .A(n[445]), .B(n28964), .Z(n28966) );
  XNOR U31015 ( .A(n28964), .B(n24414), .Z(n28965) );
  XOR U31016 ( .A(n28967), .B(n28968), .Z(n28964) );
  AND U31017 ( .A(n28969), .B(n28970), .Z(n28967) );
  XOR U31018 ( .A(n[444]), .B(n28968), .Z(n28970) );
  XNOR U31019 ( .A(n28968), .B(n24419), .Z(n28969) );
  XOR U31020 ( .A(n28971), .B(n28972), .Z(n28968) );
  AND U31021 ( .A(n28973), .B(n28974), .Z(n28971) );
  XOR U31022 ( .A(n[443]), .B(n28972), .Z(n28974) );
  XNOR U31023 ( .A(n28972), .B(n24424), .Z(n28973) );
  XOR U31024 ( .A(n28975), .B(n28976), .Z(n28972) );
  AND U31025 ( .A(n28977), .B(n28978), .Z(n28975) );
  XOR U31026 ( .A(n[442]), .B(n28976), .Z(n28978) );
  XNOR U31027 ( .A(n28976), .B(n24429), .Z(n28977) );
  XOR U31028 ( .A(n28979), .B(n28980), .Z(n28976) );
  AND U31029 ( .A(n28981), .B(n28982), .Z(n28979) );
  XOR U31030 ( .A(n[441]), .B(n28980), .Z(n28982) );
  XNOR U31031 ( .A(n28980), .B(n24434), .Z(n28981) );
  XOR U31032 ( .A(n28983), .B(n28984), .Z(n28980) );
  AND U31033 ( .A(n28985), .B(n28986), .Z(n28983) );
  XOR U31034 ( .A(n[440]), .B(n28984), .Z(n28986) );
  XNOR U31035 ( .A(n28984), .B(n24439), .Z(n28985) );
  XOR U31036 ( .A(n28987), .B(n28988), .Z(n28984) );
  AND U31037 ( .A(n28989), .B(n28990), .Z(n28987) );
  XOR U31038 ( .A(n[439]), .B(n28988), .Z(n28990) );
  XNOR U31039 ( .A(n28988), .B(n24444), .Z(n28989) );
  XOR U31040 ( .A(n28991), .B(n28992), .Z(n28988) );
  AND U31041 ( .A(n28993), .B(n28994), .Z(n28991) );
  XOR U31042 ( .A(n[438]), .B(n28992), .Z(n28994) );
  XNOR U31043 ( .A(n28992), .B(n24449), .Z(n28993) );
  XOR U31044 ( .A(n28995), .B(n28996), .Z(n28992) );
  AND U31045 ( .A(n28997), .B(n28998), .Z(n28995) );
  XOR U31046 ( .A(n[437]), .B(n28996), .Z(n28998) );
  XNOR U31047 ( .A(n28996), .B(n24454), .Z(n28997) );
  XOR U31048 ( .A(n28999), .B(n29000), .Z(n28996) );
  AND U31049 ( .A(n29001), .B(n29002), .Z(n28999) );
  XOR U31050 ( .A(n[436]), .B(n29000), .Z(n29002) );
  XNOR U31051 ( .A(n29000), .B(n24459), .Z(n29001) );
  XOR U31052 ( .A(n29003), .B(n29004), .Z(n29000) );
  AND U31053 ( .A(n29005), .B(n29006), .Z(n29003) );
  XOR U31054 ( .A(n[435]), .B(n29004), .Z(n29006) );
  XNOR U31055 ( .A(n29004), .B(n24464), .Z(n29005) );
  XOR U31056 ( .A(n29007), .B(n29008), .Z(n29004) );
  AND U31057 ( .A(n29009), .B(n29010), .Z(n29007) );
  XOR U31058 ( .A(n[434]), .B(n29008), .Z(n29010) );
  XNOR U31059 ( .A(n29008), .B(n24469), .Z(n29009) );
  XOR U31060 ( .A(n29011), .B(n29012), .Z(n29008) );
  AND U31061 ( .A(n29013), .B(n29014), .Z(n29011) );
  XOR U31062 ( .A(n[433]), .B(n29012), .Z(n29014) );
  XNOR U31063 ( .A(n29012), .B(n24474), .Z(n29013) );
  XOR U31064 ( .A(n29015), .B(n29016), .Z(n29012) );
  AND U31065 ( .A(n29017), .B(n29018), .Z(n29015) );
  XOR U31066 ( .A(n[432]), .B(n29016), .Z(n29018) );
  XNOR U31067 ( .A(n29016), .B(n24479), .Z(n29017) );
  XOR U31068 ( .A(n29019), .B(n29020), .Z(n29016) );
  AND U31069 ( .A(n29021), .B(n29022), .Z(n29019) );
  XOR U31070 ( .A(n[431]), .B(n29020), .Z(n29022) );
  XNOR U31071 ( .A(n29020), .B(n24484), .Z(n29021) );
  XOR U31072 ( .A(n29023), .B(n29024), .Z(n29020) );
  AND U31073 ( .A(n29025), .B(n29026), .Z(n29023) );
  XOR U31074 ( .A(n[430]), .B(n29024), .Z(n29026) );
  XNOR U31075 ( .A(n29024), .B(n24489), .Z(n29025) );
  XOR U31076 ( .A(n29027), .B(n29028), .Z(n29024) );
  AND U31077 ( .A(n29029), .B(n29030), .Z(n29027) );
  XOR U31078 ( .A(n[429]), .B(n29028), .Z(n29030) );
  XNOR U31079 ( .A(n29028), .B(n24494), .Z(n29029) );
  XOR U31080 ( .A(n29031), .B(n29032), .Z(n29028) );
  AND U31081 ( .A(n29033), .B(n29034), .Z(n29031) );
  XOR U31082 ( .A(n[428]), .B(n29032), .Z(n29034) );
  XNOR U31083 ( .A(n29032), .B(n24499), .Z(n29033) );
  XOR U31084 ( .A(n29035), .B(n29036), .Z(n29032) );
  AND U31085 ( .A(n29037), .B(n29038), .Z(n29035) );
  XOR U31086 ( .A(n[427]), .B(n29036), .Z(n29038) );
  XNOR U31087 ( .A(n29036), .B(n24504), .Z(n29037) );
  XOR U31088 ( .A(n29039), .B(n29040), .Z(n29036) );
  AND U31089 ( .A(n29041), .B(n29042), .Z(n29039) );
  XOR U31090 ( .A(n[426]), .B(n29040), .Z(n29042) );
  XNOR U31091 ( .A(n29040), .B(n24509), .Z(n29041) );
  XOR U31092 ( .A(n29043), .B(n29044), .Z(n29040) );
  AND U31093 ( .A(n29045), .B(n29046), .Z(n29043) );
  XOR U31094 ( .A(n[425]), .B(n29044), .Z(n29046) );
  XNOR U31095 ( .A(n29044), .B(n24514), .Z(n29045) );
  XOR U31096 ( .A(n29047), .B(n29048), .Z(n29044) );
  AND U31097 ( .A(n29049), .B(n29050), .Z(n29047) );
  XOR U31098 ( .A(n[424]), .B(n29048), .Z(n29050) );
  XNOR U31099 ( .A(n29048), .B(n24519), .Z(n29049) );
  XOR U31100 ( .A(n29051), .B(n29052), .Z(n29048) );
  AND U31101 ( .A(n29053), .B(n29054), .Z(n29051) );
  XOR U31102 ( .A(n[423]), .B(n29052), .Z(n29054) );
  XNOR U31103 ( .A(n29052), .B(n24524), .Z(n29053) );
  XOR U31104 ( .A(n29055), .B(n29056), .Z(n29052) );
  AND U31105 ( .A(n29057), .B(n29058), .Z(n29055) );
  XOR U31106 ( .A(n[422]), .B(n29056), .Z(n29058) );
  XNOR U31107 ( .A(n29056), .B(n24529), .Z(n29057) );
  XOR U31108 ( .A(n29059), .B(n29060), .Z(n29056) );
  AND U31109 ( .A(n29061), .B(n29062), .Z(n29059) );
  XOR U31110 ( .A(n[421]), .B(n29060), .Z(n29062) );
  XNOR U31111 ( .A(n29060), .B(n24534), .Z(n29061) );
  XOR U31112 ( .A(n29063), .B(n29064), .Z(n29060) );
  AND U31113 ( .A(n29065), .B(n29066), .Z(n29063) );
  XOR U31114 ( .A(n[420]), .B(n29064), .Z(n29066) );
  XNOR U31115 ( .A(n29064), .B(n24539), .Z(n29065) );
  XOR U31116 ( .A(n29067), .B(n29068), .Z(n29064) );
  AND U31117 ( .A(n29069), .B(n29070), .Z(n29067) );
  XOR U31118 ( .A(n[419]), .B(n29068), .Z(n29070) );
  XNOR U31119 ( .A(n29068), .B(n24544), .Z(n29069) );
  XOR U31120 ( .A(n29071), .B(n29072), .Z(n29068) );
  AND U31121 ( .A(n29073), .B(n29074), .Z(n29071) );
  XOR U31122 ( .A(n[418]), .B(n29072), .Z(n29074) );
  XNOR U31123 ( .A(n29072), .B(n24549), .Z(n29073) );
  XOR U31124 ( .A(n29075), .B(n29076), .Z(n29072) );
  AND U31125 ( .A(n29077), .B(n29078), .Z(n29075) );
  XOR U31126 ( .A(n[417]), .B(n29076), .Z(n29078) );
  XNOR U31127 ( .A(n29076), .B(n24554), .Z(n29077) );
  XOR U31128 ( .A(n29079), .B(n29080), .Z(n29076) );
  AND U31129 ( .A(n29081), .B(n29082), .Z(n29079) );
  XOR U31130 ( .A(n[416]), .B(n29080), .Z(n29082) );
  XNOR U31131 ( .A(n29080), .B(n24559), .Z(n29081) );
  XOR U31132 ( .A(n29083), .B(n29084), .Z(n29080) );
  AND U31133 ( .A(n29085), .B(n29086), .Z(n29083) );
  XOR U31134 ( .A(n[415]), .B(n29084), .Z(n29086) );
  XNOR U31135 ( .A(n29084), .B(n24564), .Z(n29085) );
  XOR U31136 ( .A(n29087), .B(n29088), .Z(n29084) );
  AND U31137 ( .A(n29089), .B(n29090), .Z(n29087) );
  XOR U31138 ( .A(n[414]), .B(n29088), .Z(n29090) );
  XNOR U31139 ( .A(n29088), .B(n24569), .Z(n29089) );
  XOR U31140 ( .A(n29091), .B(n29092), .Z(n29088) );
  AND U31141 ( .A(n29093), .B(n29094), .Z(n29091) );
  XOR U31142 ( .A(n[413]), .B(n29092), .Z(n29094) );
  XNOR U31143 ( .A(n29092), .B(n24574), .Z(n29093) );
  XOR U31144 ( .A(n29095), .B(n29096), .Z(n29092) );
  AND U31145 ( .A(n29097), .B(n29098), .Z(n29095) );
  XOR U31146 ( .A(n[412]), .B(n29096), .Z(n29098) );
  XNOR U31147 ( .A(n29096), .B(n24579), .Z(n29097) );
  XOR U31148 ( .A(n29099), .B(n29100), .Z(n29096) );
  AND U31149 ( .A(n29101), .B(n29102), .Z(n29099) );
  XOR U31150 ( .A(n[411]), .B(n29100), .Z(n29102) );
  XNOR U31151 ( .A(n29100), .B(n24584), .Z(n29101) );
  XOR U31152 ( .A(n29103), .B(n29104), .Z(n29100) );
  AND U31153 ( .A(n29105), .B(n29106), .Z(n29103) );
  XOR U31154 ( .A(n[410]), .B(n29104), .Z(n29106) );
  XNOR U31155 ( .A(n29104), .B(n24589), .Z(n29105) );
  XOR U31156 ( .A(n29107), .B(n29108), .Z(n29104) );
  AND U31157 ( .A(n29109), .B(n29110), .Z(n29107) );
  XOR U31158 ( .A(n[409]), .B(n29108), .Z(n29110) );
  XNOR U31159 ( .A(n29108), .B(n24594), .Z(n29109) );
  XOR U31160 ( .A(n29111), .B(n29112), .Z(n29108) );
  AND U31161 ( .A(n29113), .B(n29114), .Z(n29111) );
  XOR U31162 ( .A(n[408]), .B(n29112), .Z(n29114) );
  XNOR U31163 ( .A(n29112), .B(n24599), .Z(n29113) );
  XOR U31164 ( .A(n29115), .B(n29116), .Z(n29112) );
  AND U31165 ( .A(n29117), .B(n29118), .Z(n29115) );
  XOR U31166 ( .A(n[407]), .B(n29116), .Z(n29118) );
  XNOR U31167 ( .A(n29116), .B(n24604), .Z(n29117) );
  XOR U31168 ( .A(n29119), .B(n29120), .Z(n29116) );
  AND U31169 ( .A(n29121), .B(n29122), .Z(n29119) );
  XOR U31170 ( .A(n[406]), .B(n29120), .Z(n29122) );
  XNOR U31171 ( .A(n29120), .B(n24609), .Z(n29121) );
  XOR U31172 ( .A(n29123), .B(n29124), .Z(n29120) );
  AND U31173 ( .A(n29125), .B(n29126), .Z(n29123) );
  XOR U31174 ( .A(n[405]), .B(n29124), .Z(n29126) );
  XNOR U31175 ( .A(n29124), .B(n24614), .Z(n29125) );
  XOR U31176 ( .A(n29127), .B(n29128), .Z(n29124) );
  AND U31177 ( .A(n29129), .B(n29130), .Z(n29127) );
  XOR U31178 ( .A(n[404]), .B(n29128), .Z(n29130) );
  XNOR U31179 ( .A(n29128), .B(n24619), .Z(n29129) );
  XOR U31180 ( .A(n29131), .B(n29132), .Z(n29128) );
  AND U31181 ( .A(n29133), .B(n29134), .Z(n29131) );
  XOR U31182 ( .A(n[403]), .B(n29132), .Z(n29134) );
  XNOR U31183 ( .A(n29132), .B(n24624), .Z(n29133) );
  XOR U31184 ( .A(n29135), .B(n29136), .Z(n29132) );
  AND U31185 ( .A(n29137), .B(n29138), .Z(n29135) );
  XOR U31186 ( .A(n[402]), .B(n29136), .Z(n29138) );
  XNOR U31187 ( .A(n29136), .B(n24629), .Z(n29137) );
  XOR U31188 ( .A(n29139), .B(n29140), .Z(n29136) );
  AND U31189 ( .A(n29141), .B(n29142), .Z(n29139) );
  XOR U31190 ( .A(n[401]), .B(n29140), .Z(n29142) );
  XNOR U31191 ( .A(n29140), .B(n24634), .Z(n29141) );
  XOR U31192 ( .A(n29143), .B(n29144), .Z(n29140) );
  AND U31193 ( .A(n29145), .B(n29146), .Z(n29143) );
  XOR U31194 ( .A(n[400]), .B(n29144), .Z(n29146) );
  XNOR U31195 ( .A(n29144), .B(n24639), .Z(n29145) );
  XOR U31196 ( .A(n29147), .B(n29148), .Z(n29144) );
  AND U31197 ( .A(n29149), .B(n29150), .Z(n29147) );
  XOR U31198 ( .A(n[399]), .B(n29148), .Z(n29150) );
  XNOR U31199 ( .A(n29148), .B(n24644), .Z(n29149) );
  XOR U31200 ( .A(n29151), .B(n29152), .Z(n29148) );
  AND U31201 ( .A(n29153), .B(n29154), .Z(n29151) );
  XOR U31202 ( .A(n[398]), .B(n29152), .Z(n29154) );
  XNOR U31203 ( .A(n29152), .B(n24649), .Z(n29153) );
  XOR U31204 ( .A(n29155), .B(n29156), .Z(n29152) );
  AND U31205 ( .A(n29157), .B(n29158), .Z(n29155) );
  XOR U31206 ( .A(n[397]), .B(n29156), .Z(n29158) );
  XNOR U31207 ( .A(n29156), .B(n24654), .Z(n29157) );
  XOR U31208 ( .A(n29159), .B(n29160), .Z(n29156) );
  AND U31209 ( .A(n29161), .B(n29162), .Z(n29159) );
  XOR U31210 ( .A(n[396]), .B(n29160), .Z(n29162) );
  XNOR U31211 ( .A(n29160), .B(n24659), .Z(n29161) );
  XOR U31212 ( .A(n29163), .B(n29164), .Z(n29160) );
  AND U31213 ( .A(n29165), .B(n29166), .Z(n29163) );
  XOR U31214 ( .A(n[395]), .B(n29164), .Z(n29166) );
  XNOR U31215 ( .A(n29164), .B(n24664), .Z(n29165) );
  XOR U31216 ( .A(n29167), .B(n29168), .Z(n29164) );
  AND U31217 ( .A(n29169), .B(n29170), .Z(n29167) );
  XOR U31218 ( .A(n[394]), .B(n29168), .Z(n29170) );
  XNOR U31219 ( .A(n29168), .B(n24669), .Z(n29169) );
  XOR U31220 ( .A(n29171), .B(n29172), .Z(n29168) );
  AND U31221 ( .A(n29173), .B(n29174), .Z(n29171) );
  XOR U31222 ( .A(n[393]), .B(n29172), .Z(n29174) );
  XNOR U31223 ( .A(n29172), .B(n24674), .Z(n29173) );
  XOR U31224 ( .A(n29175), .B(n29176), .Z(n29172) );
  AND U31225 ( .A(n29177), .B(n29178), .Z(n29175) );
  XOR U31226 ( .A(n[392]), .B(n29176), .Z(n29178) );
  XNOR U31227 ( .A(n29176), .B(n24679), .Z(n29177) );
  XOR U31228 ( .A(n29179), .B(n29180), .Z(n29176) );
  AND U31229 ( .A(n29181), .B(n29182), .Z(n29179) );
  XOR U31230 ( .A(n[391]), .B(n29180), .Z(n29182) );
  XNOR U31231 ( .A(n29180), .B(n24684), .Z(n29181) );
  XOR U31232 ( .A(n29183), .B(n29184), .Z(n29180) );
  AND U31233 ( .A(n29185), .B(n29186), .Z(n29183) );
  XOR U31234 ( .A(n[390]), .B(n29184), .Z(n29186) );
  XNOR U31235 ( .A(n29184), .B(n24689), .Z(n29185) );
  XOR U31236 ( .A(n29187), .B(n29188), .Z(n29184) );
  AND U31237 ( .A(n29189), .B(n29190), .Z(n29187) );
  XOR U31238 ( .A(n[389]), .B(n29188), .Z(n29190) );
  XNOR U31239 ( .A(n29188), .B(n24694), .Z(n29189) );
  XOR U31240 ( .A(n29191), .B(n29192), .Z(n29188) );
  AND U31241 ( .A(n29193), .B(n29194), .Z(n29191) );
  XOR U31242 ( .A(n[388]), .B(n29192), .Z(n29194) );
  XNOR U31243 ( .A(n29192), .B(n24699), .Z(n29193) );
  XOR U31244 ( .A(n29195), .B(n29196), .Z(n29192) );
  AND U31245 ( .A(n29197), .B(n29198), .Z(n29195) );
  XOR U31246 ( .A(n[387]), .B(n29196), .Z(n29198) );
  XNOR U31247 ( .A(n29196), .B(n24704), .Z(n29197) );
  XOR U31248 ( .A(n29199), .B(n29200), .Z(n29196) );
  AND U31249 ( .A(n29201), .B(n29202), .Z(n29199) );
  XOR U31250 ( .A(n[386]), .B(n29200), .Z(n29202) );
  XNOR U31251 ( .A(n29200), .B(n24709), .Z(n29201) );
  XOR U31252 ( .A(n29203), .B(n29204), .Z(n29200) );
  AND U31253 ( .A(n29205), .B(n29206), .Z(n29203) );
  XOR U31254 ( .A(n[385]), .B(n29204), .Z(n29206) );
  XNOR U31255 ( .A(n29204), .B(n24714), .Z(n29205) );
  XOR U31256 ( .A(n29207), .B(n29208), .Z(n29204) );
  AND U31257 ( .A(n29209), .B(n29210), .Z(n29207) );
  XOR U31258 ( .A(n[384]), .B(n29208), .Z(n29210) );
  XNOR U31259 ( .A(n29208), .B(n24719), .Z(n29209) );
  XOR U31260 ( .A(n29211), .B(n29212), .Z(n29208) );
  AND U31261 ( .A(n29213), .B(n29214), .Z(n29211) );
  XOR U31262 ( .A(n[383]), .B(n29212), .Z(n29214) );
  XNOR U31263 ( .A(n29212), .B(n24724), .Z(n29213) );
  XOR U31264 ( .A(n29215), .B(n29216), .Z(n29212) );
  AND U31265 ( .A(n29217), .B(n29218), .Z(n29215) );
  XOR U31266 ( .A(n[382]), .B(n29216), .Z(n29218) );
  XNOR U31267 ( .A(n29216), .B(n24729), .Z(n29217) );
  XOR U31268 ( .A(n29219), .B(n29220), .Z(n29216) );
  AND U31269 ( .A(n29221), .B(n29222), .Z(n29219) );
  XOR U31270 ( .A(n[381]), .B(n29220), .Z(n29222) );
  XNOR U31271 ( .A(n29220), .B(n24734), .Z(n29221) );
  XOR U31272 ( .A(n29223), .B(n29224), .Z(n29220) );
  AND U31273 ( .A(n29225), .B(n29226), .Z(n29223) );
  XOR U31274 ( .A(n[380]), .B(n29224), .Z(n29226) );
  XNOR U31275 ( .A(n29224), .B(n24739), .Z(n29225) );
  XOR U31276 ( .A(n29227), .B(n29228), .Z(n29224) );
  AND U31277 ( .A(n29229), .B(n29230), .Z(n29227) );
  XOR U31278 ( .A(n[379]), .B(n29228), .Z(n29230) );
  XNOR U31279 ( .A(n29228), .B(n24744), .Z(n29229) );
  XOR U31280 ( .A(n29231), .B(n29232), .Z(n29228) );
  AND U31281 ( .A(n29233), .B(n29234), .Z(n29231) );
  XOR U31282 ( .A(n[378]), .B(n29232), .Z(n29234) );
  XNOR U31283 ( .A(n29232), .B(n24749), .Z(n29233) );
  XOR U31284 ( .A(n29235), .B(n29236), .Z(n29232) );
  AND U31285 ( .A(n29237), .B(n29238), .Z(n29235) );
  XOR U31286 ( .A(n[377]), .B(n29236), .Z(n29238) );
  XNOR U31287 ( .A(n29236), .B(n24754), .Z(n29237) );
  XOR U31288 ( .A(n29239), .B(n29240), .Z(n29236) );
  AND U31289 ( .A(n29241), .B(n29242), .Z(n29239) );
  XOR U31290 ( .A(n[376]), .B(n29240), .Z(n29242) );
  XNOR U31291 ( .A(n29240), .B(n24759), .Z(n29241) );
  XOR U31292 ( .A(n29243), .B(n29244), .Z(n29240) );
  AND U31293 ( .A(n29245), .B(n29246), .Z(n29243) );
  XOR U31294 ( .A(n[375]), .B(n29244), .Z(n29246) );
  XNOR U31295 ( .A(n29244), .B(n24764), .Z(n29245) );
  XOR U31296 ( .A(n29247), .B(n29248), .Z(n29244) );
  AND U31297 ( .A(n29249), .B(n29250), .Z(n29247) );
  XOR U31298 ( .A(n[374]), .B(n29248), .Z(n29250) );
  XNOR U31299 ( .A(n29248), .B(n24769), .Z(n29249) );
  XOR U31300 ( .A(n29251), .B(n29252), .Z(n29248) );
  AND U31301 ( .A(n29253), .B(n29254), .Z(n29251) );
  XOR U31302 ( .A(n[373]), .B(n29252), .Z(n29254) );
  XNOR U31303 ( .A(n29252), .B(n24774), .Z(n29253) );
  XOR U31304 ( .A(n29255), .B(n29256), .Z(n29252) );
  AND U31305 ( .A(n29257), .B(n29258), .Z(n29255) );
  XOR U31306 ( .A(n[372]), .B(n29256), .Z(n29258) );
  XNOR U31307 ( .A(n29256), .B(n24779), .Z(n29257) );
  XOR U31308 ( .A(n29259), .B(n29260), .Z(n29256) );
  AND U31309 ( .A(n29261), .B(n29262), .Z(n29259) );
  XOR U31310 ( .A(n[371]), .B(n29260), .Z(n29262) );
  XNOR U31311 ( .A(n29260), .B(n24784), .Z(n29261) );
  XOR U31312 ( .A(n29263), .B(n29264), .Z(n29260) );
  AND U31313 ( .A(n29265), .B(n29266), .Z(n29263) );
  XOR U31314 ( .A(n[370]), .B(n29264), .Z(n29266) );
  XNOR U31315 ( .A(n29264), .B(n24789), .Z(n29265) );
  XOR U31316 ( .A(n29267), .B(n29268), .Z(n29264) );
  AND U31317 ( .A(n29269), .B(n29270), .Z(n29267) );
  XOR U31318 ( .A(n[369]), .B(n29268), .Z(n29270) );
  XNOR U31319 ( .A(n29268), .B(n24794), .Z(n29269) );
  XOR U31320 ( .A(n29271), .B(n29272), .Z(n29268) );
  AND U31321 ( .A(n29273), .B(n29274), .Z(n29271) );
  XOR U31322 ( .A(n[368]), .B(n29272), .Z(n29274) );
  XNOR U31323 ( .A(n29272), .B(n24799), .Z(n29273) );
  XOR U31324 ( .A(n29275), .B(n29276), .Z(n29272) );
  AND U31325 ( .A(n29277), .B(n29278), .Z(n29275) );
  XOR U31326 ( .A(n[367]), .B(n29276), .Z(n29278) );
  XNOR U31327 ( .A(n29276), .B(n24804), .Z(n29277) );
  XOR U31328 ( .A(n29279), .B(n29280), .Z(n29276) );
  AND U31329 ( .A(n29281), .B(n29282), .Z(n29279) );
  XOR U31330 ( .A(n[366]), .B(n29280), .Z(n29282) );
  XNOR U31331 ( .A(n29280), .B(n24809), .Z(n29281) );
  XOR U31332 ( .A(n29283), .B(n29284), .Z(n29280) );
  AND U31333 ( .A(n29285), .B(n29286), .Z(n29283) );
  XOR U31334 ( .A(n[365]), .B(n29284), .Z(n29286) );
  XNOR U31335 ( .A(n29284), .B(n24814), .Z(n29285) );
  XOR U31336 ( .A(n29287), .B(n29288), .Z(n29284) );
  AND U31337 ( .A(n29289), .B(n29290), .Z(n29287) );
  XOR U31338 ( .A(n[364]), .B(n29288), .Z(n29290) );
  XNOR U31339 ( .A(n29288), .B(n24819), .Z(n29289) );
  XOR U31340 ( .A(n29291), .B(n29292), .Z(n29288) );
  AND U31341 ( .A(n29293), .B(n29294), .Z(n29291) );
  XOR U31342 ( .A(n[363]), .B(n29292), .Z(n29294) );
  XNOR U31343 ( .A(n29292), .B(n24824), .Z(n29293) );
  XOR U31344 ( .A(n29295), .B(n29296), .Z(n29292) );
  AND U31345 ( .A(n29297), .B(n29298), .Z(n29295) );
  XOR U31346 ( .A(n[362]), .B(n29296), .Z(n29298) );
  XNOR U31347 ( .A(n29296), .B(n24829), .Z(n29297) );
  XOR U31348 ( .A(n29299), .B(n29300), .Z(n29296) );
  AND U31349 ( .A(n29301), .B(n29302), .Z(n29299) );
  XOR U31350 ( .A(n[361]), .B(n29300), .Z(n29302) );
  XNOR U31351 ( .A(n29300), .B(n24834), .Z(n29301) );
  XOR U31352 ( .A(n29303), .B(n29304), .Z(n29300) );
  AND U31353 ( .A(n29305), .B(n29306), .Z(n29303) );
  XOR U31354 ( .A(n[360]), .B(n29304), .Z(n29306) );
  XNOR U31355 ( .A(n29304), .B(n24839), .Z(n29305) );
  XOR U31356 ( .A(n29307), .B(n29308), .Z(n29304) );
  AND U31357 ( .A(n29309), .B(n29310), .Z(n29307) );
  XOR U31358 ( .A(n[359]), .B(n29308), .Z(n29310) );
  XNOR U31359 ( .A(n29308), .B(n24844), .Z(n29309) );
  XOR U31360 ( .A(n29311), .B(n29312), .Z(n29308) );
  AND U31361 ( .A(n29313), .B(n29314), .Z(n29311) );
  XOR U31362 ( .A(n[358]), .B(n29312), .Z(n29314) );
  XNOR U31363 ( .A(n29312), .B(n24849), .Z(n29313) );
  XOR U31364 ( .A(n29315), .B(n29316), .Z(n29312) );
  AND U31365 ( .A(n29317), .B(n29318), .Z(n29315) );
  XOR U31366 ( .A(n[357]), .B(n29316), .Z(n29318) );
  XNOR U31367 ( .A(n29316), .B(n24854), .Z(n29317) );
  XOR U31368 ( .A(n29319), .B(n29320), .Z(n29316) );
  AND U31369 ( .A(n29321), .B(n29322), .Z(n29319) );
  XOR U31370 ( .A(n[356]), .B(n29320), .Z(n29322) );
  XNOR U31371 ( .A(n29320), .B(n24859), .Z(n29321) );
  XOR U31372 ( .A(n29323), .B(n29324), .Z(n29320) );
  AND U31373 ( .A(n29325), .B(n29326), .Z(n29323) );
  XOR U31374 ( .A(n[355]), .B(n29324), .Z(n29326) );
  XNOR U31375 ( .A(n29324), .B(n24864), .Z(n29325) );
  XOR U31376 ( .A(n29327), .B(n29328), .Z(n29324) );
  AND U31377 ( .A(n29329), .B(n29330), .Z(n29327) );
  XOR U31378 ( .A(n[354]), .B(n29328), .Z(n29330) );
  XNOR U31379 ( .A(n29328), .B(n24869), .Z(n29329) );
  XOR U31380 ( .A(n29331), .B(n29332), .Z(n29328) );
  AND U31381 ( .A(n29333), .B(n29334), .Z(n29331) );
  XOR U31382 ( .A(n[353]), .B(n29332), .Z(n29334) );
  XNOR U31383 ( .A(n29332), .B(n24874), .Z(n29333) );
  XOR U31384 ( .A(n29335), .B(n29336), .Z(n29332) );
  AND U31385 ( .A(n29337), .B(n29338), .Z(n29335) );
  XOR U31386 ( .A(n[352]), .B(n29336), .Z(n29338) );
  XNOR U31387 ( .A(n29336), .B(n24879), .Z(n29337) );
  XOR U31388 ( .A(n29339), .B(n29340), .Z(n29336) );
  AND U31389 ( .A(n29341), .B(n29342), .Z(n29339) );
  XOR U31390 ( .A(n[351]), .B(n29340), .Z(n29342) );
  XNOR U31391 ( .A(n29340), .B(n24884), .Z(n29341) );
  XOR U31392 ( .A(n29343), .B(n29344), .Z(n29340) );
  AND U31393 ( .A(n29345), .B(n29346), .Z(n29343) );
  XOR U31394 ( .A(n[350]), .B(n29344), .Z(n29346) );
  XNOR U31395 ( .A(n29344), .B(n24889), .Z(n29345) );
  XOR U31396 ( .A(n29347), .B(n29348), .Z(n29344) );
  AND U31397 ( .A(n29349), .B(n29350), .Z(n29347) );
  XOR U31398 ( .A(n[349]), .B(n29348), .Z(n29350) );
  XNOR U31399 ( .A(n29348), .B(n24894), .Z(n29349) );
  XOR U31400 ( .A(n29351), .B(n29352), .Z(n29348) );
  AND U31401 ( .A(n29353), .B(n29354), .Z(n29351) );
  XOR U31402 ( .A(n[348]), .B(n29352), .Z(n29354) );
  XNOR U31403 ( .A(n29352), .B(n24899), .Z(n29353) );
  XOR U31404 ( .A(n29355), .B(n29356), .Z(n29352) );
  AND U31405 ( .A(n29357), .B(n29358), .Z(n29355) );
  XOR U31406 ( .A(n[347]), .B(n29356), .Z(n29358) );
  XNOR U31407 ( .A(n29356), .B(n24904), .Z(n29357) );
  XOR U31408 ( .A(n29359), .B(n29360), .Z(n29356) );
  AND U31409 ( .A(n29361), .B(n29362), .Z(n29359) );
  XOR U31410 ( .A(n[346]), .B(n29360), .Z(n29362) );
  XNOR U31411 ( .A(n29360), .B(n24909), .Z(n29361) );
  XOR U31412 ( .A(n29363), .B(n29364), .Z(n29360) );
  AND U31413 ( .A(n29365), .B(n29366), .Z(n29363) );
  XOR U31414 ( .A(n[345]), .B(n29364), .Z(n29366) );
  XNOR U31415 ( .A(n29364), .B(n24914), .Z(n29365) );
  XOR U31416 ( .A(n29367), .B(n29368), .Z(n29364) );
  AND U31417 ( .A(n29369), .B(n29370), .Z(n29367) );
  XOR U31418 ( .A(n[344]), .B(n29368), .Z(n29370) );
  XNOR U31419 ( .A(n29368), .B(n24919), .Z(n29369) );
  XOR U31420 ( .A(n29371), .B(n29372), .Z(n29368) );
  AND U31421 ( .A(n29373), .B(n29374), .Z(n29371) );
  XOR U31422 ( .A(n[343]), .B(n29372), .Z(n29374) );
  XNOR U31423 ( .A(n29372), .B(n24924), .Z(n29373) );
  XOR U31424 ( .A(n29375), .B(n29376), .Z(n29372) );
  AND U31425 ( .A(n29377), .B(n29378), .Z(n29375) );
  XOR U31426 ( .A(n[342]), .B(n29376), .Z(n29378) );
  XNOR U31427 ( .A(n29376), .B(n24929), .Z(n29377) );
  XOR U31428 ( .A(n29379), .B(n29380), .Z(n29376) );
  AND U31429 ( .A(n29381), .B(n29382), .Z(n29379) );
  XOR U31430 ( .A(n[341]), .B(n29380), .Z(n29382) );
  XNOR U31431 ( .A(n29380), .B(n24934), .Z(n29381) );
  XOR U31432 ( .A(n29383), .B(n29384), .Z(n29380) );
  AND U31433 ( .A(n29385), .B(n29386), .Z(n29383) );
  XOR U31434 ( .A(n[340]), .B(n29384), .Z(n29386) );
  XNOR U31435 ( .A(n29384), .B(n24939), .Z(n29385) );
  XOR U31436 ( .A(n29387), .B(n29388), .Z(n29384) );
  AND U31437 ( .A(n29389), .B(n29390), .Z(n29387) );
  XOR U31438 ( .A(n[339]), .B(n29388), .Z(n29390) );
  XNOR U31439 ( .A(n29388), .B(n24944), .Z(n29389) );
  XOR U31440 ( .A(n29391), .B(n29392), .Z(n29388) );
  AND U31441 ( .A(n29393), .B(n29394), .Z(n29391) );
  XOR U31442 ( .A(n[338]), .B(n29392), .Z(n29394) );
  XNOR U31443 ( .A(n29392), .B(n24949), .Z(n29393) );
  XOR U31444 ( .A(n29395), .B(n29396), .Z(n29392) );
  AND U31445 ( .A(n29397), .B(n29398), .Z(n29395) );
  XOR U31446 ( .A(n[337]), .B(n29396), .Z(n29398) );
  XNOR U31447 ( .A(n29396), .B(n24954), .Z(n29397) );
  XOR U31448 ( .A(n29399), .B(n29400), .Z(n29396) );
  AND U31449 ( .A(n29401), .B(n29402), .Z(n29399) );
  XOR U31450 ( .A(n[336]), .B(n29400), .Z(n29402) );
  XNOR U31451 ( .A(n29400), .B(n24959), .Z(n29401) );
  XOR U31452 ( .A(n29403), .B(n29404), .Z(n29400) );
  AND U31453 ( .A(n29405), .B(n29406), .Z(n29403) );
  XOR U31454 ( .A(n[335]), .B(n29404), .Z(n29406) );
  XNOR U31455 ( .A(n29404), .B(n24964), .Z(n29405) );
  XOR U31456 ( .A(n29407), .B(n29408), .Z(n29404) );
  AND U31457 ( .A(n29409), .B(n29410), .Z(n29407) );
  XOR U31458 ( .A(n[334]), .B(n29408), .Z(n29410) );
  XNOR U31459 ( .A(n29408), .B(n24969), .Z(n29409) );
  XOR U31460 ( .A(n29411), .B(n29412), .Z(n29408) );
  AND U31461 ( .A(n29413), .B(n29414), .Z(n29411) );
  XOR U31462 ( .A(n[333]), .B(n29412), .Z(n29414) );
  XNOR U31463 ( .A(n29412), .B(n24974), .Z(n29413) );
  XOR U31464 ( .A(n29415), .B(n29416), .Z(n29412) );
  AND U31465 ( .A(n29417), .B(n29418), .Z(n29415) );
  XOR U31466 ( .A(n[332]), .B(n29416), .Z(n29418) );
  XNOR U31467 ( .A(n29416), .B(n24979), .Z(n29417) );
  XOR U31468 ( .A(n29419), .B(n29420), .Z(n29416) );
  AND U31469 ( .A(n29421), .B(n29422), .Z(n29419) );
  XOR U31470 ( .A(n[331]), .B(n29420), .Z(n29422) );
  XNOR U31471 ( .A(n29420), .B(n24984), .Z(n29421) );
  XOR U31472 ( .A(n29423), .B(n29424), .Z(n29420) );
  AND U31473 ( .A(n29425), .B(n29426), .Z(n29423) );
  XOR U31474 ( .A(n[330]), .B(n29424), .Z(n29426) );
  XNOR U31475 ( .A(n29424), .B(n24989), .Z(n29425) );
  XOR U31476 ( .A(n29427), .B(n29428), .Z(n29424) );
  AND U31477 ( .A(n29429), .B(n29430), .Z(n29427) );
  XOR U31478 ( .A(n[329]), .B(n29428), .Z(n29430) );
  XNOR U31479 ( .A(n29428), .B(n24994), .Z(n29429) );
  XOR U31480 ( .A(n29431), .B(n29432), .Z(n29428) );
  AND U31481 ( .A(n29433), .B(n29434), .Z(n29431) );
  XOR U31482 ( .A(n[328]), .B(n29432), .Z(n29434) );
  XNOR U31483 ( .A(n29432), .B(n24999), .Z(n29433) );
  XOR U31484 ( .A(n29435), .B(n29436), .Z(n29432) );
  AND U31485 ( .A(n29437), .B(n29438), .Z(n29435) );
  XOR U31486 ( .A(n[327]), .B(n29436), .Z(n29438) );
  XNOR U31487 ( .A(n29436), .B(n25004), .Z(n29437) );
  XOR U31488 ( .A(n29439), .B(n29440), .Z(n29436) );
  AND U31489 ( .A(n29441), .B(n29442), .Z(n29439) );
  XOR U31490 ( .A(n[326]), .B(n29440), .Z(n29442) );
  XNOR U31491 ( .A(n29440), .B(n25009), .Z(n29441) );
  XOR U31492 ( .A(n29443), .B(n29444), .Z(n29440) );
  AND U31493 ( .A(n29445), .B(n29446), .Z(n29443) );
  XOR U31494 ( .A(n[325]), .B(n29444), .Z(n29446) );
  XNOR U31495 ( .A(n29444), .B(n25014), .Z(n29445) );
  XOR U31496 ( .A(n29447), .B(n29448), .Z(n29444) );
  AND U31497 ( .A(n29449), .B(n29450), .Z(n29447) );
  XOR U31498 ( .A(n[324]), .B(n29448), .Z(n29450) );
  XNOR U31499 ( .A(n29448), .B(n25019), .Z(n29449) );
  XOR U31500 ( .A(n29451), .B(n29452), .Z(n29448) );
  AND U31501 ( .A(n29453), .B(n29454), .Z(n29451) );
  XOR U31502 ( .A(n[323]), .B(n29452), .Z(n29454) );
  XNOR U31503 ( .A(n29452), .B(n25024), .Z(n29453) );
  XOR U31504 ( .A(n29455), .B(n29456), .Z(n29452) );
  AND U31505 ( .A(n29457), .B(n29458), .Z(n29455) );
  XOR U31506 ( .A(n[322]), .B(n29456), .Z(n29458) );
  XNOR U31507 ( .A(n29456), .B(n25029), .Z(n29457) );
  XOR U31508 ( .A(n29459), .B(n29460), .Z(n29456) );
  AND U31509 ( .A(n29461), .B(n29462), .Z(n29459) );
  XOR U31510 ( .A(n[321]), .B(n29460), .Z(n29462) );
  XNOR U31511 ( .A(n29460), .B(n25034), .Z(n29461) );
  XOR U31512 ( .A(n29463), .B(n29464), .Z(n29460) );
  AND U31513 ( .A(n29465), .B(n29466), .Z(n29463) );
  XOR U31514 ( .A(n[320]), .B(n29464), .Z(n29466) );
  XNOR U31515 ( .A(n29464), .B(n25039), .Z(n29465) );
  XOR U31516 ( .A(n29467), .B(n29468), .Z(n29464) );
  AND U31517 ( .A(n29469), .B(n29470), .Z(n29467) );
  XOR U31518 ( .A(n[319]), .B(n29468), .Z(n29470) );
  XNOR U31519 ( .A(n29468), .B(n25044), .Z(n29469) );
  XOR U31520 ( .A(n29471), .B(n29472), .Z(n29468) );
  AND U31521 ( .A(n29473), .B(n29474), .Z(n29471) );
  XOR U31522 ( .A(n[318]), .B(n29472), .Z(n29474) );
  XNOR U31523 ( .A(n29472), .B(n25049), .Z(n29473) );
  XOR U31524 ( .A(n29475), .B(n29476), .Z(n29472) );
  AND U31525 ( .A(n29477), .B(n29478), .Z(n29475) );
  XOR U31526 ( .A(n[317]), .B(n29476), .Z(n29478) );
  XNOR U31527 ( .A(n29476), .B(n25054), .Z(n29477) );
  XOR U31528 ( .A(n29479), .B(n29480), .Z(n29476) );
  AND U31529 ( .A(n29481), .B(n29482), .Z(n29479) );
  XOR U31530 ( .A(n[316]), .B(n29480), .Z(n29482) );
  XNOR U31531 ( .A(n29480), .B(n25059), .Z(n29481) );
  XOR U31532 ( .A(n29483), .B(n29484), .Z(n29480) );
  AND U31533 ( .A(n29485), .B(n29486), .Z(n29483) );
  XOR U31534 ( .A(n[315]), .B(n29484), .Z(n29486) );
  XNOR U31535 ( .A(n29484), .B(n25064), .Z(n29485) );
  XOR U31536 ( .A(n29487), .B(n29488), .Z(n29484) );
  AND U31537 ( .A(n29489), .B(n29490), .Z(n29487) );
  XOR U31538 ( .A(n[314]), .B(n29488), .Z(n29490) );
  XNOR U31539 ( .A(n29488), .B(n25069), .Z(n29489) );
  XOR U31540 ( .A(n29491), .B(n29492), .Z(n29488) );
  AND U31541 ( .A(n29493), .B(n29494), .Z(n29491) );
  XOR U31542 ( .A(n[313]), .B(n29492), .Z(n29494) );
  XNOR U31543 ( .A(n29492), .B(n25074), .Z(n29493) );
  XOR U31544 ( .A(n29495), .B(n29496), .Z(n29492) );
  AND U31545 ( .A(n29497), .B(n29498), .Z(n29495) );
  XOR U31546 ( .A(n[312]), .B(n29496), .Z(n29498) );
  XNOR U31547 ( .A(n29496), .B(n25079), .Z(n29497) );
  XOR U31548 ( .A(n29499), .B(n29500), .Z(n29496) );
  AND U31549 ( .A(n29501), .B(n29502), .Z(n29499) );
  XOR U31550 ( .A(n[311]), .B(n29500), .Z(n29502) );
  XNOR U31551 ( .A(n29500), .B(n25084), .Z(n29501) );
  XOR U31552 ( .A(n29503), .B(n29504), .Z(n29500) );
  AND U31553 ( .A(n29505), .B(n29506), .Z(n29503) );
  XOR U31554 ( .A(n[310]), .B(n29504), .Z(n29506) );
  XNOR U31555 ( .A(n29504), .B(n25089), .Z(n29505) );
  XOR U31556 ( .A(n29507), .B(n29508), .Z(n29504) );
  AND U31557 ( .A(n29509), .B(n29510), .Z(n29507) );
  XOR U31558 ( .A(n[309]), .B(n29508), .Z(n29510) );
  XNOR U31559 ( .A(n29508), .B(n25094), .Z(n29509) );
  XOR U31560 ( .A(n29511), .B(n29512), .Z(n29508) );
  AND U31561 ( .A(n29513), .B(n29514), .Z(n29511) );
  XOR U31562 ( .A(n[308]), .B(n29512), .Z(n29514) );
  XNOR U31563 ( .A(n29512), .B(n25099), .Z(n29513) );
  XOR U31564 ( .A(n29515), .B(n29516), .Z(n29512) );
  AND U31565 ( .A(n29517), .B(n29518), .Z(n29515) );
  XOR U31566 ( .A(n[307]), .B(n29516), .Z(n29518) );
  XNOR U31567 ( .A(n29516), .B(n25104), .Z(n29517) );
  XOR U31568 ( .A(n29519), .B(n29520), .Z(n29516) );
  AND U31569 ( .A(n29521), .B(n29522), .Z(n29519) );
  XOR U31570 ( .A(n[306]), .B(n29520), .Z(n29522) );
  XNOR U31571 ( .A(n29520), .B(n25109), .Z(n29521) );
  XOR U31572 ( .A(n29523), .B(n29524), .Z(n29520) );
  AND U31573 ( .A(n29525), .B(n29526), .Z(n29523) );
  XOR U31574 ( .A(n[305]), .B(n29524), .Z(n29526) );
  XNOR U31575 ( .A(n29524), .B(n25114), .Z(n29525) );
  XOR U31576 ( .A(n29527), .B(n29528), .Z(n29524) );
  AND U31577 ( .A(n29529), .B(n29530), .Z(n29527) );
  XOR U31578 ( .A(n[304]), .B(n29528), .Z(n29530) );
  XNOR U31579 ( .A(n29528), .B(n25119), .Z(n29529) );
  XOR U31580 ( .A(n29531), .B(n29532), .Z(n29528) );
  AND U31581 ( .A(n29533), .B(n29534), .Z(n29531) );
  XOR U31582 ( .A(n[303]), .B(n29532), .Z(n29534) );
  XNOR U31583 ( .A(n29532), .B(n25124), .Z(n29533) );
  XOR U31584 ( .A(n29535), .B(n29536), .Z(n29532) );
  AND U31585 ( .A(n29537), .B(n29538), .Z(n29535) );
  XOR U31586 ( .A(n[302]), .B(n29536), .Z(n29538) );
  XNOR U31587 ( .A(n29536), .B(n25129), .Z(n29537) );
  XOR U31588 ( .A(n29539), .B(n29540), .Z(n29536) );
  AND U31589 ( .A(n29541), .B(n29542), .Z(n29539) );
  XOR U31590 ( .A(n[301]), .B(n29540), .Z(n29542) );
  XNOR U31591 ( .A(n29540), .B(n25134), .Z(n29541) );
  XOR U31592 ( .A(n29543), .B(n29544), .Z(n29540) );
  AND U31593 ( .A(n29545), .B(n29546), .Z(n29543) );
  XOR U31594 ( .A(n[300]), .B(n29544), .Z(n29546) );
  XNOR U31595 ( .A(n29544), .B(n25139), .Z(n29545) );
  XOR U31596 ( .A(n29547), .B(n29548), .Z(n29544) );
  AND U31597 ( .A(n29549), .B(n29550), .Z(n29547) );
  XOR U31598 ( .A(n[299]), .B(n29548), .Z(n29550) );
  XNOR U31599 ( .A(n29548), .B(n25144), .Z(n29549) );
  XOR U31600 ( .A(n29551), .B(n29552), .Z(n29548) );
  AND U31601 ( .A(n29553), .B(n29554), .Z(n29551) );
  XOR U31602 ( .A(n[298]), .B(n29552), .Z(n29554) );
  XNOR U31603 ( .A(n29552), .B(n25149), .Z(n29553) );
  XOR U31604 ( .A(n29555), .B(n29556), .Z(n29552) );
  AND U31605 ( .A(n29557), .B(n29558), .Z(n29555) );
  XOR U31606 ( .A(n[297]), .B(n29556), .Z(n29558) );
  XNOR U31607 ( .A(n29556), .B(n25154), .Z(n29557) );
  XOR U31608 ( .A(n29559), .B(n29560), .Z(n29556) );
  AND U31609 ( .A(n29561), .B(n29562), .Z(n29559) );
  XOR U31610 ( .A(n[296]), .B(n29560), .Z(n29562) );
  XNOR U31611 ( .A(n29560), .B(n25159), .Z(n29561) );
  XOR U31612 ( .A(n29563), .B(n29564), .Z(n29560) );
  AND U31613 ( .A(n29565), .B(n29566), .Z(n29563) );
  XOR U31614 ( .A(n[295]), .B(n29564), .Z(n29566) );
  XNOR U31615 ( .A(n29564), .B(n25164), .Z(n29565) );
  XOR U31616 ( .A(n29567), .B(n29568), .Z(n29564) );
  AND U31617 ( .A(n29569), .B(n29570), .Z(n29567) );
  XOR U31618 ( .A(n[294]), .B(n29568), .Z(n29570) );
  XNOR U31619 ( .A(n29568), .B(n25169), .Z(n29569) );
  XOR U31620 ( .A(n29571), .B(n29572), .Z(n29568) );
  AND U31621 ( .A(n29573), .B(n29574), .Z(n29571) );
  XOR U31622 ( .A(n[293]), .B(n29572), .Z(n29574) );
  XNOR U31623 ( .A(n29572), .B(n25174), .Z(n29573) );
  XOR U31624 ( .A(n29575), .B(n29576), .Z(n29572) );
  AND U31625 ( .A(n29577), .B(n29578), .Z(n29575) );
  XOR U31626 ( .A(n[292]), .B(n29576), .Z(n29578) );
  XNOR U31627 ( .A(n29576), .B(n25179), .Z(n29577) );
  XOR U31628 ( .A(n29579), .B(n29580), .Z(n29576) );
  AND U31629 ( .A(n29581), .B(n29582), .Z(n29579) );
  XOR U31630 ( .A(n[291]), .B(n29580), .Z(n29582) );
  XNOR U31631 ( .A(n29580), .B(n25184), .Z(n29581) );
  XOR U31632 ( .A(n29583), .B(n29584), .Z(n29580) );
  AND U31633 ( .A(n29585), .B(n29586), .Z(n29583) );
  XOR U31634 ( .A(n[290]), .B(n29584), .Z(n29586) );
  XNOR U31635 ( .A(n29584), .B(n25189), .Z(n29585) );
  XOR U31636 ( .A(n29587), .B(n29588), .Z(n29584) );
  AND U31637 ( .A(n29589), .B(n29590), .Z(n29587) );
  XOR U31638 ( .A(n[289]), .B(n29588), .Z(n29590) );
  XNOR U31639 ( .A(n29588), .B(n25194), .Z(n29589) );
  XOR U31640 ( .A(n29591), .B(n29592), .Z(n29588) );
  AND U31641 ( .A(n29593), .B(n29594), .Z(n29591) );
  XOR U31642 ( .A(n[288]), .B(n29592), .Z(n29594) );
  XNOR U31643 ( .A(n29592), .B(n25199), .Z(n29593) );
  XOR U31644 ( .A(n29595), .B(n29596), .Z(n29592) );
  AND U31645 ( .A(n29597), .B(n29598), .Z(n29595) );
  XOR U31646 ( .A(n[287]), .B(n29596), .Z(n29598) );
  XNOR U31647 ( .A(n29596), .B(n25204), .Z(n29597) );
  XOR U31648 ( .A(n29599), .B(n29600), .Z(n29596) );
  AND U31649 ( .A(n29601), .B(n29602), .Z(n29599) );
  XOR U31650 ( .A(n[286]), .B(n29600), .Z(n29602) );
  XNOR U31651 ( .A(n29600), .B(n25209), .Z(n29601) );
  XOR U31652 ( .A(n29603), .B(n29604), .Z(n29600) );
  AND U31653 ( .A(n29605), .B(n29606), .Z(n29603) );
  XOR U31654 ( .A(n[285]), .B(n29604), .Z(n29606) );
  XNOR U31655 ( .A(n29604), .B(n25214), .Z(n29605) );
  XOR U31656 ( .A(n29607), .B(n29608), .Z(n29604) );
  AND U31657 ( .A(n29609), .B(n29610), .Z(n29607) );
  XOR U31658 ( .A(n[284]), .B(n29608), .Z(n29610) );
  XNOR U31659 ( .A(n29608), .B(n25219), .Z(n29609) );
  XOR U31660 ( .A(n29611), .B(n29612), .Z(n29608) );
  AND U31661 ( .A(n29613), .B(n29614), .Z(n29611) );
  XOR U31662 ( .A(n[283]), .B(n29612), .Z(n29614) );
  XNOR U31663 ( .A(n29612), .B(n25224), .Z(n29613) );
  XOR U31664 ( .A(n29615), .B(n29616), .Z(n29612) );
  AND U31665 ( .A(n29617), .B(n29618), .Z(n29615) );
  XOR U31666 ( .A(n[282]), .B(n29616), .Z(n29618) );
  XNOR U31667 ( .A(n29616), .B(n25229), .Z(n29617) );
  XOR U31668 ( .A(n29619), .B(n29620), .Z(n29616) );
  AND U31669 ( .A(n29621), .B(n29622), .Z(n29619) );
  XOR U31670 ( .A(n[281]), .B(n29620), .Z(n29622) );
  XNOR U31671 ( .A(n29620), .B(n25234), .Z(n29621) );
  XOR U31672 ( .A(n29623), .B(n29624), .Z(n29620) );
  AND U31673 ( .A(n29625), .B(n29626), .Z(n29623) );
  XOR U31674 ( .A(n[280]), .B(n29624), .Z(n29626) );
  XNOR U31675 ( .A(n29624), .B(n25239), .Z(n29625) );
  XOR U31676 ( .A(n29627), .B(n29628), .Z(n29624) );
  AND U31677 ( .A(n29629), .B(n29630), .Z(n29627) );
  XOR U31678 ( .A(n[279]), .B(n29628), .Z(n29630) );
  XNOR U31679 ( .A(n29628), .B(n25244), .Z(n29629) );
  XOR U31680 ( .A(n29631), .B(n29632), .Z(n29628) );
  AND U31681 ( .A(n29633), .B(n29634), .Z(n29631) );
  XOR U31682 ( .A(n[278]), .B(n29632), .Z(n29634) );
  XNOR U31683 ( .A(n29632), .B(n25249), .Z(n29633) );
  XOR U31684 ( .A(n29635), .B(n29636), .Z(n29632) );
  AND U31685 ( .A(n29637), .B(n29638), .Z(n29635) );
  XOR U31686 ( .A(n[277]), .B(n29636), .Z(n29638) );
  XNOR U31687 ( .A(n29636), .B(n25254), .Z(n29637) );
  XOR U31688 ( .A(n29639), .B(n29640), .Z(n29636) );
  AND U31689 ( .A(n29641), .B(n29642), .Z(n29639) );
  XOR U31690 ( .A(n[276]), .B(n29640), .Z(n29642) );
  XNOR U31691 ( .A(n29640), .B(n25259), .Z(n29641) );
  XOR U31692 ( .A(n29643), .B(n29644), .Z(n29640) );
  AND U31693 ( .A(n29645), .B(n29646), .Z(n29643) );
  XOR U31694 ( .A(n[275]), .B(n29644), .Z(n29646) );
  XNOR U31695 ( .A(n29644), .B(n25264), .Z(n29645) );
  XOR U31696 ( .A(n29647), .B(n29648), .Z(n29644) );
  AND U31697 ( .A(n29649), .B(n29650), .Z(n29647) );
  XOR U31698 ( .A(n[274]), .B(n29648), .Z(n29650) );
  XNOR U31699 ( .A(n29648), .B(n25269), .Z(n29649) );
  XOR U31700 ( .A(n29651), .B(n29652), .Z(n29648) );
  AND U31701 ( .A(n29653), .B(n29654), .Z(n29651) );
  XOR U31702 ( .A(n[273]), .B(n29652), .Z(n29654) );
  XNOR U31703 ( .A(n29652), .B(n25274), .Z(n29653) );
  XOR U31704 ( .A(n29655), .B(n29656), .Z(n29652) );
  AND U31705 ( .A(n29657), .B(n29658), .Z(n29655) );
  XOR U31706 ( .A(n[272]), .B(n29656), .Z(n29658) );
  XNOR U31707 ( .A(n29656), .B(n25279), .Z(n29657) );
  XOR U31708 ( .A(n29659), .B(n29660), .Z(n29656) );
  AND U31709 ( .A(n29661), .B(n29662), .Z(n29659) );
  XOR U31710 ( .A(n[271]), .B(n29660), .Z(n29662) );
  XNOR U31711 ( .A(n29660), .B(n25284), .Z(n29661) );
  XOR U31712 ( .A(n29663), .B(n29664), .Z(n29660) );
  AND U31713 ( .A(n29665), .B(n29666), .Z(n29663) );
  XOR U31714 ( .A(n[270]), .B(n29664), .Z(n29666) );
  XNOR U31715 ( .A(n29664), .B(n25289), .Z(n29665) );
  XOR U31716 ( .A(n29667), .B(n29668), .Z(n29664) );
  AND U31717 ( .A(n29669), .B(n29670), .Z(n29667) );
  XOR U31718 ( .A(n[269]), .B(n29668), .Z(n29670) );
  XNOR U31719 ( .A(n29668), .B(n25294), .Z(n29669) );
  XOR U31720 ( .A(n29671), .B(n29672), .Z(n29668) );
  AND U31721 ( .A(n29673), .B(n29674), .Z(n29671) );
  XOR U31722 ( .A(n[268]), .B(n29672), .Z(n29674) );
  XNOR U31723 ( .A(n29672), .B(n25299), .Z(n29673) );
  XOR U31724 ( .A(n29675), .B(n29676), .Z(n29672) );
  AND U31725 ( .A(n29677), .B(n29678), .Z(n29675) );
  XOR U31726 ( .A(n[267]), .B(n29676), .Z(n29678) );
  XNOR U31727 ( .A(n29676), .B(n25304), .Z(n29677) );
  XOR U31728 ( .A(n29679), .B(n29680), .Z(n29676) );
  AND U31729 ( .A(n29681), .B(n29682), .Z(n29679) );
  XOR U31730 ( .A(n[266]), .B(n29680), .Z(n29682) );
  XNOR U31731 ( .A(n29680), .B(n25309), .Z(n29681) );
  XOR U31732 ( .A(n29683), .B(n29684), .Z(n29680) );
  AND U31733 ( .A(n29685), .B(n29686), .Z(n29683) );
  XOR U31734 ( .A(n[265]), .B(n29684), .Z(n29686) );
  XNOR U31735 ( .A(n29684), .B(n25314), .Z(n29685) );
  XOR U31736 ( .A(n29687), .B(n29688), .Z(n29684) );
  AND U31737 ( .A(n29689), .B(n29690), .Z(n29687) );
  XOR U31738 ( .A(n[264]), .B(n29688), .Z(n29690) );
  XNOR U31739 ( .A(n29688), .B(n25319), .Z(n29689) );
  XOR U31740 ( .A(n29691), .B(n29692), .Z(n29688) );
  AND U31741 ( .A(n29693), .B(n29694), .Z(n29691) );
  XOR U31742 ( .A(n[263]), .B(n29692), .Z(n29694) );
  XNOR U31743 ( .A(n29692), .B(n25324), .Z(n29693) );
  XOR U31744 ( .A(n29695), .B(n29696), .Z(n29692) );
  AND U31745 ( .A(n29697), .B(n29698), .Z(n29695) );
  XOR U31746 ( .A(n[262]), .B(n29696), .Z(n29698) );
  XNOR U31747 ( .A(n29696), .B(n25329), .Z(n29697) );
  XOR U31748 ( .A(n29699), .B(n29700), .Z(n29696) );
  AND U31749 ( .A(n29701), .B(n29702), .Z(n29699) );
  XOR U31750 ( .A(n[261]), .B(n29700), .Z(n29702) );
  XNOR U31751 ( .A(n29700), .B(n25334), .Z(n29701) );
  XOR U31752 ( .A(n29703), .B(n29704), .Z(n29700) );
  AND U31753 ( .A(n29705), .B(n29706), .Z(n29703) );
  XOR U31754 ( .A(n[260]), .B(n29704), .Z(n29706) );
  XNOR U31755 ( .A(n29704), .B(n25339), .Z(n29705) );
  XOR U31756 ( .A(n29707), .B(n29708), .Z(n29704) );
  AND U31757 ( .A(n29709), .B(n29710), .Z(n29707) );
  XOR U31758 ( .A(n[259]), .B(n29708), .Z(n29710) );
  XNOR U31759 ( .A(n29708), .B(n25344), .Z(n29709) );
  XOR U31760 ( .A(n29711), .B(n29712), .Z(n29708) );
  AND U31761 ( .A(n29713), .B(n29714), .Z(n29711) );
  XOR U31762 ( .A(n[258]), .B(n29712), .Z(n29714) );
  XNOR U31763 ( .A(n29712), .B(n25349), .Z(n29713) );
  XOR U31764 ( .A(n29715), .B(n29716), .Z(n29712) );
  AND U31765 ( .A(n29717), .B(n29718), .Z(n29715) );
  XOR U31766 ( .A(n[257]), .B(n29716), .Z(n29718) );
  XNOR U31767 ( .A(n29716), .B(n25354), .Z(n29717) );
  XOR U31768 ( .A(n29719), .B(n29720), .Z(n29716) );
  AND U31769 ( .A(n29721), .B(n29722), .Z(n29719) );
  XOR U31770 ( .A(n[256]), .B(n29720), .Z(n29722) );
  XNOR U31771 ( .A(n29720), .B(n25359), .Z(n29721) );
  XOR U31772 ( .A(n29723), .B(n29724), .Z(n29720) );
  AND U31773 ( .A(n29725), .B(n29726), .Z(n29723) );
  XOR U31774 ( .A(n[255]), .B(n29724), .Z(n29726) );
  XNOR U31775 ( .A(n29724), .B(n25364), .Z(n29725) );
  XOR U31776 ( .A(n29727), .B(n29728), .Z(n29724) );
  AND U31777 ( .A(n29729), .B(n29730), .Z(n29727) );
  XOR U31778 ( .A(n[254]), .B(n29728), .Z(n29730) );
  XNOR U31779 ( .A(n29728), .B(n25369), .Z(n29729) );
  XOR U31780 ( .A(n29731), .B(n29732), .Z(n29728) );
  AND U31781 ( .A(n29733), .B(n29734), .Z(n29731) );
  XOR U31782 ( .A(n[253]), .B(n29732), .Z(n29734) );
  XNOR U31783 ( .A(n29732), .B(n25374), .Z(n29733) );
  XOR U31784 ( .A(n29735), .B(n29736), .Z(n29732) );
  AND U31785 ( .A(n29737), .B(n29738), .Z(n29735) );
  XOR U31786 ( .A(n[252]), .B(n29736), .Z(n29738) );
  XNOR U31787 ( .A(n29736), .B(n25379), .Z(n29737) );
  XOR U31788 ( .A(n29739), .B(n29740), .Z(n29736) );
  AND U31789 ( .A(n29741), .B(n29742), .Z(n29739) );
  XOR U31790 ( .A(n[251]), .B(n29740), .Z(n29742) );
  XNOR U31791 ( .A(n29740), .B(n25384), .Z(n29741) );
  XOR U31792 ( .A(n29743), .B(n29744), .Z(n29740) );
  AND U31793 ( .A(n29745), .B(n29746), .Z(n29743) );
  XOR U31794 ( .A(n[250]), .B(n29744), .Z(n29746) );
  XNOR U31795 ( .A(n29744), .B(n25389), .Z(n29745) );
  XOR U31796 ( .A(n29747), .B(n29748), .Z(n29744) );
  AND U31797 ( .A(n29749), .B(n29750), .Z(n29747) );
  XOR U31798 ( .A(n[249]), .B(n29748), .Z(n29750) );
  XNOR U31799 ( .A(n29748), .B(n25394), .Z(n29749) );
  XOR U31800 ( .A(n29751), .B(n29752), .Z(n29748) );
  AND U31801 ( .A(n29753), .B(n29754), .Z(n29751) );
  XOR U31802 ( .A(n[248]), .B(n29752), .Z(n29754) );
  XNOR U31803 ( .A(n29752), .B(n25399), .Z(n29753) );
  XOR U31804 ( .A(n29755), .B(n29756), .Z(n29752) );
  AND U31805 ( .A(n29757), .B(n29758), .Z(n29755) );
  XOR U31806 ( .A(n[247]), .B(n29756), .Z(n29758) );
  XNOR U31807 ( .A(n29756), .B(n25404), .Z(n29757) );
  XOR U31808 ( .A(n29759), .B(n29760), .Z(n29756) );
  AND U31809 ( .A(n29761), .B(n29762), .Z(n29759) );
  XOR U31810 ( .A(n[246]), .B(n29760), .Z(n29762) );
  XNOR U31811 ( .A(n29760), .B(n25409), .Z(n29761) );
  XOR U31812 ( .A(n29763), .B(n29764), .Z(n29760) );
  AND U31813 ( .A(n29765), .B(n29766), .Z(n29763) );
  XOR U31814 ( .A(n[245]), .B(n29764), .Z(n29766) );
  XNOR U31815 ( .A(n29764), .B(n25414), .Z(n29765) );
  XOR U31816 ( .A(n29767), .B(n29768), .Z(n29764) );
  AND U31817 ( .A(n29769), .B(n29770), .Z(n29767) );
  XOR U31818 ( .A(n[244]), .B(n29768), .Z(n29770) );
  XNOR U31819 ( .A(n29768), .B(n25419), .Z(n29769) );
  XOR U31820 ( .A(n29771), .B(n29772), .Z(n29768) );
  AND U31821 ( .A(n29773), .B(n29774), .Z(n29771) );
  XOR U31822 ( .A(n[243]), .B(n29772), .Z(n29774) );
  XNOR U31823 ( .A(n29772), .B(n25424), .Z(n29773) );
  XOR U31824 ( .A(n29775), .B(n29776), .Z(n29772) );
  AND U31825 ( .A(n29777), .B(n29778), .Z(n29775) );
  XOR U31826 ( .A(n[242]), .B(n29776), .Z(n29778) );
  XNOR U31827 ( .A(n29776), .B(n25429), .Z(n29777) );
  XOR U31828 ( .A(n29779), .B(n29780), .Z(n29776) );
  AND U31829 ( .A(n29781), .B(n29782), .Z(n29779) );
  XOR U31830 ( .A(n[241]), .B(n29780), .Z(n29782) );
  XNOR U31831 ( .A(n29780), .B(n25434), .Z(n29781) );
  XOR U31832 ( .A(n29783), .B(n29784), .Z(n29780) );
  AND U31833 ( .A(n29785), .B(n29786), .Z(n29783) );
  XOR U31834 ( .A(n[240]), .B(n29784), .Z(n29786) );
  XNOR U31835 ( .A(n29784), .B(n25439), .Z(n29785) );
  XOR U31836 ( .A(n29787), .B(n29788), .Z(n29784) );
  AND U31837 ( .A(n29789), .B(n29790), .Z(n29787) );
  XOR U31838 ( .A(n[239]), .B(n29788), .Z(n29790) );
  XNOR U31839 ( .A(n29788), .B(n25444), .Z(n29789) );
  XOR U31840 ( .A(n29791), .B(n29792), .Z(n29788) );
  AND U31841 ( .A(n29793), .B(n29794), .Z(n29791) );
  XOR U31842 ( .A(n[238]), .B(n29792), .Z(n29794) );
  XNOR U31843 ( .A(n29792), .B(n25449), .Z(n29793) );
  XOR U31844 ( .A(n29795), .B(n29796), .Z(n29792) );
  AND U31845 ( .A(n29797), .B(n29798), .Z(n29795) );
  XOR U31846 ( .A(n[237]), .B(n29796), .Z(n29798) );
  XNOR U31847 ( .A(n29796), .B(n25454), .Z(n29797) );
  XOR U31848 ( .A(n29799), .B(n29800), .Z(n29796) );
  AND U31849 ( .A(n29801), .B(n29802), .Z(n29799) );
  XOR U31850 ( .A(n[236]), .B(n29800), .Z(n29802) );
  XNOR U31851 ( .A(n29800), .B(n25459), .Z(n29801) );
  XOR U31852 ( .A(n29803), .B(n29804), .Z(n29800) );
  AND U31853 ( .A(n29805), .B(n29806), .Z(n29803) );
  XOR U31854 ( .A(n[235]), .B(n29804), .Z(n29806) );
  XNOR U31855 ( .A(n29804), .B(n25464), .Z(n29805) );
  XOR U31856 ( .A(n29807), .B(n29808), .Z(n29804) );
  AND U31857 ( .A(n29809), .B(n29810), .Z(n29807) );
  XOR U31858 ( .A(n[234]), .B(n29808), .Z(n29810) );
  XNOR U31859 ( .A(n29808), .B(n25469), .Z(n29809) );
  XOR U31860 ( .A(n29811), .B(n29812), .Z(n29808) );
  AND U31861 ( .A(n29813), .B(n29814), .Z(n29811) );
  XOR U31862 ( .A(n[233]), .B(n29812), .Z(n29814) );
  XNOR U31863 ( .A(n29812), .B(n25474), .Z(n29813) );
  XOR U31864 ( .A(n29815), .B(n29816), .Z(n29812) );
  AND U31865 ( .A(n29817), .B(n29818), .Z(n29815) );
  XOR U31866 ( .A(n[232]), .B(n29816), .Z(n29818) );
  XNOR U31867 ( .A(n29816), .B(n25479), .Z(n29817) );
  XOR U31868 ( .A(n29819), .B(n29820), .Z(n29816) );
  AND U31869 ( .A(n29821), .B(n29822), .Z(n29819) );
  XOR U31870 ( .A(n[231]), .B(n29820), .Z(n29822) );
  XNOR U31871 ( .A(n29820), .B(n25484), .Z(n29821) );
  XOR U31872 ( .A(n29823), .B(n29824), .Z(n29820) );
  AND U31873 ( .A(n29825), .B(n29826), .Z(n29823) );
  XOR U31874 ( .A(n[230]), .B(n29824), .Z(n29826) );
  XNOR U31875 ( .A(n29824), .B(n25489), .Z(n29825) );
  XOR U31876 ( .A(n29827), .B(n29828), .Z(n29824) );
  AND U31877 ( .A(n29829), .B(n29830), .Z(n29827) );
  XOR U31878 ( .A(n[229]), .B(n29828), .Z(n29830) );
  XNOR U31879 ( .A(n29828), .B(n25494), .Z(n29829) );
  XOR U31880 ( .A(n29831), .B(n29832), .Z(n29828) );
  AND U31881 ( .A(n29833), .B(n29834), .Z(n29831) );
  XOR U31882 ( .A(n[228]), .B(n29832), .Z(n29834) );
  XNOR U31883 ( .A(n29832), .B(n25499), .Z(n29833) );
  XOR U31884 ( .A(n29835), .B(n29836), .Z(n29832) );
  AND U31885 ( .A(n29837), .B(n29838), .Z(n29835) );
  XOR U31886 ( .A(n[227]), .B(n29836), .Z(n29838) );
  XNOR U31887 ( .A(n29836), .B(n25504), .Z(n29837) );
  XOR U31888 ( .A(n29839), .B(n29840), .Z(n29836) );
  AND U31889 ( .A(n29841), .B(n29842), .Z(n29839) );
  XOR U31890 ( .A(n[226]), .B(n29840), .Z(n29842) );
  XNOR U31891 ( .A(n29840), .B(n25509), .Z(n29841) );
  XOR U31892 ( .A(n29843), .B(n29844), .Z(n29840) );
  AND U31893 ( .A(n29845), .B(n29846), .Z(n29843) );
  XOR U31894 ( .A(n[225]), .B(n29844), .Z(n29846) );
  XNOR U31895 ( .A(n29844), .B(n25514), .Z(n29845) );
  XOR U31896 ( .A(n29847), .B(n29848), .Z(n29844) );
  AND U31897 ( .A(n29849), .B(n29850), .Z(n29847) );
  XOR U31898 ( .A(n[224]), .B(n29848), .Z(n29850) );
  XNOR U31899 ( .A(n29848), .B(n25519), .Z(n29849) );
  XOR U31900 ( .A(n29851), .B(n29852), .Z(n29848) );
  AND U31901 ( .A(n29853), .B(n29854), .Z(n29851) );
  XOR U31902 ( .A(n[223]), .B(n29852), .Z(n29854) );
  XNOR U31903 ( .A(n29852), .B(n25524), .Z(n29853) );
  XOR U31904 ( .A(n29855), .B(n29856), .Z(n29852) );
  AND U31905 ( .A(n29857), .B(n29858), .Z(n29855) );
  XOR U31906 ( .A(n[222]), .B(n29856), .Z(n29858) );
  XNOR U31907 ( .A(n29856), .B(n25529), .Z(n29857) );
  XOR U31908 ( .A(n29859), .B(n29860), .Z(n29856) );
  AND U31909 ( .A(n29861), .B(n29862), .Z(n29859) );
  XOR U31910 ( .A(n[221]), .B(n29860), .Z(n29862) );
  XNOR U31911 ( .A(n29860), .B(n25534), .Z(n29861) );
  XOR U31912 ( .A(n29863), .B(n29864), .Z(n29860) );
  AND U31913 ( .A(n29865), .B(n29866), .Z(n29863) );
  XOR U31914 ( .A(n[220]), .B(n29864), .Z(n29866) );
  XNOR U31915 ( .A(n29864), .B(n25539), .Z(n29865) );
  XOR U31916 ( .A(n29867), .B(n29868), .Z(n29864) );
  AND U31917 ( .A(n29869), .B(n29870), .Z(n29867) );
  XOR U31918 ( .A(n[219]), .B(n29868), .Z(n29870) );
  XNOR U31919 ( .A(n29868), .B(n25544), .Z(n29869) );
  XOR U31920 ( .A(n29871), .B(n29872), .Z(n29868) );
  AND U31921 ( .A(n29873), .B(n29874), .Z(n29871) );
  XOR U31922 ( .A(n[218]), .B(n29872), .Z(n29874) );
  XNOR U31923 ( .A(n29872), .B(n25549), .Z(n29873) );
  XOR U31924 ( .A(n29875), .B(n29876), .Z(n29872) );
  AND U31925 ( .A(n29877), .B(n29878), .Z(n29875) );
  XOR U31926 ( .A(n[217]), .B(n29876), .Z(n29878) );
  XNOR U31927 ( .A(n29876), .B(n25554), .Z(n29877) );
  XOR U31928 ( .A(n29879), .B(n29880), .Z(n29876) );
  AND U31929 ( .A(n29881), .B(n29882), .Z(n29879) );
  XOR U31930 ( .A(n[216]), .B(n29880), .Z(n29882) );
  XNOR U31931 ( .A(n29880), .B(n25559), .Z(n29881) );
  XOR U31932 ( .A(n29883), .B(n29884), .Z(n29880) );
  AND U31933 ( .A(n29885), .B(n29886), .Z(n29883) );
  XOR U31934 ( .A(n[215]), .B(n29884), .Z(n29886) );
  XNOR U31935 ( .A(n29884), .B(n25564), .Z(n29885) );
  XOR U31936 ( .A(n29887), .B(n29888), .Z(n29884) );
  AND U31937 ( .A(n29889), .B(n29890), .Z(n29887) );
  XOR U31938 ( .A(n[214]), .B(n29888), .Z(n29890) );
  XNOR U31939 ( .A(n29888), .B(n25569), .Z(n29889) );
  XOR U31940 ( .A(n29891), .B(n29892), .Z(n29888) );
  AND U31941 ( .A(n29893), .B(n29894), .Z(n29891) );
  XOR U31942 ( .A(n[213]), .B(n29892), .Z(n29894) );
  XNOR U31943 ( .A(n29892), .B(n25574), .Z(n29893) );
  XOR U31944 ( .A(n29895), .B(n29896), .Z(n29892) );
  AND U31945 ( .A(n29897), .B(n29898), .Z(n29895) );
  XOR U31946 ( .A(n[212]), .B(n29896), .Z(n29898) );
  XNOR U31947 ( .A(n29896), .B(n25579), .Z(n29897) );
  XOR U31948 ( .A(n29899), .B(n29900), .Z(n29896) );
  AND U31949 ( .A(n29901), .B(n29902), .Z(n29899) );
  XOR U31950 ( .A(n[211]), .B(n29900), .Z(n29902) );
  XNOR U31951 ( .A(n29900), .B(n25584), .Z(n29901) );
  XOR U31952 ( .A(n29903), .B(n29904), .Z(n29900) );
  AND U31953 ( .A(n29905), .B(n29906), .Z(n29903) );
  XOR U31954 ( .A(n[210]), .B(n29904), .Z(n29906) );
  XNOR U31955 ( .A(n29904), .B(n25589), .Z(n29905) );
  XOR U31956 ( .A(n29907), .B(n29908), .Z(n29904) );
  AND U31957 ( .A(n29909), .B(n29910), .Z(n29907) );
  XOR U31958 ( .A(n[209]), .B(n29908), .Z(n29910) );
  XNOR U31959 ( .A(n29908), .B(n25594), .Z(n29909) );
  XOR U31960 ( .A(n29911), .B(n29912), .Z(n29908) );
  AND U31961 ( .A(n29913), .B(n29914), .Z(n29911) );
  XOR U31962 ( .A(n[208]), .B(n29912), .Z(n29914) );
  XNOR U31963 ( .A(n29912), .B(n25599), .Z(n29913) );
  XOR U31964 ( .A(n29915), .B(n29916), .Z(n29912) );
  AND U31965 ( .A(n29917), .B(n29918), .Z(n29915) );
  XOR U31966 ( .A(n[207]), .B(n29916), .Z(n29918) );
  XNOR U31967 ( .A(n29916), .B(n25604), .Z(n29917) );
  XOR U31968 ( .A(n29919), .B(n29920), .Z(n29916) );
  AND U31969 ( .A(n29921), .B(n29922), .Z(n29919) );
  XOR U31970 ( .A(n[206]), .B(n29920), .Z(n29922) );
  XNOR U31971 ( .A(n29920), .B(n25609), .Z(n29921) );
  XOR U31972 ( .A(n29923), .B(n29924), .Z(n29920) );
  AND U31973 ( .A(n29925), .B(n29926), .Z(n29923) );
  XOR U31974 ( .A(n[205]), .B(n29924), .Z(n29926) );
  XNOR U31975 ( .A(n29924), .B(n25614), .Z(n29925) );
  XOR U31976 ( .A(n29927), .B(n29928), .Z(n29924) );
  AND U31977 ( .A(n29929), .B(n29930), .Z(n29927) );
  XOR U31978 ( .A(n[204]), .B(n29928), .Z(n29930) );
  XNOR U31979 ( .A(n29928), .B(n25619), .Z(n29929) );
  XOR U31980 ( .A(n29931), .B(n29932), .Z(n29928) );
  AND U31981 ( .A(n29933), .B(n29934), .Z(n29931) );
  XOR U31982 ( .A(n[203]), .B(n29932), .Z(n29934) );
  XNOR U31983 ( .A(n29932), .B(n25624), .Z(n29933) );
  XOR U31984 ( .A(n29935), .B(n29936), .Z(n29932) );
  AND U31985 ( .A(n29937), .B(n29938), .Z(n29935) );
  XOR U31986 ( .A(n[202]), .B(n29936), .Z(n29938) );
  XNOR U31987 ( .A(n29936), .B(n25629), .Z(n29937) );
  XOR U31988 ( .A(n29939), .B(n29940), .Z(n29936) );
  AND U31989 ( .A(n29941), .B(n29942), .Z(n29939) );
  XOR U31990 ( .A(n[201]), .B(n29940), .Z(n29942) );
  XNOR U31991 ( .A(n29940), .B(n25634), .Z(n29941) );
  XOR U31992 ( .A(n29943), .B(n29944), .Z(n29940) );
  AND U31993 ( .A(n29945), .B(n29946), .Z(n29943) );
  XOR U31994 ( .A(n[200]), .B(n29944), .Z(n29946) );
  XNOR U31995 ( .A(n29944), .B(n25639), .Z(n29945) );
  XOR U31996 ( .A(n29947), .B(n29948), .Z(n29944) );
  AND U31997 ( .A(n29949), .B(n29950), .Z(n29947) );
  XOR U31998 ( .A(n[199]), .B(n29948), .Z(n29950) );
  XNOR U31999 ( .A(n29948), .B(n25644), .Z(n29949) );
  XOR U32000 ( .A(n29951), .B(n29952), .Z(n29948) );
  AND U32001 ( .A(n29953), .B(n29954), .Z(n29951) );
  XOR U32002 ( .A(n[198]), .B(n29952), .Z(n29954) );
  XNOR U32003 ( .A(n29952), .B(n25649), .Z(n29953) );
  XOR U32004 ( .A(n29955), .B(n29956), .Z(n29952) );
  AND U32005 ( .A(n29957), .B(n29958), .Z(n29955) );
  XOR U32006 ( .A(n[197]), .B(n29956), .Z(n29958) );
  XNOR U32007 ( .A(n29956), .B(n25654), .Z(n29957) );
  XOR U32008 ( .A(n29959), .B(n29960), .Z(n29956) );
  AND U32009 ( .A(n29961), .B(n29962), .Z(n29959) );
  XOR U32010 ( .A(n[196]), .B(n29960), .Z(n29962) );
  XNOR U32011 ( .A(n29960), .B(n25659), .Z(n29961) );
  XOR U32012 ( .A(n29963), .B(n29964), .Z(n29960) );
  AND U32013 ( .A(n29965), .B(n29966), .Z(n29963) );
  XOR U32014 ( .A(n[195]), .B(n29964), .Z(n29966) );
  XNOR U32015 ( .A(n29964), .B(n25664), .Z(n29965) );
  XOR U32016 ( .A(n29967), .B(n29968), .Z(n29964) );
  AND U32017 ( .A(n29969), .B(n29970), .Z(n29967) );
  XOR U32018 ( .A(n[194]), .B(n29968), .Z(n29970) );
  XNOR U32019 ( .A(n29968), .B(n25669), .Z(n29969) );
  XOR U32020 ( .A(n29971), .B(n29972), .Z(n29968) );
  AND U32021 ( .A(n29973), .B(n29974), .Z(n29971) );
  XOR U32022 ( .A(n[193]), .B(n29972), .Z(n29974) );
  XNOR U32023 ( .A(n29972), .B(n25674), .Z(n29973) );
  XOR U32024 ( .A(n29975), .B(n29976), .Z(n29972) );
  AND U32025 ( .A(n29977), .B(n29978), .Z(n29975) );
  XOR U32026 ( .A(n[192]), .B(n29976), .Z(n29978) );
  XNOR U32027 ( .A(n29976), .B(n25679), .Z(n29977) );
  XOR U32028 ( .A(n29979), .B(n29980), .Z(n29976) );
  AND U32029 ( .A(n29981), .B(n29982), .Z(n29979) );
  XOR U32030 ( .A(n[191]), .B(n29980), .Z(n29982) );
  XNOR U32031 ( .A(n29980), .B(n25684), .Z(n29981) );
  XOR U32032 ( .A(n29983), .B(n29984), .Z(n29980) );
  AND U32033 ( .A(n29985), .B(n29986), .Z(n29983) );
  XOR U32034 ( .A(n[190]), .B(n29984), .Z(n29986) );
  XNOR U32035 ( .A(n29984), .B(n25689), .Z(n29985) );
  XOR U32036 ( .A(n29987), .B(n29988), .Z(n29984) );
  AND U32037 ( .A(n29989), .B(n29990), .Z(n29987) );
  XOR U32038 ( .A(n[189]), .B(n29988), .Z(n29990) );
  XNOR U32039 ( .A(n29988), .B(n25694), .Z(n29989) );
  XOR U32040 ( .A(n29991), .B(n29992), .Z(n29988) );
  AND U32041 ( .A(n29993), .B(n29994), .Z(n29991) );
  XOR U32042 ( .A(n[188]), .B(n29992), .Z(n29994) );
  XNOR U32043 ( .A(n29992), .B(n25699), .Z(n29993) );
  XOR U32044 ( .A(n29995), .B(n29996), .Z(n29992) );
  AND U32045 ( .A(n29997), .B(n29998), .Z(n29995) );
  XOR U32046 ( .A(n[187]), .B(n29996), .Z(n29998) );
  XNOR U32047 ( .A(n29996), .B(n25704), .Z(n29997) );
  XOR U32048 ( .A(n29999), .B(n30000), .Z(n29996) );
  AND U32049 ( .A(n30001), .B(n30002), .Z(n29999) );
  XOR U32050 ( .A(n[186]), .B(n30000), .Z(n30002) );
  XNOR U32051 ( .A(n30000), .B(n25709), .Z(n30001) );
  XOR U32052 ( .A(n30003), .B(n30004), .Z(n30000) );
  AND U32053 ( .A(n30005), .B(n30006), .Z(n30003) );
  XOR U32054 ( .A(n[185]), .B(n30004), .Z(n30006) );
  XNOR U32055 ( .A(n30004), .B(n25714), .Z(n30005) );
  XOR U32056 ( .A(n30007), .B(n30008), .Z(n30004) );
  AND U32057 ( .A(n30009), .B(n30010), .Z(n30007) );
  XOR U32058 ( .A(n[184]), .B(n30008), .Z(n30010) );
  XNOR U32059 ( .A(n30008), .B(n25719), .Z(n30009) );
  XOR U32060 ( .A(n30011), .B(n30012), .Z(n30008) );
  AND U32061 ( .A(n30013), .B(n30014), .Z(n30011) );
  XOR U32062 ( .A(n[183]), .B(n30012), .Z(n30014) );
  XNOR U32063 ( .A(n30012), .B(n25724), .Z(n30013) );
  XOR U32064 ( .A(n30015), .B(n30016), .Z(n30012) );
  AND U32065 ( .A(n30017), .B(n30018), .Z(n30015) );
  XOR U32066 ( .A(n[182]), .B(n30016), .Z(n30018) );
  XNOR U32067 ( .A(n30016), .B(n25729), .Z(n30017) );
  XOR U32068 ( .A(n30019), .B(n30020), .Z(n30016) );
  AND U32069 ( .A(n30021), .B(n30022), .Z(n30019) );
  XOR U32070 ( .A(n[181]), .B(n30020), .Z(n30022) );
  XNOR U32071 ( .A(n30020), .B(n25734), .Z(n30021) );
  XOR U32072 ( .A(n30023), .B(n30024), .Z(n30020) );
  AND U32073 ( .A(n30025), .B(n30026), .Z(n30023) );
  XOR U32074 ( .A(n[180]), .B(n30024), .Z(n30026) );
  XNOR U32075 ( .A(n30024), .B(n25739), .Z(n30025) );
  XOR U32076 ( .A(n30027), .B(n30028), .Z(n30024) );
  AND U32077 ( .A(n30029), .B(n30030), .Z(n30027) );
  XOR U32078 ( .A(n[179]), .B(n30028), .Z(n30030) );
  XNOR U32079 ( .A(n30028), .B(n25744), .Z(n30029) );
  XOR U32080 ( .A(n30031), .B(n30032), .Z(n30028) );
  AND U32081 ( .A(n30033), .B(n30034), .Z(n30031) );
  XOR U32082 ( .A(n[178]), .B(n30032), .Z(n30034) );
  XNOR U32083 ( .A(n30032), .B(n25749), .Z(n30033) );
  XOR U32084 ( .A(n30035), .B(n30036), .Z(n30032) );
  AND U32085 ( .A(n30037), .B(n30038), .Z(n30035) );
  XOR U32086 ( .A(n[177]), .B(n30036), .Z(n30038) );
  XNOR U32087 ( .A(n30036), .B(n25754), .Z(n30037) );
  XOR U32088 ( .A(n30039), .B(n30040), .Z(n30036) );
  AND U32089 ( .A(n30041), .B(n30042), .Z(n30039) );
  XOR U32090 ( .A(n[176]), .B(n30040), .Z(n30042) );
  XNOR U32091 ( .A(n30040), .B(n25759), .Z(n30041) );
  XOR U32092 ( .A(n30043), .B(n30044), .Z(n30040) );
  AND U32093 ( .A(n30045), .B(n30046), .Z(n30043) );
  XOR U32094 ( .A(n[175]), .B(n30044), .Z(n30046) );
  XNOR U32095 ( .A(n30044), .B(n25764), .Z(n30045) );
  XOR U32096 ( .A(n30047), .B(n30048), .Z(n30044) );
  AND U32097 ( .A(n30049), .B(n30050), .Z(n30047) );
  XOR U32098 ( .A(n[174]), .B(n30048), .Z(n30050) );
  XNOR U32099 ( .A(n30048), .B(n25769), .Z(n30049) );
  XOR U32100 ( .A(n30051), .B(n30052), .Z(n30048) );
  AND U32101 ( .A(n30053), .B(n30054), .Z(n30051) );
  XOR U32102 ( .A(n[173]), .B(n30052), .Z(n30054) );
  XNOR U32103 ( .A(n30052), .B(n25774), .Z(n30053) );
  XOR U32104 ( .A(n30055), .B(n30056), .Z(n30052) );
  AND U32105 ( .A(n30057), .B(n30058), .Z(n30055) );
  XOR U32106 ( .A(n[172]), .B(n30056), .Z(n30058) );
  XNOR U32107 ( .A(n30056), .B(n25779), .Z(n30057) );
  XOR U32108 ( .A(n30059), .B(n30060), .Z(n30056) );
  AND U32109 ( .A(n30061), .B(n30062), .Z(n30059) );
  XOR U32110 ( .A(n[171]), .B(n30060), .Z(n30062) );
  XNOR U32111 ( .A(n30060), .B(n25784), .Z(n30061) );
  XOR U32112 ( .A(n30063), .B(n30064), .Z(n30060) );
  AND U32113 ( .A(n30065), .B(n30066), .Z(n30063) );
  XOR U32114 ( .A(n[170]), .B(n30064), .Z(n30066) );
  XNOR U32115 ( .A(n30064), .B(n25789), .Z(n30065) );
  XOR U32116 ( .A(n30067), .B(n30068), .Z(n30064) );
  AND U32117 ( .A(n30069), .B(n30070), .Z(n30067) );
  XOR U32118 ( .A(n[169]), .B(n30068), .Z(n30070) );
  XNOR U32119 ( .A(n30068), .B(n25794), .Z(n30069) );
  XOR U32120 ( .A(n30071), .B(n30072), .Z(n30068) );
  AND U32121 ( .A(n30073), .B(n30074), .Z(n30071) );
  XOR U32122 ( .A(n[168]), .B(n30072), .Z(n30074) );
  XNOR U32123 ( .A(n30072), .B(n25799), .Z(n30073) );
  XOR U32124 ( .A(n30075), .B(n30076), .Z(n30072) );
  AND U32125 ( .A(n30077), .B(n30078), .Z(n30075) );
  XOR U32126 ( .A(n[167]), .B(n30076), .Z(n30078) );
  XNOR U32127 ( .A(n30076), .B(n25804), .Z(n30077) );
  XOR U32128 ( .A(n30079), .B(n30080), .Z(n30076) );
  AND U32129 ( .A(n30081), .B(n30082), .Z(n30079) );
  XOR U32130 ( .A(n[166]), .B(n30080), .Z(n30082) );
  XNOR U32131 ( .A(n30080), .B(n25809), .Z(n30081) );
  XOR U32132 ( .A(n30083), .B(n30084), .Z(n30080) );
  AND U32133 ( .A(n30085), .B(n30086), .Z(n30083) );
  XOR U32134 ( .A(n[165]), .B(n30084), .Z(n30086) );
  XNOR U32135 ( .A(n30084), .B(n25814), .Z(n30085) );
  XOR U32136 ( .A(n30087), .B(n30088), .Z(n30084) );
  AND U32137 ( .A(n30089), .B(n30090), .Z(n30087) );
  XOR U32138 ( .A(n[164]), .B(n30088), .Z(n30090) );
  XNOR U32139 ( .A(n30088), .B(n25819), .Z(n30089) );
  XOR U32140 ( .A(n30091), .B(n30092), .Z(n30088) );
  AND U32141 ( .A(n30093), .B(n30094), .Z(n30091) );
  XOR U32142 ( .A(n[163]), .B(n30092), .Z(n30094) );
  XNOR U32143 ( .A(n30092), .B(n25824), .Z(n30093) );
  XOR U32144 ( .A(n30095), .B(n30096), .Z(n30092) );
  AND U32145 ( .A(n30097), .B(n30098), .Z(n30095) );
  XOR U32146 ( .A(n[162]), .B(n30096), .Z(n30098) );
  XNOR U32147 ( .A(n30096), .B(n25829), .Z(n30097) );
  XOR U32148 ( .A(n30099), .B(n30100), .Z(n30096) );
  AND U32149 ( .A(n30101), .B(n30102), .Z(n30099) );
  XOR U32150 ( .A(n[161]), .B(n30100), .Z(n30102) );
  XNOR U32151 ( .A(n30100), .B(n25834), .Z(n30101) );
  XOR U32152 ( .A(n30103), .B(n30104), .Z(n30100) );
  AND U32153 ( .A(n30105), .B(n30106), .Z(n30103) );
  XOR U32154 ( .A(n[160]), .B(n30104), .Z(n30106) );
  XNOR U32155 ( .A(n30104), .B(n25839), .Z(n30105) );
  XOR U32156 ( .A(n30107), .B(n30108), .Z(n30104) );
  AND U32157 ( .A(n30109), .B(n30110), .Z(n30107) );
  XOR U32158 ( .A(n[159]), .B(n30108), .Z(n30110) );
  XNOR U32159 ( .A(n30108), .B(n25844), .Z(n30109) );
  XOR U32160 ( .A(n30111), .B(n30112), .Z(n30108) );
  AND U32161 ( .A(n30113), .B(n30114), .Z(n30111) );
  XOR U32162 ( .A(n[158]), .B(n30112), .Z(n30114) );
  XNOR U32163 ( .A(n30112), .B(n25849), .Z(n30113) );
  XOR U32164 ( .A(n30115), .B(n30116), .Z(n30112) );
  AND U32165 ( .A(n30117), .B(n30118), .Z(n30115) );
  XOR U32166 ( .A(n[157]), .B(n30116), .Z(n30118) );
  XNOR U32167 ( .A(n30116), .B(n25854), .Z(n30117) );
  XOR U32168 ( .A(n30119), .B(n30120), .Z(n30116) );
  AND U32169 ( .A(n30121), .B(n30122), .Z(n30119) );
  XOR U32170 ( .A(n[156]), .B(n30120), .Z(n30122) );
  XNOR U32171 ( .A(n30120), .B(n25859), .Z(n30121) );
  XOR U32172 ( .A(n30123), .B(n30124), .Z(n30120) );
  AND U32173 ( .A(n30125), .B(n30126), .Z(n30123) );
  XOR U32174 ( .A(n[155]), .B(n30124), .Z(n30126) );
  XNOR U32175 ( .A(n30124), .B(n25864), .Z(n30125) );
  XOR U32176 ( .A(n30127), .B(n30128), .Z(n30124) );
  AND U32177 ( .A(n30129), .B(n30130), .Z(n30127) );
  XOR U32178 ( .A(n[154]), .B(n30128), .Z(n30130) );
  XNOR U32179 ( .A(n30128), .B(n25869), .Z(n30129) );
  XOR U32180 ( .A(n30131), .B(n30132), .Z(n30128) );
  AND U32181 ( .A(n30133), .B(n30134), .Z(n30131) );
  XOR U32182 ( .A(n[153]), .B(n30132), .Z(n30134) );
  XNOR U32183 ( .A(n30132), .B(n25874), .Z(n30133) );
  XOR U32184 ( .A(n30135), .B(n30136), .Z(n30132) );
  AND U32185 ( .A(n30137), .B(n30138), .Z(n30135) );
  XOR U32186 ( .A(n[152]), .B(n30136), .Z(n30138) );
  XNOR U32187 ( .A(n30136), .B(n25879), .Z(n30137) );
  XOR U32188 ( .A(n30139), .B(n30140), .Z(n30136) );
  AND U32189 ( .A(n30141), .B(n30142), .Z(n30139) );
  XOR U32190 ( .A(n[151]), .B(n30140), .Z(n30142) );
  XNOR U32191 ( .A(n30140), .B(n25884), .Z(n30141) );
  XOR U32192 ( .A(n30143), .B(n30144), .Z(n30140) );
  AND U32193 ( .A(n30145), .B(n30146), .Z(n30143) );
  XOR U32194 ( .A(n[150]), .B(n30144), .Z(n30146) );
  XNOR U32195 ( .A(n30144), .B(n25889), .Z(n30145) );
  XOR U32196 ( .A(n30147), .B(n30148), .Z(n30144) );
  AND U32197 ( .A(n30149), .B(n30150), .Z(n30147) );
  XOR U32198 ( .A(n[149]), .B(n30148), .Z(n30150) );
  XNOR U32199 ( .A(n30148), .B(n25894), .Z(n30149) );
  XOR U32200 ( .A(n30151), .B(n30152), .Z(n30148) );
  AND U32201 ( .A(n30153), .B(n30154), .Z(n30151) );
  XOR U32202 ( .A(n[148]), .B(n30152), .Z(n30154) );
  XNOR U32203 ( .A(n30152), .B(n25899), .Z(n30153) );
  XOR U32204 ( .A(n30155), .B(n30156), .Z(n30152) );
  AND U32205 ( .A(n30157), .B(n30158), .Z(n30155) );
  XOR U32206 ( .A(n[147]), .B(n30156), .Z(n30158) );
  XNOR U32207 ( .A(n30156), .B(n25904), .Z(n30157) );
  XOR U32208 ( .A(n30159), .B(n30160), .Z(n30156) );
  AND U32209 ( .A(n30161), .B(n30162), .Z(n30159) );
  XOR U32210 ( .A(n[146]), .B(n30160), .Z(n30162) );
  XNOR U32211 ( .A(n30160), .B(n25909), .Z(n30161) );
  XOR U32212 ( .A(n30163), .B(n30164), .Z(n30160) );
  AND U32213 ( .A(n30165), .B(n30166), .Z(n30163) );
  XOR U32214 ( .A(n[145]), .B(n30164), .Z(n30166) );
  XNOR U32215 ( .A(n30164), .B(n25914), .Z(n30165) );
  XOR U32216 ( .A(n30167), .B(n30168), .Z(n30164) );
  AND U32217 ( .A(n30169), .B(n30170), .Z(n30167) );
  XOR U32218 ( .A(n[144]), .B(n30168), .Z(n30170) );
  XNOR U32219 ( .A(n30168), .B(n25919), .Z(n30169) );
  XOR U32220 ( .A(n30171), .B(n30172), .Z(n30168) );
  AND U32221 ( .A(n30173), .B(n30174), .Z(n30171) );
  XOR U32222 ( .A(n[143]), .B(n30172), .Z(n30174) );
  XNOR U32223 ( .A(n30172), .B(n25924), .Z(n30173) );
  XOR U32224 ( .A(n30175), .B(n30176), .Z(n30172) );
  AND U32225 ( .A(n30177), .B(n30178), .Z(n30175) );
  XOR U32226 ( .A(n[142]), .B(n30176), .Z(n30178) );
  XNOR U32227 ( .A(n30176), .B(n25929), .Z(n30177) );
  XOR U32228 ( .A(n30179), .B(n30180), .Z(n30176) );
  AND U32229 ( .A(n30181), .B(n30182), .Z(n30179) );
  XOR U32230 ( .A(n[141]), .B(n30180), .Z(n30182) );
  XNOR U32231 ( .A(n30180), .B(n25934), .Z(n30181) );
  XOR U32232 ( .A(n30183), .B(n30184), .Z(n30180) );
  AND U32233 ( .A(n30185), .B(n30186), .Z(n30183) );
  XOR U32234 ( .A(n[140]), .B(n30184), .Z(n30186) );
  XNOR U32235 ( .A(n30184), .B(n25939), .Z(n30185) );
  XOR U32236 ( .A(n30187), .B(n30188), .Z(n30184) );
  AND U32237 ( .A(n30189), .B(n30190), .Z(n30187) );
  XOR U32238 ( .A(n[139]), .B(n30188), .Z(n30190) );
  XNOR U32239 ( .A(n30188), .B(n25944), .Z(n30189) );
  XOR U32240 ( .A(n30191), .B(n30192), .Z(n30188) );
  AND U32241 ( .A(n30193), .B(n30194), .Z(n30191) );
  XOR U32242 ( .A(n[138]), .B(n30192), .Z(n30194) );
  XNOR U32243 ( .A(n30192), .B(n25949), .Z(n30193) );
  XOR U32244 ( .A(n30195), .B(n30196), .Z(n30192) );
  AND U32245 ( .A(n30197), .B(n30198), .Z(n30195) );
  XOR U32246 ( .A(n[137]), .B(n30196), .Z(n30198) );
  XNOR U32247 ( .A(n30196), .B(n25954), .Z(n30197) );
  XOR U32248 ( .A(n30199), .B(n30200), .Z(n30196) );
  AND U32249 ( .A(n30201), .B(n30202), .Z(n30199) );
  XOR U32250 ( .A(n[136]), .B(n30200), .Z(n30202) );
  XNOR U32251 ( .A(n30200), .B(n25959), .Z(n30201) );
  XOR U32252 ( .A(n30203), .B(n30204), .Z(n30200) );
  AND U32253 ( .A(n30205), .B(n30206), .Z(n30203) );
  XOR U32254 ( .A(n[135]), .B(n30204), .Z(n30206) );
  XNOR U32255 ( .A(n30204), .B(n25964), .Z(n30205) );
  XOR U32256 ( .A(n30207), .B(n30208), .Z(n30204) );
  AND U32257 ( .A(n30209), .B(n30210), .Z(n30207) );
  XOR U32258 ( .A(n[134]), .B(n30208), .Z(n30210) );
  XNOR U32259 ( .A(n30208), .B(n25969), .Z(n30209) );
  XOR U32260 ( .A(n30211), .B(n30212), .Z(n30208) );
  AND U32261 ( .A(n30213), .B(n30214), .Z(n30211) );
  XOR U32262 ( .A(n[133]), .B(n30212), .Z(n30214) );
  XNOR U32263 ( .A(n30212), .B(n25974), .Z(n30213) );
  XOR U32264 ( .A(n30215), .B(n30216), .Z(n30212) );
  AND U32265 ( .A(n30217), .B(n30218), .Z(n30215) );
  XOR U32266 ( .A(n[132]), .B(n30216), .Z(n30218) );
  XNOR U32267 ( .A(n30216), .B(n25979), .Z(n30217) );
  XOR U32268 ( .A(n30219), .B(n30220), .Z(n30216) );
  AND U32269 ( .A(n30221), .B(n30222), .Z(n30219) );
  XOR U32270 ( .A(n[131]), .B(n30220), .Z(n30222) );
  XNOR U32271 ( .A(n30220), .B(n25984), .Z(n30221) );
  XOR U32272 ( .A(n30223), .B(n30224), .Z(n30220) );
  AND U32273 ( .A(n30225), .B(n30226), .Z(n30223) );
  XOR U32274 ( .A(n[130]), .B(n30224), .Z(n30226) );
  XNOR U32275 ( .A(n30224), .B(n25989), .Z(n30225) );
  XOR U32276 ( .A(n30227), .B(n30228), .Z(n30224) );
  AND U32277 ( .A(n30229), .B(n30230), .Z(n30227) );
  XOR U32278 ( .A(n[129]), .B(n30228), .Z(n30230) );
  XNOR U32279 ( .A(n30228), .B(n25994), .Z(n30229) );
  XOR U32280 ( .A(n30231), .B(n30232), .Z(n30228) );
  AND U32281 ( .A(n30233), .B(n30234), .Z(n30231) );
  XOR U32282 ( .A(n[128]), .B(n30232), .Z(n30234) );
  XNOR U32283 ( .A(n30232), .B(n25999), .Z(n30233) );
  XOR U32284 ( .A(n30235), .B(n30236), .Z(n30232) );
  AND U32285 ( .A(n30237), .B(n30238), .Z(n30235) );
  XOR U32286 ( .A(n[127]), .B(n30236), .Z(n30238) );
  XNOR U32287 ( .A(n30236), .B(n26004), .Z(n30237) );
  XOR U32288 ( .A(n30239), .B(n30240), .Z(n30236) );
  AND U32289 ( .A(n30241), .B(n30242), .Z(n30239) );
  XOR U32290 ( .A(n[126]), .B(n30240), .Z(n30242) );
  XNOR U32291 ( .A(n30240), .B(n26009), .Z(n30241) );
  XOR U32292 ( .A(n30243), .B(n30244), .Z(n30240) );
  AND U32293 ( .A(n30245), .B(n30246), .Z(n30243) );
  XOR U32294 ( .A(n[125]), .B(n30244), .Z(n30246) );
  XNOR U32295 ( .A(n30244), .B(n26014), .Z(n30245) );
  XOR U32296 ( .A(n30247), .B(n30248), .Z(n30244) );
  AND U32297 ( .A(n30249), .B(n30250), .Z(n30247) );
  XOR U32298 ( .A(n[124]), .B(n30248), .Z(n30250) );
  XNOR U32299 ( .A(n30248), .B(n26019), .Z(n30249) );
  XOR U32300 ( .A(n30251), .B(n30252), .Z(n30248) );
  AND U32301 ( .A(n30253), .B(n30254), .Z(n30251) );
  XOR U32302 ( .A(n[123]), .B(n30252), .Z(n30254) );
  XNOR U32303 ( .A(n30252), .B(n26024), .Z(n30253) );
  XOR U32304 ( .A(n30255), .B(n30256), .Z(n30252) );
  AND U32305 ( .A(n30257), .B(n30258), .Z(n30255) );
  XOR U32306 ( .A(n[122]), .B(n30256), .Z(n30258) );
  XNOR U32307 ( .A(n30256), .B(n26029), .Z(n30257) );
  XOR U32308 ( .A(n30259), .B(n30260), .Z(n30256) );
  AND U32309 ( .A(n30261), .B(n30262), .Z(n30259) );
  XOR U32310 ( .A(n[121]), .B(n30260), .Z(n30262) );
  XNOR U32311 ( .A(n30260), .B(n26034), .Z(n30261) );
  XOR U32312 ( .A(n30263), .B(n30264), .Z(n30260) );
  AND U32313 ( .A(n30265), .B(n30266), .Z(n30263) );
  XOR U32314 ( .A(n[120]), .B(n30264), .Z(n30266) );
  XNOR U32315 ( .A(n30264), .B(n26039), .Z(n30265) );
  XOR U32316 ( .A(n30267), .B(n30268), .Z(n30264) );
  AND U32317 ( .A(n30269), .B(n30270), .Z(n30267) );
  XOR U32318 ( .A(n[119]), .B(n30268), .Z(n30270) );
  XNOR U32319 ( .A(n30268), .B(n26044), .Z(n30269) );
  XOR U32320 ( .A(n30271), .B(n30272), .Z(n30268) );
  AND U32321 ( .A(n30273), .B(n30274), .Z(n30271) );
  XOR U32322 ( .A(n[118]), .B(n30272), .Z(n30274) );
  XNOR U32323 ( .A(n30272), .B(n26049), .Z(n30273) );
  XOR U32324 ( .A(n30275), .B(n30276), .Z(n30272) );
  AND U32325 ( .A(n30277), .B(n30278), .Z(n30275) );
  XOR U32326 ( .A(n[117]), .B(n30276), .Z(n30278) );
  XNOR U32327 ( .A(n30276), .B(n26054), .Z(n30277) );
  XOR U32328 ( .A(n30279), .B(n30280), .Z(n30276) );
  AND U32329 ( .A(n30281), .B(n30282), .Z(n30279) );
  XOR U32330 ( .A(n[116]), .B(n30280), .Z(n30282) );
  XNOR U32331 ( .A(n30280), .B(n26059), .Z(n30281) );
  XOR U32332 ( .A(n30283), .B(n30284), .Z(n30280) );
  AND U32333 ( .A(n30285), .B(n30286), .Z(n30283) );
  XOR U32334 ( .A(n[115]), .B(n30284), .Z(n30286) );
  XNOR U32335 ( .A(n30284), .B(n26064), .Z(n30285) );
  XOR U32336 ( .A(n30287), .B(n30288), .Z(n30284) );
  AND U32337 ( .A(n30289), .B(n30290), .Z(n30287) );
  XOR U32338 ( .A(n[114]), .B(n30288), .Z(n30290) );
  XNOR U32339 ( .A(n30288), .B(n26069), .Z(n30289) );
  XOR U32340 ( .A(n30291), .B(n30292), .Z(n30288) );
  AND U32341 ( .A(n30293), .B(n30294), .Z(n30291) );
  XOR U32342 ( .A(n[113]), .B(n30292), .Z(n30294) );
  XNOR U32343 ( .A(n30292), .B(n26074), .Z(n30293) );
  XOR U32344 ( .A(n30295), .B(n30296), .Z(n30292) );
  AND U32345 ( .A(n30297), .B(n30298), .Z(n30295) );
  XOR U32346 ( .A(n[112]), .B(n30296), .Z(n30298) );
  XNOR U32347 ( .A(n30296), .B(n26079), .Z(n30297) );
  XOR U32348 ( .A(n30299), .B(n30300), .Z(n30296) );
  AND U32349 ( .A(n30301), .B(n30302), .Z(n30299) );
  XOR U32350 ( .A(n[111]), .B(n30300), .Z(n30302) );
  XNOR U32351 ( .A(n30300), .B(n26084), .Z(n30301) );
  XOR U32352 ( .A(n30303), .B(n30304), .Z(n30300) );
  AND U32353 ( .A(n30305), .B(n30306), .Z(n30303) );
  XOR U32354 ( .A(n[110]), .B(n30304), .Z(n30306) );
  XNOR U32355 ( .A(n30304), .B(n26089), .Z(n30305) );
  XOR U32356 ( .A(n30307), .B(n30308), .Z(n30304) );
  AND U32357 ( .A(n30309), .B(n30310), .Z(n30307) );
  XOR U32358 ( .A(n[109]), .B(n30308), .Z(n30310) );
  XNOR U32359 ( .A(n30308), .B(n26094), .Z(n30309) );
  XOR U32360 ( .A(n30311), .B(n30312), .Z(n30308) );
  AND U32361 ( .A(n30313), .B(n30314), .Z(n30311) );
  XOR U32362 ( .A(n[108]), .B(n30312), .Z(n30314) );
  XNOR U32363 ( .A(n30312), .B(n26099), .Z(n30313) );
  XOR U32364 ( .A(n30315), .B(n30316), .Z(n30312) );
  AND U32365 ( .A(n30317), .B(n30318), .Z(n30315) );
  XOR U32366 ( .A(n[107]), .B(n30316), .Z(n30318) );
  XNOR U32367 ( .A(n30316), .B(n26104), .Z(n30317) );
  XOR U32368 ( .A(n30319), .B(n30320), .Z(n30316) );
  AND U32369 ( .A(n30321), .B(n30322), .Z(n30319) );
  XOR U32370 ( .A(n[106]), .B(n30320), .Z(n30322) );
  XNOR U32371 ( .A(n30320), .B(n26109), .Z(n30321) );
  XOR U32372 ( .A(n30323), .B(n30324), .Z(n30320) );
  AND U32373 ( .A(n30325), .B(n30326), .Z(n30323) );
  XOR U32374 ( .A(n[105]), .B(n30324), .Z(n30326) );
  XNOR U32375 ( .A(n30324), .B(n26114), .Z(n30325) );
  XOR U32376 ( .A(n30327), .B(n30328), .Z(n30324) );
  AND U32377 ( .A(n30329), .B(n30330), .Z(n30327) );
  XOR U32378 ( .A(n[104]), .B(n30328), .Z(n30330) );
  XNOR U32379 ( .A(n30328), .B(n26119), .Z(n30329) );
  XOR U32380 ( .A(n30331), .B(n30332), .Z(n30328) );
  AND U32381 ( .A(n30333), .B(n30334), .Z(n30331) );
  XOR U32382 ( .A(n[103]), .B(n30332), .Z(n30334) );
  XNOR U32383 ( .A(n30332), .B(n26124), .Z(n30333) );
  XOR U32384 ( .A(n30335), .B(n30336), .Z(n30332) );
  AND U32385 ( .A(n30337), .B(n30338), .Z(n30335) );
  XOR U32386 ( .A(n[102]), .B(n30336), .Z(n30338) );
  XNOR U32387 ( .A(n30336), .B(n26129), .Z(n30337) );
  XOR U32388 ( .A(n30339), .B(n30340), .Z(n30336) );
  AND U32389 ( .A(n30341), .B(n30342), .Z(n30339) );
  XOR U32390 ( .A(n[101]), .B(n30340), .Z(n30342) );
  XNOR U32391 ( .A(n30340), .B(n26134), .Z(n30341) );
  XOR U32392 ( .A(n30343), .B(n30344), .Z(n30340) );
  AND U32393 ( .A(n30345), .B(n30346), .Z(n30343) );
  XOR U32394 ( .A(n[100]), .B(n30344), .Z(n30346) );
  XNOR U32395 ( .A(n30344), .B(n26139), .Z(n30345) );
  XOR U32396 ( .A(n30347), .B(n30348), .Z(n30344) );
  AND U32397 ( .A(n30349), .B(n30350), .Z(n30347) );
  XOR U32398 ( .A(n[99]), .B(n30348), .Z(n30350) );
  XNOR U32399 ( .A(n30348), .B(n26144), .Z(n30349) );
  XOR U32400 ( .A(n30351), .B(n30352), .Z(n30348) );
  AND U32401 ( .A(n30353), .B(n30354), .Z(n30351) );
  XOR U32402 ( .A(n[98]), .B(n30352), .Z(n30354) );
  XNOR U32403 ( .A(n30352), .B(n26149), .Z(n30353) );
  XOR U32404 ( .A(n30355), .B(n30356), .Z(n30352) );
  AND U32405 ( .A(n30357), .B(n30358), .Z(n30355) );
  XOR U32406 ( .A(n[97]), .B(n30356), .Z(n30358) );
  XNOR U32407 ( .A(n30356), .B(n26154), .Z(n30357) );
  XOR U32408 ( .A(n30359), .B(n30360), .Z(n30356) );
  AND U32409 ( .A(n30361), .B(n30362), .Z(n30359) );
  XOR U32410 ( .A(n[96]), .B(n30360), .Z(n30362) );
  XNOR U32411 ( .A(n30360), .B(n26159), .Z(n30361) );
  XOR U32412 ( .A(n30363), .B(n30364), .Z(n30360) );
  AND U32413 ( .A(n30365), .B(n30366), .Z(n30363) );
  XOR U32414 ( .A(n[95]), .B(n30364), .Z(n30366) );
  XNOR U32415 ( .A(n30364), .B(n26164), .Z(n30365) );
  XOR U32416 ( .A(n30367), .B(n30368), .Z(n30364) );
  AND U32417 ( .A(n30369), .B(n30370), .Z(n30367) );
  XOR U32418 ( .A(n[94]), .B(n30368), .Z(n30370) );
  XNOR U32419 ( .A(n30368), .B(n26169), .Z(n30369) );
  XOR U32420 ( .A(n30371), .B(n30372), .Z(n30368) );
  AND U32421 ( .A(n30373), .B(n30374), .Z(n30371) );
  XOR U32422 ( .A(n[93]), .B(n30372), .Z(n30374) );
  XNOR U32423 ( .A(n30372), .B(n26174), .Z(n30373) );
  XOR U32424 ( .A(n30375), .B(n30376), .Z(n30372) );
  AND U32425 ( .A(n30377), .B(n30378), .Z(n30375) );
  XOR U32426 ( .A(n[92]), .B(n30376), .Z(n30378) );
  XNOR U32427 ( .A(n30376), .B(n26179), .Z(n30377) );
  XOR U32428 ( .A(n30379), .B(n30380), .Z(n30376) );
  AND U32429 ( .A(n30381), .B(n30382), .Z(n30379) );
  XOR U32430 ( .A(n[91]), .B(n30380), .Z(n30382) );
  XNOR U32431 ( .A(n30380), .B(n26184), .Z(n30381) );
  XOR U32432 ( .A(n30383), .B(n30384), .Z(n30380) );
  AND U32433 ( .A(n30385), .B(n30386), .Z(n30383) );
  XOR U32434 ( .A(n[90]), .B(n30384), .Z(n30386) );
  XNOR U32435 ( .A(n30384), .B(n26189), .Z(n30385) );
  XOR U32436 ( .A(n30387), .B(n30388), .Z(n30384) );
  AND U32437 ( .A(n30389), .B(n30390), .Z(n30387) );
  XOR U32438 ( .A(n[89]), .B(n30388), .Z(n30390) );
  XNOR U32439 ( .A(n30388), .B(n26194), .Z(n30389) );
  XOR U32440 ( .A(n30391), .B(n30392), .Z(n30388) );
  AND U32441 ( .A(n30393), .B(n30394), .Z(n30391) );
  XOR U32442 ( .A(n[88]), .B(n30392), .Z(n30394) );
  XNOR U32443 ( .A(n30392), .B(n26199), .Z(n30393) );
  XOR U32444 ( .A(n30395), .B(n30396), .Z(n30392) );
  AND U32445 ( .A(n30397), .B(n30398), .Z(n30395) );
  XOR U32446 ( .A(n[87]), .B(n30396), .Z(n30398) );
  XNOR U32447 ( .A(n30396), .B(n26204), .Z(n30397) );
  XOR U32448 ( .A(n30399), .B(n30400), .Z(n30396) );
  AND U32449 ( .A(n30401), .B(n30402), .Z(n30399) );
  XOR U32450 ( .A(n[86]), .B(n30400), .Z(n30402) );
  XNOR U32451 ( .A(n30400), .B(n26209), .Z(n30401) );
  XOR U32452 ( .A(n30403), .B(n30404), .Z(n30400) );
  AND U32453 ( .A(n30405), .B(n30406), .Z(n30403) );
  XOR U32454 ( .A(n[85]), .B(n30404), .Z(n30406) );
  XNOR U32455 ( .A(n30404), .B(n26214), .Z(n30405) );
  XOR U32456 ( .A(n30407), .B(n30408), .Z(n30404) );
  AND U32457 ( .A(n30409), .B(n30410), .Z(n30407) );
  XOR U32458 ( .A(n[84]), .B(n30408), .Z(n30410) );
  XNOR U32459 ( .A(n30408), .B(n26219), .Z(n30409) );
  XOR U32460 ( .A(n30411), .B(n30412), .Z(n30408) );
  AND U32461 ( .A(n30413), .B(n30414), .Z(n30411) );
  XOR U32462 ( .A(n[83]), .B(n30412), .Z(n30414) );
  XNOR U32463 ( .A(n30412), .B(n26224), .Z(n30413) );
  XOR U32464 ( .A(n30415), .B(n30416), .Z(n30412) );
  AND U32465 ( .A(n30417), .B(n30418), .Z(n30415) );
  XOR U32466 ( .A(n[82]), .B(n30416), .Z(n30418) );
  XNOR U32467 ( .A(n30416), .B(n26229), .Z(n30417) );
  XOR U32468 ( .A(n30419), .B(n30420), .Z(n30416) );
  AND U32469 ( .A(n30421), .B(n30422), .Z(n30419) );
  XOR U32470 ( .A(n[81]), .B(n30420), .Z(n30422) );
  XNOR U32471 ( .A(n30420), .B(n26234), .Z(n30421) );
  XOR U32472 ( .A(n30423), .B(n30424), .Z(n30420) );
  AND U32473 ( .A(n30425), .B(n30426), .Z(n30423) );
  XOR U32474 ( .A(n[80]), .B(n30424), .Z(n30426) );
  XNOR U32475 ( .A(n30424), .B(n26239), .Z(n30425) );
  XOR U32476 ( .A(n30427), .B(n30428), .Z(n30424) );
  AND U32477 ( .A(n30429), .B(n30430), .Z(n30427) );
  XOR U32478 ( .A(n[79]), .B(n30428), .Z(n30430) );
  XNOR U32479 ( .A(n30428), .B(n26244), .Z(n30429) );
  XOR U32480 ( .A(n30431), .B(n30432), .Z(n30428) );
  AND U32481 ( .A(n30433), .B(n30434), .Z(n30431) );
  XOR U32482 ( .A(n[78]), .B(n30432), .Z(n30434) );
  XNOR U32483 ( .A(n30432), .B(n26249), .Z(n30433) );
  XOR U32484 ( .A(n30435), .B(n30436), .Z(n30432) );
  AND U32485 ( .A(n30437), .B(n30438), .Z(n30435) );
  XOR U32486 ( .A(n[77]), .B(n30436), .Z(n30438) );
  XNOR U32487 ( .A(n30436), .B(n26254), .Z(n30437) );
  XOR U32488 ( .A(n30439), .B(n30440), .Z(n30436) );
  AND U32489 ( .A(n30441), .B(n30442), .Z(n30439) );
  XOR U32490 ( .A(n[76]), .B(n30440), .Z(n30442) );
  XNOR U32491 ( .A(n30440), .B(n26259), .Z(n30441) );
  XOR U32492 ( .A(n30443), .B(n30444), .Z(n30440) );
  AND U32493 ( .A(n30445), .B(n30446), .Z(n30443) );
  XOR U32494 ( .A(n[75]), .B(n30444), .Z(n30446) );
  XNOR U32495 ( .A(n30444), .B(n26264), .Z(n30445) );
  XOR U32496 ( .A(n30447), .B(n30448), .Z(n30444) );
  AND U32497 ( .A(n30449), .B(n30450), .Z(n30447) );
  XOR U32498 ( .A(n[74]), .B(n30448), .Z(n30450) );
  XNOR U32499 ( .A(n30448), .B(n26269), .Z(n30449) );
  XOR U32500 ( .A(n30451), .B(n30452), .Z(n30448) );
  AND U32501 ( .A(n30453), .B(n30454), .Z(n30451) );
  XOR U32502 ( .A(n[73]), .B(n30452), .Z(n30454) );
  XNOR U32503 ( .A(n30452), .B(n26274), .Z(n30453) );
  XOR U32504 ( .A(n30455), .B(n30456), .Z(n30452) );
  AND U32505 ( .A(n30457), .B(n30458), .Z(n30455) );
  XOR U32506 ( .A(n[72]), .B(n30456), .Z(n30458) );
  XNOR U32507 ( .A(n30456), .B(n26279), .Z(n30457) );
  XOR U32508 ( .A(n30459), .B(n30460), .Z(n30456) );
  AND U32509 ( .A(n30461), .B(n30462), .Z(n30459) );
  XOR U32510 ( .A(n[71]), .B(n30460), .Z(n30462) );
  XNOR U32511 ( .A(n30460), .B(n26284), .Z(n30461) );
  XOR U32512 ( .A(n30463), .B(n30464), .Z(n30460) );
  AND U32513 ( .A(n30465), .B(n30466), .Z(n30463) );
  XOR U32514 ( .A(n[70]), .B(n30464), .Z(n30466) );
  XNOR U32515 ( .A(n30464), .B(n26289), .Z(n30465) );
  XOR U32516 ( .A(n30467), .B(n30468), .Z(n30464) );
  AND U32517 ( .A(n30469), .B(n30470), .Z(n30467) );
  XOR U32518 ( .A(n[69]), .B(n30468), .Z(n30470) );
  XNOR U32519 ( .A(n30468), .B(n26294), .Z(n30469) );
  XOR U32520 ( .A(n30471), .B(n30472), .Z(n30468) );
  AND U32521 ( .A(n30473), .B(n30474), .Z(n30471) );
  XOR U32522 ( .A(n[68]), .B(n30472), .Z(n30474) );
  XNOR U32523 ( .A(n30472), .B(n26299), .Z(n30473) );
  XOR U32524 ( .A(n30475), .B(n30476), .Z(n30472) );
  AND U32525 ( .A(n30477), .B(n30478), .Z(n30475) );
  XOR U32526 ( .A(n[67]), .B(n30476), .Z(n30478) );
  XNOR U32527 ( .A(n30476), .B(n26304), .Z(n30477) );
  XOR U32528 ( .A(n30479), .B(n30480), .Z(n30476) );
  AND U32529 ( .A(n30481), .B(n30482), .Z(n30479) );
  XOR U32530 ( .A(n[66]), .B(n30480), .Z(n30482) );
  XNOR U32531 ( .A(n30480), .B(n26309), .Z(n30481) );
  XOR U32532 ( .A(n30483), .B(n30484), .Z(n30480) );
  AND U32533 ( .A(n30485), .B(n30486), .Z(n30483) );
  XOR U32534 ( .A(n[65]), .B(n30484), .Z(n30486) );
  XNOR U32535 ( .A(n30484), .B(n26314), .Z(n30485) );
  XOR U32536 ( .A(n30487), .B(n30488), .Z(n30484) );
  AND U32537 ( .A(n30489), .B(n30490), .Z(n30487) );
  XOR U32538 ( .A(n[64]), .B(n30488), .Z(n30490) );
  XNOR U32539 ( .A(n30488), .B(n26319), .Z(n30489) );
  XOR U32540 ( .A(n30491), .B(n30492), .Z(n30488) );
  AND U32541 ( .A(n30493), .B(n30494), .Z(n30491) );
  XOR U32542 ( .A(n[63]), .B(n30492), .Z(n30494) );
  XNOR U32543 ( .A(n30492), .B(n26324), .Z(n30493) );
  XOR U32544 ( .A(n30495), .B(n30496), .Z(n30492) );
  AND U32545 ( .A(n30497), .B(n30498), .Z(n30495) );
  XOR U32546 ( .A(n[62]), .B(n30496), .Z(n30498) );
  XNOR U32547 ( .A(n30496), .B(n26329), .Z(n30497) );
  XOR U32548 ( .A(n30499), .B(n30500), .Z(n30496) );
  AND U32549 ( .A(n30501), .B(n30502), .Z(n30499) );
  XOR U32550 ( .A(n[61]), .B(n30500), .Z(n30502) );
  XNOR U32551 ( .A(n30500), .B(n26334), .Z(n30501) );
  XOR U32552 ( .A(n30503), .B(n30504), .Z(n30500) );
  AND U32553 ( .A(n30505), .B(n30506), .Z(n30503) );
  XOR U32554 ( .A(n[60]), .B(n30504), .Z(n30506) );
  XNOR U32555 ( .A(n30504), .B(n26339), .Z(n30505) );
  XOR U32556 ( .A(n30507), .B(n30508), .Z(n30504) );
  AND U32557 ( .A(n30509), .B(n30510), .Z(n30507) );
  XOR U32558 ( .A(n[59]), .B(n30508), .Z(n30510) );
  XNOR U32559 ( .A(n30508), .B(n26344), .Z(n30509) );
  XOR U32560 ( .A(n30511), .B(n30512), .Z(n30508) );
  AND U32561 ( .A(n30513), .B(n30514), .Z(n30511) );
  XOR U32562 ( .A(n[58]), .B(n30512), .Z(n30514) );
  XNOR U32563 ( .A(n30512), .B(n26349), .Z(n30513) );
  XOR U32564 ( .A(n30515), .B(n30516), .Z(n30512) );
  AND U32565 ( .A(n30517), .B(n30518), .Z(n30515) );
  XOR U32566 ( .A(n[57]), .B(n30516), .Z(n30518) );
  XNOR U32567 ( .A(n30516), .B(n26354), .Z(n30517) );
  XOR U32568 ( .A(n30519), .B(n30520), .Z(n30516) );
  AND U32569 ( .A(n30521), .B(n30522), .Z(n30519) );
  XOR U32570 ( .A(n[56]), .B(n30520), .Z(n30522) );
  XNOR U32571 ( .A(n30520), .B(n26359), .Z(n30521) );
  XOR U32572 ( .A(n30523), .B(n30524), .Z(n30520) );
  AND U32573 ( .A(n30525), .B(n30526), .Z(n30523) );
  XOR U32574 ( .A(n[55]), .B(n30524), .Z(n30526) );
  XNOR U32575 ( .A(n30524), .B(n26364), .Z(n30525) );
  XOR U32576 ( .A(n30527), .B(n30528), .Z(n30524) );
  AND U32577 ( .A(n30529), .B(n30530), .Z(n30527) );
  XOR U32578 ( .A(n[54]), .B(n30528), .Z(n30530) );
  XNOR U32579 ( .A(n30528), .B(n26369), .Z(n30529) );
  XOR U32580 ( .A(n30531), .B(n30532), .Z(n30528) );
  AND U32581 ( .A(n30533), .B(n30534), .Z(n30531) );
  XOR U32582 ( .A(n[53]), .B(n30532), .Z(n30534) );
  XNOR U32583 ( .A(n30532), .B(n26374), .Z(n30533) );
  XOR U32584 ( .A(n30535), .B(n30536), .Z(n30532) );
  AND U32585 ( .A(n30537), .B(n30538), .Z(n30535) );
  XOR U32586 ( .A(n[52]), .B(n30536), .Z(n30538) );
  XNOR U32587 ( .A(n30536), .B(n26379), .Z(n30537) );
  XOR U32588 ( .A(n30539), .B(n30540), .Z(n30536) );
  AND U32589 ( .A(n30541), .B(n30542), .Z(n30539) );
  XOR U32590 ( .A(n[51]), .B(n30540), .Z(n30542) );
  XNOR U32591 ( .A(n30540), .B(n26384), .Z(n30541) );
  XOR U32592 ( .A(n30543), .B(n30544), .Z(n30540) );
  AND U32593 ( .A(n30545), .B(n30546), .Z(n30543) );
  XOR U32594 ( .A(n[50]), .B(n30544), .Z(n30546) );
  XNOR U32595 ( .A(n30544), .B(n26389), .Z(n30545) );
  XOR U32596 ( .A(n30547), .B(n30548), .Z(n30544) );
  AND U32597 ( .A(n30549), .B(n30550), .Z(n30547) );
  XOR U32598 ( .A(n[49]), .B(n30548), .Z(n30550) );
  XNOR U32599 ( .A(n30548), .B(n26394), .Z(n30549) );
  XOR U32600 ( .A(n30551), .B(n30552), .Z(n30548) );
  AND U32601 ( .A(n30553), .B(n30554), .Z(n30551) );
  XOR U32602 ( .A(n[48]), .B(n30552), .Z(n30554) );
  XNOR U32603 ( .A(n30552), .B(n26399), .Z(n30553) );
  XOR U32604 ( .A(n30555), .B(n30556), .Z(n30552) );
  AND U32605 ( .A(n30557), .B(n30558), .Z(n30555) );
  XOR U32606 ( .A(n[47]), .B(n30556), .Z(n30558) );
  XNOR U32607 ( .A(n30556), .B(n26404), .Z(n30557) );
  XOR U32608 ( .A(n30559), .B(n30560), .Z(n30556) );
  AND U32609 ( .A(n30561), .B(n30562), .Z(n30559) );
  XOR U32610 ( .A(n[46]), .B(n30560), .Z(n30562) );
  XNOR U32611 ( .A(n30560), .B(n26409), .Z(n30561) );
  XOR U32612 ( .A(n30563), .B(n30564), .Z(n30560) );
  AND U32613 ( .A(n30565), .B(n30566), .Z(n30563) );
  XOR U32614 ( .A(n[45]), .B(n30564), .Z(n30566) );
  XNOR U32615 ( .A(n30564), .B(n26414), .Z(n30565) );
  XOR U32616 ( .A(n30567), .B(n30568), .Z(n30564) );
  AND U32617 ( .A(n30569), .B(n30570), .Z(n30567) );
  XOR U32618 ( .A(n[44]), .B(n30568), .Z(n30570) );
  XNOR U32619 ( .A(n30568), .B(n26419), .Z(n30569) );
  XOR U32620 ( .A(n30571), .B(n30572), .Z(n30568) );
  AND U32621 ( .A(n30573), .B(n30574), .Z(n30571) );
  XOR U32622 ( .A(n[43]), .B(n30572), .Z(n30574) );
  XNOR U32623 ( .A(n30572), .B(n26424), .Z(n30573) );
  XOR U32624 ( .A(n30575), .B(n30576), .Z(n30572) );
  AND U32625 ( .A(n30577), .B(n30578), .Z(n30575) );
  XOR U32626 ( .A(n[42]), .B(n30576), .Z(n30578) );
  XNOR U32627 ( .A(n30576), .B(n26429), .Z(n30577) );
  XOR U32628 ( .A(n30579), .B(n30580), .Z(n30576) );
  AND U32629 ( .A(n30581), .B(n30582), .Z(n30579) );
  XOR U32630 ( .A(n[41]), .B(n30580), .Z(n30582) );
  XNOR U32631 ( .A(n30580), .B(n26434), .Z(n30581) );
  XOR U32632 ( .A(n30583), .B(n30584), .Z(n30580) );
  AND U32633 ( .A(n30585), .B(n30586), .Z(n30583) );
  XOR U32634 ( .A(n[40]), .B(n30584), .Z(n30586) );
  XNOR U32635 ( .A(n30584), .B(n26439), .Z(n30585) );
  XOR U32636 ( .A(n30587), .B(n30588), .Z(n30584) );
  AND U32637 ( .A(n30589), .B(n30590), .Z(n30587) );
  XOR U32638 ( .A(n[39]), .B(n30588), .Z(n30590) );
  XNOR U32639 ( .A(n30588), .B(n26444), .Z(n30589) );
  XOR U32640 ( .A(n30591), .B(n30592), .Z(n30588) );
  AND U32641 ( .A(n30593), .B(n30594), .Z(n30591) );
  XOR U32642 ( .A(n[38]), .B(n30592), .Z(n30594) );
  XNOR U32643 ( .A(n30592), .B(n26449), .Z(n30593) );
  XOR U32644 ( .A(n30595), .B(n30596), .Z(n30592) );
  AND U32645 ( .A(n30597), .B(n30598), .Z(n30595) );
  XOR U32646 ( .A(n[37]), .B(n30596), .Z(n30598) );
  XNOR U32647 ( .A(n30596), .B(n26454), .Z(n30597) );
  XOR U32648 ( .A(n30599), .B(n30600), .Z(n30596) );
  AND U32649 ( .A(n30601), .B(n30602), .Z(n30599) );
  XOR U32650 ( .A(n[36]), .B(n30600), .Z(n30602) );
  XNOR U32651 ( .A(n30600), .B(n26459), .Z(n30601) );
  XOR U32652 ( .A(n30603), .B(n30604), .Z(n30600) );
  AND U32653 ( .A(n30605), .B(n30606), .Z(n30603) );
  XOR U32654 ( .A(n[35]), .B(n30604), .Z(n30606) );
  XNOR U32655 ( .A(n30604), .B(n26464), .Z(n30605) );
  XOR U32656 ( .A(n30607), .B(n30608), .Z(n30604) );
  AND U32657 ( .A(n30609), .B(n30610), .Z(n30607) );
  XOR U32658 ( .A(n[34]), .B(n30608), .Z(n30610) );
  XNOR U32659 ( .A(n30608), .B(n26469), .Z(n30609) );
  XOR U32660 ( .A(n30611), .B(n30612), .Z(n30608) );
  AND U32661 ( .A(n30613), .B(n30614), .Z(n30611) );
  XOR U32662 ( .A(n[33]), .B(n30612), .Z(n30614) );
  XNOR U32663 ( .A(n30612), .B(n26474), .Z(n30613) );
  XOR U32664 ( .A(n30615), .B(n30616), .Z(n30612) );
  AND U32665 ( .A(n30617), .B(n30618), .Z(n30615) );
  XOR U32666 ( .A(n[32]), .B(n30616), .Z(n30618) );
  XNOR U32667 ( .A(n30616), .B(n26479), .Z(n30617) );
  XOR U32668 ( .A(n30619), .B(n30620), .Z(n30616) );
  AND U32669 ( .A(n30621), .B(n30622), .Z(n30619) );
  XOR U32670 ( .A(n[31]), .B(n30620), .Z(n30622) );
  XNOR U32671 ( .A(n30620), .B(n26484), .Z(n30621) );
  XOR U32672 ( .A(n30623), .B(n30624), .Z(n30620) );
  AND U32673 ( .A(n30625), .B(n30626), .Z(n30623) );
  XOR U32674 ( .A(n[30]), .B(n30624), .Z(n30626) );
  XNOR U32675 ( .A(n30624), .B(n26489), .Z(n30625) );
  XOR U32676 ( .A(n30627), .B(n30628), .Z(n30624) );
  AND U32677 ( .A(n30629), .B(n30630), .Z(n30627) );
  XOR U32678 ( .A(n[29]), .B(n30628), .Z(n30630) );
  XNOR U32679 ( .A(n30628), .B(n26494), .Z(n30629) );
  XOR U32680 ( .A(n30631), .B(n30632), .Z(n30628) );
  AND U32681 ( .A(n30633), .B(n30634), .Z(n30631) );
  XOR U32682 ( .A(n[28]), .B(n30632), .Z(n30634) );
  XNOR U32683 ( .A(n30632), .B(n26499), .Z(n30633) );
  XOR U32684 ( .A(n30635), .B(n30636), .Z(n30632) );
  AND U32685 ( .A(n30637), .B(n30638), .Z(n30635) );
  XOR U32686 ( .A(n[27]), .B(n30636), .Z(n30638) );
  XNOR U32687 ( .A(n30636), .B(n26504), .Z(n30637) );
  XOR U32688 ( .A(n30639), .B(n30640), .Z(n30636) );
  AND U32689 ( .A(n30641), .B(n30642), .Z(n30639) );
  XOR U32690 ( .A(n[26]), .B(n30640), .Z(n30642) );
  XNOR U32691 ( .A(n30640), .B(n26509), .Z(n30641) );
  XOR U32692 ( .A(n30643), .B(n30644), .Z(n30640) );
  AND U32693 ( .A(n30645), .B(n30646), .Z(n30643) );
  XOR U32694 ( .A(n[25]), .B(n30644), .Z(n30646) );
  XNOR U32695 ( .A(n30644), .B(n26514), .Z(n30645) );
  XOR U32696 ( .A(n30647), .B(n30648), .Z(n30644) );
  AND U32697 ( .A(n30649), .B(n30650), .Z(n30647) );
  XOR U32698 ( .A(n[24]), .B(n30648), .Z(n30650) );
  XNOR U32699 ( .A(n30648), .B(n26519), .Z(n30649) );
  XOR U32700 ( .A(n30651), .B(n30652), .Z(n30648) );
  AND U32701 ( .A(n30653), .B(n30654), .Z(n30651) );
  XOR U32702 ( .A(n[23]), .B(n30652), .Z(n30654) );
  XNOR U32703 ( .A(n30652), .B(n26524), .Z(n30653) );
  XOR U32704 ( .A(n30655), .B(n30656), .Z(n30652) );
  AND U32705 ( .A(n30657), .B(n30658), .Z(n30655) );
  XOR U32706 ( .A(n[22]), .B(n30656), .Z(n30658) );
  XNOR U32707 ( .A(n30656), .B(n26529), .Z(n30657) );
  XOR U32708 ( .A(n30659), .B(n30660), .Z(n30656) );
  AND U32709 ( .A(n30661), .B(n30662), .Z(n30659) );
  XOR U32710 ( .A(n[21]), .B(n30660), .Z(n30662) );
  XNOR U32711 ( .A(n30660), .B(n26534), .Z(n30661) );
  XOR U32712 ( .A(n30663), .B(n30664), .Z(n30660) );
  AND U32713 ( .A(n30665), .B(n30666), .Z(n30663) );
  XOR U32714 ( .A(n[20]), .B(n30664), .Z(n30666) );
  XNOR U32715 ( .A(n30664), .B(n26539), .Z(n30665) );
  XOR U32716 ( .A(n30667), .B(n30668), .Z(n30664) );
  AND U32717 ( .A(n30669), .B(n30670), .Z(n30667) );
  XOR U32718 ( .A(n[19]), .B(n30668), .Z(n30670) );
  XNOR U32719 ( .A(n30668), .B(n26544), .Z(n30669) );
  XOR U32720 ( .A(n30671), .B(n30672), .Z(n30668) );
  AND U32721 ( .A(n30673), .B(n30674), .Z(n30671) );
  XOR U32722 ( .A(n[18]), .B(n30672), .Z(n30674) );
  XNOR U32723 ( .A(n30672), .B(n26549), .Z(n30673) );
  XOR U32724 ( .A(n30675), .B(n30676), .Z(n30672) );
  AND U32725 ( .A(n30677), .B(n30678), .Z(n30675) );
  XOR U32726 ( .A(n[17]), .B(n30676), .Z(n30678) );
  XNOR U32727 ( .A(n30676), .B(n26554), .Z(n30677) );
  XOR U32728 ( .A(n30679), .B(n30680), .Z(n30676) );
  AND U32729 ( .A(n30681), .B(n30682), .Z(n30679) );
  XOR U32730 ( .A(n[16]), .B(n30680), .Z(n30682) );
  XNOR U32731 ( .A(n30680), .B(n26559), .Z(n30681) );
  XOR U32732 ( .A(n30683), .B(n30684), .Z(n30680) );
  AND U32733 ( .A(n30685), .B(n30686), .Z(n30683) );
  XOR U32734 ( .A(n[15]), .B(n30684), .Z(n30686) );
  XNOR U32735 ( .A(n30684), .B(n26564), .Z(n30685) );
  XOR U32736 ( .A(n30687), .B(n30688), .Z(n30684) );
  AND U32737 ( .A(n30689), .B(n30690), .Z(n30687) );
  XOR U32738 ( .A(n[14]), .B(n30688), .Z(n30690) );
  XNOR U32739 ( .A(n30688), .B(n26569), .Z(n30689) );
  XOR U32740 ( .A(n30691), .B(n30692), .Z(n30688) );
  AND U32741 ( .A(n30693), .B(n30694), .Z(n30691) );
  XOR U32742 ( .A(n[13]), .B(n30692), .Z(n30694) );
  XNOR U32743 ( .A(n30692), .B(n26574), .Z(n30693) );
  XOR U32744 ( .A(n30695), .B(n30696), .Z(n30692) );
  AND U32745 ( .A(n30697), .B(n30698), .Z(n30695) );
  XOR U32746 ( .A(n[12]), .B(n30696), .Z(n30698) );
  XNOR U32747 ( .A(n30696), .B(n26579), .Z(n30697) );
  XOR U32748 ( .A(n30699), .B(n30700), .Z(n30696) );
  AND U32749 ( .A(n30701), .B(n30702), .Z(n30699) );
  XOR U32750 ( .A(n[11]), .B(n30700), .Z(n30702) );
  XNOR U32751 ( .A(n30700), .B(n26584), .Z(n30701) );
  XOR U32752 ( .A(n30703), .B(n30704), .Z(n30700) );
  AND U32753 ( .A(n30705), .B(n30706), .Z(n30703) );
  XOR U32754 ( .A(n[10]), .B(n30704), .Z(n30706) );
  XNOR U32755 ( .A(n30704), .B(n26589), .Z(n30705) );
  XOR U32756 ( .A(n30707), .B(n30708), .Z(n30704) );
  AND U32757 ( .A(n30709), .B(n30710), .Z(n30707) );
  XOR U32758 ( .A(n[9]), .B(n30708), .Z(n30710) );
  XNOR U32759 ( .A(n30708), .B(n26594), .Z(n30709) );
  XOR U32760 ( .A(n30711), .B(n30712), .Z(n30708) );
  AND U32761 ( .A(n30713), .B(n30714), .Z(n30711) );
  XOR U32762 ( .A(n[8]), .B(n30712), .Z(n30714) );
  XNOR U32763 ( .A(n30712), .B(n26599), .Z(n30713) );
  XOR U32764 ( .A(n30715), .B(n30716), .Z(n30712) );
  AND U32765 ( .A(n30717), .B(n30718), .Z(n30715) );
  XOR U32766 ( .A(n[7]), .B(n30716), .Z(n30718) );
  XNOR U32767 ( .A(n30716), .B(n26604), .Z(n30717) );
  XOR U32768 ( .A(n30719), .B(n30720), .Z(n30716) );
  AND U32769 ( .A(n30721), .B(n30722), .Z(n30719) );
  XOR U32770 ( .A(n[6]), .B(n30720), .Z(n30722) );
  XNOR U32771 ( .A(n30720), .B(n26609), .Z(n30721) );
  XOR U32772 ( .A(n30723), .B(n30724), .Z(n30720) );
  AND U32773 ( .A(n30725), .B(n30726), .Z(n30723) );
  XOR U32774 ( .A(n[5]), .B(n30724), .Z(n30726) );
  XNOR U32775 ( .A(n30724), .B(n26614), .Z(n30725) );
  XOR U32776 ( .A(n30727), .B(n30728), .Z(n30724) );
  AND U32777 ( .A(n30729), .B(n30730), .Z(n30727) );
  XOR U32778 ( .A(n[4]), .B(n30728), .Z(n30730) );
  XNOR U32779 ( .A(n30728), .B(n26619), .Z(n30729) );
  XOR U32780 ( .A(n30731), .B(n30732), .Z(n30728) );
  AND U32781 ( .A(n30733), .B(n30734), .Z(n30731) );
  XOR U32782 ( .A(n[3]), .B(n30732), .Z(n30734) );
  XNOR U32783 ( .A(n30732), .B(n26624), .Z(n30733) );
  XNOR U32784 ( .A(n30735), .B(n30736), .Z(n30732) );
  AND U32785 ( .A(n30737), .B(n30738), .Z(n30735) );
  XNOR U32786 ( .A(n[2]), .B(n30736), .Z(n30738) );
  XNOR U32787 ( .A(n30736), .B(n26629), .Z(n30737) );
  XNOR U32788 ( .A(n30739), .B(n30740), .Z(n30736) );
  NAND U32789 ( .A(n30741), .B(n30742), .Z(n30740) );
  XOR U32790 ( .A(n[1]), .B(n30743), .Z(n30742) );
  XOR U32791 ( .A(n30739), .B(n26634), .Z(n30741) );
  XNOR U32792 ( .A(\modmult_1/zin[0][0] ), .B(n30744), .Z(n26634) );
  IV U32793 ( .A(n30743), .Z(n30739) );
  ANDN U32794 ( .B(n[0]), .A(n21514), .Z(n30743) );
  XOR U32795 ( .A(n30745), .B(n30746), .Z(n21514) );
  ANDN U32796 ( .B(\modmult_1/xin[1023] ), .A(n30747), .Z(n30745) );
  IV U32797 ( .A(n30746), .Z(n30747) );
  XNOR U32798 ( .A(m[0]), .B(n30748), .Z(n30746) );
  NAND U32799 ( .A(n30749), .B(mul_pow), .Z(n30748) );
  XOR U32800 ( .A(m[0]), .B(c[0]), .Z(n30749) );
  XOR U32801 ( .A(n30750), .B(n30751), .Z(n26629) );
  XOR U32802 ( .A(n30752), .B(n30753), .Z(n26624) );
  XOR U32803 ( .A(n30754), .B(n30755), .Z(n26619) );
  XOR U32804 ( .A(n30756), .B(n30757), .Z(n26614) );
  XOR U32805 ( .A(n30758), .B(n30759), .Z(n26609) );
  XOR U32806 ( .A(n30760), .B(n30761), .Z(n26604) );
  XOR U32807 ( .A(n30762), .B(n30763), .Z(n26599) );
  XOR U32808 ( .A(n30764), .B(n30765), .Z(n26594) );
  XOR U32809 ( .A(n30766), .B(n30767), .Z(n26589) );
  XOR U32810 ( .A(n30768), .B(n30769), .Z(n26584) );
  XOR U32811 ( .A(n30770), .B(n30771), .Z(n26579) );
  XOR U32812 ( .A(n30772), .B(n30773), .Z(n26574) );
  XOR U32813 ( .A(n30774), .B(n30775), .Z(n26569) );
  XOR U32814 ( .A(n30776), .B(n30777), .Z(n26564) );
  XOR U32815 ( .A(n30778), .B(n30779), .Z(n26559) );
  XOR U32816 ( .A(n30780), .B(n30781), .Z(n26554) );
  XOR U32817 ( .A(n30782), .B(n30783), .Z(n26549) );
  XOR U32818 ( .A(n30784), .B(n30785), .Z(n26544) );
  XOR U32819 ( .A(n30786), .B(n30787), .Z(n26539) );
  XOR U32820 ( .A(n30788), .B(n30789), .Z(n26534) );
  XOR U32821 ( .A(n30790), .B(n30791), .Z(n26529) );
  XOR U32822 ( .A(n30792), .B(n30793), .Z(n26524) );
  XOR U32823 ( .A(n30794), .B(n30795), .Z(n26519) );
  XOR U32824 ( .A(n30796), .B(n30797), .Z(n26514) );
  XOR U32825 ( .A(n30798), .B(n30799), .Z(n26509) );
  XOR U32826 ( .A(n30800), .B(n30801), .Z(n26504) );
  XOR U32827 ( .A(n30802), .B(n30803), .Z(n26499) );
  XOR U32828 ( .A(n30804), .B(n30805), .Z(n26494) );
  XOR U32829 ( .A(n30806), .B(n30807), .Z(n26489) );
  XOR U32830 ( .A(n30808), .B(n30809), .Z(n26484) );
  XOR U32831 ( .A(n30810), .B(n30811), .Z(n26479) );
  XOR U32832 ( .A(n30812), .B(n30813), .Z(n26474) );
  XOR U32833 ( .A(n30814), .B(n30815), .Z(n26469) );
  XOR U32834 ( .A(n30816), .B(n30817), .Z(n26464) );
  XOR U32835 ( .A(n30818), .B(n30819), .Z(n26459) );
  XOR U32836 ( .A(n30820), .B(n30821), .Z(n26454) );
  XOR U32837 ( .A(n30822), .B(n30823), .Z(n26449) );
  XOR U32838 ( .A(n30824), .B(n30825), .Z(n26444) );
  XOR U32839 ( .A(n30826), .B(n30827), .Z(n26439) );
  XOR U32840 ( .A(n30828), .B(n30829), .Z(n26434) );
  XOR U32841 ( .A(n30830), .B(n30831), .Z(n26429) );
  XOR U32842 ( .A(n30832), .B(n30833), .Z(n26424) );
  XOR U32843 ( .A(n30834), .B(n30835), .Z(n26419) );
  XOR U32844 ( .A(n30836), .B(n30837), .Z(n26414) );
  XOR U32845 ( .A(n30838), .B(n30839), .Z(n26409) );
  XOR U32846 ( .A(n30840), .B(n30841), .Z(n26404) );
  XOR U32847 ( .A(n30842), .B(n30843), .Z(n26399) );
  XOR U32848 ( .A(n30844), .B(n30845), .Z(n26394) );
  XOR U32849 ( .A(n30846), .B(n30847), .Z(n26389) );
  XOR U32850 ( .A(n30848), .B(n30849), .Z(n26384) );
  XOR U32851 ( .A(n30850), .B(n30851), .Z(n26379) );
  XOR U32852 ( .A(n30852), .B(n30853), .Z(n26374) );
  XOR U32853 ( .A(n30854), .B(n30855), .Z(n26369) );
  XOR U32854 ( .A(n30856), .B(n30857), .Z(n26364) );
  XOR U32855 ( .A(n30858), .B(n30859), .Z(n26359) );
  XOR U32856 ( .A(n30860), .B(n30861), .Z(n26354) );
  XOR U32857 ( .A(n30862), .B(n30863), .Z(n26349) );
  XOR U32858 ( .A(n30864), .B(n30865), .Z(n26344) );
  XOR U32859 ( .A(n30866), .B(n30867), .Z(n26339) );
  XOR U32860 ( .A(n30868), .B(n30869), .Z(n26334) );
  XOR U32861 ( .A(n30870), .B(n30871), .Z(n26329) );
  XOR U32862 ( .A(n30872), .B(n30873), .Z(n26324) );
  XOR U32863 ( .A(n30874), .B(n30875), .Z(n26319) );
  XOR U32864 ( .A(n30876), .B(n30877), .Z(n26314) );
  XOR U32865 ( .A(n30878), .B(n30879), .Z(n26309) );
  XOR U32866 ( .A(n30880), .B(n30881), .Z(n26304) );
  XOR U32867 ( .A(n30882), .B(n30883), .Z(n26299) );
  XOR U32868 ( .A(n30884), .B(n30885), .Z(n26294) );
  XOR U32869 ( .A(n30886), .B(n30887), .Z(n26289) );
  XOR U32870 ( .A(n30888), .B(n30889), .Z(n26284) );
  XOR U32871 ( .A(n30890), .B(n30891), .Z(n26279) );
  XOR U32872 ( .A(n30892), .B(n30893), .Z(n26274) );
  XOR U32873 ( .A(n30894), .B(n30895), .Z(n26269) );
  XOR U32874 ( .A(n30896), .B(n30897), .Z(n26264) );
  XOR U32875 ( .A(n30898), .B(n30899), .Z(n26259) );
  XOR U32876 ( .A(n30900), .B(n30901), .Z(n26254) );
  XOR U32877 ( .A(n30902), .B(n30903), .Z(n26249) );
  XOR U32878 ( .A(n30904), .B(n30905), .Z(n26244) );
  XOR U32879 ( .A(n30906), .B(n30907), .Z(n26239) );
  XOR U32880 ( .A(n30908), .B(n30909), .Z(n26234) );
  XOR U32881 ( .A(n30910), .B(n30911), .Z(n26229) );
  XOR U32882 ( .A(n30912), .B(n30913), .Z(n26224) );
  XOR U32883 ( .A(n30914), .B(n30915), .Z(n26219) );
  XOR U32884 ( .A(n30916), .B(n30917), .Z(n26214) );
  XOR U32885 ( .A(n30918), .B(n30919), .Z(n26209) );
  XOR U32886 ( .A(n30920), .B(n30921), .Z(n26204) );
  XOR U32887 ( .A(n30922), .B(n30923), .Z(n26199) );
  XOR U32888 ( .A(n30924), .B(n30925), .Z(n26194) );
  XOR U32889 ( .A(n30926), .B(n30927), .Z(n26189) );
  XOR U32890 ( .A(n30928), .B(n30929), .Z(n26184) );
  XOR U32891 ( .A(n30930), .B(n30931), .Z(n26179) );
  XOR U32892 ( .A(n30932), .B(n30933), .Z(n26174) );
  XOR U32893 ( .A(n30934), .B(n30935), .Z(n26169) );
  XOR U32894 ( .A(n30936), .B(n30937), .Z(n26164) );
  XOR U32895 ( .A(n30938), .B(n30939), .Z(n26159) );
  XOR U32896 ( .A(n30940), .B(n30941), .Z(n26154) );
  XOR U32897 ( .A(n30942), .B(n30943), .Z(n26149) );
  XOR U32898 ( .A(n30944), .B(n30945), .Z(n26144) );
  XOR U32899 ( .A(n30946), .B(n30947), .Z(n26139) );
  XOR U32900 ( .A(n30948), .B(n30949), .Z(n26134) );
  XOR U32901 ( .A(n30950), .B(n30951), .Z(n26129) );
  XOR U32902 ( .A(n30952), .B(n30953), .Z(n26124) );
  XOR U32903 ( .A(n30954), .B(n30955), .Z(n26119) );
  XOR U32904 ( .A(n30956), .B(n30957), .Z(n26114) );
  XOR U32905 ( .A(n30958), .B(n30959), .Z(n26109) );
  XOR U32906 ( .A(n30960), .B(n30961), .Z(n26104) );
  XOR U32907 ( .A(n30962), .B(n30963), .Z(n26099) );
  XOR U32908 ( .A(n30964), .B(n30965), .Z(n26094) );
  XOR U32909 ( .A(n30966), .B(n30967), .Z(n26089) );
  XOR U32910 ( .A(n30968), .B(n30969), .Z(n26084) );
  XOR U32911 ( .A(n30970), .B(n30971), .Z(n26079) );
  XOR U32912 ( .A(n30972), .B(n30973), .Z(n26074) );
  XOR U32913 ( .A(n30974), .B(n30975), .Z(n26069) );
  XOR U32914 ( .A(n30976), .B(n30977), .Z(n26064) );
  XOR U32915 ( .A(n30978), .B(n30979), .Z(n26059) );
  XOR U32916 ( .A(n30980), .B(n30981), .Z(n26054) );
  XOR U32917 ( .A(n30982), .B(n30983), .Z(n26049) );
  XOR U32918 ( .A(n30984), .B(n30985), .Z(n26044) );
  XOR U32919 ( .A(n30986), .B(n30987), .Z(n26039) );
  XOR U32920 ( .A(n30988), .B(n30989), .Z(n26034) );
  XOR U32921 ( .A(n30990), .B(n30991), .Z(n26029) );
  XOR U32922 ( .A(n30992), .B(n30993), .Z(n26024) );
  XOR U32923 ( .A(n30994), .B(n30995), .Z(n26019) );
  XOR U32924 ( .A(n30996), .B(n30997), .Z(n26014) );
  XOR U32925 ( .A(n30998), .B(n30999), .Z(n26009) );
  XOR U32926 ( .A(n31000), .B(n31001), .Z(n26004) );
  XOR U32927 ( .A(n31002), .B(n31003), .Z(n25999) );
  XOR U32928 ( .A(n31004), .B(n31005), .Z(n25994) );
  XOR U32929 ( .A(n31006), .B(n31007), .Z(n25989) );
  XOR U32930 ( .A(n31008), .B(n31009), .Z(n25984) );
  XOR U32931 ( .A(n31010), .B(n31011), .Z(n25979) );
  XOR U32932 ( .A(n31012), .B(n31013), .Z(n25974) );
  XOR U32933 ( .A(n31014), .B(n31015), .Z(n25969) );
  XOR U32934 ( .A(n31016), .B(n31017), .Z(n25964) );
  XOR U32935 ( .A(n31018), .B(n31019), .Z(n25959) );
  XOR U32936 ( .A(n31020), .B(n31021), .Z(n25954) );
  XOR U32937 ( .A(n31022), .B(n31023), .Z(n25949) );
  XOR U32938 ( .A(n31024), .B(n31025), .Z(n25944) );
  XOR U32939 ( .A(n31026), .B(n31027), .Z(n25939) );
  XOR U32940 ( .A(n31028), .B(n31029), .Z(n25934) );
  XOR U32941 ( .A(n31030), .B(n31031), .Z(n25929) );
  XOR U32942 ( .A(n31032), .B(n31033), .Z(n25924) );
  XOR U32943 ( .A(n31034), .B(n31035), .Z(n25919) );
  XOR U32944 ( .A(n31036), .B(n31037), .Z(n25914) );
  XOR U32945 ( .A(n31038), .B(n31039), .Z(n25909) );
  XOR U32946 ( .A(n31040), .B(n31041), .Z(n25904) );
  XOR U32947 ( .A(n31042), .B(n31043), .Z(n25899) );
  XOR U32948 ( .A(n31044), .B(n31045), .Z(n25894) );
  XOR U32949 ( .A(n31046), .B(n31047), .Z(n25889) );
  XOR U32950 ( .A(n31048), .B(n31049), .Z(n25884) );
  XOR U32951 ( .A(n31050), .B(n31051), .Z(n25879) );
  XOR U32952 ( .A(n31052), .B(n31053), .Z(n25874) );
  XOR U32953 ( .A(n31054), .B(n31055), .Z(n25869) );
  XOR U32954 ( .A(n31056), .B(n31057), .Z(n25864) );
  XOR U32955 ( .A(n31058), .B(n31059), .Z(n25859) );
  XOR U32956 ( .A(n31060), .B(n31061), .Z(n25854) );
  XOR U32957 ( .A(n31062), .B(n31063), .Z(n25849) );
  XOR U32958 ( .A(n31064), .B(n31065), .Z(n25844) );
  XOR U32959 ( .A(n31066), .B(n31067), .Z(n25839) );
  XOR U32960 ( .A(n31068), .B(n31069), .Z(n25834) );
  XOR U32961 ( .A(n31070), .B(n31071), .Z(n25829) );
  XOR U32962 ( .A(n31072), .B(n31073), .Z(n25824) );
  XOR U32963 ( .A(n31074), .B(n31075), .Z(n25819) );
  XOR U32964 ( .A(n31076), .B(n31077), .Z(n25814) );
  XOR U32965 ( .A(n31078), .B(n31079), .Z(n25809) );
  XOR U32966 ( .A(n31080), .B(n31081), .Z(n25804) );
  XOR U32967 ( .A(n31082), .B(n31083), .Z(n25799) );
  XOR U32968 ( .A(n31084), .B(n31085), .Z(n25794) );
  XOR U32969 ( .A(n31086), .B(n31087), .Z(n25789) );
  XOR U32970 ( .A(n31088), .B(n31089), .Z(n25784) );
  XOR U32971 ( .A(n31090), .B(n31091), .Z(n25779) );
  XOR U32972 ( .A(n31092), .B(n31093), .Z(n25774) );
  XOR U32973 ( .A(n31094), .B(n31095), .Z(n25769) );
  XOR U32974 ( .A(n31096), .B(n31097), .Z(n25764) );
  XOR U32975 ( .A(n31098), .B(n31099), .Z(n25759) );
  XOR U32976 ( .A(n31100), .B(n31101), .Z(n25754) );
  XOR U32977 ( .A(n31102), .B(n31103), .Z(n25749) );
  XOR U32978 ( .A(n31104), .B(n31105), .Z(n25744) );
  XOR U32979 ( .A(n31106), .B(n31107), .Z(n25739) );
  XOR U32980 ( .A(n31108), .B(n31109), .Z(n25734) );
  XOR U32981 ( .A(n31110), .B(n31111), .Z(n25729) );
  XOR U32982 ( .A(n31112), .B(n31113), .Z(n25724) );
  XOR U32983 ( .A(n31114), .B(n31115), .Z(n25719) );
  XOR U32984 ( .A(n31116), .B(n31117), .Z(n25714) );
  XOR U32985 ( .A(n31118), .B(n31119), .Z(n25709) );
  XOR U32986 ( .A(n31120), .B(n31121), .Z(n25704) );
  XOR U32987 ( .A(n31122), .B(n31123), .Z(n25699) );
  XOR U32988 ( .A(n31124), .B(n31125), .Z(n25694) );
  XOR U32989 ( .A(n31126), .B(n31127), .Z(n25689) );
  XOR U32990 ( .A(n31128), .B(n31129), .Z(n25684) );
  XOR U32991 ( .A(n31130), .B(n31131), .Z(n25679) );
  XOR U32992 ( .A(n31132), .B(n31133), .Z(n25674) );
  XOR U32993 ( .A(n31134), .B(n31135), .Z(n25669) );
  XOR U32994 ( .A(n31136), .B(n31137), .Z(n25664) );
  XOR U32995 ( .A(n31138), .B(n31139), .Z(n25659) );
  XOR U32996 ( .A(n31140), .B(n31141), .Z(n25654) );
  XOR U32997 ( .A(n31142), .B(n31143), .Z(n25649) );
  XOR U32998 ( .A(n31144), .B(n31145), .Z(n25644) );
  XOR U32999 ( .A(n31146), .B(n31147), .Z(n25639) );
  XOR U33000 ( .A(n31148), .B(n31149), .Z(n25634) );
  XOR U33001 ( .A(n31150), .B(n31151), .Z(n25629) );
  XOR U33002 ( .A(n31152), .B(n31153), .Z(n25624) );
  XOR U33003 ( .A(n31154), .B(n31155), .Z(n25619) );
  XOR U33004 ( .A(n31156), .B(n31157), .Z(n25614) );
  XOR U33005 ( .A(n31158), .B(n31159), .Z(n25609) );
  XOR U33006 ( .A(n31160), .B(n31161), .Z(n25604) );
  XOR U33007 ( .A(n31162), .B(n31163), .Z(n25599) );
  XOR U33008 ( .A(n31164), .B(n31165), .Z(n25594) );
  XOR U33009 ( .A(n31166), .B(n31167), .Z(n25589) );
  XOR U33010 ( .A(n31168), .B(n31169), .Z(n25584) );
  XOR U33011 ( .A(n31170), .B(n31171), .Z(n25579) );
  XOR U33012 ( .A(n31172), .B(n31173), .Z(n25574) );
  XOR U33013 ( .A(n31174), .B(n31175), .Z(n25569) );
  XOR U33014 ( .A(n31176), .B(n31177), .Z(n25564) );
  XOR U33015 ( .A(n31178), .B(n31179), .Z(n25559) );
  XOR U33016 ( .A(n31180), .B(n31181), .Z(n25554) );
  XOR U33017 ( .A(n31182), .B(n31183), .Z(n25549) );
  XOR U33018 ( .A(n31184), .B(n31185), .Z(n25544) );
  XOR U33019 ( .A(n31186), .B(n31187), .Z(n25539) );
  XOR U33020 ( .A(n31188), .B(n31189), .Z(n25534) );
  XOR U33021 ( .A(n31190), .B(n31191), .Z(n25529) );
  XOR U33022 ( .A(n31192), .B(n31193), .Z(n25524) );
  XOR U33023 ( .A(n31194), .B(n31195), .Z(n25519) );
  XOR U33024 ( .A(n31196), .B(n31197), .Z(n25514) );
  XOR U33025 ( .A(n31198), .B(n31199), .Z(n25509) );
  XOR U33026 ( .A(n31200), .B(n31201), .Z(n25504) );
  XOR U33027 ( .A(n31202), .B(n31203), .Z(n25499) );
  XOR U33028 ( .A(n31204), .B(n31205), .Z(n25494) );
  XOR U33029 ( .A(n31206), .B(n31207), .Z(n25489) );
  XOR U33030 ( .A(n31208), .B(n31209), .Z(n25484) );
  XOR U33031 ( .A(n31210), .B(n31211), .Z(n25479) );
  XOR U33032 ( .A(n31212), .B(n31213), .Z(n25474) );
  XOR U33033 ( .A(n31214), .B(n31215), .Z(n25469) );
  XOR U33034 ( .A(n31216), .B(n31217), .Z(n25464) );
  XOR U33035 ( .A(n31218), .B(n31219), .Z(n25459) );
  XOR U33036 ( .A(n31220), .B(n31221), .Z(n25454) );
  XOR U33037 ( .A(n31222), .B(n31223), .Z(n25449) );
  XOR U33038 ( .A(n31224), .B(n31225), .Z(n25444) );
  XOR U33039 ( .A(n31226), .B(n31227), .Z(n25439) );
  XOR U33040 ( .A(n31228), .B(n31229), .Z(n25434) );
  XOR U33041 ( .A(n31230), .B(n31231), .Z(n25429) );
  XOR U33042 ( .A(n31232), .B(n31233), .Z(n25424) );
  XOR U33043 ( .A(n31234), .B(n31235), .Z(n25419) );
  XOR U33044 ( .A(n31236), .B(n31237), .Z(n25414) );
  XOR U33045 ( .A(n31238), .B(n31239), .Z(n25409) );
  XOR U33046 ( .A(n31240), .B(n31241), .Z(n25404) );
  XOR U33047 ( .A(n31242), .B(n31243), .Z(n25399) );
  XOR U33048 ( .A(n31244), .B(n31245), .Z(n25394) );
  XOR U33049 ( .A(n31246), .B(n31247), .Z(n25389) );
  XOR U33050 ( .A(n31248), .B(n31249), .Z(n25384) );
  XOR U33051 ( .A(n31250), .B(n31251), .Z(n25379) );
  XOR U33052 ( .A(n31252), .B(n31253), .Z(n25374) );
  XOR U33053 ( .A(n31254), .B(n31255), .Z(n25369) );
  XOR U33054 ( .A(n31256), .B(n31257), .Z(n25364) );
  XOR U33055 ( .A(n31258), .B(n31259), .Z(n25359) );
  XOR U33056 ( .A(n31260), .B(n31261), .Z(n25354) );
  XOR U33057 ( .A(n31262), .B(n31263), .Z(n25349) );
  XOR U33058 ( .A(n31264), .B(n31265), .Z(n25344) );
  XOR U33059 ( .A(n31266), .B(n31267), .Z(n25339) );
  XOR U33060 ( .A(n31268), .B(n31269), .Z(n25334) );
  XOR U33061 ( .A(n31270), .B(n31271), .Z(n25329) );
  XOR U33062 ( .A(n31272), .B(n31273), .Z(n25324) );
  XOR U33063 ( .A(n31274), .B(n31275), .Z(n25319) );
  XOR U33064 ( .A(n31276), .B(n31277), .Z(n25314) );
  XOR U33065 ( .A(n31278), .B(n31279), .Z(n25309) );
  XOR U33066 ( .A(n31280), .B(n31281), .Z(n25304) );
  XOR U33067 ( .A(n31282), .B(n31283), .Z(n25299) );
  XOR U33068 ( .A(n31284), .B(n31285), .Z(n25294) );
  XOR U33069 ( .A(n31286), .B(n31287), .Z(n25289) );
  XOR U33070 ( .A(n31288), .B(n31289), .Z(n25284) );
  XOR U33071 ( .A(n31290), .B(n31291), .Z(n25279) );
  XOR U33072 ( .A(n31292), .B(n31293), .Z(n25274) );
  XOR U33073 ( .A(n31294), .B(n31295), .Z(n25269) );
  XOR U33074 ( .A(n31296), .B(n31297), .Z(n25264) );
  XOR U33075 ( .A(n31298), .B(n31299), .Z(n25259) );
  XOR U33076 ( .A(n31300), .B(n31301), .Z(n25254) );
  XOR U33077 ( .A(n31302), .B(n31303), .Z(n25249) );
  XOR U33078 ( .A(n31304), .B(n31305), .Z(n25244) );
  XOR U33079 ( .A(n31306), .B(n31307), .Z(n25239) );
  XOR U33080 ( .A(n31308), .B(n31309), .Z(n25234) );
  XOR U33081 ( .A(n31310), .B(n31311), .Z(n25229) );
  XOR U33082 ( .A(n31312), .B(n31313), .Z(n25224) );
  XOR U33083 ( .A(n31314), .B(n31315), .Z(n25219) );
  XOR U33084 ( .A(n31316), .B(n31317), .Z(n25214) );
  XOR U33085 ( .A(n31318), .B(n31319), .Z(n25209) );
  XOR U33086 ( .A(n31320), .B(n31321), .Z(n25204) );
  XOR U33087 ( .A(n31322), .B(n31323), .Z(n25199) );
  XOR U33088 ( .A(n31324), .B(n31325), .Z(n25194) );
  XOR U33089 ( .A(n31326), .B(n31327), .Z(n25189) );
  XOR U33090 ( .A(n31328), .B(n31329), .Z(n25184) );
  XOR U33091 ( .A(n31330), .B(n31331), .Z(n25179) );
  XOR U33092 ( .A(n31332), .B(n31333), .Z(n25174) );
  XOR U33093 ( .A(n31334), .B(n31335), .Z(n25169) );
  XOR U33094 ( .A(n31336), .B(n31337), .Z(n25164) );
  XOR U33095 ( .A(n31338), .B(n31339), .Z(n25159) );
  XOR U33096 ( .A(n31340), .B(n31341), .Z(n25154) );
  XOR U33097 ( .A(n31342), .B(n31343), .Z(n25149) );
  XOR U33098 ( .A(n31344), .B(n31345), .Z(n25144) );
  XOR U33099 ( .A(n31346), .B(n31347), .Z(n25139) );
  XOR U33100 ( .A(n31348), .B(n31349), .Z(n25134) );
  XOR U33101 ( .A(n31350), .B(n31351), .Z(n25129) );
  XOR U33102 ( .A(n31352), .B(n31353), .Z(n25124) );
  XOR U33103 ( .A(n31354), .B(n31355), .Z(n25119) );
  XOR U33104 ( .A(n31356), .B(n31357), .Z(n25114) );
  XOR U33105 ( .A(n31358), .B(n31359), .Z(n25109) );
  XOR U33106 ( .A(n31360), .B(n31361), .Z(n25104) );
  XOR U33107 ( .A(n31362), .B(n31363), .Z(n25099) );
  XOR U33108 ( .A(n31364), .B(n31365), .Z(n25094) );
  XOR U33109 ( .A(n31366), .B(n31367), .Z(n25089) );
  XOR U33110 ( .A(n31368), .B(n31369), .Z(n25084) );
  XOR U33111 ( .A(n31370), .B(n31371), .Z(n25079) );
  XOR U33112 ( .A(n31372), .B(n31373), .Z(n25074) );
  XOR U33113 ( .A(n31374), .B(n31375), .Z(n25069) );
  XOR U33114 ( .A(n31376), .B(n31377), .Z(n25064) );
  XOR U33115 ( .A(n31378), .B(n31379), .Z(n25059) );
  XOR U33116 ( .A(n31380), .B(n31381), .Z(n25054) );
  XOR U33117 ( .A(n31382), .B(n31383), .Z(n25049) );
  XOR U33118 ( .A(n31384), .B(n31385), .Z(n25044) );
  XOR U33119 ( .A(n31386), .B(n31387), .Z(n25039) );
  XOR U33120 ( .A(n31388), .B(n31389), .Z(n25034) );
  XOR U33121 ( .A(n31390), .B(n31391), .Z(n25029) );
  XOR U33122 ( .A(n31392), .B(n31393), .Z(n25024) );
  XOR U33123 ( .A(n31394), .B(n31395), .Z(n25019) );
  XOR U33124 ( .A(n31396), .B(n31397), .Z(n25014) );
  XOR U33125 ( .A(n31398), .B(n31399), .Z(n25009) );
  XOR U33126 ( .A(n31400), .B(n31401), .Z(n25004) );
  XOR U33127 ( .A(n31402), .B(n31403), .Z(n24999) );
  XOR U33128 ( .A(n31404), .B(n31405), .Z(n24994) );
  XOR U33129 ( .A(n31406), .B(n31407), .Z(n24989) );
  XOR U33130 ( .A(n31408), .B(n31409), .Z(n24984) );
  XOR U33131 ( .A(n31410), .B(n31411), .Z(n24979) );
  XOR U33132 ( .A(n31412), .B(n31413), .Z(n24974) );
  XOR U33133 ( .A(n31414), .B(n31415), .Z(n24969) );
  XOR U33134 ( .A(n31416), .B(n31417), .Z(n24964) );
  XOR U33135 ( .A(n31418), .B(n31419), .Z(n24959) );
  XOR U33136 ( .A(n31420), .B(n31421), .Z(n24954) );
  XOR U33137 ( .A(n31422), .B(n31423), .Z(n24949) );
  XOR U33138 ( .A(n31424), .B(n31425), .Z(n24944) );
  XOR U33139 ( .A(n31426), .B(n31427), .Z(n24939) );
  XOR U33140 ( .A(n31428), .B(n31429), .Z(n24934) );
  XOR U33141 ( .A(n31430), .B(n31431), .Z(n24929) );
  XOR U33142 ( .A(n31432), .B(n31433), .Z(n24924) );
  XOR U33143 ( .A(n31434), .B(n31435), .Z(n24919) );
  XOR U33144 ( .A(n31436), .B(n31437), .Z(n24914) );
  XOR U33145 ( .A(n31438), .B(n31439), .Z(n24909) );
  XOR U33146 ( .A(n31440), .B(n31441), .Z(n24904) );
  XOR U33147 ( .A(n31442), .B(n31443), .Z(n24899) );
  XOR U33148 ( .A(n31444), .B(n31445), .Z(n24894) );
  XOR U33149 ( .A(n31446), .B(n31447), .Z(n24889) );
  XOR U33150 ( .A(n31448), .B(n31449), .Z(n24884) );
  XOR U33151 ( .A(n31450), .B(n31451), .Z(n24879) );
  XOR U33152 ( .A(n31452), .B(n31453), .Z(n24874) );
  XOR U33153 ( .A(n31454), .B(n31455), .Z(n24869) );
  XOR U33154 ( .A(n31456), .B(n31457), .Z(n24864) );
  XOR U33155 ( .A(n31458), .B(n31459), .Z(n24859) );
  XOR U33156 ( .A(n31460), .B(n31461), .Z(n24854) );
  XOR U33157 ( .A(n31462), .B(n31463), .Z(n24849) );
  XOR U33158 ( .A(n31464), .B(n31465), .Z(n24844) );
  XOR U33159 ( .A(n31466), .B(n31467), .Z(n24839) );
  XOR U33160 ( .A(n31468), .B(n31469), .Z(n24834) );
  XOR U33161 ( .A(n31470), .B(n31471), .Z(n24829) );
  XOR U33162 ( .A(n31472), .B(n31473), .Z(n24824) );
  XOR U33163 ( .A(n31474), .B(n31475), .Z(n24819) );
  XOR U33164 ( .A(n31476), .B(n31477), .Z(n24814) );
  XOR U33165 ( .A(n31478), .B(n31479), .Z(n24809) );
  XOR U33166 ( .A(n31480), .B(n31481), .Z(n24804) );
  XOR U33167 ( .A(n31482), .B(n31483), .Z(n24799) );
  XOR U33168 ( .A(n31484), .B(n31485), .Z(n24794) );
  XOR U33169 ( .A(n31486), .B(n31487), .Z(n24789) );
  XOR U33170 ( .A(n31488), .B(n31489), .Z(n24784) );
  XOR U33171 ( .A(n31490), .B(n31491), .Z(n24779) );
  XOR U33172 ( .A(n31492), .B(n31493), .Z(n24774) );
  XOR U33173 ( .A(n31494), .B(n31495), .Z(n24769) );
  XOR U33174 ( .A(n31496), .B(n31497), .Z(n24764) );
  XOR U33175 ( .A(n31498), .B(n31499), .Z(n24759) );
  XOR U33176 ( .A(n31500), .B(n31501), .Z(n24754) );
  XOR U33177 ( .A(n31502), .B(n31503), .Z(n24749) );
  XOR U33178 ( .A(n31504), .B(n31505), .Z(n24744) );
  XOR U33179 ( .A(n31506), .B(n31507), .Z(n24739) );
  XOR U33180 ( .A(n31508), .B(n31509), .Z(n24734) );
  XOR U33181 ( .A(n31510), .B(n31511), .Z(n24729) );
  XOR U33182 ( .A(n31512), .B(n31513), .Z(n24724) );
  XOR U33183 ( .A(n31514), .B(n31515), .Z(n24719) );
  XOR U33184 ( .A(n31516), .B(n31517), .Z(n24714) );
  XOR U33185 ( .A(n31518), .B(n31519), .Z(n24709) );
  XOR U33186 ( .A(n31520), .B(n31521), .Z(n24704) );
  XOR U33187 ( .A(n31522), .B(n31523), .Z(n24699) );
  XOR U33188 ( .A(n31524), .B(n31525), .Z(n24694) );
  XOR U33189 ( .A(n31526), .B(n31527), .Z(n24689) );
  XOR U33190 ( .A(n31528), .B(n31529), .Z(n24684) );
  XOR U33191 ( .A(n31530), .B(n31531), .Z(n24679) );
  XOR U33192 ( .A(n31532), .B(n31533), .Z(n24674) );
  XOR U33193 ( .A(n31534), .B(n31535), .Z(n24669) );
  XOR U33194 ( .A(n31536), .B(n31537), .Z(n24664) );
  XOR U33195 ( .A(n31538), .B(n31539), .Z(n24659) );
  XOR U33196 ( .A(n31540), .B(n31541), .Z(n24654) );
  XOR U33197 ( .A(n31542), .B(n31543), .Z(n24649) );
  XOR U33198 ( .A(n31544), .B(n31545), .Z(n24644) );
  XOR U33199 ( .A(n31546), .B(n31547), .Z(n24639) );
  XOR U33200 ( .A(n31548), .B(n31549), .Z(n24634) );
  XOR U33201 ( .A(n31550), .B(n31551), .Z(n24629) );
  XOR U33202 ( .A(n31552), .B(n31553), .Z(n24624) );
  XOR U33203 ( .A(n31554), .B(n31555), .Z(n24619) );
  XOR U33204 ( .A(n31556), .B(n31557), .Z(n24614) );
  XOR U33205 ( .A(n31558), .B(n31559), .Z(n24609) );
  XOR U33206 ( .A(n31560), .B(n31561), .Z(n24604) );
  XOR U33207 ( .A(n31562), .B(n31563), .Z(n24599) );
  XOR U33208 ( .A(n31564), .B(n31565), .Z(n24594) );
  XOR U33209 ( .A(n31566), .B(n31567), .Z(n24589) );
  XOR U33210 ( .A(n31568), .B(n31569), .Z(n24584) );
  XOR U33211 ( .A(n31570), .B(n31571), .Z(n24579) );
  XOR U33212 ( .A(n31572), .B(n31573), .Z(n24574) );
  XOR U33213 ( .A(n31574), .B(n31575), .Z(n24569) );
  XOR U33214 ( .A(n31576), .B(n31577), .Z(n24564) );
  XOR U33215 ( .A(n31578), .B(n31579), .Z(n24559) );
  XOR U33216 ( .A(n31580), .B(n31581), .Z(n24554) );
  XOR U33217 ( .A(n31582), .B(n31583), .Z(n24549) );
  XOR U33218 ( .A(n31584), .B(n31585), .Z(n24544) );
  XOR U33219 ( .A(n31586), .B(n31587), .Z(n24539) );
  XOR U33220 ( .A(n31588), .B(n31589), .Z(n24534) );
  XOR U33221 ( .A(n31590), .B(n31591), .Z(n24529) );
  XOR U33222 ( .A(n31592), .B(n31593), .Z(n24524) );
  XOR U33223 ( .A(n31594), .B(n31595), .Z(n24519) );
  XOR U33224 ( .A(n31596), .B(n31597), .Z(n24514) );
  XOR U33225 ( .A(n31598), .B(n31599), .Z(n24509) );
  XOR U33226 ( .A(n31600), .B(n31601), .Z(n24504) );
  XOR U33227 ( .A(n31602), .B(n31603), .Z(n24499) );
  XOR U33228 ( .A(n31604), .B(n31605), .Z(n24494) );
  XOR U33229 ( .A(n31606), .B(n31607), .Z(n24489) );
  XOR U33230 ( .A(n31608), .B(n31609), .Z(n24484) );
  XOR U33231 ( .A(n31610), .B(n31611), .Z(n24479) );
  XOR U33232 ( .A(n31612), .B(n31613), .Z(n24474) );
  XOR U33233 ( .A(n31614), .B(n31615), .Z(n24469) );
  XOR U33234 ( .A(n31616), .B(n31617), .Z(n24464) );
  XOR U33235 ( .A(n31618), .B(n31619), .Z(n24459) );
  XOR U33236 ( .A(n31620), .B(n31621), .Z(n24454) );
  XOR U33237 ( .A(n31622), .B(n31623), .Z(n24449) );
  XOR U33238 ( .A(n31624), .B(n31625), .Z(n24444) );
  XOR U33239 ( .A(n31626), .B(n31627), .Z(n24439) );
  XOR U33240 ( .A(n31628), .B(n31629), .Z(n24434) );
  XOR U33241 ( .A(n31630), .B(n31631), .Z(n24429) );
  XOR U33242 ( .A(n31632), .B(n31633), .Z(n24424) );
  XOR U33243 ( .A(n31634), .B(n31635), .Z(n24419) );
  XOR U33244 ( .A(n31636), .B(n31637), .Z(n24414) );
  XOR U33245 ( .A(n31638), .B(n31639), .Z(n24409) );
  XOR U33246 ( .A(n31640), .B(n31641), .Z(n24404) );
  XOR U33247 ( .A(n31642), .B(n31643), .Z(n24399) );
  XOR U33248 ( .A(n31644), .B(n31645), .Z(n24394) );
  XOR U33249 ( .A(n31646), .B(n31647), .Z(n24389) );
  XOR U33250 ( .A(n31648), .B(n31649), .Z(n24384) );
  XOR U33251 ( .A(n31650), .B(n31651), .Z(n24379) );
  XOR U33252 ( .A(n31652), .B(n31653), .Z(n24374) );
  XOR U33253 ( .A(n31654), .B(n31655), .Z(n24369) );
  XOR U33254 ( .A(n31656), .B(n31657), .Z(n24364) );
  XOR U33255 ( .A(n31658), .B(n31659), .Z(n24359) );
  XOR U33256 ( .A(n31660), .B(n31661), .Z(n24354) );
  XOR U33257 ( .A(n31662), .B(n31663), .Z(n24349) );
  XOR U33258 ( .A(n31664), .B(n31665), .Z(n24344) );
  XOR U33259 ( .A(n31666), .B(n31667), .Z(n24339) );
  XOR U33260 ( .A(n31668), .B(n31669), .Z(n24334) );
  XOR U33261 ( .A(n31670), .B(n31671), .Z(n24329) );
  XOR U33262 ( .A(n31672), .B(n31673), .Z(n24324) );
  XOR U33263 ( .A(n31674), .B(n31675), .Z(n24319) );
  XOR U33264 ( .A(n31676), .B(n31677), .Z(n24314) );
  XOR U33265 ( .A(n31678), .B(n31679), .Z(n24309) );
  XOR U33266 ( .A(n31680), .B(n31681), .Z(n24304) );
  XOR U33267 ( .A(n31682), .B(n31683), .Z(n24299) );
  XOR U33268 ( .A(n31684), .B(n31685), .Z(n24294) );
  XOR U33269 ( .A(n31686), .B(n31687), .Z(n24289) );
  XOR U33270 ( .A(n31688), .B(n31689), .Z(n24284) );
  XOR U33271 ( .A(n31690), .B(n31691), .Z(n24279) );
  XOR U33272 ( .A(n31692), .B(n31693), .Z(n24274) );
  XOR U33273 ( .A(n31694), .B(n31695), .Z(n24269) );
  XOR U33274 ( .A(n31696), .B(n31697), .Z(n24264) );
  XOR U33275 ( .A(n31698), .B(n31699), .Z(n24259) );
  XOR U33276 ( .A(n31700), .B(n31701), .Z(n24254) );
  XOR U33277 ( .A(n31702), .B(n31703), .Z(n24249) );
  XOR U33278 ( .A(n31704), .B(n31705), .Z(n24244) );
  XOR U33279 ( .A(n31706), .B(n31707), .Z(n24239) );
  XOR U33280 ( .A(n31708), .B(n31709), .Z(n24234) );
  XOR U33281 ( .A(n31710), .B(n31711), .Z(n24229) );
  XOR U33282 ( .A(n31712), .B(n31713), .Z(n24224) );
  XOR U33283 ( .A(n31714), .B(n31715), .Z(n24219) );
  XOR U33284 ( .A(n31716), .B(n31717), .Z(n24214) );
  XOR U33285 ( .A(n31718), .B(n31719), .Z(n24209) );
  XOR U33286 ( .A(n31720), .B(n31721), .Z(n24204) );
  XOR U33287 ( .A(n31722), .B(n31723), .Z(n24199) );
  XOR U33288 ( .A(n31724), .B(n31725), .Z(n24194) );
  XOR U33289 ( .A(n31726), .B(n31727), .Z(n24189) );
  XOR U33290 ( .A(n31728), .B(n31729), .Z(n24184) );
  XOR U33291 ( .A(n31730), .B(n31731), .Z(n24179) );
  XOR U33292 ( .A(n31732), .B(n31733), .Z(n24174) );
  XOR U33293 ( .A(n31734), .B(n31735), .Z(n24169) );
  XOR U33294 ( .A(n31736), .B(n31737), .Z(n24164) );
  XOR U33295 ( .A(n31738), .B(n31739), .Z(n24159) );
  XOR U33296 ( .A(n31740), .B(n31741), .Z(n24154) );
  XOR U33297 ( .A(n31742), .B(n31743), .Z(n24149) );
  XOR U33298 ( .A(n31744), .B(n31745), .Z(n24144) );
  XOR U33299 ( .A(n31746), .B(n31747), .Z(n24139) );
  XOR U33300 ( .A(n31748), .B(n31749), .Z(n24134) );
  XOR U33301 ( .A(n31750), .B(n31751), .Z(n24129) );
  XOR U33302 ( .A(n31752), .B(n31753), .Z(n24124) );
  XOR U33303 ( .A(n31754), .B(n31755), .Z(n24119) );
  XOR U33304 ( .A(n31756), .B(n31757), .Z(n24114) );
  XOR U33305 ( .A(n31758), .B(n31759), .Z(n24109) );
  XOR U33306 ( .A(n31760), .B(n31761), .Z(n24104) );
  XOR U33307 ( .A(n31762), .B(n31763), .Z(n24099) );
  XOR U33308 ( .A(n31764), .B(n31765), .Z(n24094) );
  XOR U33309 ( .A(n31766), .B(n31767), .Z(n24089) );
  XOR U33310 ( .A(n31768), .B(n31769), .Z(n24084) );
  XOR U33311 ( .A(n31770), .B(n31771), .Z(n24079) );
  XOR U33312 ( .A(n31772), .B(n31773), .Z(n24074) );
  XOR U33313 ( .A(n31774), .B(n31775), .Z(n24069) );
  XOR U33314 ( .A(n31776), .B(n31777), .Z(n24064) );
  XOR U33315 ( .A(n31778), .B(n31779), .Z(n24059) );
  XOR U33316 ( .A(n31780), .B(n31781), .Z(n24054) );
  XOR U33317 ( .A(n31782), .B(n31783), .Z(n24049) );
  XOR U33318 ( .A(n31784), .B(n31785), .Z(n24044) );
  XOR U33319 ( .A(n31786), .B(n31787), .Z(n24039) );
  XOR U33320 ( .A(n31788), .B(n31789), .Z(n24034) );
  XOR U33321 ( .A(n31790), .B(n31791), .Z(n24029) );
  XOR U33322 ( .A(n31792), .B(n31793), .Z(n24024) );
  XOR U33323 ( .A(n31794), .B(n31795), .Z(n24019) );
  XOR U33324 ( .A(n31796), .B(n31797), .Z(n24014) );
  XOR U33325 ( .A(n31798), .B(n31799), .Z(n24009) );
  XOR U33326 ( .A(n31800), .B(n31801), .Z(n24004) );
  XOR U33327 ( .A(n31802), .B(n31803), .Z(n23999) );
  XOR U33328 ( .A(n31804), .B(n31805), .Z(n23994) );
  XOR U33329 ( .A(n31806), .B(n31807), .Z(n23989) );
  XOR U33330 ( .A(n31808), .B(n31809), .Z(n23984) );
  XOR U33331 ( .A(n31810), .B(n31811), .Z(n23979) );
  XOR U33332 ( .A(n31812), .B(n31813), .Z(n23974) );
  XOR U33333 ( .A(n31814), .B(n31815), .Z(n23969) );
  XOR U33334 ( .A(n31816), .B(n31817), .Z(n23964) );
  XOR U33335 ( .A(n31818), .B(n31819), .Z(n23959) );
  XOR U33336 ( .A(n31820), .B(n31821), .Z(n23954) );
  XOR U33337 ( .A(n31822), .B(n31823), .Z(n23949) );
  XOR U33338 ( .A(n31824), .B(n31825), .Z(n23944) );
  XOR U33339 ( .A(n31826), .B(n31827), .Z(n23939) );
  XOR U33340 ( .A(n31828), .B(n31829), .Z(n23934) );
  XOR U33341 ( .A(n31830), .B(n31831), .Z(n23929) );
  XOR U33342 ( .A(n31832), .B(n31833), .Z(n23924) );
  XOR U33343 ( .A(n31834), .B(n31835), .Z(n23919) );
  XOR U33344 ( .A(n31836), .B(n31837), .Z(n23914) );
  XOR U33345 ( .A(n31838), .B(n31839), .Z(n23909) );
  XOR U33346 ( .A(n31840), .B(n31841), .Z(n23904) );
  XOR U33347 ( .A(n31842), .B(n31843), .Z(n23899) );
  XOR U33348 ( .A(n31844), .B(n31845), .Z(n23894) );
  XOR U33349 ( .A(n31846), .B(n31847), .Z(n23889) );
  XOR U33350 ( .A(n31848), .B(n31849), .Z(n23884) );
  XOR U33351 ( .A(n31850), .B(n31851), .Z(n23879) );
  XOR U33352 ( .A(n31852), .B(n31853), .Z(n23874) );
  XOR U33353 ( .A(n31854), .B(n31855), .Z(n23869) );
  XOR U33354 ( .A(n31856), .B(n31857), .Z(n23864) );
  XOR U33355 ( .A(n31858), .B(n31859), .Z(n23859) );
  XOR U33356 ( .A(n31860), .B(n31861), .Z(n23854) );
  XOR U33357 ( .A(n31862), .B(n31863), .Z(n23849) );
  XOR U33358 ( .A(n31864), .B(n31865), .Z(n23844) );
  XOR U33359 ( .A(n31866), .B(n31867), .Z(n23839) );
  XOR U33360 ( .A(n31868), .B(n31869), .Z(n23834) );
  XOR U33361 ( .A(n31870), .B(n31871), .Z(n23829) );
  XOR U33362 ( .A(n31872), .B(n31873), .Z(n23824) );
  XOR U33363 ( .A(n31874), .B(n31875), .Z(n23819) );
  XOR U33364 ( .A(n31876), .B(n31877), .Z(n23814) );
  XOR U33365 ( .A(n31878), .B(n31879), .Z(n23809) );
  XOR U33366 ( .A(n31880), .B(n31881), .Z(n23804) );
  XOR U33367 ( .A(n31882), .B(n31883), .Z(n23799) );
  XOR U33368 ( .A(n31884), .B(n31885), .Z(n23794) );
  XOR U33369 ( .A(n31886), .B(n31887), .Z(n23789) );
  XOR U33370 ( .A(n31888), .B(n31889), .Z(n23784) );
  XOR U33371 ( .A(n31890), .B(n31891), .Z(n23779) );
  XOR U33372 ( .A(n31892), .B(n31893), .Z(n23774) );
  XOR U33373 ( .A(n31894), .B(n31895), .Z(n23769) );
  XOR U33374 ( .A(n31896), .B(n31897), .Z(n23764) );
  XOR U33375 ( .A(n31898), .B(n31899), .Z(n23759) );
  XOR U33376 ( .A(n31900), .B(n31901), .Z(n23754) );
  XOR U33377 ( .A(n31902), .B(n31903), .Z(n23749) );
  XOR U33378 ( .A(n31904), .B(n31905), .Z(n23744) );
  XOR U33379 ( .A(n31906), .B(n31907), .Z(n23739) );
  XOR U33380 ( .A(n31908), .B(n31909), .Z(n23734) );
  XOR U33381 ( .A(n31910), .B(n31911), .Z(n23729) );
  XOR U33382 ( .A(n31912), .B(n31913), .Z(n23724) );
  XOR U33383 ( .A(n31914), .B(n31915), .Z(n23719) );
  XOR U33384 ( .A(n31916), .B(n31917), .Z(n23714) );
  XOR U33385 ( .A(n31918), .B(n31919), .Z(n23709) );
  XOR U33386 ( .A(n31920), .B(n31921), .Z(n23704) );
  XOR U33387 ( .A(n31922), .B(n31923), .Z(n23699) );
  XOR U33388 ( .A(n31924), .B(n31925), .Z(n23694) );
  XOR U33389 ( .A(n31926), .B(n31927), .Z(n23689) );
  XOR U33390 ( .A(n31928), .B(n31929), .Z(n23684) );
  XOR U33391 ( .A(n31930), .B(n31931), .Z(n23679) );
  XOR U33392 ( .A(n31932), .B(n31933), .Z(n23674) );
  XOR U33393 ( .A(n31934), .B(n31935), .Z(n23669) );
  XOR U33394 ( .A(n31936), .B(n31937), .Z(n23664) );
  XOR U33395 ( .A(n31938), .B(n31939), .Z(n23659) );
  XOR U33396 ( .A(n31940), .B(n31941), .Z(n23654) );
  XOR U33397 ( .A(n31942), .B(n31943), .Z(n23649) );
  XOR U33398 ( .A(n31944), .B(n31945), .Z(n23644) );
  XOR U33399 ( .A(n31946), .B(n31947), .Z(n23639) );
  XOR U33400 ( .A(n31948), .B(n31949), .Z(n23634) );
  XOR U33401 ( .A(n31950), .B(n31951), .Z(n23629) );
  XOR U33402 ( .A(n31952), .B(n31953), .Z(n23624) );
  XOR U33403 ( .A(n31954), .B(n31955), .Z(n23619) );
  XOR U33404 ( .A(n31956), .B(n31957), .Z(n23614) );
  XOR U33405 ( .A(n31958), .B(n31959), .Z(n23609) );
  XOR U33406 ( .A(n31960), .B(n31961), .Z(n23604) );
  XOR U33407 ( .A(n31962), .B(n31963), .Z(n23599) );
  XOR U33408 ( .A(n31964), .B(n31965), .Z(n23594) );
  XOR U33409 ( .A(n31966), .B(n31967), .Z(n23589) );
  XOR U33410 ( .A(n31968), .B(n31969), .Z(n23584) );
  XOR U33411 ( .A(n31970), .B(n31971), .Z(n23579) );
  XOR U33412 ( .A(n31972), .B(n31973), .Z(n23574) );
  XOR U33413 ( .A(n31974), .B(n31975), .Z(n23569) );
  XOR U33414 ( .A(n31976), .B(n31977), .Z(n23564) );
  XOR U33415 ( .A(n31978), .B(n31979), .Z(n23559) );
  XOR U33416 ( .A(n31980), .B(n31981), .Z(n23554) );
  XOR U33417 ( .A(n31982), .B(n31983), .Z(n23549) );
  XOR U33418 ( .A(n31984), .B(n31985), .Z(n23544) );
  XOR U33419 ( .A(n31986), .B(n31987), .Z(n23539) );
  XOR U33420 ( .A(n31988), .B(n31989), .Z(n23534) );
  XOR U33421 ( .A(n31990), .B(n31991), .Z(n23529) );
  XOR U33422 ( .A(n31992), .B(n31993), .Z(n23524) );
  XOR U33423 ( .A(n31994), .B(n31995), .Z(n23519) );
  XOR U33424 ( .A(n31996), .B(n31997), .Z(n23514) );
  XOR U33425 ( .A(n31998), .B(n31999), .Z(n23509) );
  XOR U33426 ( .A(n32000), .B(n32001), .Z(n23504) );
  XOR U33427 ( .A(n32002), .B(n32003), .Z(n23499) );
  XOR U33428 ( .A(n32004), .B(n32005), .Z(n23494) );
  XOR U33429 ( .A(n32006), .B(n32007), .Z(n23489) );
  XOR U33430 ( .A(n32008), .B(n32009), .Z(n23484) );
  XOR U33431 ( .A(n32010), .B(n32011), .Z(n23479) );
  XOR U33432 ( .A(n32012), .B(n32013), .Z(n23474) );
  XOR U33433 ( .A(n32014), .B(n32015), .Z(n23469) );
  XOR U33434 ( .A(n32016), .B(n32017), .Z(n23464) );
  XOR U33435 ( .A(n32018), .B(n32019), .Z(n23459) );
  XOR U33436 ( .A(n32020), .B(n32021), .Z(n23454) );
  XOR U33437 ( .A(n32022), .B(n32023), .Z(n23449) );
  XOR U33438 ( .A(n32024), .B(n32025), .Z(n23444) );
  XOR U33439 ( .A(n32026), .B(n32027), .Z(n23439) );
  XOR U33440 ( .A(n32028), .B(n32029), .Z(n23434) );
  XOR U33441 ( .A(n32030), .B(n32031), .Z(n23429) );
  XOR U33442 ( .A(n32032), .B(n32033), .Z(n23424) );
  XOR U33443 ( .A(n32034), .B(n32035), .Z(n23419) );
  XOR U33444 ( .A(n32036), .B(n32037), .Z(n23414) );
  XOR U33445 ( .A(n32038), .B(n32039), .Z(n23409) );
  XOR U33446 ( .A(n32040), .B(n32041), .Z(n23404) );
  XOR U33447 ( .A(n32042), .B(n32043), .Z(n23399) );
  XOR U33448 ( .A(n32044), .B(n32045), .Z(n23394) );
  XOR U33449 ( .A(n32046), .B(n32047), .Z(n23389) );
  XOR U33450 ( .A(n32048), .B(n32049), .Z(n23384) );
  XOR U33451 ( .A(n32050), .B(n32051), .Z(n23379) );
  XOR U33452 ( .A(n32052), .B(n32053), .Z(n23374) );
  XOR U33453 ( .A(n32054), .B(n32055), .Z(n23369) );
  XOR U33454 ( .A(n32056), .B(n32057), .Z(n23364) );
  XOR U33455 ( .A(n32058), .B(n32059), .Z(n23359) );
  XOR U33456 ( .A(n32060), .B(n32061), .Z(n23354) );
  XOR U33457 ( .A(n32062), .B(n32063), .Z(n23349) );
  XOR U33458 ( .A(n32064), .B(n32065), .Z(n23344) );
  XOR U33459 ( .A(n32066), .B(n32067), .Z(n23339) );
  XOR U33460 ( .A(n32068), .B(n32069), .Z(n23334) );
  XOR U33461 ( .A(n32070), .B(n32071), .Z(n23329) );
  XOR U33462 ( .A(n32072), .B(n32073), .Z(n23324) );
  XOR U33463 ( .A(n32074), .B(n32075), .Z(n23319) );
  XOR U33464 ( .A(n32076), .B(n32077), .Z(n23314) );
  XOR U33465 ( .A(n32078), .B(n32079), .Z(n23309) );
  XOR U33466 ( .A(n32080), .B(n32081), .Z(n23304) );
  XOR U33467 ( .A(n32082), .B(n32083), .Z(n23299) );
  XOR U33468 ( .A(n32084), .B(n32085), .Z(n23294) );
  XOR U33469 ( .A(n32086), .B(n32087), .Z(n23289) );
  XOR U33470 ( .A(n32088), .B(n32089), .Z(n23284) );
  XOR U33471 ( .A(n32090), .B(n32091), .Z(n23279) );
  XOR U33472 ( .A(n32092), .B(n32093), .Z(n23274) );
  XOR U33473 ( .A(n32094), .B(n32095), .Z(n23269) );
  XOR U33474 ( .A(n32096), .B(n32097), .Z(n23264) );
  XOR U33475 ( .A(n32098), .B(n32099), .Z(n23259) );
  XOR U33476 ( .A(n32100), .B(n32101), .Z(n23254) );
  XOR U33477 ( .A(n32102), .B(n32103), .Z(n23249) );
  XOR U33478 ( .A(n32104), .B(n32105), .Z(n23244) );
  XOR U33479 ( .A(n32106), .B(n32107), .Z(n23239) );
  XOR U33480 ( .A(n32108), .B(n32109), .Z(n23234) );
  XOR U33481 ( .A(n32110), .B(n32111), .Z(n23229) );
  XOR U33482 ( .A(n32112), .B(n32113), .Z(n23224) );
  XOR U33483 ( .A(n32114), .B(n32115), .Z(n23219) );
  XOR U33484 ( .A(n32116), .B(n32117), .Z(n23214) );
  XOR U33485 ( .A(n32118), .B(n32119), .Z(n23209) );
  XOR U33486 ( .A(n32120), .B(n32121), .Z(n23204) );
  XOR U33487 ( .A(n32122), .B(n32123), .Z(n23199) );
  XOR U33488 ( .A(n32124), .B(n32125), .Z(n23194) );
  XOR U33489 ( .A(n32126), .B(n32127), .Z(n23189) );
  XOR U33490 ( .A(n32128), .B(n32129), .Z(n23184) );
  XOR U33491 ( .A(n32130), .B(n32131), .Z(n23179) );
  XOR U33492 ( .A(n32132), .B(n32133), .Z(n23174) );
  XOR U33493 ( .A(n32134), .B(n32135), .Z(n23169) );
  XOR U33494 ( .A(n32136), .B(n32137), .Z(n23164) );
  XOR U33495 ( .A(n32138), .B(n32139), .Z(n23159) );
  XOR U33496 ( .A(n32140), .B(n32141), .Z(n23154) );
  XOR U33497 ( .A(n32142), .B(n32143), .Z(n23149) );
  XOR U33498 ( .A(n32144), .B(n32145), .Z(n23144) );
  XOR U33499 ( .A(n32146), .B(n32147), .Z(n23139) );
  XOR U33500 ( .A(n32148), .B(n32149), .Z(n23134) );
  XOR U33501 ( .A(n32150), .B(n32151), .Z(n23129) );
  XOR U33502 ( .A(n32152), .B(n32153), .Z(n23124) );
  XOR U33503 ( .A(n32154), .B(n32155), .Z(n23119) );
  XOR U33504 ( .A(n32156), .B(n32157), .Z(n23114) );
  XOR U33505 ( .A(n32158), .B(n32159), .Z(n23109) );
  XOR U33506 ( .A(n32160), .B(n32161), .Z(n23104) );
  XOR U33507 ( .A(n32162), .B(n32163), .Z(n23099) );
  XOR U33508 ( .A(n32164), .B(n32165), .Z(n23094) );
  XOR U33509 ( .A(n32166), .B(n32167), .Z(n23089) );
  XOR U33510 ( .A(n32168), .B(n32169), .Z(n23084) );
  XOR U33511 ( .A(n32170), .B(n32171), .Z(n23079) );
  XOR U33512 ( .A(n32172), .B(n32173), .Z(n23074) );
  XOR U33513 ( .A(n32174), .B(n32175), .Z(n23069) );
  XOR U33514 ( .A(n32176), .B(n32177), .Z(n23064) );
  XOR U33515 ( .A(n32178), .B(n32179), .Z(n23059) );
  XOR U33516 ( .A(n32180), .B(n32181), .Z(n23054) );
  XOR U33517 ( .A(n32182), .B(n32183), .Z(n23049) );
  XOR U33518 ( .A(n32184), .B(n32185), .Z(n23044) );
  XOR U33519 ( .A(n32186), .B(n32187), .Z(n23039) );
  XOR U33520 ( .A(n32188), .B(n32189), .Z(n23034) );
  XOR U33521 ( .A(n32190), .B(n32191), .Z(n23029) );
  XOR U33522 ( .A(n32192), .B(n32193), .Z(n23024) );
  XOR U33523 ( .A(n32194), .B(n32195), .Z(n23019) );
  XOR U33524 ( .A(n32196), .B(n32197), .Z(n23014) );
  XOR U33525 ( .A(n32198), .B(n32199), .Z(n23009) );
  XOR U33526 ( .A(n32200), .B(n32201), .Z(n23004) );
  XOR U33527 ( .A(n32202), .B(n32203), .Z(n22999) );
  XOR U33528 ( .A(n32204), .B(n32205), .Z(n22994) );
  XOR U33529 ( .A(n32206), .B(n32207), .Z(n22989) );
  XOR U33530 ( .A(n32208), .B(n32209), .Z(n22984) );
  XOR U33531 ( .A(n32210), .B(n32211), .Z(n22979) );
  XOR U33532 ( .A(n32212), .B(n32213), .Z(n22974) );
  XOR U33533 ( .A(n32214), .B(n32215), .Z(n22969) );
  XOR U33534 ( .A(n32216), .B(n32217), .Z(n22964) );
  XOR U33535 ( .A(n32218), .B(n32219), .Z(n22959) );
  XOR U33536 ( .A(n32220), .B(n32221), .Z(n22954) );
  XOR U33537 ( .A(n32222), .B(n32223), .Z(n22949) );
  XOR U33538 ( .A(n32224), .B(n32225), .Z(n22944) );
  XOR U33539 ( .A(n32226), .B(n32227), .Z(n22939) );
  XOR U33540 ( .A(n32228), .B(n32229), .Z(n22934) );
  XOR U33541 ( .A(n32230), .B(n32231), .Z(n22929) );
  XOR U33542 ( .A(n32232), .B(n32233), .Z(n22924) );
  XOR U33543 ( .A(n32234), .B(n32235), .Z(n22919) );
  XOR U33544 ( .A(n32236), .B(n32237), .Z(n22914) );
  XOR U33545 ( .A(n32238), .B(n32239), .Z(n22909) );
  XOR U33546 ( .A(n32240), .B(n32241), .Z(n22904) );
  XOR U33547 ( .A(n32242), .B(n32243), .Z(n22899) );
  XOR U33548 ( .A(n32244), .B(n32245), .Z(n22894) );
  XOR U33549 ( .A(n32246), .B(n32247), .Z(n22889) );
  XOR U33550 ( .A(n32248), .B(n32249), .Z(n22884) );
  XOR U33551 ( .A(n32250), .B(n32251), .Z(n22879) );
  XOR U33552 ( .A(n32252), .B(n32253), .Z(n22874) );
  XOR U33553 ( .A(n32254), .B(n32255), .Z(n22869) );
  XOR U33554 ( .A(n32256), .B(n32257), .Z(n22864) );
  XOR U33555 ( .A(n32258), .B(n32259), .Z(n22859) );
  XOR U33556 ( .A(n32260), .B(n32261), .Z(n22854) );
  XOR U33557 ( .A(n32262), .B(n32263), .Z(n22849) );
  XOR U33558 ( .A(n32264), .B(n32265), .Z(n22844) );
  XOR U33559 ( .A(n32266), .B(n32267), .Z(n22839) );
  XOR U33560 ( .A(n32268), .B(n32269), .Z(n22834) );
  XOR U33561 ( .A(n32270), .B(n32271), .Z(n22829) );
  XOR U33562 ( .A(n32272), .B(n32273), .Z(n22824) );
  XOR U33563 ( .A(n32274), .B(n32275), .Z(n22819) );
  XOR U33564 ( .A(n32276), .B(n32277), .Z(n22814) );
  XOR U33565 ( .A(n32278), .B(n32279), .Z(n22809) );
  XOR U33566 ( .A(n32280), .B(n32281), .Z(n22804) );
  XOR U33567 ( .A(n32282), .B(n32283), .Z(n22799) );
  XOR U33568 ( .A(n32284), .B(n32285), .Z(n22794) );
  XOR U33569 ( .A(n32286), .B(n32287), .Z(n22789) );
  XOR U33570 ( .A(n32288), .B(n32289), .Z(n22784) );
  XOR U33571 ( .A(n32290), .B(n32291), .Z(n22779) );
  XOR U33572 ( .A(n32292), .B(n32293), .Z(n22774) );
  XOR U33573 ( .A(n32294), .B(n32295), .Z(n22769) );
  XOR U33574 ( .A(n32296), .B(n32297), .Z(n22764) );
  XOR U33575 ( .A(n32298), .B(n32299), .Z(n22759) );
  XOR U33576 ( .A(n32300), .B(n32301), .Z(n22754) );
  XOR U33577 ( .A(n32302), .B(n32303), .Z(n22749) );
  XOR U33578 ( .A(n32304), .B(n32305), .Z(n22744) );
  XOR U33579 ( .A(n32306), .B(n32307), .Z(n22739) );
  XOR U33580 ( .A(n32308), .B(n32309), .Z(n22734) );
  XOR U33581 ( .A(n32310), .B(n32311), .Z(n22729) );
  XOR U33582 ( .A(n32312), .B(n32313), .Z(n22724) );
  XOR U33583 ( .A(n32314), .B(n32315), .Z(n22719) );
  XOR U33584 ( .A(n32316), .B(n32317), .Z(n22714) );
  XOR U33585 ( .A(n32318), .B(n32319), .Z(n22709) );
  XOR U33586 ( .A(n32320), .B(n32321), .Z(n22704) );
  XOR U33587 ( .A(n32322), .B(n32323), .Z(n22699) );
  XOR U33588 ( .A(n32324), .B(n32325), .Z(n22694) );
  XOR U33589 ( .A(n32326), .B(n32327), .Z(n22689) );
  XOR U33590 ( .A(n32328), .B(n32329), .Z(n22684) );
  XOR U33591 ( .A(n32330), .B(n32331), .Z(n22679) );
  XOR U33592 ( .A(n32332), .B(n32333), .Z(n22674) );
  XOR U33593 ( .A(n32334), .B(n32335), .Z(n22669) );
  XOR U33594 ( .A(n32336), .B(n32337), .Z(n22664) );
  XOR U33595 ( .A(n32338), .B(n32339), .Z(n22659) );
  XOR U33596 ( .A(n32340), .B(n32341), .Z(n22654) );
  XOR U33597 ( .A(n32342), .B(n32343), .Z(n22649) );
  XOR U33598 ( .A(n32344), .B(n32345), .Z(n22644) );
  XOR U33599 ( .A(n32346), .B(n32347), .Z(n22639) );
  XOR U33600 ( .A(n32348), .B(n32349), .Z(n22634) );
  XOR U33601 ( .A(n32350), .B(n32351), .Z(n22629) );
  XOR U33602 ( .A(n32352), .B(n32353), .Z(n22624) );
  XOR U33603 ( .A(n32354), .B(n32355), .Z(n22619) );
  XOR U33604 ( .A(n32356), .B(n32357), .Z(n22614) );
  XOR U33605 ( .A(n32358), .B(n32359), .Z(n22609) );
  XOR U33606 ( .A(n32360), .B(n32361), .Z(n22604) );
  XOR U33607 ( .A(n32362), .B(n32363), .Z(n22599) );
  XOR U33608 ( .A(n32364), .B(n32365), .Z(n22594) );
  XOR U33609 ( .A(n32366), .B(n32367), .Z(n22589) );
  XOR U33610 ( .A(n32368), .B(n32369), .Z(n22584) );
  XOR U33611 ( .A(n32370), .B(n32371), .Z(n22579) );
  XOR U33612 ( .A(n32372), .B(n32373), .Z(n22574) );
  XOR U33613 ( .A(n32374), .B(n32375), .Z(n22569) );
  XOR U33614 ( .A(n32376), .B(n32377), .Z(n22564) );
  XOR U33615 ( .A(n32378), .B(n32379), .Z(n22559) );
  XOR U33616 ( .A(n32380), .B(n32381), .Z(n22554) );
  XOR U33617 ( .A(n32382), .B(n32383), .Z(n22549) );
  XOR U33618 ( .A(n32384), .B(n32385), .Z(n22544) );
  XOR U33619 ( .A(n32386), .B(n32387), .Z(n22539) );
  XOR U33620 ( .A(n32388), .B(n32389), .Z(n22534) );
  XOR U33621 ( .A(n32390), .B(n32391), .Z(n22529) );
  XOR U33622 ( .A(n32392), .B(n32393), .Z(n22524) );
  XOR U33623 ( .A(n32394), .B(n32395), .Z(n22519) );
  XOR U33624 ( .A(n32396), .B(n32397), .Z(n22514) );
  XOR U33625 ( .A(n32398), .B(n32399), .Z(n22509) );
  XOR U33626 ( .A(n32400), .B(n32401), .Z(n22504) );
  XOR U33627 ( .A(n32402), .B(n32403), .Z(n22499) );
  XOR U33628 ( .A(n32404), .B(n32405), .Z(n22494) );
  XOR U33629 ( .A(n32406), .B(n32407), .Z(n22489) );
  XOR U33630 ( .A(n32408), .B(n32409), .Z(n22484) );
  XOR U33631 ( .A(n32410), .B(n32411), .Z(n22479) );
  XOR U33632 ( .A(n32412), .B(n32413), .Z(n22474) );
  XOR U33633 ( .A(n32414), .B(n32415), .Z(n22469) );
  XOR U33634 ( .A(n32416), .B(n32417), .Z(n22464) );
  XOR U33635 ( .A(n32418), .B(n32419), .Z(n22459) );
  XOR U33636 ( .A(n32420), .B(n32421), .Z(n22454) );
  XOR U33637 ( .A(n32422), .B(n32423), .Z(n22449) );
  XOR U33638 ( .A(n32424), .B(n32425), .Z(n22444) );
  XOR U33639 ( .A(n32426), .B(n32427), .Z(n22439) );
  XOR U33640 ( .A(n32428), .B(n32429), .Z(n22434) );
  XOR U33641 ( .A(n32430), .B(n32431), .Z(n22429) );
  XOR U33642 ( .A(n32432), .B(n32433), .Z(n22424) );
  XOR U33643 ( .A(n32434), .B(n32435), .Z(n22419) );
  XOR U33644 ( .A(n32436), .B(n32437), .Z(n22414) );
  XOR U33645 ( .A(n32438), .B(n32439), .Z(n22409) );
  XOR U33646 ( .A(n32440), .B(n32441), .Z(n22404) );
  XOR U33647 ( .A(n32442), .B(n32443), .Z(n22399) );
  XOR U33648 ( .A(n32444), .B(n32445), .Z(n22394) );
  XOR U33649 ( .A(n32446), .B(n32447), .Z(n22389) );
  XOR U33650 ( .A(n32448), .B(n32449), .Z(n22384) );
  XOR U33651 ( .A(n32450), .B(n32451), .Z(n22379) );
  XOR U33652 ( .A(n32452), .B(n32453), .Z(n22374) );
  XOR U33653 ( .A(n32454), .B(n32455), .Z(n22369) );
  XOR U33654 ( .A(n32456), .B(n32457), .Z(n22364) );
  XOR U33655 ( .A(n32458), .B(n32459), .Z(n22359) );
  XOR U33656 ( .A(n32460), .B(n32461), .Z(n22354) );
  XOR U33657 ( .A(n32462), .B(n32463), .Z(n22349) );
  XOR U33658 ( .A(n32464), .B(n32465), .Z(n22344) );
  XOR U33659 ( .A(n32466), .B(n32467), .Z(n22339) );
  XOR U33660 ( .A(n32468), .B(n32469), .Z(n22334) );
  XOR U33661 ( .A(n32470), .B(n32471), .Z(n22329) );
  XOR U33662 ( .A(n32472), .B(n32473), .Z(n22324) );
  XOR U33663 ( .A(n32474), .B(n32475), .Z(n22319) );
  XOR U33664 ( .A(n32476), .B(n32477), .Z(n22314) );
  XOR U33665 ( .A(n32478), .B(n32479), .Z(n22309) );
  XOR U33666 ( .A(n32480), .B(n32481), .Z(n22304) );
  XOR U33667 ( .A(n32482), .B(n32483), .Z(n22299) );
  XOR U33668 ( .A(n32484), .B(n32485), .Z(n22294) );
  XOR U33669 ( .A(n32486), .B(n32487), .Z(n22289) );
  XOR U33670 ( .A(n32488), .B(n32489), .Z(n22284) );
  XOR U33671 ( .A(n32490), .B(n32491), .Z(n22279) );
  XOR U33672 ( .A(n32492), .B(n32493), .Z(n22274) );
  XOR U33673 ( .A(n32494), .B(n32495), .Z(n22269) );
  XOR U33674 ( .A(n32496), .B(n32497), .Z(n22264) );
  XOR U33675 ( .A(n32498), .B(n32499), .Z(n22259) );
  XOR U33676 ( .A(n32500), .B(n32501), .Z(n22254) );
  XOR U33677 ( .A(n32502), .B(n32503), .Z(n22249) );
  XOR U33678 ( .A(n32504), .B(n32505), .Z(n22244) );
  XOR U33679 ( .A(n32506), .B(n32507), .Z(n22239) );
  XOR U33680 ( .A(n32508), .B(n32509), .Z(n22234) );
  XOR U33681 ( .A(n32510), .B(n32511), .Z(n22229) );
  XOR U33682 ( .A(n32512), .B(n32513), .Z(n22224) );
  XOR U33683 ( .A(n32514), .B(n32515), .Z(n22219) );
  XOR U33684 ( .A(n32516), .B(n32517), .Z(n22214) );
  XOR U33685 ( .A(n32518), .B(n32519), .Z(n22209) );
  XOR U33686 ( .A(n32520), .B(n32521), .Z(n22204) );
  XOR U33687 ( .A(n32522), .B(n32523), .Z(n22199) );
  XOR U33688 ( .A(n32524), .B(n32525), .Z(n22194) );
  XOR U33689 ( .A(n32526), .B(n32527), .Z(n22189) );
  XOR U33690 ( .A(n32528), .B(n32529), .Z(n22184) );
  XOR U33691 ( .A(n32530), .B(n32531), .Z(n22179) );
  XOR U33692 ( .A(n32532), .B(n32533), .Z(n22174) );
  XOR U33693 ( .A(n32534), .B(n32535), .Z(n22169) );
  XOR U33694 ( .A(n32536), .B(n32537), .Z(n22164) );
  XOR U33695 ( .A(n32538), .B(n32539), .Z(n22159) );
  XOR U33696 ( .A(n32540), .B(n32541), .Z(n22154) );
  XOR U33697 ( .A(n32542), .B(n32543), .Z(n22149) );
  XOR U33698 ( .A(n32544), .B(n32545), .Z(n22144) );
  XOR U33699 ( .A(n32546), .B(n32547), .Z(n22139) );
  XOR U33700 ( .A(n32548), .B(n32549), .Z(n22134) );
  XOR U33701 ( .A(n32550), .B(n32551), .Z(n22129) );
  XOR U33702 ( .A(n32552), .B(n32553), .Z(n22124) );
  XOR U33703 ( .A(n32554), .B(n32555), .Z(n22119) );
  XOR U33704 ( .A(n32556), .B(n32557), .Z(n22114) );
  XOR U33705 ( .A(n32558), .B(n32559), .Z(n22109) );
  XOR U33706 ( .A(n32560), .B(n32561), .Z(n22104) );
  XOR U33707 ( .A(n32562), .B(n32563), .Z(n22099) );
  XOR U33708 ( .A(n32564), .B(n32565), .Z(n22094) );
  XOR U33709 ( .A(n32566), .B(n32567), .Z(n22089) );
  XOR U33710 ( .A(n32568), .B(n32569), .Z(n22084) );
  XOR U33711 ( .A(n32570), .B(n32571), .Z(n22079) );
  XOR U33712 ( .A(n32572), .B(n32573), .Z(n22074) );
  XOR U33713 ( .A(n32574), .B(n32575), .Z(n22069) );
  XOR U33714 ( .A(n32576), .B(n32577), .Z(n22064) );
  XOR U33715 ( .A(n32578), .B(n32579), .Z(n22059) );
  XOR U33716 ( .A(n32580), .B(n32581), .Z(n22054) );
  XOR U33717 ( .A(n32582), .B(n32583), .Z(n22049) );
  XOR U33718 ( .A(n32584), .B(n32585), .Z(n22044) );
  XOR U33719 ( .A(n32586), .B(n32587), .Z(n22039) );
  XOR U33720 ( .A(n32588), .B(n32589), .Z(n22034) );
  XOR U33721 ( .A(n32590), .B(n32591), .Z(n22029) );
  XOR U33722 ( .A(n32592), .B(n32593), .Z(n22024) );
  XOR U33723 ( .A(n32594), .B(n32595), .Z(n22019) );
  XOR U33724 ( .A(n32596), .B(n32597), .Z(n22014) );
  XOR U33725 ( .A(n32598), .B(n32599), .Z(n22009) );
  XOR U33726 ( .A(n32600), .B(n32601), .Z(n22004) );
  XOR U33727 ( .A(n32602), .B(n32603), .Z(n21999) );
  XOR U33728 ( .A(n32604), .B(n32605), .Z(n21994) );
  XOR U33729 ( .A(n32606), .B(n32607), .Z(n21989) );
  XOR U33730 ( .A(n32608), .B(n32609), .Z(n21984) );
  XOR U33731 ( .A(n32610), .B(n32611), .Z(n21979) );
  XOR U33732 ( .A(n32612), .B(n32613), .Z(n21974) );
  XOR U33733 ( .A(n32614), .B(n32615), .Z(n21969) );
  XOR U33734 ( .A(n32616), .B(n32617), .Z(n21964) );
  XOR U33735 ( .A(n32618), .B(n32619), .Z(n21959) );
  XOR U33736 ( .A(n32620), .B(n32621), .Z(n21954) );
  XOR U33737 ( .A(n32622), .B(n32623), .Z(n21949) );
  XOR U33738 ( .A(n32624), .B(n32625), .Z(n21944) );
  XOR U33739 ( .A(n32626), .B(n32627), .Z(n21939) );
  XOR U33740 ( .A(n32628), .B(n32629), .Z(n21934) );
  XOR U33741 ( .A(n32630), .B(n32631), .Z(n21929) );
  XOR U33742 ( .A(n32632), .B(n32633), .Z(n21924) );
  XOR U33743 ( .A(n32634), .B(n32635), .Z(n21919) );
  XOR U33744 ( .A(n32636), .B(n32637), .Z(n21914) );
  XOR U33745 ( .A(n32638), .B(n32639), .Z(n21909) );
  XOR U33746 ( .A(n32640), .B(n32641), .Z(n21904) );
  XOR U33747 ( .A(n32642), .B(n32643), .Z(n21899) );
  XOR U33748 ( .A(n32644), .B(n32645), .Z(n21894) );
  XOR U33749 ( .A(n32646), .B(n32647), .Z(n21889) );
  XOR U33750 ( .A(n32648), .B(n32649), .Z(n21884) );
  XOR U33751 ( .A(n32650), .B(n32651), .Z(n21879) );
  XOR U33752 ( .A(n32652), .B(n32653), .Z(n21874) );
  XOR U33753 ( .A(n32654), .B(n32655), .Z(n21869) );
  XOR U33754 ( .A(n32656), .B(n32657), .Z(n21864) );
  XOR U33755 ( .A(n32658), .B(n32659), .Z(n21859) );
  XOR U33756 ( .A(n32660), .B(n32661), .Z(n21854) );
  XOR U33757 ( .A(n32662), .B(n32663), .Z(n21849) );
  XOR U33758 ( .A(n32664), .B(n32665), .Z(n21844) );
  XOR U33759 ( .A(n32666), .B(n32667), .Z(n21839) );
  XOR U33760 ( .A(n32668), .B(n32669), .Z(n21834) );
  XOR U33761 ( .A(n32670), .B(n32671), .Z(n21829) );
  XOR U33762 ( .A(n32672), .B(n32673), .Z(n21824) );
  XOR U33763 ( .A(n32674), .B(n32675), .Z(n21819) );
  XOR U33764 ( .A(n32676), .B(n32677), .Z(n21814) );
  XOR U33765 ( .A(n32678), .B(n32679), .Z(n21809) );
  XOR U33766 ( .A(n32680), .B(n32681), .Z(n21804) );
  XOR U33767 ( .A(n32682), .B(n32683), .Z(n21799) );
  XOR U33768 ( .A(n32684), .B(n32685), .Z(n21794) );
  XOR U33769 ( .A(n32686), .B(n32687), .Z(n21789) );
  XOR U33770 ( .A(n32688), .B(n32689), .Z(n21784) );
  XOR U33771 ( .A(n32690), .B(n32691), .Z(n21779) );
  XOR U33772 ( .A(n32692), .B(n32693), .Z(n21774) );
  XOR U33773 ( .A(n32694), .B(n32695), .Z(n21769) );
  XOR U33774 ( .A(n32696), .B(n32697), .Z(n21764) );
  XOR U33775 ( .A(n32698), .B(n32699), .Z(n21759) );
  XOR U33776 ( .A(n32700), .B(n32701), .Z(n21754) );
  XOR U33777 ( .A(n32702), .B(n32703), .Z(n21749) );
  XOR U33778 ( .A(n32704), .B(n32705), .Z(n21744) );
  XOR U33779 ( .A(n32706), .B(n32707), .Z(n21739) );
  XOR U33780 ( .A(n32708), .B(n32709), .Z(n21734) );
  XOR U33781 ( .A(n32710), .B(n32711), .Z(n21729) );
  XOR U33782 ( .A(n32712), .B(n32713), .Z(n21724) );
  XOR U33783 ( .A(n32714), .B(n32715), .Z(n21719) );
  XOR U33784 ( .A(n32716), .B(n32717), .Z(n21714) );
  XOR U33785 ( .A(n32718), .B(n32719), .Z(n21709) );
  XOR U33786 ( .A(n32720), .B(n32721), .Z(n21704) );
  XOR U33787 ( .A(n32722), .B(n32723), .Z(n21699) );
  XOR U33788 ( .A(n32724), .B(n32725), .Z(n21694) );
  XOR U33789 ( .A(n32726), .B(n32727), .Z(n21689) );
  XOR U33790 ( .A(n32728), .B(n32729), .Z(n21684) );
  XOR U33791 ( .A(n32730), .B(n32731), .Z(n21679) );
  XOR U33792 ( .A(n32732), .B(n32733), .Z(n21674) );
  XOR U33793 ( .A(n32734), .B(n32735), .Z(n21669) );
  XOR U33794 ( .A(n32736), .B(n32737), .Z(n21664) );
  XOR U33795 ( .A(n32738), .B(n32739), .Z(n21659) );
  XOR U33796 ( .A(n32740), .B(n32741), .Z(n21654) );
  XOR U33797 ( .A(n32742), .B(n32743), .Z(n21649) );
  XOR U33798 ( .A(n32744), .B(n32745), .Z(n21644) );
  XOR U33799 ( .A(n32746), .B(n32747), .Z(n21639) );
  XOR U33800 ( .A(n32748), .B(n32749), .Z(n21634) );
  XOR U33801 ( .A(n32750), .B(n32751), .Z(n21629) );
  XOR U33802 ( .A(n32752), .B(n32753), .Z(n21624) );
  XOR U33803 ( .A(n32754), .B(n32755), .Z(n21619) );
  XOR U33804 ( .A(n32756), .B(n32757), .Z(n21614) );
  XOR U33805 ( .A(n32758), .B(n32759), .Z(n21609) );
  XOR U33806 ( .A(n32760), .B(n32761), .Z(n21604) );
  XOR U33807 ( .A(n32762), .B(n32763), .Z(n21599) );
  XOR U33808 ( .A(n32764), .B(n32765), .Z(n21594) );
  XOR U33809 ( .A(n32766), .B(n32767), .Z(n21589) );
  XOR U33810 ( .A(n32768), .B(n32769), .Z(n21584) );
  XOR U33811 ( .A(n32770), .B(n32771), .Z(n21579) );
  XOR U33812 ( .A(n32772), .B(n32773), .Z(n21574) );
  XOR U33813 ( .A(n32774), .B(n32775), .Z(n21569) );
  XOR U33814 ( .A(n32776), .B(n32777), .Z(n21564) );
  XOR U33815 ( .A(n32778), .B(n32779), .Z(n21559) );
  XOR U33816 ( .A(n32780), .B(n32781), .Z(n21554) );
  XOR U33817 ( .A(n32782), .B(n32783), .Z(n21549) );
  XOR U33818 ( .A(n32784), .B(n32785), .Z(n21544) );
  XOR U33819 ( .A(n32786), .B(n32787), .Z(n21539) );
  XOR U33820 ( .A(n32788), .B(n32789), .Z(n21534) );
  XOR U33821 ( .A(n32790), .B(n32791), .Z(n21529) );
  XOR U33822 ( .A(n26649), .B(n26650), .Z(n21524) );
  XOR U33823 ( .A(n32792), .B(n32793), .Z(n26650) );
  ANDN U33824 ( .B(\modmult_1/xin[1023] ), .A(n32793), .Z(n32792) );
  XOR U33825 ( .A(m[1023]), .B(n32794), .Z(n32793) );
  NAND U33826 ( .A(n32795), .B(mul_pow), .Z(n32794) );
  XOR U33827 ( .A(m[1023]), .B(c[1023]), .Z(n32795) );
  XNOR U33828 ( .A(\modmult_1/zin[0][1022] ), .B(n32796), .Z(n26649) );
  IV U33829 ( .A(n26647), .Z(n32796) );
  XOR U33830 ( .A(n32797), .B(n32798), .Z(n26647) );
  ANDN U33831 ( .B(n32799), .A(n32790), .Z(n32797) );
  XNOR U33832 ( .A(\modmult_1/zin[0][1021] ), .B(n32800), .Z(n32790) );
  IV U33833 ( .A(n32798), .Z(n32800) );
  XOR U33834 ( .A(n32798), .B(n32791), .Z(n32799) );
  XNOR U33835 ( .A(n32801), .B(n32802), .Z(n32791) );
  ANDN U33836 ( .B(\modmult_1/xin[1023] ), .A(n32803), .Z(n32801) );
  IV U33837 ( .A(n32802), .Z(n32803) );
  XNOR U33838 ( .A(m[1022]), .B(n32804), .Z(n32802) );
  NAND U33839 ( .A(n32805), .B(mul_pow), .Z(n32804) );
  XOR U33840 ( .A(m[1022]), .B(c[1022]), .Z(n32805) );
  XOR U33841 ( .A(n32806), .B(n32807), .Z(n32798) );
  ANDN U33842 ( .B(n32808), .A(n32788), .Z(n32806) );
  XNOR U33843 ( .A(\modmult_1/zin[0][1020] ), .B(n32809), .Z(n32788) );
  IV U33844 ( .A(n32807), .Z(n32809) );
  XOR U33845 ( .A(n32807), .B(n32789), .Z(n32808) );
  XNOR U33846 ( .A(n32810), .B(n32811), .Z(n32789) );
  ANDN U33847 ( .B(\modmult_1/xin[1023] ), .A(n32812), .Z(n32810) );
  IV U33848 ( .A(n32811), .Z(n32812) );
  XNOR U33849 ( .A(m[1021]), .B(n32813), .Z(n32811) );
  NAND U33850 ( .A(n32814), .B(mul_pow), .Z(n32813) );
  XOR U33851 ( .A(m[1021]), .B(c[1021]), .Z(n32814) );
  XOR U33852 ( .A(n32815), .B(n32816), .Z(n32807) );
  ANDN U33853 ( .B(n32817), .A(n32786), .Z(n32815) );
  XNOR U33854 ( .A(\modmult_1/zin[0][1019] ), .B(n32818), .Z(n32786) );
  IV U33855 ( .A(n32816), .Z(n32818) );
  XOR U33856 ( .A(n32816), .B(n32787), .Z(n32817) );
  XNOR U33857 ( .A(n32819), .B(n32820), .Z(n32787) );
  ANDN U33858 ( .B(\modmult_1/xin[1023] ), .A(n32821), .Z(n32819) );
  IV U33859 ( .A(n32820), .Z(n32821) );
  XNOR U33860 ( .A(m[1020]), .B(n32822), .Z(n32820) );
  NAND U33861 ( .A(n32823), .B(mul_pow), .Z(n32822) );
  XOR U33862 ( .A(m[1020]), .B(c[1020]), .Z(n32823) );
  XOR U33863 ( .A(n32824), .B(n32825), .Z(n32816) );
  ANDN U33864 ( .B(n32826), .A(n32784), .Z(n32824) );
  XNOR U33865 ( .A(\modmult_1/zin[0][1018] ), .B(n32827), .Z(n32784) );
  IV U33866 ( .A(n32825), .Z(n32827) );
  XOR U33867 ( .A(n32825), .B(n32785), .Z(n32826) );
  XNOR U33868 ( .A(n32828), .B(n32829), .Z(n32785) );
  ANDN U33869 ( .B(\modmult_1/xin[1023] ), .A(n32830), .Z(n32828) );
  IV U33870 ( .A(n32829), .Z(n32830) );
  XNOR U33871 ( .A(m[1019]), .B(n32831), .Z(n32829) );
  NAND U33872 ( .A(n32832), .B(mul_pow), .Z(n32831) );
  XOR U33873 ( .A(m[1019]), .B(c[1019]), .Z(n32832) );
  XOR U33874 ( .A(n32833), .B(n32834), .Z(n32825) );
  ANDN U33875 ( .B(n32835), .A(n32782), .Z(n32833) );
  XNOR U33876 ( .A(\modmult_1/zin[0][1017] ), .B(n32836), .Z(n32782) );
  IV U33877 ( .A(n32834), .Z(n32836) );
  XOR U33878 ( .A(n32834), .B(n32783), .Z(n32835) );
  XNOR U33879 ( .A(n32837), .B(n32838), .Z(n32783) );
  ANDN U33880 ( .B(\modmult_1/xin[1023] ), .A(n32839), .Z(n32837) );
  IV U33881 ( .A(n32838), .Z(n32839) );
  XNOR U33882 ( .A(m[1018]), .B(n32840), .Z(n32838) );
  NAND U33883 ( .A(n32841), .B(mul_pow), .Z(n32840) );
  XOR U33884 ( .A(m[1018]), .B(c[1018]), .Z(n32841) );
  XOR U33885 ( .A(n32842), .B(n32843), .Z(n32834) );
  ANDN U33886 ( .B(n32844), .A(n32780), .Z(n32842) );
  XNOR U33887 ( .A(\modmult_1/zin[0][1016] ), .B(n32845), .Z(n32780) );
  IV U33888 ( .A(n32843), .Z(n32845) );
  XOR U33889 ( .A(n32843), .B(n32781), .Z(n32844) );
  XNOR U33890 ( .A(n32846), .B(n32847), .Z(n32781) );
  ANDN U33891 ( .B(\modmult_1/xin[1023] ), .A(n32848), .Z(n32846) );
  IV U33892 ( .A(n32847), .Z(n32848) );
  XNOR U33893 ( .A(m[1017]), .B(n32849), .Z(n32847) );
  NAND U33894 ( .A(n32850), .B(mul_pow), .Z(n32849) );
  XOR U33895 ( .A(m[1017]), .B(c[1017]), .Z(n32850) );
  XOR U33896 ( .A(n32851), .B(n32852), .Z(n32843) );
  ANDN U33897 ( .B(n32853), .A(n32778), .Z(n32851) );
  XNOR U33898 ( .A(\modmult_1/zin[0][1015] ), .B(n32854), .Z(n32778) );
  IV U33899 ( .A(n32852), .Z(n32854) );
  XOR U33900 ( .A(n32852), .B(n32779), .Z(n32853) );
  XNOR U33901 ( .A(n32855), .B(n32856), .Z(n32779) );
  ANDN U33902 ( .B(\modmult_1/xin[1023] ), .A(n32857), .Z(n32855) );
  IV U33903 ( .A(n32856), .Z(n32857) );
  XNOR U33904 ( .A(m[1016]), .B(n32858), .Z(n32856) );
  NAND U33905 ( .A(n32859), .B(mul_pow), .Z(n32858) );
  XOR U33906 ( .A(m[1016]), .B(c[1016]), .Z(n32859) );
  XOR U33907 ( .A(n32860), .B(n32861), .Z(n32852) );
  ANDN U33908 ( .B(n32862), .A(n32776), .Z(n32860) );
  XNOR U33909 ( .A(\modmult_1/zin[0][1014] ), .B(n32863), .Z(n32776) );
  IV U33910 ( .A(n32861), .Z(n32863) );
  XOR U33911 ( .A(n32861), .B(n32777), .Z(n32862) );
  XNOR U33912 ( .A(n32864), .B(n32865), .Z(n32777) );
  ANDN U33913 ( .B(\modmult_1/xin[1023] ), .A(n32866), .Z(n32864) );
  IV U33914 ( .A(n32865), .Z(n32866) );
  XNOR U33915 ( .A(m[1015]), .B(n32867), .Z(n32865) );
  NAND U33916 ( .A(n32868), .B(mul_pow), .Z(n32867) );
  XOR U33917 ( .A(m[1015]), .B(c[1015]), .Z(n32868) );
  XOR U33918 ( .A(n32869), .B(n32870), .Z(n32861) );
  ANDN U33919 ( .B(n32871), .A(n32774), .Z(n32869) );
  XNOR U33920 ( .A(\modmult_1/zin[0][1013] ), .B(n32872), .Z(n32774) );
  IV U33921 ( .A(n32870), .Z(n32872) );
  XOR U33922 ( .A(n32870), .B(n32775), .Z(n32871) );
  XNOR U33923 ( .A(n32873), .B(n32874), .Z(n32775) );
  ANDN U33924 ( .B(\modmult_1/xin[1023] ), .A(n32875), .Z(n32873) );
  IV U33925 ( .A(n32874), .Z(n32875) );
  XNOR U33926 ( .A(m[1014]), .B(n32876), .Z(n32874) );
  NAND U33927 ( .A(n32877), .B(mul_pow), .Z(n32876) );
  XOR U33928 ( .A(m[1014]), .B(c[1014]), .Z(n32877) );
  XOR U33929 ( .A(n32878), .B(n32879), .Z(n32870) );
  ANDN U33930 ( .B(n32880), .A(n32772), .Z(n32878) );
  XNOR U33931 ( .A(\modmult_1/zin[0][1012] ), .B(n32881), .Z(n32772) );
  IV U33932 ( .A(n32879), .Z(n32881) );
  XOR U33933 ( .A(n32879), .B(n32773), .Z(n32880) );
  XNOR U33934 ( .A(n32882), .B(n32883), .Z(n32773) );
  ANDN U33935 ( .B(\modmult_1/xin[1023] ), .A(n32884), .Z(n32882) );
  IV U33936 ( .A(n32883), .Z(n32884) );
  XNOR U33937 ( .A(m[1013]), .B(n32885), .Z(n32883) );
  NAND U33938 ( .A(n32886), .B(mul_pow), .Z(n32885) );
  XOR U33939 ( .A(m[1013]), .B(c[1013]), .Z(n32886) );
  XOR U33940 ( .A(n32887), .B(n32888), .Z(n32879) );
  ANDN U33941 ( .B(n32889), .A(n32770), .Z(n32887) );
  XNOR U33942 ( .A(\modmult_1/zin[0][1011] ), .B(n32890), .Z(n32770) );
  IV U33943 ( .A(n32888), .Z(n32890) );
  XOR U33944 ( .A(n32888), .B(n32771), .Z(n32889) );
  XNOR U33945 ( .A(n32891), .B(n32892), .Z(n32771) );
  ANDN U33946 ( .B(\modmult_1/xin[1023] ), .A(n32893), .Z(n32891) );
  IV U33947 ( .A(n32892), .Z(n32893) );
  XNOR U33948 ( .A(m[1012]), .B(n32894), .Z(n32892) );
  NAND U33949 ( .A(n32895), .B(mul_pow), .Z(n32894) );
  XOR U33950 ( .A(m[1012]), .B(c[1012]), .Z(n32895) );
  XOR U33951 ( .A(n32896), .B(n32897), .Z(n32888) );
  ANDN U33952 ( .B(n32898), .A(n32768), .Z(n32896) );
  XNOR U33953 ( .A(\modmult_1/zin[0][1010] ), .B(n32899), .Z(n32768) );
  IV U33954 ( .A(n32897), .Z(n32899) );
  XOR U33955 ( .A(n32897), .B(n32769), .Z(n32898) );
  XNOR U33956 ( .A(n32900), .B(n32901), .Z(n32769) );
  ANDN U33957 ( .B(\modmult_1/xin[1023] ), .A(n32902), .Z(n32900) );
  IV U33958 ( .A(n32901), .Z(n32902) );
  XNOR U33959 ( .A(m[1011]), .B(n32903), .Z(n32901) );
  NAND U33960 ( .A(n32904), .B(mul_pow), .Z(n32903) );
  XOR U33961 ( .A(m[1011]), .B(c[1011]), .Z(n32904) );
  XOR U33962 ( .A(n32905), .B(n32906), .Z(n32897) );
  ANDN U33963 ( .B(n32907), .A(n32766), .Z(n32905) );
  XNOR U33964 ( .A(\modmult_1/zin[0][1009] ), .B(n32908), .Z(n32766) );
  IV U33965 ( .A(n32906), .Z(n32908) );
  XOR U33966 ( .A(n32906), .B(n32767), .Z(n32907) );
  XNOR U33967 ( .A(n32909), .B(n32910), .Z(n32767) );
  ANDN U33968 ( .B(\modmult_1/xin[1023] ), .A(n32911), .Z(n32909) );
  IV U33969 ( .A(n32910), .Z(n32911) );
  XNOR U33970 ( .A(m[1010]), .B(n32912), .Z(n32910) );
  NAND U33971 ( .A(n32913), .B(mul_pow), .Z(n32912) );
  XOR U33972 ( .A(m[1010]), .B(c[1010]), .Z(n32913) );
  XOR U33973 ( .A(n32914), .B(n32915), .Z(n32906) );
  ANDN U33974 ( .B(n32916), .A(n32764), .Z(n32914) );
  XNOR U33975 ( .A(\modmult_1/zin[0][1008] ), .B(n32917), .Z(n32764) );
  IV U33976 ( .A(n32915), .Z(n32917) );
  XOR U33977 ( .A(n32915), .B(n32765), .Z(n32916) );
  XNOR U33978 ( .A(n32918), .B(n32919), .Z(n32765) );
  ANDN U33979 ( .B(\modmult_1/xin[1023] ), .A(n32920), .Z(n32918) );
  IV U33980 ( .A(n32919), .Z(n32920) );
  XNOR U33981 ( .A(m[1009]), .B(n32921), .Z(n32919) );
  NAND U33982 ( .A(n32922), .B(mul_pow), .Z(n32921) );
  XOR U33983 ( .A(m[1009]), .B(c[1009]), .Z(n32922) );
  XOR U33984 ( .A(n32923), .B(n32924), .Z(n32915) );
  ANDN U33985 ( .B(n32925), .A(n32762), .Z(n32923) );
  XNOR U33986 ( .A(\modmult_1/zin[0][1007] ), .B(n32926), .Z(n32762) );
  IV U33987 ( .A(n32924), .Z(n32926) );
  XOR U33988 ( .A(n32924), .B(n32763), .Z(n32925) );
  XNOR U33989 ( .A(n32927), .B(n32928), .Z(n32763) );
  ANDN U33990 ( .B(\modmult_1/xin[1023] ), .A(n32929), .Z(n32927) );
  IV U33991 ( .A(n32928), .Z(n32929) );
  XNOR U33992 ( .A(m[1008]), .B(n32930), .Z(n32928) );
  NAND U33993 ( .A(n32931), .B(mul_pow), .Z(n32930) );
  XOR U33994 ( .A(m[1008]), .B(c[1008]), .Z(n32931) );
  XOR U33995 ( .A(n32932), .B(n32933), .Z(n32924) );
  ANDN U33996 ( .B(n32934), .A(n32760), .Z(n32932) );
  XNOR U33997 ( .A(\modmult_1/zin[0][1006] ), .B(n32935), .Z(n32760) );
  IV U33998 ( .A(n32933), .Z(n32935) );
  XOR U33999 ( .A(n32933), .B(n32761), .Z(n32934) );
  XNOR U34000 ( .A(n32936), .B(n32937), .Z(n32761) );
  ANDN U34001 ( .B(\modmult_1/xin[1023] ), .A(n32938), .Z(n32936) );
  IV U34002 ( .A(n32937), .Z(n32938) );
  XNOR U34003 ( .A(m[1007]), .B(n32939), .Z(n32937) );
  NAND U34004 ( .A(n32940), .B(mul_pow), .Z(n32939) );
  XOR U34005 ( .A(m[1007]), .B(c[1007]), .Z(n32940) );
  XOR U34006 ( .A(n32941), .B(n32942), .Z(n32933) );
  ANDN U34007 ( .B(n32943), .A(n32758), .Z(n32941) );
  XNOR U34008 ( .A(\modmult_1/zin[0][1005] ), .B(n32944), .Z(n32758) );
  IV U34009 ( .A(n32942), .Z(n32944) );
  XOR U34010 ( .A(n32942), .B(n32759), .Z(n32943) );
  XNOR U34011 ( .A(n32945), .B(n32946), .Z(n32759) );
  ANDN U34012 ( .B(\modmult_1/xin[1023] ), .A(n32947), .Z(n32945) );
  IV U34013 ( .A(n32946), .Z(n32947) );
  XNOR U34014 ( .A(m[1006]), .B(n32948), .Z(n32946) );
  NAND U34015 ( .A(n32949), .B(mul_pow), .Z(n32948) );
  XOR U34016 ( .A(m[1006]), .B(c[1006]), .Z(n32949) );
  XOR U34017 ( .A(n32950), .B(n32951), .Z(n32942) );
  ANDN U34018 ( .B(n32952), .A(n32756), .Z(n32950) );
  XNOR U34019 ( .A(\modmult_1/zin[0][1004] ), .B(n32953), .Z(n32756) );
  IV U34020 ( .A(n32951), .Z(n32953) );
  XOR U34021 ( .A(n32951), .B(n32757), .Z(n32952) );
  XNOR U34022 ( .A(n32954), .B(n32955), .Z(n32757) );
  ANDN U34023 ( .B(\modmult_1/xin[1023] ), .A(n32956), .Z(n32954) );
  IV U34024 ( .A(n32955), .Z(n32956) );
  XNOR U34025 ( .A(m[1005]), .B(n32957), .Z(n32955) );
  NAND U34026 ( .A(n32958), .B(mul_pow), .Z(n32957) );
  XOR U34027 ( .A(m[1005]), .B(c[1005]), .Z(n32958) );
  XOR U34028 ( .A(n32959), .B(n32960), .Z(n32951) );
  ANDN U34029 ( .B(n32961), .A(n32754), .Z(n32959) );
  XNOR U34030 ( .A(\modmult_1/zin[0][1003] ), .B(n32962), .Z(n32754) );
  IV U34031 ( .A(n32960), .Z(n32962) );
  XOR U34032 ( .A(n32960), .B(n32755), .Z(n32961) );
  XNOR U34033 ( .A(n32963), .B(n32964), .Z(n32755) );
  ANDN U34034 ( .B(\modmult_1/xin[1023] ), .A(n32965), .Z(n32963) );
  IV U34035 ( .A(n32964), .Z(n32965) );
  XNOR U34036 ( .A(m[1004]), .B(n32966), .Z(n32964) );
  NAND U34037 ( .A(n32967), .B(mul_pow), .Z(n32966) );
  XOR U34038 ( .A(m[1004]), .B(c[1004]), .Z(n32967) );
  XOR U34039 ( .A(n32968), .B(n32969), .Z(n32960) );
  ANDN U34040 ( .B(n32970), .A(n32752), .Z(n32968) );
  XNOR U34041 ( .A(\modmult_1/zin[0][1002] ), .B(n32971), .Z(n32752) );
  IV U34042 ( .A(n32969), .Z(n32971) );
  XOR U34043 ( .A(n32969), .B(n32753), .Z(n32970) );
  XNOR U34044 ( .A(n32972), .B(n32973), .Z(n32753) );
  ANDN U34045 ( .B(\modmult_1/xin[1023] ), .A(n32974), .Z(n32972) );
  IV U34046 ( .A(n32973), .Z(n32974) );
  XNOR U34047 ( .A(m[1003]), .B(n32975), .Z(n32973) );
  NAND U34048 ( .A(n32976), .B(mul_pow), .Z(n32975) );
  XOR U34049 ( .A(m[1003]), .B(c[1003]), .Z(n32976) );
  XOR U34050 ( .A(n32977), .B(n32978), .Z(n32969) );
  ANDN U34051 ( .B(n32979), .A(n32750), .Z(n32977) );
  XNOR U34052 ( .A(\modmult_1/zin[0][1001] ), .B(n32980), .Z(n32750) );
  IV U34053 ( .A(n32978), .Z(n32980) );
  XOR U34054 ( .A(n32978), .B(n32751), .Z(n32979) );
  XNOR U34055 ( .A(n32981), .B(n32982), .Z(n32751) );
  ANDN U34056 ( .B(\modmult_1/xin[1023] ), .A(n32983), .Z(n32981) );
  IV U34057 ( .A(n32982), .Z(n32983) );
  XNOR U34058 ( .A(m[1002]), .B(n32984), .Z(n32982) );
  NAND U34059 ( .A(n32985), .B(mul_pow), .Z(n32984) );
  XOR U34060 ( .A(m[1002]), .B(c[1002]), .Z(n32985) );
  XOR U34061 ( .A(n32986), .B(n32987), .Z(n32978) );
  ANDN U34062 ( .B(n32988), .A(n32748), .Z(n32986) );
  XNOR U34063 ( .A(\modmult_1/zin[0][1000] ), .B(n32989), .Z(n32748) );
  IV U34064 ( .A(n32987), .Z(n32989) );
  XOR U34065 ( .A(n32987), .B(n32749), .Z(n32988) );
  XNOR U34066 ( .A(n32990), .B(n32991), .Z(n32749) );
  ANDN U34067 ( .B(\modmult_1/xin[1023] ), .A(n32992), .Z(n32990) );
  IV U34068 ( .A(n32991), .Z(n32992) );
  XNOR U34069 ( .A(m[1001]), .B(n32993), .Z(n32991) );
  NAND U34070 ( .A(n32994), .B(mul_pow), .Z(n32993) );
  XOR U34071 ( .A(m[1001]), .B(c[1001]), .Z(n32994) );
  XOR U34072 ( .A(n32995), .B(n32996), .Z(n32987) );
  ANDN U34073 ( .B(n32997), .A(n32746), .Z(n32995) );
  XNOR U34074 ( .A(\modmult_1/zin[0][999] ), .B(n32998), .Z(n32746) );
  IV U34075 ( .A(n32996), .Z(n32998) );
  XOR U34076 ( .A(n32996), .B(n32747), .Z(n32997) );
  XNOR U34077 ( .A(n32999), .B(n33000), .Z(n32747) );
  ANDN U34078 ( .B(\modmult_1/xin[1023] ), .A(n33001), .Z(n32999) );
  IV U34079 ( .A(n33000), .Z(n33001) );
  XNOR U34080 ( .A(m[1000]), .B(n33002), .Z(n33000) );
  NAND U34081 ( .A(n33003), .B(mul_pow), .Z(n33002) );
  XOR U34082 ( .A(m[1000]), .B(c[1000]), .Z(n33003) );
  XOR U34083 ( .A(n33004), .B(n33005), .Z(n32996) );
  ANDN U34084 ( .B(n33006), .A(n32744), .Z(n33004) );
  XNOR U34085 ( .A(\modmult_1/zin[0][998] ), .B(n33007), .Z(n32744) );
  IV U34086 ( .A(n33005), .Z(n33007) );
  XOR U34087 ( .A(n33005), .B(n32745), .Z(n33006) );
  XNOR U34088 ( .A(n33008), .B(n33009), .Z(n32745) );
  ANDN U34089 ( .B(\modmult_1/xin[1023] ), .A(n33010), .Z(n33008) );
  IV U34090 ( .A(n33009), .Z(n33010) );
  XNOR U34091 ( .A(m[999]), .B(n33011), .Z(n33009) );
  NAND U34092 ( .A(n33012), .B(mul_pow), .Z(n33011) );
  XOR U34093 ( .A(m[999]), .B(c[999]), .Z(n33012) );
  XOR U34094 ( .A(n33013), .B(n33014), .Z(n33005) );
  ANDN U34095 ( .B(n33015), .A(n32742), .Z(n33013) );
  XNOR U34096 ( .A(\modmult_1/zin[0][997] ), .B(n33016), .Z(n32742) );
  IV U34097 ( .A(n33014), .Z(n33016) );
  XOR U34098 ( .A(n33014), .B(n32743), .Z(n33015) );
  XNOR U34099 ( .A(n33017), .B(n33018), .Z(n32743) );
  ANDN U34100 ( .B(\modmult_1/xin[1023] ), .A(n33019), .Z(n33017) );
  IV U34101 ( .A(n33018), .Z(n33019) );
  XNOR U34102 ( .A(m[998]), .B(n33020), .Z(n33018) );
  NAND U34103 ( .A(n33021), .B(mul_pow), .Z(n33020) );
  XOR U34104 ( .A(m[998]), .B(c[998]), .Z(n33021) );
  XOR U34105 ( .A(n33022), .B(n33023), .Z(n33014) );
  ANDN U34106 ( .B(n33024), .A(n32740), .Z(n33022) );
  XNOR U34107 ( .A(\modmult_1/zin[0][996] ), .B(n33025), .Z(n32740) );
  IV U34108 ( .A(n33023), .Z(n33025) );
  XOR U34109 ( .A(n33023), .B(n32741), .Z(n33024) );
  XNOR U34110 ( .A(n33026), .B(n33027), .Z(n32741) );
  ANDN U34111 ( .B(\modmult_1/xin[1023] ), .A(n33028), .Z(n33026) );
  IV U34112 ( .A(n33027), .Z(n33028) );
  XNOR U34113 ( .A(m[997]), .B(n33029), .Z(n33027) );
  NAND U34114 ( .A(n33030), .B(mul_pow), .Z(n33029) );
  XOR U34115 ( .A(m[997]), .B(c[997]), .Z(n33030) );
  XOR U34116 ( .A(n33031), .B(n33032), .Z(n33023) );
  ANDN U34117 ( .B(n33033), .A(n32738), .Z(n33031) );
  XNOR U34118 ( .A(\modmult_1/zin[0][995] ), .B(n33034), .Z(n32738) );
  IV U34119 ( .A(n33032), .Z(n33034) );
  XOR U34120 ( .A(n33032), .B(n32739), .Z(n33033) );
  XNOR U34121 ( .A(n33035), .B(n33036), .Z(n32739) );
  ANDN U34122 ( .B(\modmult_1/xin[1023] ), .A(n33037), .Z(n33035) );
  IV U34123 ( .A(n33036), .Z(n33037) );
  XNOR U34124 ( .A(m[996]), .B(n33038), .Z(n33036) );
  NAND U34125 ( .A(n33039), .B(mul_pow), .Z(n33038) );
  XOR U34126 ( .A(m[996]), .B(c[996]), .Z(n33039) );
  XOR U34127 ( .A(n33040), .B(n33041), .Z(n33032) );
  ANDN U34128 ( .B(n33042), .A(n32736), .Z(n33040) );
  XNOR U34129 ( .A(\modmult_1/zin[0][994] ), .B(n33043), .Z(n32736) );
  IV U34130 ( .A(n33041), .Z(n33043) );
  XOR U34131 ( .A(n33041), .B(n32737), .Z(n33042) );
  XNOR U34132 ( .A(n33044), .B(n33045), .Z(n32737) );
  ANDN U34133 ( .B(\modmult_1/xin[1023] ), .A(n33046), .Z(n33044) );
  IV U34134 ( .A(n33045), .Z(n33046) );
  XNOR U34135 ( .A(m[995]), .B(n33047), .Z(n33045) );
  NAND U34136 ( .A(n33048), .B(mul_pow), .Z(n33047) );
  XOR U34137 ( .A(m[995]), .B(c[995]), .Z(n33048) );
  XOR U34138 ( .A(n33049), .B(n33050), .Z(n33041) );
  ANDN U34139 ( .B(n33051), .A(n32734), .Z(n33049) );
  XNOR U34140 ( .A(\modmult_1/zin[0][993] ), .B(n33052), .Z(n32734) );
  IV U34141 ( .A(n33050), .Z(n33052) );
  XOR U34142 ( .A(n33050), .B(n32735), .Z(n33051) );
  XNOR U34143 ( .A(n33053), .B(n33054), .Z(n32735) );
  ANDN U34144 ( .B(\modmult_1/xin[1023] ), .A(n33055), .Z(n33053) );
  IV U34145 ( .A(n33054), .Z(n33055) );
  XNOR U34146 ( .A(m[994]), .B(n33056), .Z(n33054) );
  NAND U34147 ( .A(n33057), .B(mul_pow), .Z(n33056) );
  XOR U34148 ( .A(m[994]), .B(c[994]), .Z(n33057) );
  XOR U34149 ( .A(n33058), .B(n33059), .Z(n33050) );
  ANDN U34150 ( .B(n33060), .A(n32732), .Z(n33058) );
  XNOR U34151 ( .A(\modmult_1/zin[0][992] ), .B(n33061), .Z(n32732) );
  IV U34152 ( .A(n33059), .Z(n33061) );
  XOR U34153 ( .A(n33059), .B(n32733), .Z(n33060) );
  XNOR U34154 ( .A(n33062), .B(n33063), .Z(n32733) );
  ANDN U34155 ( .B(\modmult_1/xin[1023] ), .A(n33064), .Z(n33062) );
  IV U34156 ( .A(n33063), .Z(n33064) );
  XNOR U34157 ( .A(m[993]), .B(n33065), .Z(n33063) );
  NAND U34158 ( .A(n33066), .B(mul_pow), .Z(n33065) );
  XOR U34159 ( .A(m[993]), .B(c[993]), .Z(n33066) );
  XOR U34160 ( .A(n33067), .B(n33068), .Z(n33059) );
  ANDN U34161 ( .B(n33069), .A(n32730), .Z(n33067) );
  XNOR U34162 ( .A(\modmult_1/zin[0][991] ), .B(n33070), .Z(n32730) );
  IV U34163 ( .A(n33068), .Z(n33070) );
  XOR U34164 ( .A(n33068), .B(n32731), .Z(n33069) );
  XNOR U34165 ( .A(n33071), .B(n33072), .Z(n32731) );
  ANDN U34166 ( .B(\modmult_1/xin[1023] ), .A(n33073), .Z(n33071) );
  IV U34167 ( .A(n33072), .Z(n33073) );
  XNOR U34168 ( .A(m[992]), .B(n33074), .Z(n33072) );
  NAND U34169 ( .A(n33075), .B(mul_pow), .Z(n33074) );
  XOR U34170 ( .A(m[992]), .B(c[992]), .Z(n33075) );
  XOR U34171 ( .A(n33076), .B(n33077), .Z(n33068) );
  ANDN U34172 ( .B(n33078), .A(n32728), .Z(n33076) );
  XNOR U34173 ( .A(\modmult_1/zin[0][990] ), .B(n33079), .Z(n32728) );
  IV U34174 ( .A(n33077), .Z(n33079) );
  XOR U34175 ( .A(n33077), .B(n32729), .Z(n33078) );
  XNOR U34176 ( .A(n33080), .B(n33081), .Z(n32729) );
  ANDN U34177 ( .B(\modmult_1/xin[1023] ), .A(n33082), .Z(n33080) );
  IV U34178 ( .A(n33081), .Z(n33082) );
  XNOR U34179 ( .A(m[991]), .B(n33083), .Z(n33081) );
  NAND U34180 ( .A(n33084), .B(mul_pow), .Z(n33083) );
  XOR U34181 ( .A(m[991]), .B(c[991]), .Z(n33084) );
  XOR U34182 ( .A(n33085), .B(n33086), .Z(n33077) );
  ANDN U34183 ( .B(n33087), .A(n32726), .Z(n33085) );
  XNOR U34184 ( .A(\modmult_1/zin[0][989] ), .B(n33088), .Z(n32726) );
  IV U34185 ( .A(n33086), .Z(n33088) );
  XOR U34186 ( .A(n33086), .B(n32727), .Z(n33087) );
  XNOR U34187 ( .A(n33089), .B(n33090), .Z(n32727) );
  ANDN U34188 ( .B(\modmult_1/xin[1023] ), .A(n33091), .Z(n33089) );
  IV U34189 ( .A(n33090), .Z(n33091) );
  XNOR U34190 ( .A(m[990]), .B(n33092), .Z(n33090) );
  NAND U34191 ( .A(n33093), .B(mul_pow), .Z(n33092) );
  XOR U34192 ( .A(m[990]), .B(c[990]), .Z(n33093) );
  XOR U34193 ( .A(n33094), .B(n33095), .Z(n33086) );
  ANDN U34194 ( .B(n33096), .A(n32724), .Z(n33094) );
  XNOR U34195 ( .A(\modmult_1/zin[0][988] ), .B(n33097), .Z(n32724) );
  IV U34196 ( .A(n33095), .Z(n33097) );
  XOR U34197 ( .A(n33095), .B(n32725), .Z(n33096) );
  XNOR U34198 ( .A(n33098), .B(n33099), .Z(n32725) );
  ANDN U34199 ( .B(\modmult_1/xin[1023] ), .A(n33100), .Z(n33098) );
  IV U34200 ( .A(n33099), .Z(n33100) );
  XNOR U34201 ( .A(m[989]), .B(n33101), .Z(n33099) );
  NAND U34202 ( .A(n33102), .B(mul_pow), .Z(n33101) );
  XOR U34203 ( .A(m[989]), .B(c[989]), .Z(n33102) );
  XOR U34204 ( .A(n33103), .B(n33104), .Z(n33095) );
  ANDN U34205 ( .B(n33105), .A(n32722), .Z(n33103) );
  XNOR U34206 ( .A(\modmult_1/zin[0][987] ), .B(n33106), .Z(n32722) );
  IV U34207 ( .A(n33104), .Z(n33106) );
  XOR U34208 ( .A(n33104), .B(n32723), .Z(n33105) );
  XNOR U34209 ( .A(n33107), .B(n33108), .Z(n32723) );
  ANDN U34210 ( .B(\modmult_1/xin[1023] ), .A(n33109), .Z(n33107) );
  IV U34211 ( .A(n33108), .Z(n33109) );
  XNOR U34212 ( .A(m[988]), .B(n33110), .Z(n33108) );
  NAND U34213 ( .A(n33111), .B(mul_pow), .Z(n33110) );
  XOR U34214 ( .A(m[988]), .B(c[988]), .Z(n33111) );
  XOR U34215 ( .A(n33112), .B(n33113), .Z(n33104) );
  ANDN U34216 ( .B(n33114), .A(n32720), .Z(n33112) );
  XNOR U34217 ( .A(\modmult_1/zin[0][986] ), .B(n33115), .Z(n32720) );
  IV U34218 ( .A(n33113), .Z(n33115) );
  XOR U34219 ( .A(n33113), .B(n32721), .Z(n33114) );
  XNOR U34220 ( .A(n33116), .B(n33117), .Z(n32721) );
  ANDN U34221 ( .B(\modmult_1/xin[1023] ), .A(n33118), .Z(n33116) );
  IV U34222 ( .A(n33117), .Z(n33118) );
  XNOR U34223 ( .A(m[987]), .B(n33119), .Z(n33117) );
  NAND U34224 ( .A(n33120), .B(mul_pow), .Z(n33119) );
  XOR U34225 ( .A(m[987]), .B(c[987]), .Z(n33120) );
  XOR U34226 ( .A(n33121), .B(n33122), .Z(n33113) );
  ANDN U34227 ( .B(n33123), .A(n32718), .Z(n33121) );
  XNOR U34228 ( .A(\modmult_1/zin[0][985] ), .B(n33124), .Z(n32718) );
  IV U34229 ( .A(n33122), .Z(n33124) );
  XOR U34230 ( .A(n33122), .B(n32719), .Z(n33123) );
  XNOR U34231 ( .A(n33125), .B(n33126), .Z(n32719) );
  ANDN U34232 ( .B(\modmult_1/xin[1023] ), .A(n33127), .Z(n33125) );
  IV U34233 ( .A(n33126), .Z(n33127) );
  XNOR U34234 ( .A(m[986]), .B(n33128), .Z(n33126) );
  NAND U34235 ( .A(n33129), .B(mul_pow), .Z(n33128) );
  XOR U34236 ( .A(m[986]), .B(c[986]), .Z(n33129) );
  XOR U34237 ( .A(n33130), .B(n33131), .Z(n33122) );
  ANDN U34238 ( .B(n33132), .A(n32716), .Z(n33130) );
  XNOR U34239 ( .A(\modmult_1/zin[0][984] ), .B(n33133), .Z(n32716) );
  IV U34240 ( .A(n33131), .Z(n33133) );
  XOR U34241 ( .A(n33131), .B(n32717), .Z(n33132) );
  XNOR U34242 ( .A(n33134), .B(n33135), .Z(n32717) );
  ANDN U34243 ( .B(\modmult_1/xin[1023] ), .A(n33136), .Z(n33134) );
  IV U34244 ( .A(n33135), .Z(n33136) );
  XNOR U34245 ( .A(m[985]), .B(n33137), .Z(n33135) );
  NAND U34246 ( .A(n33138), .B(mul_pow), .Z(n33137) );
  XOR U34247 ( .A(m[985]), .B(c[985]), .Z(n33138) );
  XOR U34248 ( .A(n33139), .B(n33140), .Z(n33131) );
  ANDN U34249 ( .B(n33141), .A(n32714), .Z(n33139) );
  XNOR U34250 ( .A(\modmult_1/zin[0][983] ), .B(n33142), .Z(n32714) );
  IV U34251 ( .A(n33140), .Z(n33142) );
  XOR U34252 ( .A(n33140), .B(n32715), .Z(n33141) );
  XNOR U34253 ( .A(n33143), .B(n33144), .Z(n32715) );
  ANDN U34254 ( .B(\modmult_1/xin[1023] ), .A(n33145), .Z(n33143) );
  IV U34255 ( .A(n33144), .Z(n33145) );
  XNOR U34256 ( .A(m[984]), .B(n33146), .Z(n33144) );
  NAND U34257 ( .A(n33147), .B(mul_pow), .Z(n33146) );
  XOR U34258 ( .A(m[984]), .B(c[984]), .Z(n33147) );
  XOR U34259 ( .A(n33148), .B(n33149), .Z(n33140) );
  ANDN U34260 ( .B(n33150), .A(n32712), .Z(n33148) );
  XNOR U34261 ( .A(\modmult_1/zin[0][982] ), .B(n33151), .Z(n32712) );
  IV U34262 ( .A(n33149), .Z(n33151) );
  XOR U34263 ( .A(n33149), .B(n32713), .Z(n33150) );
  XNOR U34264 ( .A(n33152), .B(n33153), .Z(n32713) );
  ANDN U34265 ( .B(\modmult_1/xin[1023] ), .A(n33154), .Z(n33152) );
  IV U34266 ( .A(n33153), .Z(n33154) );
  XNOR U34267 ( .A(m[983]), .B(n33155), .Z(n33153) );
  NAND U34268 ( .A(n33156), .B(mul_pow), .Z(n33155) );
  XOR U34269 ( .A(m[983]), .B(c[983]), .Z(n33156) );
  XOR U34270 ( .A(n33157), .B(n33158), .Z(n33149) );
  ANDN U34271 ( .B(n33159), .A(n32710), .Z(n33157) );
  XNOR U34272 ( .A(\modmult_1/zin[0][981] ), .B(n33160), .Z(n32710) );
  IV U34273 ( .A(n33158), .Z(n33160) );
  XOR U34274 ( .A(n33158), .B(n32711), .Z(n33159) );
  XNOR U34275 ( .A(n33161), .B(n33162), .Z(n32711) );
  ANDN U34276 ( .B(\modmult_1/xin[1023] ), .A(n33163), .Z(n33161) );
  IV U34277 ( .A(n33162), .Z(n33163) );
  XNOR U34278 ( .A(m[982]), .B(n33164), .Z(n33162) );
  NAND U34279 ( .A(n33165), .B(mul_pow), .Z(n33164) );
  XOR U34280 ( .A(m[982]), .B(c[982]), .Z(n33165) );
  XOR U34281 ( .A(n33166), .B(n33167), .Z(n33158) );
  ANDN U34282 ( .B(n33168), .A(n32708), .Z(n33166) );
  XNOR U34283 ( .A(\modmult_1/zin[0][980] ), .B(n33169), .Z(n32708) );
  IV U34284 ( .A(n33167), .Z(n33169) );
  XOR U34285 ( .A(n33167), .B(n32709), .Z(n33168) );
  XNOR U34286 ( .A(n33170), .B(n33171), .Z(n32709) );
  ANDN U34287 ( .B(\modmult_1/xin[1023] ), .A(n33172), .Z(n33170) );
  IV U34288 ( .A(n33171), .Z(n33172) );
  XNOR U34289 ( .A(m[981]), .B(n33173), .Z(n33171) );
  NAND U34290 ( .A(n33174), .B(mul_pow), .Z(n33173) );
  XOR U34291 ( .A(m[981]), .B(c[981]), .Z(n33174) );
  XOR U34292 ( .A(n33175), .B(n33176), .Z(n33167) );
  ANDN U34293 ( .B(n33177), .A(n32706), .Z(n33175) );
  XNOR U34294 ( .A(\modmult_1/zin[0][979] ), .B(n33178), .Z(n32706) );
  IV U34295 ( .A(n33176), .Z(n33178) );
  XOR U34296 ( .A(n33176), .B(n32707), .Z(n33177) );
  XNOR U34297 ( .A(n33179), .B(n33180), .Z(n32707) );
  ANDN U34298 ( .B(\modmult_1/xin[1023] ), .A(n33181), .Z(n33179) );
  IV U34299 ( .A(n33180), .Z(n33181) );
  XNOR U34300 ( .A(m[980]), .B(n33182), .Z(n33180) );
  NAND U34301 ( .A(n33183), .B(mul_pow), .Z(n33182) );
  XOR U34302 ( .A(m[980]), .B(c[980]), .Z(n33183) );
  XOR U34303 ( .A(n33184), .B(n33185), .Z(n33176) );
  ANDN U34304 ( .B(n33186), .A(n32704), .Z(n33184) );
  XNOR U34305 ( .A(\modmult_1/zin[0][978] ), .B(n33187), .Z(n32704) );
  IV U34306 ( .A(n33185), .Z(n33187) );
  XOR U34307 ( .A(n33185), .B(n32705), .Z(n33186) );
  XNOR U34308 ( .A(n33188), .B(n33189), .Z(n32705) );
  ANDN U34309 ( .B(\modmult_1/xin[1023] ), .A(n33190), .Z(n33188) );
  IV U34310 ( .A(n33189), .Z(n33190) );
  XNOR U34311 ( .A(m[979]), .B(n33191), .Z(n33189) );
  NAND U34312 ( .A(n33192), .B(mul_pow), .Z(n33191) );
  XOR U34313 ( .A(m[979]), .B(c[979]), .Z(n33192) );
  XOR U34314 ( .A(n33193), .B(n33194), .Z(n33185) );
  ANDN U34315 ( .B(n33195), .A(n32702), .Z(n33193) );
  XNOR U34316 ( .A(\modmult_1/zin[0][977] ), .B(n33196), .Z(n32702) );
  IV U34317 ( .A(n33194), .Z(n33196) );
  XOR U34318 ( .A(n33194), .B(n32703), .Z(n33195) );
  XNOR U34319 ( .A(n33197), .B(n33198), .Z(n32703) );
  ANDN U34320 ( .B(\modmult_1/xin[1023] ), .A(n33199), .Z(n33197) );
  IV U34321 ( .A(n33198), .Z(n33199) );
  XNOR U34322 ( .A(m[978]), .B(n33200), .Z(n33198) );
  NAND U34323 ( .A(n33201), .B(mul_pow), .Z(n33200) );
  XOR U34324 ( .A(m[978]), .B(c[978]), .Z(n33201) );
  XOR U34325 ( .A(n33202), .B(n33203), .Z(n33194) );
  ANDN U34326 ( .B(n33204), .A(n32700), .Z(n33202) );
  XNOR U34327 ( .A(\modmult_1/zin[0][976] ), .B(n33205), .Z(n32700) );
  IV U34328 ( .A(n33203), .Z(n33205) );
  XOR U34329 ( .A(n33203), .B(n32701), .Z(n33204) );
  XNOR U34330 ( .A(n33206), .B(n33207), .Z(n32701) );
  ANDN U34331 ( .B(\modmult_1/xin[1023] ), .A(n33208), .Z(n33206) );
  IV U34332 ( .A(n33207), .Z(n33208) );
  XNOR U34333 ( .A(m[977]), .B(n33209), .Z(n33207) );
  NAND U34334 ( .A(n33210), .B(mul_pow), .Z(n33209) );
  XOR U34335 ( .A(m[977]), .B(c[977]), .Z(n33210) );
  XOR U34336 ( .A(n33211), .B(n33212), .Z(n33203) );
  ANDN U34337 ( .B(n33213), .A(n32698), .Z(n33211) );
  XNOR U34338 ( .A(\modmult_1/zin[0][975] ), .B(n33214), .Z(n32698) );
  IV U34339 ( .A(n33212), .Z(n33214) );
  XOR U34340 ( .A(n33212), .B(n32699), .Z(n33213) );
  XNOR U34341 ( .A(n33215), .B(n33216), .Z(n32699) );
  ANDN U34342 ( .B(\modmult_1/xin[1023] ), .A(n33217), .Z(n33215) );
  IV U34343 ( .A(n33216), .Z(n33217) );
  XNOR U34344 ( .A(m[976]), .B(n33218), .Z(n33216) );
  NAND U34345 ( .A(n33219), .B(mul_pow), .Z(n33218) );
  XOR U34346 ( .A(m[976]), .B(c[976]), .Z(n33219) );
  XOR U34347 ( .A(n33220), .B(n33221), .Z(n33212) );
  ANDN U34348 ( .B(n33222), .A(n32696), .Z(n33220) );
  XNOR U34349 ( .A(\modmult_1/zin[0][974] ), .B(n33223), .Z(n32696) );
  IV U34350 ( .A(n33221), .Z(n33223) );
  XOR U34351 ( .A(n33221), .B(n32697), .Z(n33222) );
  XNOR U34352 ( .A(n33224), .B(n33225), .Z(n32697) );
  ANDN U34353 ( .B(\modmult_1/xin[1023] ), .A(n33226), .Z(n33224) );
  IV U34354 ( .A(n33225), .Z(n33226) );
  XNOR U34355 ( .A(m[975]), .B(n33227), .Z(n33225) );
  NAND U34356 ( .A(n33228), .B(mul_pow), .Z(n33227) );
  XOR U34357 ( .A(m[975]), .B(c[975]), .Z(n33228) );
  XOR U34358 ( .A(n33229), .B(n33230), .Z(n33221) );
  ANDN U34359 ( .B(n33231), .A(n32694), .Z(n33229) );
  XNOR U34360 ( .A(\modmult_1/zin[0][973] ), .B(n33232), .Z(n32694) );
  IV U34361 ( .A(n33230), .Z(n33232) );
  XOR U34362 ( .A(n33230), .B(n32695), .Z(n33231) );
  XNOR U34363 ( .A(n33233), .B(n33234), .Z(n32695) );
  ANDN U34364 ( .B(\modmult_1/xin[1023] ), .A(n33235), .Z(n33233) );
  IV U34365 ( .A(n33234), .Z(n33235) );
  XNOR U34366 ( .A(m[974]), .B(n33236), .Z(n33234) );
  NAND U34367 ( .A(n33237), .B(mul_pow), .Z(n33236) );
  XOR U34368 ( .A(m[974]), .B(c[974]), .Z(n33237) );
  XOR U34369 ( .A(n33238), .B(n33239), .Z(n33230) );
  ANDN U34370 ( .B(n33240), .A(n32692), .Z(n33238) );
  XNOR U34371 ( .A(\modmult_1/zin[0][972] ), .B(n33241), .Z(n32692) );
  IV U34372 ( .A(n33239), .Z(n33241) );
  XOR U34373 ( .A(n33239), .B(n32693), .Z(n33240) );
  XNOR U34374 ( .A(n33242), .B(n33243), .Z(n32693) );
  ANDN U34375 ( .B(\modmult_1/xin[1023] ), .A(n33244), .Z(n33242) );
  IV U34376 ( .A(n33243), .Z(n33244) );
  XNOR U34377 ( .A(m[973]), .B(n33245), .Z(n33243) );
  NAND U34378 ( .A(n33246), .B(mul_pow), .Z(n33245) );
  XOR U34379 ( .A(m[973]), .B(c[973]), .Z(n33246) );
  XOR U34380 ( .A(n33247), .B(n33248), .Z(n33239) );
  ANDN U34381 ( .B(n33249), .A(n32690), .Z(n33247) );
  XNOR U34382 ( .A(\modmult_1/zin[0][971] ), .B(n33250), .Z(n32690) );
  IV U34383 ( .A(n33248), .Z(n33250) );
  XOR U34384 ( .A(n33248), .B(n32691), .Z(n33249) );
  XNOR U34385 ( .A(n33251), .B(n33252), .Z(n32691) );
  ANDN U34386 ( .B(\modmult_1/xin[1023] ), .A(n33253), .Z(n33251) );
  IV U34387 ( .A(n33252), .Z(n33253) );
  XNOR U34388 ( .A(m[972]), .B(n33254), .Z(n33252) );
  NAND U34389 ( .A(n33255), .B(mul_pow), .Z(n33254) );
  XOR U34390 ( .A(m[972]), .B(c[972]), .Z(n33255) );
  XOR U34391 ( .A(n33256), .B(n33257), .Z(n33248) );
  ANDN U34392 ( .B(n33258), .A(n32688), .Z(n33256) );
  XNOR U34393 ( .A(\modmult_1/zin[0][970] ), .B(n33259), .Z(n32688) );
  IV U34394 ( .A(n33257), .Z(n33259) );
  XOR U34395 ( .A(n33257), .B(n32689), .Z(n33258) );
  XNOR U34396 ( .A(n33260), .B(n33261), .Z(n32689) );
  ANDN U34397 ( .B(\modmult_1/xin[1023] ), .A(n33262), .Z(n33260) );
  IV U34398 ( .A(n33261), .Z(n33262) );
  XNOR U34399 ( .A(m[971]), .B(n33263), .Z(n33261) );
  NAND U34400 ( .A(n33264), .B(mul_pow), .Z(n33263) );
  XOR U34401 ( .A(m[971]), .B(c[971]), .Z(n33264) );
  XOR U34402 ( .A(n33265), .B(n33266), .Z(n33257) );
  ANDN U34403 ( .B(n33267), .A(n32686), .Z(n33265) );
  XNOR U34404 ( .A(\modmult_1/zin[0][969] ), .B(n33268), .Z(n32686) );
  IV U34405 ( .A(n33266), .Z(n33268) );
  XOR U34406 ( .A(n33266), .B(n32687), .Z(n33267) );
  XNOR U34407 ( .A(n33269), .B(n33270), .Z(n32687) );
  ANDN U34408 ( .B(\modmult_1/xin[1023] ), .A(n33271), .Z(n33269) );
  IV U34409 ( .A(n33270), .Z(n33271) );
  XNOR U34410 ( .A(m[970]), .B(n33272), .Z(n33270) );
  NAND U34411 ( .A(n33273), .B(mul_pow), .Z(n33272) );
  XOR U34412 ( .A(m[970]), .B(c[970]), .Z(n33273) );
  XOR U34413 ( .A(n33274), .B(n33275), .Z(n33266) );
  ANDN U34414 ( .B(n33276), .A(n32684), .Z(n33274) );
  XNOR U34415 ( .A(\modmult_1/zin[0][968] ), .B(n33277), .Z(n32684) );
  IV U34416 ( .A(n33275), .Z(n33277) );
  XOR U34417 ( .A(n33275), .B(n32685), .Z(n33276) );
  XNOR U34418 ( .A(n33278), .B(n33279), .Z(n32685) );
  ANDN U34419 ( .B(\modmult_1/xin[1023] ), .A(n33280), .Z(n33278) );
  IV U34420 ( .A(n33279), .Z(n33280) );
  XNOR U34421 ( .A(m[969]), .B(n33281), .Z(n33279) );
  NAND U34422 ( .A(n33282), .B(mul_pow), .Z(n33281) );
  XOR U34423 ( .A(m[969]), .B(c[969]), .Z(n33282) );
  XOR U34424 ( .A(n33283), .B(n33284), .Z(n33275) );
  ANDN U34425 ( .B(n33285), .A(n32682), .Z(n33283) );
  XNOR U34426 ( .A(\modmult_1/zin[0][967] ), .B(n33286), .Z(n32682) );
  IV U34427 ( .A(n33284), .Z(n33286) );
  XOR U34428 ( .A(n33284), .B(n32683), .Z(n33285) );
  XNOR U34429 ( .A(n33287), .B(n33288), .Z(n32683) );
  ANDN U34430 ( .B(\modmult_1/xin[1023] ), .A(n33289), .Z(n33287) );
  IV U34431 ( .A(n33288), .Z(n33289) );
  XNOR U34432 ( .A(m[968]), .B(n33290), .Z(n33288) );
  NAND U34433 ( .A(n33291), .B(mul_pow), .Z(n33290) );
  XOR U34434 ( .A(m[968]), .B(c[968]), .Z(n33291) );
  XOR U34435 ( .A(n33292), .B(n33293), .Z(n33284) );
  ANDN U34436 ( .B(n33294), .A(n32680), .Z(n33292) );
  XNOR U34437 ( .A(\modmult_1/zin[0][966] ), .B(n33295), .Z(n32680) );
  IV U34438 ( .A(n33293), .Z(n33295) );
  XOR U34439 ( .A(n33293), .B(n32681), .Z(n33294) );
  XNOR U34440 ( .A(n33296), .B(n33297), .Z(n32681) );
  ANDN U34441 ( .B(\modmult_1/xin[1023] ), .A(n33298), .Z(n33296) );
  IV U34442 ( .A(n33297), .Z(n33298) );
  XNOR U34443 ( .A(m[967]), .B(n33299), .Z(n33297) );
  NAND U34444 ( .A(n33300), .B(mul_pow), .Z(n33299) );
  XOR U34445 ( .A(m[967]), .B(c[967]), .Z(n33300) );
  XOR U34446 ( .A(n33301), .B(n33302), .Z(n33293) );
  ANDN U34447 ( .B(n33303), .A(n32678), .Z(n33301) );
  XNOR U34448 ( .A(\modmult_1/zin[0][965] ), .B(n33304), .Z(n32678) );
  IV U34449 ( .A(n33302), .Z(n33304) );
  XOR U34450 ( .A(n33302), .B(n32679), .Z(n33303) );
  XNOR U34451 ( .A(n33305), .B(n33306), .Z(n32679) );
  ANDN U34452 ( .B(\modmult_1/xin[1023] ), .A(n33307), .Z(n33305) );
  IV U34453 ( .A(n33306), .Z(n33307) );
  XNOR U34454 ( .A(m[966]), .B(n33308), .Z(n33306) );
  NAND U34455 ( .A(n33309), .B(mul_pow), .Z(n33308) );
  XOR U34456 ( .A(m[966]), .B(c[966]), .Z(n33309) );
  XOR U34457 ( .A(n33310), .B(n33311), .Z(n33302) );
  ANDN U34458 ( .B(n33312), .A(n32676), .Z(n33310) );
  XNOR U34459 ( .A(\modmult_1/zin[0][964] ), .B(n33313), .Z(n32676) );
  IV U34460 ( .A(n33311), .Z(n33313) );
  XOR U34461 ( .A(n33311), .B(n32677), .Z(n33312) );
  XNOR U34462 ( .A(n33314), .B(n33315), .Z(n32677) );
  ANDN U34463 ( .B(\modmult_1/xin[1023] ), .A(n33316), .Z(n33314) );
  IV U34464 ( .A(n33315), .Z(n33316) );
  XNOR U34465 ( .A(m[965]), .B(n33317), .Z(n33315) );
  NAND U34466 ( .A(n33318), .B(mul_pow), .Z(n33317) );
  XOR U34467 ( .A(m[965]), .B(c[965]), .Z(n33318) );
  XOR U34468 ( .A(n33319), .B(n33320), .Z(n33311) );
  ANDN U34469 ( .B(n33321), .A(n32674), .Z(n33319) );
  XNOR U34470 ( .A(\modmult_1/zin[0][963] ), .B(n33322), .Z(n32674) );
  IV U34471 ( .A(n33320), .Z(n33322) );
  XOR U34472 ( .A(n33320), .B(n32675), .Z(n33321) );
  XNOR U34473 ( .A(n33323), .B(n33324), .Z(n32675) );
  ANDN U34474 ( .B(\modmult_1/xin[1023] ), .A(n33325), .Z(n33323) );
  IV U34475 ( .A(n33324), .Z(n33325) );
  XNOR U34476 ( .A(m[964]), .B(n33326), .Z(n33324) );
  NAND U34477 ( .A(n33327), .B(mul_pow), .Z(n33326) );
  XOR U34478 ( .A(m[964]), .B(c[964]), .Z(n33327) );
  XOR U34479 ( .A(n33328), .B(n33329), .Z(n33320) );
  ANDN U34480 ( .B(n33330), .A(n32672), .Z(n33328) );
  XNOR U34481 ( .A(\modmult_1/zin[0][962] ), .B(n33331), .Z(n32672) );
  IV U34482 ( .A(n33329), .Z(n33331) );
  XOR U34483 ( .A(n33329), .B(n32673), .Z(n33330) );
  XNOR U34484 ( .A(n33332), .B(n33333), .Z(n32673) );
  ANDN U34485 ( .B(\modmult_1/xin[1023] ), .A(n33334), .Z(n33332) );
  IV U34486 ( .A(n33333), .Z(n33334) );
  XNOR U34487 ( .A(m[963]), .B(n33335), .Z(n33333) );
  NAND U34488 ( .A(n33336), .B(mul_pow), .Z(n33335) );
  XOR U34489 ( .A(m[963]), .B(c[963]), .Z(n33336) );
  XOR U34490 ( .A(n33337), .B(n33338), .Z(n33329) );
  ANDN U34491 ( .B(n33339), .A(n32670), .Z(n33337) );
  XNOR U34492 ( .A(\modmult_1/zin[0][961] ), .B(n33340), .Z(n32670) );
  IV U34493 ( .A(n33338), .Z(n33340) );
  XOR U34494 ( .A(n33338), .B(n32671), .Z(n33339) );
  XNOR U34495 ( .A(n33341), .B(n33342), .Z(n32671) );
  ANDN U34496 ( .B(\modmult_1/xin[1023] ), .A(n33343), .Z(n33341) );
  IV U34497 ( .A(n33342), .Z(n33343) );
  XNOR U34498 ( .A(m[962]), .B(n33344), .Z(n33342) );
  NAND U34499 ( .A(n33345), .B(mul_pow), .Z(n33344) );
  XOR U34500 ( .A(m[962]), .B(c[962]), .Z(n33345) );
  XOR U34501 ( .A(n33346), .B(n33347), .Z(n33338) );
  ANDN U34502 ( .B(n33348), .A(n32668), .Z(n33346) );
  XNOR U34503 ( .A(\modmult_1/zin[0][960] ), .B(n33349), .Z(n32668) );
  IV U34504 ( .A(n33347), .Z(n33349) );
  XOR U34505 ( .A(n33347), .B(n32669), .Z(n33348) );
  XNOR U34506 ( .A(n33350), .B(n33351), .Z(n32669) );
  ANDN U34507 ( .B(\modmult_1/xin[1023] ), .A(n33352), .Z(n33350) );
  IV U34508 ( .A(n33351), .Z(n33352) );
  XNOR U34509 ( .A(m[961]), .B(n33353), .Z(n33351) );
  NAND U34510 ( .A(n33354), .B(mul_pow), .Z(n33353) );
  XOR U34511 ( .A(m[961]), .B(c[961]), .Z(n33354) );
  XOR U34512 ( .A(n33355), .B(n33356), .Z(n33347) );
  ANDN U34513 ( .B(n33357), .A(n32666), .Z(n33355) );
  XNOR U34514 ( .A(\modmult_1/zin[0][959] ), .B(n33358), .Z(n32666) );
  IV U34515 ( .A(n33356), .Z(n33358) );
  XOR U34516 ( .A(n33356), .B(n32667), .Z(n33357) );
  XNOR U34517 ( .A(n33359), .B(n33360), .Z(n32667) );
  ANDN U34518 ( .B(\modmult_1/xin[1023] ), .A(n33361), .Z(n33359) );
  IV U34519 ( .A(n33360), .Z(n33361) );
  XNOR U34520 ( .A(m[960]), .B(n33362), .Z(n33360) );
  NAND U34521 ( .A(n33363), .B(mul_pow), .Z(n33362) );
  XOR U34522 ( .A(m[960]), .B(c[960]), .Z(n33363) );
  XOR U34523 ( .A(n33364), .B(n33365), .Z(n33356) );
  ANDN U34524 ( .B(n33366), .A(n32664), .Z(n33364) );
  XNOR U34525 ( .A(\modmult_1/zin[0][958] ), .B(n33367), .Z(n32664) );
  IV U34526 ( .A(n33365), .Z(n33367) );
  XOR U34527 ( .A(n33365), .B(n32665), .Z(n33366) );
  XNOR U34528 ( .A(n33368), .B(n33369), .Z(n32665) );
  ANDN U34529 ( .B(\modmult_1/xin[1023] ), .A(n33370), .Z(n33368) );
  IV U34530 ( .A(n33369), .Z(n33370) );
  XNOR U34531 ( .A(m[959]), .B(n33371), .Z(n33369) );
  NAND U34532 ( .A(n33372), .B(mul_pow), .Z(n33371) );
  XOR U34533 ( .A(m[959]), .B(c[959]), .Z(n33372) );
  XOR U34534 ( .A(n33373), .B(n33374), .Z(n33365) );
  ANDN U34535 ( .B(n33375), .A(n32662), .Z(n33373) );
  XNOR U34536 ( .A(\modmult_1/zin[0][957] ), .B(n33376), .Z(n32662) );
  IV U34537 ( .A(n33374), .Z(n33376) );
  XOR U34538 ( .A(n33374), .B(n32663), .Z(n33375) );
  XNOR U34539 ( .A(n33377), .B(n33378), .Z(n32663) );
  ANDN U34540 ( .B(\modmult_1/xin[1023] ), .A(n33379), .Z(n33377) );
  IV U34541 ( .A(n33378), .Z(n33379) );
  XNOR U34542 ( .A(m[958]), .B(n33380), .Z(n33378) );
  NAND U34543 ( .A(n33381), .B(mul_pow), .Z(n33380) );
  XOR U34544 ( .A(m[958]), .B(c[958]), .Z(n33381) );
  XOR U34545 ( .A(n33382), .B(n33383), .Z(n33374) );
  ANDN U34546 ( .B(n33384), .A(n32660), .Z(n33382) );
  XNOR U34547 ( .A(\modmult_1/zin[0][956] ), .B(n33385), .Z(n32660) );
  IV U34548 ( .A(n33383), .Z(n33385) );
  XOR U34549 ( .A(n33383), .B(n32661), .Z(n33384) );
  XNOR U34550 ( .A(n33386), .B(n33387), .Z(n32661) );
  ANDN U34551 ( .B(\modmult_1/xin[1023] ), .A(n33388), .Z(n33386) );
  IV U34552 ( .A(n33387), .Z(n33388) );
  XNOR U34553 ( .A(m[957]), .B(n33389), .Z(n33387) );
  NAND U34554 ( .A(n33390), .B(mul_pow), .Z(n33389) );
  XOR U34555 ( .A(m[957]), .B(c[957]), .Z(n33390) );
  XOR U34556 ( .A(n33391), .B(n33392), .Z(n33383) );
  ANDN U34557 ( .B(n33393), .A(n32658), .Z(n33391) );
  XNOR U34558 ( .A(\modmult_1/zin[0][955] ), .B(n33394), .Z(n32658) );
  IV U34559 ( .A(n33392), .Z(n33394) );
  XOR U34560 ( .A(n33392), .B(n32659), .Z(n33393) );
  XNOR U34561 ( .A(n33395), .B(n33396), .Z(n32659) );
  ANDN U34562 ( .B(\modmult_1/xin[1023] ), .A(n33397), .Z(n33395) );
  IV U34563 ( .A(n33396), .Z(n33397) );
  XNOR U34564 ( .A(m[956]), .B(n33398), .Z(n33396) );
  NAND U34565 ( .A(n33399), .B(mul_pow), .Z(n33398) );
  XOR U34566 ( .A(m[956]), .B(c[956]), .Z(n33399) );
  XOR U34567 ( .A(n33400), .B(n33401), .Z(n33392) );
  ANDN U34568 ( .B(n33402), .A(n32656), .Z(n33400) );
  XNOR U34569 ( .A(\modmult_1/zin[0][954] ), .B(n33403), .Z(n32656) );
  IV U34570 ( .A(n33401), .Z(n33403) );
  XOR U34571 ( .A(n33401), .B(n32657), .Z(n33402) );
  XNOR U34572 ( .A(n33404), .B(n33405), .Z(n32657) );
  ANDN U34573 ( .B(\modmult_1/xin[1023] ), .A(n33406), .Z(n33404) );
  IV U34574 ( .A(n33405), .Z(n33406) );
  XNOR U34575 ( .A(m[955]), .B(n33407), .Z(n33405) );
  NAND U34576 ( .A(n33408), .B(mul_pow), .Z(n33407) );
  XOR U34577 ( .A(m[955]), .B(c[955]), .Z(n33408) );
  XOR U34578 ( .A(n33409), .B(n33410), .Z(n33401) );
  ANDN U34579 ( .B(n33411), .A(n32654), .Z(n33409) );
  XNOR U34580 ( .A(\modmult_1/zin[0][953] ), .B(n33412), .Z(n32654) );
  IV U34581 ( .A(n33410), .Z(n33412) );
  XOR U34582 ( .A(n33410), .B(n32655), .Z(n33411) );
  XNOR U34583 ( .A(n33413), .B(n33414), .Z(n32655) );
  ANDN U34584 ( .B(\modmult_1/xin[1023] ), .A(n33415), .Z(n33413) );
  IV U34585 ( .A(n33414), .Z(n33415) );
  XNOR U34586 ( .A(m[954]), .B(n33416), .Z(n33414) );
  NAND U34587 ( .A(n33417), .B(mul_pow), .Z(n33416) );
  XOR U34588 ( .A(m[954]), .B(c[954]), .Z(n33417) );
  XOR U34589 ( .A(n33418), .B(n33419), .Z(n33410) );
  ANDN U34590 ( .B(n33420), .A(n32652), .Z(n33418) );
  XNOR U34591 ( .A(\modmult_1/zin[0][952] ), .B(n33421), .Z(n32652) );
  IV U34592 ( .A(n33419), .Z(n33421) );
  XOR U34593 ( .A(n33419), .B(n32653), .Z(n33420) );
  XNOR U34594 ( .A(n33422), .B(n33423), .Z(n32653) );
  ANDN U34595 ( .B(\modmult_1/xin[1023] ), .A(n33424), .Z(n33422) );
  IV U34596 ( .A(n33423), .Z(n33424) );
  XNOR U34597 ( .A(m[953]), .B(n33425), .Z(n33423) );
  NAND U34598 ( .A(n33426), .B(mul_pow), .Z(n33425) );
  XOR U34599 ( .A(m[953]), .B(c[953]), .Z(n33426) );
  XOR U34600 ( .A(n33427), .B(n33428), .Z(n33419) );
  ANDN U34601 ( .B(n33429), .A(n32650), .Z(n33427) );
  XNOR U34602 ( .A(\modmult_1/zin[0][951] ), .B(n33430), .Z(n32650) );
  IV U34603 ( .A(n33428), .Z(n33430) );
  XOR U34604 ( .A(n33428), .B(n32651), .Z(n33429) );
  XNOR U34605 ( .A(n33431), .B(n33432), .Z(n32651) );
  ANDN U34606 ( .B(\modmult_1/xin[1023] ), .A(n33433), .Z(n33431) );
  IV U34607 ( .A(n33432), .Z(n33433) );
  XNOR U34608 ( .A(m[952]), .B(n33434), .Z(n33432) );
  NAND U34609 ( .A(n33435), .B(mul_pow), .Z(n33434) );
  XOR U34610 ( .A(m[952]), .B(c[952]), .Z(n33435) );
  XOR U34611 ( .A(n33436), .B(n33437), .Z(n33428) );
  ANDN U34612 ( .B(n33438), .A(n32648), .Z(n33436) );
  XNOR U34613 ( .A(\modmult_1/zin[0][950] ), .B(n33439), .Z(n32648) );
  IV U34614 ( .A(n33437), .Z(n33439) );
  XOR U34615 ( .A(n33437), .B(n32649), .Z(n33438) );
  XNOR U34616 ( .A(n33440), .B(n33441), .Z(n32649) );
  ANDN U34617 ( .B(\modmult_1/xin[1023] ), .A(n33442), .Z(n33440) );
  IV U34618 ( .A(n33441), .Z(n33442) );
  XNOR U34619 ( .A(m[951]), .B(n33443), .Z(n33441) );
  NAND U34620 ( .A(n33444), .B(mul_pow), .Z(n33443) );
  XOR U34621 ( .A(m[951]), .B(c[951]), .Z(n33444) );
  XOR U34622 ( .A(n33445), .B(n33446), .Z(n33437) );
  ANDN U34623 ( .B(n33447), .A(n32646), .Z(n33445) );
  XNOR U34624 ( .A(\modmult_1/zin[0][949] ), .B(n33448), .Z(n32646) );
  IV U34625 ( .A(n33446), .Z(n33448) );
  XOR U34626 ( .A(n33446), .B(n32647), .Z(n33447) );
  XNOR U34627 ( .A(n33449), .B(n33450), .Z(n32647) );
  ANDN U34628 ( .B(\modmult_1/xin[1023] ), .A(n33451), .Z(n33449) );
  IV U34629 ( .A(n33450), .Z(n33451) );
  XNOR U34630 ( .A(m[950]), .B(n33452), .Z(n33450) );
  NAND U34631 ( .A(n33453), .B(mul_pow), .Z(n33452) );
  XOR U34632 ( .A(m[950]), .B(c[950]), .Z(n33453) );
  XOR U34633 ( .A(n33454), .B(n33455), .Z(n33446) );
  ANDN U34634 ( .B(n33456), .A(n32644), .Z(n33454) );
  XNOR U34635 ( .A(\modmult_1/zin[0][948] ), .B(n33457), .Z(n32644) );
  IV U34636 ( .A(n33455), .Z(n33457) );
  XOR U34637 ( .A(n33455), .B(n32645), .Z(n33456) );
  XNOR U34638 ( .A(n33458), .B(n33459), .Z(n32645) );
  ANDN U34639 ( .B(\modmult_1/xin[1023] ), .A(n33460), .Z(n33458) );
  IV U34640 ( .A(n33459), .Z(n33460) );
  XNOR U34641 ( .A(m[949]), .B(n33461), .Z(n33459) );
  NAND U34642 ( .A(n33462), .B(mul_pow), .Z(n33461) );
  XOR U34643 ( .A(m[949]), .B(c[949]), .Z(n33462) );
  XOR U34644 ( .A(n33463), .B(n33464), .Z(n33455) );
  ANDN U34645 ( .B(n33465), .A(n32642), .Z(n33463) );
  XNOR U34646 ( .A(\modmult_1/zin[0][947] ), .B(n33466), .Z(n32642) );
  IV U34647 ( .A(n33464), .Z(n33466) );
  XOR U34648 ( .A(n33464), .B(n32643), .Z(n33465) );
  XNOR U34649 ( .A(n33467), .B(n33468), .Z(n32643) );
  ANDN U34650 ( .B(\modmult_1/xin[1023] ), .A(n33469), .Z(n33467) );
  IV U34651 ( .A(n33468), .Z(n33469) );
  XNOR U34652 ( .A(m[948]), .B(n33470), .Z(n33468) );
  NAND U34653 ( .A(n33471), .B(mul_pow), .Z(n33470) );
  XOR U34654 ( .A(m[948]), .B(c[948]), .Z(n33471) );
  XOR U34655 ( .A(n33472), .B(n33473), .Z(n33464) );
  ANDN U34656 ( .B(n33474), .A(n32640), .Z(n33472) );
  XNOR U34657 ( .A(\modmult_1/zin[0][946] ), .B(n33475), .Z(n32640) );
  IV U34658 ( .A(n33473), .Z(n33475) );
  XOR U34659 ( .A(n33473), .B(n32641), .Z(n33474) );
  XNOR U34660 ( .A(n33476), .B(n33477), .Z(n32641) );
  ANDN U34661 ( .B(\modmult_1/xin[1023] ), .A(n33478), .Z(n33476) );
  IV U34662 ( .A(n33477), .Z(n33478) );
  XNOR U34663 ( .A(m[947]), .B(n33479), .Z(n33477) );
  NAND U34664 ( .A(n33480), .B(mul_pow), .Z(n33479) );
  XOR U34665 ( .A(m[947]), .B(c[947]), .Z(n33480) );
  XOR U34666 ( .A(n33481), .B(n33482), .Z(n33473) );
  ANDN U34667 ( .B(n33483), .A(n32638), .Z(n33481) );
  XNOR U34668 ( .A(\modmult_1/zin[0][945] ), .B(n33484), .Z(n32638) );
  IV U34669 ( .A(n33482), .Z(n33484) );
  XOR U34670 ( .A(n33482), .B(n32639), .Z(n33483) );
  XNOR U34671 ( .A(n33485), .B(n33486), .Z(n32639) );
  ANDN U34672 ( .B(\modmult_1/xin[1023] ), .A(n33487), .Z(n33485) );
  IV U34673 ( .A(n33486), .Z(n33487) );
  XNOR U34674 ( .A(m[946]), .B(n33488), .Z(n33486) );
  NAND U34675 ( .A(n33489), .B(mul_pow), .Z(n33488) );
  XOR U34676 ( .A(m[946]), .B(c[946]), .Z(n33489) );
  XOR U34677 ( .A(n33490), .B(n33491), .Z(n33482) );
  ANDN U34678 ( .B(n33492), .A(n32636), .Z(n33490) );
  XNOR U34679 ( .A(\modmult_1/zin[0][944] ), .B(n33493), .Z(n32636) );
  IV U34680 ( .A(n33491), .Z(n33493) );
  XOR U34681 ( .A(n33491), .B(n32637), .Z(n33492) );
  XNOR U34682 ( .A(n33494), .B(n33495), .Z(n32637) );
  ANDN U34683 ( .B(\modmult_1/xin[1023] ), .A(n33496), .Z(n33494) );
  IV U34684 ( .A(n33495), .Z(n33496) );
  XNOR U34685 ( .A(m[945]), .B(n33497), .Z(n33495) );
  NAND U34686 ( .A(n33498), .B(mul_pow), .Z(n33497) );
  XOR U34687 ( .A(m[945]), .B(c[945]), .Z(n33498) );
  XOR U34688 ( .A(n33499), .B(n33500), .Z(n33491) );
  ANDN U34689 ( .B(n33501), .A(n32634), .Z(n33499) );
  XNOR U34690 ( .A(\modmult_1/zin[0][943] ), .B(n33502), .Z(n32634) );
  IV U34691 ( .A(n33500), .Z(n33502) );
  XOR U34692 ( .A(n33500), .B(n32635), .Z(n33501) );
  XNOR U34693 ( .A(n33503), .B(n33504), .Z(n32635) );
  ANDN U34694 ( .B(\modmult_1/xin[1023] ), .A(n33505), .Z(n33503) );
  IV U34695 ( .A(n33504), .Z(n33505) );
  XNOR U34696 ( .A(m[944]), .B(n33506), .Z(n33504) );
  NAND U34697 ( .A(n33507), .B(mul_pow), .Z(n33506) );
  XOR U34698 ( .A(m[944]), .B(c[944]), .Z(n33507) );
  XOR U34699 ( .A(n33508), .B(n33509), .Z(n33500) );
  ANDN U34700 ( .B(n33510), .A(n32632), .Z(n33508) );
  XNOR U34701 ( .A(\modmult_1/zin[0][942] ), .B(n33511), .Z(n32632) );
  IV U34702 ( .A(n33509), .Z(n33511) );
  XOR U34703 ( .A(n33509), .B(n32633), .Z(n33510) );
  XNOR U34704 ( .A(n33512), .B(n33513), .Z(n32633) );
  ANDN U34705 ( .B(\modmult_1/xin[1023] ), .A(n33514), .Z(n33512) );
  IV U34706 ( .A(n33513), .Z(n33514) );
  XNOR U34707 ( .A(m[943]), .B(n33515), .Z(n33513) );
  NAND U34708 ( .A(n33516), .B(mul_pow), .Z(n33515) );
  XOR U34709 ( .A(m[943]), .B(c[943]), .Z(n33516) );
  XOR U34710 ( .A(n33517), .B(n33518), .Z(n33509) );
  ANDN U34711 ( .B(n33519), .A(n32630), .Z(n33517) );
  XNOR U34712 ( .A(\modmult_1/zin[0][941] ), .B(n33520), .Z(n32630) );
  IV U34713 ( .A(n33518), .Z(n33520) );
  XOR U34714 ( .A(n33518), .B(n32631), .Z(n33519) );
  XNOR U34715 ( .A(n33521), .B(n33522), .Z(n32631) );
  ANDN U34716 ( .B(\modmult_1/xin[1023] ), .A(n33523), .Z(n33521) );
  IV U34717 ( .A(n33522), .Z(n33523) );
  XNOR U34718 ( .A(m[942]), .B(n33524), .Z(n33522) );
  NAND U34719 ( .A(n33525), .B(mul_pow), .Z(n33524) );
  XOR U34720 ( .A(m[942]), .B(c[942]), .Z(n33525) );
  XOR U34721 ( .A(n33526), .B(n33527), .Z(n33518) );
  ANDN U34722 ( .B(n33528), .A(n32628), .Z(n33526) );
  XNOR U34723 ( .A(\modmult_1/zin[0][940] ), .B(n33529), .Z(n32628) );
  IV U34724 ( .A(n33527), .Z(n33529) );
  XOR U34725 ( .A(n33527), .B(n32629), .Z(n33528) );
  XNOR U34726 ( .A(n33530), .B(n33531), .Z(n32629) );
  ANDN U34727 ( .B(\modmult_1/xin[1023] ), .A(n33532), .Z(n33530) );
  IV U34728 ( .A(n33531), .Z(n33532) );
  XNOR U34729 ( .A(m[941]), .B(n33533), .Z(n33531) );
  NAND U34730 ( .A(n33534), .B(mul_pow), .Z(n33533) );
  XOR U34731 ( .A(m[941]), .B(c[941]), .Z(n33534) );
  XOR U34732 ( .A(n33535), .B(n33536), .Z(n33527) );
  ANDN U34733 ( .B(n33537), .A(n32626), .Z(n33535) );
  XNOR U34734 ( .A(\modmult_1/zin[0][939] ), .B(n33538), .Z(n32626) );
  IV U34735 ( .A(n33536), .Z(n33538) );
  XOR U34736 ( .A(n33536), .B(n32627), .Z(n33537) );
  XNOR U34737 ( .A(n33539), .B(n33540), .Z(n32627) );
  ANDN U34738 ( .B(\modmult_1/xin[1023] ), .A(n33541), .Z(n33539) );
  IV U34739 ( .A(n33540), .Z(n33541) );
  XNOR U34740 ( .A(m[940]), .B(n33542), .Z(n33540) );
  NAND U34741 ( .A(n33543), .B(mul_pow), .Z(n33542) );
  XOR U34742 ( .A(m[940]), .B(c[940]), .Z(n33543) );
  XOR U34743 ( .A(n33544), .B(n33545), .Z(n33536) );
  ANDN U34744 ( .B(n33546), .A(n32624), .Z(n33544) );
  XNOR U34745 ( .A(\modmult_1/zin[0][938] ), .B(n33547), .Z(n32624) );
  IV U34746 ( .A(n33545), .Z(n33547) );
  XOR U34747 ( .A(n33545), .B(n32625), .Z(n33546) );
  XNOR U34748 ( .A(n33548), .B(n33549), .Z(n32625) );
  ANDN U34749 ( .B(\modmult_1/xin[1023] ), .A(n33550), .Z(n33548) );
  IV U34750 ( .A(n33549), .Z(n33550) );
  XNOR U34751 ( .A(m[939]), .B(n33551), .Z(n33549) );
  NAND U34752 ( .A(n33552), .B(mul_pow), .Z(n33551) );
  XOR U34753 ( .A(m[939]), .B(c[939]), .Z(n33552) );
  XOR U34754 ( .A(n33553), .B(n33554), .Z(n33545) );
  ANDN U34755 ( .B(n33555), .A(n32622), .Z(n33553) );
  XNOR U34756 ( .A(\modmult_1/zin[0][937] ), .B(n33556), .Z(n32622) );
  IV U34757 ( .A(n33554), .Z(n33556) );
  XOR U34758 ( .A(n33554), .B(n32623), .Z(n33555) );
  XNOR U34759 ( .A(n33557), .B(n33558), .Z(n32623) );
  ANDN U34760 ( .B(\modmult_1/xin[1023] ), .A(n33559), .Z(n33557) );
  IV U34761 ( .A(n33558), .Z(n33559) );
  XNOR U34762 ( .A(m[938]), .B(n33560), .Z(n33558) );
  NAND U34763 ( .A(n33561), .B(mul_pow), .Z(n33560) );
  XOR U34764 ( .A(m[938]), .B(c[938]), .Z(n33561) );
  XOR U34765 ( .A(n33562), .B(n33563), .Z(n33554) );
  ANDN U34766 ( .B(n33564), .A(n32620), .Z(n33562) );
  XNOR U34767 ( .A(\modmult_1/zin[0][936] ), .B(n33565), .Z(n32620) );
  IV U34768 ( .A(n33563), .Z(n33565) );
  XOR U34769 ( .A(n33563), .B(n32621), .Z(n33564) );
  XNOR U34770 ( .A(n33566), .B(n33567), .Z(n32621) );
  ANDN U34771 ( .B(\modmult_1/xin[1023] ), .A(n33568), .Z(n33566) );
  IV U34772 ( .A(n33567), .Z(n33568) );
  XNOR U34773 ( .A(m[937]), .B(n33569), .Z(n33567) );
  NAND U34774 ( .A(n33570), .B(mul_pow), .Z(n33569) );
  XOR U34775 ( .A(m[937]), .B(c[937]), .Z(n33570) );
  XOR U34776 ( .A(n33571), .B(n33572), .Z(n33563) );
  ANDN U34777 ( .B(n33573), .A(n32618), .Z(n33571) );
  XNOR U34778 ( .A(\modmult_1/zin[0][935] ), .B(n33574), .Z(n32618) );
  IV U34779 ( .A(n33572), .Z(n33574) );
  XOR U34780 ( .A(n33572), .B(n32619), .Z(n33573) );
  XNOR U34781 ( .A(n33575), .B(n33576), .Z(n32619) );
  ANDN U34782 ( .B(\modmult_1/xin[1023] ), .A(n33577), .Z(n33575) );
  IV U34783 ( .A(n33576), .Z(n33577) );
  XNOR U34784 ( .A(m[936]), .B(n33578), .Z(n33576) );
  NAND U34785 ( .A(n33579), .B(mul_pow), .Z(n33578) );
  XOR U34786 ( .A(m[936]), .B(c[936]), .Z(n33579) );
  XOR U34787 ( .A(n33580), .B(n33581), .Z(n33572) );
  ANDN U34788 ( .B(n33582), .A(n32616), .Z(n33580) );
  XNOR U34789 ( .A(\modmult_1/zin[0][934] ), .B(n33583), .Z(n32616) );
  IV U34790 ( .A(n33581), .Z(n33583) );
  XOR U34791 ( .A(n33581), .B(n32617), .Z(n33582) );
  XNOR U34792 ( .A(n33584), .B(n33585), .Z(n32617) );
  ANDN U34793 ( .B(\modmult_1/xin[1023] ), .A(n33586), .Z(n33584) );
  IV U34794 ( .A(n33585), .Z(n33586) );
  XNOR U34795 ( .A(m[935]), .B(n33587), .Z(n33585) );
  NAND U34796 ( .A(n33588), .B(mul_pow), .Z(n33587) );
  XOR U34797 ( .A(m[935]), .B(c[935]), .Z(n33588) );
  XOR U34798 ( .A(n33589), .B(n33590), .Z(n33581) );
  ANDN U34799 ( .B(n33591), .A(n32614), .Z(n33589) );
  XNOR U34800 ( .A(\modmult_1/zin[0][933] ), .B(n33592), .Z(n32614) );
  IV U34801 ( .A(n33590), .Z(n33592) );
  XOR U34802 ( .A(n33590), .B(n32615), .Z(n33591) );
  XNOR U34803 ( .A(n33593), .B(n33594), .Z(n32615) );
  ANDN U34804 ( .B(\modmult_1/xin[1023] ), .A(n33595), .Z(n33593) );
  IV U34805 ( .A(n33594), .Z(n33595) );
  XNOR U34806 ( .A(m[934]), .B(n33596), .Z(n33594) );
  NAND U34807 ( .A(n33597), .B(mul_pow), .Z(n33596) );
  XOR U34808 ( .A(m[934]), .B(c[934]), .Z(n33597) );
  XOR U34809 ( .A(n33598), .B(n33599), .Z(n33590) );
  ANDN U34810 ( .B(n33600), .A(n32612), .Z(n33598) );
  XNOR U34811 ( .A(\modmult_1/zin[0][932] ), .B(n33601), .Z(n32612) );
  IV U34812 ( .A(n33599), .Z(n33601) );
  XOR U34813 ( .A(n33599), .B(n32613), .Z(n33600) );
  XNOR U34814 ( .A(n33602), .B(n33603), .Z(n32613) );
  ANDN U34815 ( .B(\modmult_1/xin[1023] ), .A(n33604), .Z(n33602) );
  IV U34816 ( .A(n33603), .Z(n33604) );
  XNOR U34817 ( .A(m[933]), .B(n33605), .Z(n33603) );
  NAND U34818 ( .A(n33606), .B(mul_pow), .Z(n33605) );
  XOR U34819 ( .A(m[933]), .B(c[933]), .Z(n33606) );
  XOR U34820 ( .A(n33607), .B(n33608), .Z(n33599) );
  ANDN U34821 ( .B(n33609), .A(n32610), .Z(n33607) );
  XNOR U34822 ( .A(\modmult_1/zin[0][931] ), .B(n33610), .Z(n32610) );
  IV U34823 ( .A(n33608), .Z(n33610) );
  XOR U34824 ( .A(n33608), .B(n32611), .Z(n33609) );
  XNOR U34825 ( .A(n33611), .B(n33612), .Z(n32611) );
  ANDN U34826 ( .B(\modmult_1/xin[1023] ), .A(n33613), .Z(n33611) );
  IV U34827 ( .A(n33612), .Z(n33613) );
  XNOR U34828 ( .A(m[932]), .B(n33614), .Z(n33612) );
  NAND U34829 ( .A(n33615), .B(mul_pow), .Z(n33614) );
  XOR U34830 ( .A(m[932]), .B(c[932]), .Z(n33615) );
  XOR U34831 ( .A(n33616), .B(n33617), .Z(n33608) );
  ANDN U34832 ( .B(n33618), .A(n32608), .Z(n33616) );
  XNOR U34833 ( .A(\modmult_1/zin[0][930] ), .B(n33619), .Z(n32608) );
  IV U34834 ( .A(n33617), .Z(n33619) );
  XOR U34835 ( .A(n33617), .B(n32609), .Z(n33618) );
  XNOR U34836 ( .A(n33620), .B(n33621), .Z(n32609) );
  ANDN U34837 ( .B(\modmult_1/xin[1023] ), .A(n33622), .Z(n33620) );
  IV U34838 ( .A(n33621), .Z(n33622) );
  XNOR U34839 ( .A(m[931]), .B(n33623), .Z(n33621) );
  NAND U34840 ( .A(n33624), .B(mul_pow), .Z(n33623) );
  XOR U34841 ( .A(m[931]), .B(c[931]), .Z(n33624) );
  XOR U34842 ( .A(n33625), .B(n33626), .Z(n33617) );
  ANDN U34843 ( .B(n33627), .A(n32606), .Z(n33625) );
  XNOR U34844 ( .A(\modmult_1/zin[0][929] ), .B(n33628), .Z(n32606) );
  IV U34845 ( .A(n33626), .Z(n33628) );
  XOR U34846 ( .A(n33626), .B(n32607), .Z(n33627) );
  XNOR U34847 ( .A(n33629), .B(n33630), .Z(n32607) );
  ANDN U34848 ( .B(\modmult_1/xin[1023] ), .A(n33631), .Z(n33629) );
  IV U34849 ( .A(n33630), .Z(n33631) );
  XNOR U34850 ( .A(m[930]), .B(n33632), .Z(n33630) );
  NAND U34851 ( .A(n33633), .B(mul_pow), .Z(n33632) );
  XOR U34852 ( .A(m[930]), .B(c[930]), .Z(n33633) );
  XOR U34853 ( .A(n33634), .B(n33635), .Z(n33626) );
  ANDN U34854 ( .B(n33636), .A(n32604), .Z(n33634) );
  XNOR U34855 ( .A(\modmult_1/zin[0][928] ), .B(n33637), .Z(n32604) );
  IV U34856 ( .A(n33635), .Z(n33637) );
  XOR U34857 ( .A(n33635), .B(n32605), .Z(n33636) );
  XNOR U34858 ( .A(n33638), .B(n33639), .Z(n32605) );
  ANDN U34859 ( .B(\modmult_1/xin[1023] ), .A(n33640), .Z(n33638) );
  IV U34860 ( .A(n33639), .Z(n33640) );
  XNOR U34861 ( .A(m[929]), .B(n33641), .Z(n33639) );
  NAND U34862 ( .A(n33642), .B(mul_pow), .Z(n33641) );
  XOR U34863 ( .A(m[929]), .B(c[929]), .Z(n33642) );
  XOR U34864 ( .A(n33643), .B(n33644), .Z(n33635) );
  ANDN U34865 ( .B(n33645), .A(n32602), .Z(n33643) );
  XNOR U34866 ( .A(\modmult_1/zin[0][927] ), .B(n33646), .Z(n32602) );
  IV U34867 ( .A(n33644), .Z(n33646) );
  XOR U34868 ( .A(n33644), .B(n32603), .Z(n33645) );
  XNOR U34869 ( .A(n33647), .B(n33648), .Z(n32603) );
  ANDN U34870 ( .B(\modmult_1/xin[1023] ), .A(n33649), .Z(n33647) );
  IV U34871 ( .A(n33648), .Z(n33649) );
  XNOR U34872 ( .A(m[928]), .B(n33650), .Z(n33648) );
  NAND U34873 ( .A(n33651), .B(mul_pow), .Z(n33650) );
  XOR U34874 ( .A(m[928]), .B(c[928]), .Z(n33651) );
  XOR U34875 ( .A(n33652), .B(n33653), .Z(n33644) );
  ANDN U34876 ( .B(n33654), .A(n32600), .Z(n33652) );
  XNOR U34877 ( .A(\modmult_1/zin[0][926] ), .B(n33655), .Z(n32600) );
  IV U34878 ( .A(n33653), .Z(n33655) );
  XOR U34879 ( .A(n33653), .B(n32601), .Z(n33654) );
  XNOR U34880 ( .A(n33656), .B(n33657), .Z(n32601) );
  ANDN U34881 ( .B(\modmult_1/xin[1023] ), .A(n33658), .Z(n33656) );
  IV U34882 ( .A(n33657), .Z(n33658) );
  XNOR U34883 ( .A(m[927]), .B(n33659), .Z(n33657) );
  NAND U34884 ( .A(n33660), .B(mul_pow), .Z(n33659) );
  XOR U34885 ( .A(m[927]), .B(c[927]), .Z(n33660) );
  XOR U34886 ( .A(n33661), .B(n33662), .Z(n33653) );
  ANDN U34887 ( .B(n33663), .A(n32598), .Z(n33661) );
  XNOR U34888 ( .A(\modmult_1/zin[0][925] ), .B(n33664), .Z(n32598) );
  IV U34889 ( .A(n33662), .Z(n33664) );
  XOR U34890 ( .A(n33662), .B(n32599), .Z(n33663) );
  XNOR U34891 ( .A(n33665), .B(n33666), .Z(n32599) );
  ANDN U34892 ( .B(\modmult_1/xin[1023] ), .A(n33667), .Z(n33665) );
  IV U34893 ( .A(n33666), .Z(n33667) );
  XNOR U34894 ( .A(m[926]), .B(n33668), .Z(n33666) );
  NAND U34895 ( .A(n33669), .B(mul_pow), .Z(n33668) );
  XOR U34896 ( .A(m[926]), .B(c[926]), .Z(n33669) );
  XOR U34897 ( .A(n33670), .B(n33671), .Z(n33662) );
  ANDN U34898 ( .B(n33672), .A(n32596), .Z(n33670) );
  XNOR U34899 ( .A(\modmult_1/zin[0][924] ), .B(n33673), .Z(n32596) );
  IV U34900 ( .A(n33671), .Z(n33673) );
  XOR U34901 ( .A(n33671), .B(n32597), .Z(n33672) );
  XNOR U34902 ( .A(n33674), .B(n33675), .Z(n32597) );
  ANDN U34903 ( .B(\modmult_1/xin[1023] ), .A(n33676), .Z(n33674) );
  IV U34904 ( .A(n33675), .Z(n33676) );
  XNOR U34905 ( .A(m[925]), .B(n33677), .Z(n33675) );
  NAND U34906 ( .A(n33678), .B(mul_pow), .Z(n33677) );
  XOR U34907 ( .A(m[925]), .B(c[925]), .Z(n33678) );
  XOR U34908 ( .A(n33679), .B(n33680), .Z(n33671) );
  ANDN U34909 ( .B(n33681), .A(n32594), .Z(n33679) );
  XNOR U34910 ( .A(\modmult_1/zin[0][923] ), .B(n33682), .Z(n32594) );
  IV U34911 ( .A(n33680), .Z(n33682) );
  XOR U34912 ( .A(n33680), .B(n32595), .Z(n33681) );
  XNOR U34913 ( .A(n33683), .B(n33684), .Z(n32595) );
  ANDN U34914 ( .B(\modmult_1/xin[1023] ), .A(n33685), .Z(n33683) );
  IV U34915 ( .A(n33684), .Z(n33685) );
  XNOR U34916 ( .A(m[924]), .B(n33686), .Z(n33684) );
  NAND U34917 ( .A(n33687), .B(mul_pow), .Z(n33686) );
  XOR U34918 ( .A(m[924]), .B(c[924]), .Z(n33687) );
  XOR U34919 ( .A(n33688), .B(n33689), .Z(n33680) );
  ANDN U34920 ( .B(n33690), .A(n32592), .Z(n33688) );
  XNOR U34921 ( .A(\modmult_1/zin[0][922] ), .B(n33691), .Z(n32592) );
  IV U34922 ( .A(n33689), .Z(n33691) );
  XOR U34923 ( .A(n33689), .B(n32593), .Z(n33690) );
  XNOR U34924 ( .A(n33692), .B(n33693), .Z(n32593) );
  ANDN U34925 ( .B(\modmult_1/xin[1023] ), .A(n33694), .Z(n33692) );
  IV U34926 ( .A(n33693), .Z(n33694) );
  XNOR U34927 ( .A(m[923]), .B(n33695), .Z(n33693) );
  NAND U34928 ( .A(n33696), .B(mul_pow), .Z(n33695) );
  XOR U34929 ( .A(m[923]), .B(c[923]), .Z(n33696) );
  XOR U34930 ( .A(n33697), .B(n33698), .Z(n33689) );
  ANDN U34931 ( .B(n33699), .A(n32590), .Z(n33697) );
  XNOR U34932 ( .A(\modmult_1/zin[0][921] ), .B(n33700), .Z(n32590) );
  IV U34933 ( .A(n33698), .Z(n33700) );
  XOR U34934 ( .A(n33698), .B(n32591), .Z(n33699) );
  XNOR U34935 ( .A(n33701), .B(n33702), .Z(n32591) );
  ANDN U34936 ( .B(\modmult_1/xin[1023] ), .A(n33703), .Z(n33701) );
  IV U34937 ( .A(n33702), .Z(n33703) );
  XNOR U34938 ( .A(m[922]), .B(n33704), .Z(n33702) );
  NAND U34939 ( .A(n33705), .B(mul_pow), .Z(n33704) );
  XOR U34940 ( .A(m[922]), .B(c[922]), .Z(n33705) );
  XOR U34941 ( .A(n33706), .B(n33707), .Z(n33698) );
  ANDN U34942 ( .B(n33708), .A(n32588), .Z(n33706) );
  XNOR U34943 ( .A(\modmult_1/zin[0][920] ), .B(n33709), .Z(n32588) );
  IV U34944 ( .A(n33707), .Z(n33709) );
  XOR U34945 ( .A(n33707), .B(n32589), .Z(n33708) );
  XNOR U34946 ( .A(n33710), .B(n33711), .Z(n32589) );
  ANDN U34947 ( .B(\modmult_1/xin[1023] ), .A(n33712), .Z(n33710) );
  IV U34948 ( .A(n33711), .Z(n33712) );
  XNOR U34949 ( .A(m[921]), .B(n33713), .Z(n33711) );
  NAND U34950 ( .A(n33714), .B(mul_pow), .Z(n33713) );
  XOR U34951 ( .A(m[921]), .B(c[921]), .Z(n33714) );
  XOR U34952 ( .A(n33715), .B(n33716), .Z(n33707) );
  ANDN U34953 ( .B(n33717), .A(n32586), .Z(n33715) );
  XNOR U34954 ( .A(\modmult_1/zin[0][919] ), .B(n33718), .Z(n32586) );
  IV U34955 ( .A(n33716), .Z(n33718) );
  XOR U34956 ( .A(n33716), .B(n32587), .Z(n33717) );
  XNOR U34957 ( .A(n33719), .B(n33720), .Z(n32587) );
  ANDN U34958 ( .B(\modmult_1/xin[1023] ), .A(n33721), .Z(n33719) );
  IV U34959 ( .A(n33720), .Z(n33721) );
  XNOR U34960 ( .A(m[920]), .B(n33722), .Z(n33720) );
  NAND U34961 ( .A(n33723), .B(mul_pow), .Z(n33722) );
  XOR U34962 ( .A(m[920]), .B(c[920]), .Z(n33723) );
  XOR U34963 ( .A(n33724), .B(n33725), .Z(n33716) );
  ANDN U34964 ( .B(n33726), .A(n32584), .Z(n33724) );
  XNOR U34965 ( .A(\modmult_1/zin[0][918] ), .B(n33727), .Z(n32584) );
  IV U34966 ( .A(n33725), .Z(n33727) );
  XOR U34967 ( .A(n33725), .B(n32585), .Z(n33726) );
  XNOR U34968 ( .A(n33728), .B(n33729), .Z(n32585) );
  ANDN U34969 ( .B(\modmult_1/xin[1023] ), .A(n33730), .Z(n33728) );
  IV U34970 ( .A(n33729), .Z(n33730) );
  XNOR U34971 ( .A(m[919]), .B(n33731), .Z(n33729) );
  NAND U34972 ( .A(n33732), .B(mul_pow), .Z(n33731) );
  XOR U34973 ( .A(m[919]), .B(c[919]), .Z(n33732) );
  XOR U34974 ( .A(n33733), .B(n33734), .Z(n33725) );
  ANDN U34975 ( .B(n33735), .A(n32582), .Z(n33733) );
  XNOR U34976 ( .A(\modmult_1/zin[0][917] ), .B(n33736), .Z(n32582) );
  IV U34977 ( .A(n33734), .Z(n33736) );
  XOR U34978 ( .A(n33734), .B(n32583), .Z(n33735) );
  XNOR U34979 ( .A(n33737), .B(n33738), .Z(n32583) );
  ANDN U34980 ( .B(\modmult_1/xin[1023] ), .A(n33739), .Z(n33737) );
  IV U34981 ( .A(n33738), .Z(n33739) );
  XNOR U34982 ( .A(m[918]), .B(n33740), .Z(n33738) );
  NAND U34983 ( .A(n33741), .B(mul_pow), .Z(n33740) );
  XOR U34984 ( .A(m[918]), .B(c[918]), .Z(n33741) );
  XOR U34985 ( .A(n33742), .B(n33743), .Z(n33734) );
  ANDN U34986 ( .B(n33744), .A(n32580), .Z(n33742) );
  XNOR U34987 ( .A(\modmult_1/zin[0][916] ), .B(n33745), .Z(n32580) );
  IV U34988 ( .A(n33743), .Z(n33745) );
  XOR U34989 ( .A(n33743), .B(n32581), .Z(n33744) );
  XNOR U34990 ( .A(n33746), .B(n33747), .Z(n32581) );
  ANDN U34991 ( .B(\modmult_1/xin[1023] ), .A(n33748), .Z(n33746) );
  IV U34992 ( .A(n33747), .Z(n33748) );
  XNOR U34993 ( .A(m[917]), .B(n33749), .Z(n33747) );
  NAND U34994 ( .A(n33750), .B(mul_pow), .Z(n33749) );
  XOR U34995 ( .A(m[917]), .B(c[917]), .Z(n33750) );
  XOR U34996 ( .A(n33751), .B(n33752), .Z(n33743) );
  ANDN U34997 ( .B(n33753), .A(n32578), .Z(n33751) );
  XNOR U34998 ( .A(\modmult_1/zin[0][915] ), .B(n33754), .Z(n32578) );
  IV U34999 ( .A(n33752), .Z(n33754) );
  XOR U35000 ( .A(n33752), .B(n32579), .Z(n33753) );
  XNOR U35001 ( .A(n33755), .B(n33756), .Z(n32579) );
  ANDN U35002 ( .B(\modmult_1/xin[1023] ), .A(n33757), .Z(n33755) );
  IV U35003 ( .A(n33756), .Z(n33757) );
  XNOR U35004 ( .A(m[916]), .B(n33758), .Z(n33756) );
  NAND U35005 ( .A(n33759), .B(mul_pow), .Z(n33758) );
  XOR U35006 ( .A(m[916]), .B(c[916]), .Z(n33759) );
  XOR U35007 ( .A(n33760), .B(n33761), .Z(n33752) );
  ANDN U35008 ( .B(n33762), .A(n32576), .Z(n33760) );
  XNOR U35009 ( .A(\modmult_1/zin[0][914] ), .B(n33763), .Z(n32576) );
  IV U35010 ( .A(n33761), .Z(n33763) );
  XOR U35011 ( .A(n33761), .B(n32577), .Z(n33762) );
  XNOR U35012 ( .A(n33764), .B(n33765), .Z(n32577) );
  ANDN U35013 ( .B(\modmult_1/xin[1023] ), .A(n33766), .Z(n33764) );
  IV U35014 ( .A(n33765), .Z(n33766) );
  XNOR U35015 ( .A(m[915]), .B(n33767), .Z(n33765) );
  NAND U35016 ( .A(n33768), .B(mul_pow), .Z(n33767) );
  XOR U35017 ( .A(m[915]), .B(c[915]), .Z(n33768) );
  XOR U35018 ( .A(n33769), .B(n33770), .Z(n33761) );
  ANDN U35019 ( .B(n33771), .A(n32574), .Z(n33769) );
  XNOR U35020 ( .A(\modmult_1/zin[0][913] ), .B(n33772), .Z(n32574) );
  IV U35021 ( .A(n33770), .Z(n33772) );
  XOR U35022 ( .A(n33770), .B(n32575), .Z(n33771) );
  XNOR U35023 ( .A(n33773), .B(n33774), .Z(n32575) );
  ANDN U35024 ( .B(\modmult_1/xin[1023] ), .A(n33775), .Z(n33773) );
  IV U35025 ( .A(n33774), .Z(n33775) );
  XNOR U35026 ( .A(m[914]), .B(n33776), .Z(n33774) );
  NAND U35027 ( .A(n33777), .B(mul_pow), .Z(n33776) );
  XOR U35028 ( .A(m[914]), .B(c[914]), .Z(n33777) );
  XOR U35029 ( .A(n33778), .B(n33779), .Z(n33770) );
  ANDN U35030 ( .B(n33780), .A(n32572), .Z(n33778) );
  XNOR U35031 ( .A(\modmult_1/zin[0][912] ), .B(n33781), .Z(n32572) );
  IV U35032 ( .A(n33779), .Z(n33781) );
  XOR U35033 ( .A(n33779), .B(n32573), .Z(n33780) );
  XNOR U35034 ( .A(n33782), .B(n33783), .Z(n32573) );
  ANDN U35035 ( .B(\modmult_1/xin[1023] ), .A(n33784), .Z(n33782) );
  IV U35036 ( .A(n33783), .Z(n33784) );
  XNOR U35037 ( .A(m[913]), .B(n33785), .Z(n33783) );
  NAND U35038 ( .A(n33786), .B(mul_pow), .Z(n33785) );
  XOR U35039 ( .A(m[913]), .B(c[913]), .Z(n33786) );
  XOR U35040 ( .A(n33787), .B(n33788), .Z(n33779) );
  ANDN U35041 ( .B(n33789), .A(n32570), .Z(n33787) );
  XNOR U35042 ( .A(\modmult_1/zin[0][911] ), .B(n33790), .Z(n32570) );
  IV U35043 ( .A(n33788), .Z(n33790) );
  XOR U35044 ( .A(n33788), .B(n32571), .Z(n33789) );
  XNOR U35045 ( .A(n33791), .B(n33792), .Z(n32571) );
  ANDN U35046 ( .B(\modmult_1/xin[1023] ), .A(n33793), .Z(n33791) );
  IV U35047 ( .A(n33792), .Z(n33793) );
  XNOR U35048 ( .A(m[912]), .B(n33794), .Z(n33792) );
  NAND U35049 ( .A(n33795), .B(mul_pow), .Z(n33794) );
  XOR U35050 ( .A(m[912]), .B(c[912]), .Z(n33795) );
  XOR U35051 ( .A(n33796), .B(n33797), .Z(n33788) );
  ANDN U35052 ( .B(n33798), .A(n32568), .Z(n33796) );
  XNOR U35053 ( .A(\modmult_1/zin[0][910] ), .B(n33799), .Z(n32568) );
  IV U35054 ( .A(n33797), .Z(n33799) );
  XOR U35055 ( .A(n33797), .B(n32569), .Z(n33798) );
  XNOR U35056 ( .A(n33800), .B(n33801), .Z(n32569) );
  ANDN U35057 ( .B(\modmult_1/xin[1023] ), .A(n33802), .Z(n33800) );
  IV U35058 ( .A(n33801), .Z(n33802) );
  XNOR U35059 ( .A(m[911]), .B(n33803), .Z(n33801) );
  NAND U35060 ( .A(n33804), .B(mul_pow), .Z(n33803) );
  XOR U35061 ( .A(m[911]), .B(c[911]), .Z(n33804) );
  XOR U35062 ( .A(n33805), .B(n33806), .Z(n33797) );
  ANDN U35063 ( .B(n33807), .A(n32566), .Z(n33805) );
  XNOR U35064 ( .A(\modmult_1/zin[0][909] ), .B(n33808), .Z(n32566) );
  IV U35065 ( .A(n33806), .Z(n33808) );
  XOR U35066 ( .A(n33806), .B(n32567), .Z(n33807) );
  XNOR U35067 ( .A(n33809), .B(n33810), .Z(n32567) );
  ANDN U35068 ( .B(\modmult_1/xin[1023] ), .A(n33811), .Z(n33809) );
  IV U35069 ( .A(n33810), .Z(n33811) );
  XNOR U35070 ( .A(m[910]), .B(n33812), .Z(n33810) );
  NAND U35071 ( .A(n33813), .B(mul_pow), .Z(n33812) );
  XOR U35072 ( .A(m[910]), .B(c[910]), .Z(n33813) );
  XOR U35073 ( .A(n33814), .B(n33815), .Z(n33806) );
  ANDN U35074 ( .B(n33816), .A(n32564), .Z(n33814) );
  XNOR U35075 ( .A(\modmult_1/zin[0][908] ), .B(n33817), .Z(n32564) );
  IV U35076 ( .A(n33815), .Z(n33817) );
  XOR U35077 ( .A(n33815), .B(n32565), .Z(n33816) );
  XNOR U35078 ( .A(n33818), .B(n33819), .Z(n32565) );
  ANDN U35079 ( .B(\modmult_1/xin[1023] ), .A(n33820), .Z(n33818) );
  IV U35080 ( .A(n33819), .Z(n33820) );
  XNOR U35081 ( .A(m[909]), .B(n33821), .Z(n33819) );
  NAND U35082 ( .A(n33822), .B(mul_pow), .Z(n33821) );
  XOR U35083 ( .A(m[909]), .B(c[909]), .Z(n33822) );
  XOR U35084 ( .A(n33823), .B(n33824), .Z(n33815) );
  ANDN U35085 ( .B(n33825), .A(n32562), .Z(n33823) );
  XNOR U35086 ( .A(\modmult_1/zin[0][907] ), .B(n33826), .Z(n32562) );
  IV U35087 ( .A(n33824), .Z(n33826) );
  XOR U35088 ( .A(n33824), .B(n32563), .Z(n33825) );
  XNOR U35089 ( .A(n33827), .B(n33828), .Z(n32563) );
  ANDN U35090 ( .B(\modmult_1/xin[1023] ), .A(n33829), .Z(n33827) );
  IV U35091 ( .A(n33828), .Z(n33829) );
  XNOR U35092 ( .A(m[908]), .B(n33830), .Z(n33828) );
  NAND U35093 ( .A(n33831), .B(mul_pow), .Z(n33830) );
  XOR U35094 ( .A(m[908]), .B(c[908]), .Z(n33831) );
  XOR U35095 ( .A(n33832), .B(n33833), .Z(n33824) );
  ANDN U35096 ( .B(n33834), .A(n32560), .Z(n33832) );
  XNOR U35097 ( .A(\modmult_1/zin[0][906] ), .B(n33835), .Z(n32560) );
  IV U35098 ( .A(n33833), .Z(n33835) );
  XOR U35099 ( .A(n33833), .B(n32561), .Z(n33834) );
  XNOR U35100 ( .A(n33836), .B(n33837), .Z(n32561) );
  ANDN U35101 ( .B(\modmult_1/xin[1023] ), .A(n33838), .Z(n33836) );
  IV U35102 ( .A(n33837), .Z(n33838) );
  XNOR U35103 ( .A(m[907]), .B(n33839), .Z(n33837) );
  NAND U35104 ( .A(n33840), .B(mul_pow), .Z(n33839) );
  XOR U35105 ( .A(m[907]), .B(c[907]), .Z(n33840) );
  XOR U35106 ( .A(n33841), .B(n33842), .Z(n33833) );
  ANDN U35107 ( .B(n33843), .A(n32558), .Z(n33841) );
  XNOR U35108 ( .A(\modmult_1/zin[0][905] ), .B(n33844), .Z(n32558) );
  IV U35109 ( .A(n33842), .Z(n33844) );
  XOR U35110 ( .A(n33842), .B(n32559), .Z(n33843) );
  XNOR U35111 ( .A(n33845), .B(n33846), .Z(n32559) );
  ANDN U35112 ( .B(\modmult_1/xin[1023] ), .A(n33847), .Z(n33845) );
  IV U35113 ( .A(n33846), .Z(n33847) );
  XNOR U35114 ( .A(m[906]), .B(n33848), .Z(n33846) );
  NAND U35115 ( .A(n33849), .B(mul_pow), .Z(n33848) );
  XOR U35116 ( .A(m[906]), .B(c[906]), .Z(n33849) );
  XOR U35117 ( .A(n33850), .B(n33851), .Z(n33842) );
  ANDN U35118 ( .B(n33852), .A(n32556), .Z(n33850) );
  XNOR U35119 ( .A(\modmult_1/zin[0][904] ), .B(n33853), .Z(n32556) );
  IV U35120 ( .A(n33851), .Z(n33853) );
  XOR U35121 ( .A(n33851), .B(n32557), .Z(n33852) );
  XNOR U35122 ( .A(n33854), .B(n33855), .Z(n32557) );
  ANDN U35123 ( .B(\modmult_1/xin[1023] ), .A(n33856), .Z(n33854) );
  IV U35124 ( .A(n33855), .Z(n33856) );
  XNOR U35125 ( .A(m[905]), .B(n33857), .Z(n33855) );
  NAND U35126 ( .A(n33858), .B(mul_pow), .Z(n33857) );
  XOR U35127 ( .A(m[905]), .B(c[905]), .Z(n33858) );
  XOR U35128 ( .A(n33859), .B(n33860), .Z(n33851) );
  ANDN U35129 ( .B(n33861), .A(n32554), .Z(n33859) );
  XNOR U35130 ( .A(\modmult_1/zin[0][903] ), .B(n33862), .Z(n32554) );
  IV U35131 ( .A(n33860), .Z(n33862) );
  XOR U35132 ( .A(n33860), .B(n32555), .Z(n33861) );
  XNOR U35133 ( .A(n33863), .B(n33864), .Z(n32555) );
  ANDN U35134 ( .B(\modmult_1/xin[1023] ), .A(n33865), .Z(n33863) );
  IV U35135 ( .A(n33864), .Z(n33865) );
  XNOR U35136 ( .A(m[904]), .B(n33866), .Z(n33864) );
  NAND U35137 ( .A(n33867), .B(mul_pow), .Z(n33866) );
  XOR U35138 ( .A(m[904]), .B(c[904]), .Z(n33867) );
  XOR U35139 ( .A(n33868), .B(n33869), .Z(n33860) );
  ANDN U35140 ( .B(n33870), .A(n32552), .Z(n33868) );
  XNOR U35141 ( .A(\modmult_1/zin[0][902] ), .B(n33871), .Z(n32552) );
  IV U35142 ( .A(n33869), .Z(n33871) );
  XOR U35143 ( .A(n33869), .B(n32553), .Z(n33870) );
  XNOR U35144 ( .A(n33872), .B(n33873), .Z(n32553) );
  ANDN U35145 ( .B(\modmult_1/xin[1023] ), .A(n33874), .Z(n33872) );
  IV U35146 ( .A(n33873), .Z(n33874) );
  XNOR U35147 ( .A(m[903]), .B(n33875), .Z(n33873) );
  NAND U35148 ( .A(n33876), .B(mul_pow), .Z(n33875) );
  XOR U35149 ( .A(m[903]), .B(c[903]), .Z(n33876) );
  XOR U35150 ( .A(n33877), .B(n33878), .Z(n33869) );
  ANDN U35151 ( .B(n33879), .A(n32550), .Z(n33877) );
  XNOR U35152 ( .A(\modmult_1/zin[0][901] ), .B(n33880), .Z(n32550) );
  IV U35153 ( .A(n33878), .Z(n33880) );
  XOR U35154 ( .A(n33878), .B(n32551), .Z(n33879) );
  XNOR U35155 ( .A(n33881), .B(n33882), .Z(n32551) );
  ANDN U35156 ( .B(\modmult_1/xin[1023] ), .A(n33883), .Z(n33881) );
  IV U35157 ( .A(n33882), .Z(n33883) );
  XNOR U35158 ( .A(m[902]), .B(n33884), .Z(n33882) );
  NAND U35159 ( .A(n33885), .B(mul_pow), .Z(n33884) );
  XOR U35160 ( .A(m[902]), .B(c[902]), .Z(n33885) );
  XOR U35161 ( .A(n33886), .B(n33887), .Z(n33878) );
  ANDN U35162 ( .B(n33888), .A(n32548), .Z(n33886) );
  XNOR U35163 ( .A(\modmult_1/zin[0][900] ), .B(n33889), .Z(n32548) );
  IV U35164 ( .A(n33887), .Z(n33889) );
  XOR U35165 ( .A(n33887), .B(n32549), .Z(n33888) );
  XNOR U35166 ( .A(n33890), .B(n33891), .Z(n32549) );
  ANDN U35167 ( .B(\modmult_1/xin[1023] ), .A(n33892), .Z(n33890) );
  IV U35168 ( .A(n33891), .Z(n33892) );
  XNOR U35169 ( .A(m[901]), .B(n33893), .Z(n33891) );
  NAND U35170 ( .A(n33894), .B(mul_pow), .Z(n33893) );
  XOR U35171 ( .A(m[901]), .B(c[901]), .Z(n33894) );
  XOR U35172 ( .A(n33895), .B(n33896), .Z(n33887) );
  ANDN U35173 ( .B(n33897), .A(n32546), .Z(n33895) );
  XNOR U35174 ( .A(\modmult_1/zin[0][899] ), .B(n33898), .Z(n32546) );
  IV U35175 ( .A(n33896), .Z(n33898) );
  XOR U35176 ( .A(n33896), .B(n32547), .Z(n33897) );
  XNOR U35177 ( .A(n33899), .B(n33900), .Z(n32547) );
  ANDN U35178 ( .B(\modmult_1/xin[1023] ), .A(n33901), .Z(n33899) );
  IV U35179 ( .A(n33900), .Z(n33901) );
  XNOR U35180 ( .A(m[900]), .B(n33902), .Z(n33900) );
  NAND U35181 ( .A(n33903), .B(mul_pow), .Z(n33902) );
  XOR U35182 ( .A(m[900]), .B(c[900]), .Z(n33903) );
  XOR U35183 ( .A(n33904), .B(n33905), .Z(n33896) );
  ANDN U35184 ( .B(n33906), .A(n32544), .Z(n33904) );
  XNOR U35185 ( .A(\modmult_1/zin[0][898] ), .B(n33907), .Z(n32544) );
  IV U35186 ( .A(n33905), .Z(n33907) );
  XOR U35187 ( .A(n33905), .B(n32545), .Z(n33906) );
  XNOR U35188 ( .A(n33908), .B(n33909), .Z(n32545) );
  ANDN U35189 ( .B(\modmult_1/xin[1023] ), .A(n33910), .Z(n33908) );
  IV U35190 ( .A(n33909), .Z(n33910) );
  XNOR U35191 ( .A(m[899]), .B(n33911), .Z(n33909) );
  NAND U35192 ( .A(n33912), .B(mul_pow), .Z(n33911) );
  XOR U35193 ( .A(m[899]), .B(c[899]), .Z(n33912) );
  XOR U35194 ( .A(n33913), .B(n33914), .Z(n33905) );
  ANDN U35195 ( .B(n33915), .A(n32542), .Z(n33913) );
  XNOR U35196 ( .A(\modmult_1/zin[0][897] ), .B(n33916), .Z(n32542) );
  IV U35197 ( .A(n33914), .Z(n33916) );
  XOR U35198 ( .A(n33914), .B(n32543), .Z(n33915) );
  XNOR U35199 ( .A(n33917), .B(n33918), .Z(n32543) );
  ANDN U35200 ( .B(\modmult_1/xin[1023] ), .A(n33919), .Z(n33917) );
  IV U35201 ( .A(n33918), .Z(n33919) );
  XNOR U35202 ( .A(m[898]), .B(n33920), .Z(n33918) );
  NAND U35203 ( .A(n33921), .B(mul_pow), .Z(n33920) );
  XOR U35204 ( .A(m[898]), .B(c[898]), .Z(n33921) );
  XOR U35205 ( .A(n33922), .B(n33923), .Z(n33914) );
  ANDN U35206 ( .B(n33924), .A(n32540), .Z(n33922) );
  XNOR U35207 ( .A(\modmult_1/zin[0][896] ), .B(n33925), .Z(n32540) );
  IV U35208 ( .A(n33923), .Z(n33925) );
  XOR U35209 ( .A(n33923), .B(n32541), .Z(n33924) );
  XNOR U35210 ( .A(n33926), .B(n33927), .Z(n32541) );
  ANDN U35211 ( .B(\modmult_1/xin[1023] ), .A(n33928), .Z(n33926) );
  IV U35212 ( .A(n33927), .Z(n33928) );
  XNOR U35213 ( .A(m[897]), .B(n33929), .Z(n33927) );
  NAND U35214 ( .A(n33930), .B(mul_pow), .Z(n33929) );
  XOR U35215 ( .A(m[897]), .B(c[897]), .Z(n33930) );
  XOR U35216 ( .A(n33931), .B(n33932), .Z(n33923) );
  ANDN U35217 ( .B(n33933), .A(n32538), .Z(n33931) );
  XNOR U35218 ( .A(\modmult_1/zin[0][895] ), .B(n33934), .Z(n32538) );
  IV U35219 ( .A(n33932), .Z(n33934) );
  XOR U35220 ( .A(n33932), .B(n32539), .Z(n33933) );
  XNOR U35221 ( .A(n33935), .B(n33936), .Z(n32539) );
  ANDN U35222 ( .B(\modmult_1/xin[1023] ), .A(n33937), .Z(n33935) );
  IV U35223 ( .A(n33936), .Z(n33937) );
  XNOR U35224 ( .A(m[896]), .B(n33938), .Z(n33936) );
  NAND U35225 ( .A(n33939), .B(mul_pow), .Z(n33938) );
  XOR U35226 ( .A(m[896]), .B(c[896]), .Z(n33939) );
  XOR U35227 ( .A(n33940), .B(n33941), .Z(n33932) );
  ANDN U35228 ( .B(n33942), .A(n32536), .Z(n33940) );
  XNOR U35229 ( .A(\modmult_1/zin[0][894] ), .B(n33943), .Z(n32536) );
  IV U35230 ( .A(n33941), .Z(n33943) );
  XOR U35231 ( .A(n33941), .B(n32537), .Z(n33942) );
  XNOR U35232 ( .A(n33944), .B(n33945), .Z(n32537) );
  ANDN U35233 ( .B(\modmult_1/xin[1023] ), .A(n33946), .Z(n33944) );
  IV U35234 ( .A(n33945), .Z(n33946) );
  XNOR U35235 ( .A(m[895]), .B(n33947), .Z(n33945) );
  NAND U35236 ( .A(n33948), .B(mul_pow), .Z(n33947) );
  XOR U35237 ( .A(m[895]), .B(c[895]), .Z(n33948) );
  XOR U35238 ( .A(n33949), .B(n33950), .Z(n33941) );
  ANDN U35239 ( .B(n33951), .A(n32534), .Z(n33949) );
  XNOR U35240 ( .A(\modmult_1/zin[0][893] ), .B(n33952), .Z(n32534) );
  IV U35241 ( .A(n33950), .Z(n33952) );
  XOR U35242 ( .A(n33950), .B(n32535), .Z(n33951) );
  XNOR U35243 ( .A(n33953), .B(n33954), .Z(n32535) );
  ANDN U35244 ( .B(\modmult_1/xin[1023] ), .A(n33955), .Z(n33953) );
  IV U35245 ( .A(n33954), .Z(n33955) );
  XNOR U35246 ( .A(m[894]), .B(n33956), .Z(n33954) );
  NAND U35247 ( .A(n33957), .B(mul_pow), .Z(n33956) );
  XOR U35248 ( .A(m[894]), .B(c[894]), .Z(n33957) );
  XOR U35249 ( .A(n33958), .B(n33959), .Z(n33950) );
  ANDN U35250 ( .B(n33960), .A(n32532), .Z(n33958) );
  XNOR U35251 ( .A(\modmult_1/zin[0][892] ), .B(n33961), .Z(n32532) );
  IV U35252 ( .A(n33959), .Z(n33961) );
  XOR U35253 ( .A(n33959), .B(n32533), .Z(n33960) );
  XNOR U35254 ( .A(n33962), .B(n33963), .Z(n32533) );
  ANDN U35255 ( .B(\modmult_1/xin[1023] ), .A(n33964), .Z(n33962) );
  IV U35256 ( .A(n33963), .Z(n33964) );
  XNOR U35257 ( .A(m[893]), .B(n33965), .Z(n33963) );
  NAND U35258 ( .A(n33966), .B(mul_pow), .Z(n33965) );
  XOR U35259 ( .A(m[893]), .B(c[893]), .Z(n33966) );
  XOR U35260 ( .A(n33967), .B(n33968), .Z(n33959) );
  ANDN U35261 ( .B(n33969), .A(n32530), .Z(n33967) );
  XNOR U35262 ( .A(\modmult_1/zin[0][891] ), .B(n33970), .Z(n32530) );
  IV U35263 ( .A(n33968), .Z(n33970) );
  XOR U35264 ( .A(n33968), .B(n32531), .Z(n33969) );
  XNOR U35265 ( .A(n33971), .B(n33972), .Z(n32531) );
  ANDN U35266 ( .B(\modmult_1/xin[1023] ), .A(n33973), .Z(n33971) );
  IV U35267 ( .A(n33972), .Z(n33973) );
  XNOR U35268 ( .A(m[892]), .B(n33974), .Z(n33972) );
  NAND U35269 ( .A(n33975), .B(mul_pow), .Z(n33974) );
  XOR U35270 ( .A(m[892]), .B(c[892]), .Z(n33975) );
  XOR U35271 ( .A(n33976), .B(n33977), .Z(n33968) );
  ANDN U35272 ( .B(n33978), .A(n32528), .Z(n33976) );
  XNOR U35273 ( .A(\modmult_1/zin[0][890] ), .B(n33979), .Z(n32528) );
  IV U35274 ( .A(n33977), .Z(n33979) );
  XOR U35275 ( .A(n33977), .B(n32529), .Z(n33978) );
  XNOR U35276 ( .A(n33980), .B(n33981), .Z(n32529) );
  ANDN U35277 ( .B(\modmult_1/xin[1023] ), .A(n33982), .Z(n33980) );
  IV U35278 ( .A(n33981), .Z(n33982) );
  XNOR U35279 ( .A(m[891]), .B(n33983), .Z(n33981) );
  NAND U35280 ( .A(n33984), .B(mul_pow), .Z(n33983) );
  XOR U35281 ( .A(m[891]), .B(c[891]), .Z(n33984) );
  XOR U35282 ( .A(n33985), .B(n33986), .Z(n33977) );
  ANDN U35283 ( .B(n33987), .A(n32526), .Z(n33985) );
  XNOR U35284 ( .A(\modmult_1/zin[0][889] ), .B(n33988), .Z(n32526) );
  IV U35285 ( .A(n33986), .Z(n33988) );
  XOR U35286 ( .A(n33986), .B(n32527), .Z(n33987) );
  XNOR U35287 ( .A(n33989), .B(n33990), .Z(n32527) );
  ANDN U35288 ( .B(\modmult_1/xin[1023] ), .A(n33991), .Z(n33989) );
  IV U35289 ( .A(n33990), .Z(n33991) );
  XNOR U35290 ( .A(m[890]), .B(n33992), .Z(n33990) );
  NAND U35291 ( .A(n33993), .B(mul_pow), .Z(n33992) );
  XOR U35292 ( .A(m[890]), .B(c[890]), .Z(n33993) );
  XOR U35293 ( .A(n33994), .B(n33995), .Z(n33986) );
  ANDN U35294 ( .B(n33996), .A(n32524), .Z(n33994) );
  XNOR U35295 ( .A(\modmult_1/zin[0][888] ), .B(n33997), .Z(n32524) );
  IV U35296 ( .A(n33995), .Z(n33997) );
  XOR U35297 ( .A(n33995), .B(n32525), .Z(n33996) );
  XNOR U35298 ( .A(n33998), .B(n33999), .Z(n32525) );
  ANDN U35299 ( .B(\modmult_1/xin[1023] ), .A(n34000), .Z(n33998) );
  IV U35300 ( .A(n33999), .Z(n34000) );
  XNOR U35301 ( .A(m[889]), .B(n34001), .Z(n33999) );
  NAND U35302 ( .A(n34002), .B(mul_pow), .Z(n34001) );
  XOR U35303 ( .A(m[889]), .B(c[889]), .Z(n34002) );
  XOR U35304 ( .A(n34003), .B(n34004), .Z(n33995) );
  ANDN U35305 ( .B(n34005), .A(n32522), .Z(n34003) );
  XNOR U35306 ( .A(\modmult_1/zin[0][887] ), .B(n34006), .Z(n32522) );
  IV U35307 ( .A(n34004), .Z(n34006) );
  XOR U35308 ( .A(n34004), .B(n32523), .Z(n34005) );
  XNOR U35309 ( .A(n34007), .B(n34008), .Z(n32523) );
  ANDN U35310 ( .B(\modmult_1/xin[1023] ), .A(n34009), .Z(n34007) );
  IV U35311 ( .A(n34008), .Z(n34009) );
  XNOR U35312 ( .A(m[888]), .B(n34010), .Z(n34008) );
  NAND U35313 ( .A(n34011), .B(mul_pow), .Z(n34010) );
  XOR U35314 ( .A(m[888]), .B(c[888]), .Z(n34011) );
  XOR U35315 ( .A(n34012), .B(n34013), .Z(n34004) );
  ANDN U35316 ( .B(n34014), .A(n32520), .Z(n34012) );
  XNOR U35317 ( .A(\modmult_1/zin[0][886] ), .B(n34015), .Z(n32520) );
  IV U35318 ( .A(n34013), .Z(n34015) );
  XOR U35319 ( .A(n34013), .B(n32521), .Z(n34014) );
  XNOR U35320 ( .A(n34016), .B(n34017), .Z(n32521) );
  ANDN U35321 ( .B(\modmult_1/xin[1023] ), .A(n34018), .Z(n34016) );
  IV U35322 ( .A(n34017), .Z(n34018) );
  XNOR U35323 ( .A(m[887]), .B(n34019), .Z(n34017) );
  NAND U35324 ( .A(n34020), .B(mul_pow), .Z(n34019) );
  XOR U35325 ( .A(m[887]), .B(c[887]), .Z(n34020) );
  XOR U35326 ( .A(n34021), .B(n34022), .Z(n34013) );
  ANDN U35327 ( .B(n34023), .A(n32518), .Z(n34021) );
  XNOR U35328 ( .A(\modmult_1/zin[0][885] ), .B(n34024), .Z(n32518) );
  IV U35329 ( .A(n34022), .Z(n34024) );
  XOR U35330 ( .A(n34022), .B(n32519), .Z(n34023) );
  XNOR U35331 ( .A(n34025), .B(n34026), .Z(n32519) );
  ANDN U35332 ( .B(\modmult_1/xin[1023] ), .A(n34027), .Z(n34025) );
  IV U35333 ( .A(n34026), .Z(n34027) );
  XNOR U35334 ( .A(m[886]), .B(n34028), .Z(n34026) );
  NAND U35335 ( .A(n34029), .B(mul_pow), .Z(n34028) );
  XOR U35336 ( .A(m[886]), .B(c[886]), .Z(n34029) );
  XOR U35337 ( .A(n34030), .B(n34031), .Z(n34022) );
  ANDN U35338 ( .B(n34032), .A(n32516), .Z(n34030) );
  XNOR U35339 ( .A(\modmult_1/zin[0][884] ), .B(n34033), .Z(n32516) );
  IV U35340 ( .A(n34031), .Z(n34033) );
  XOR U35341 ( .A(n34031), .B(n32517), .Z(n34032) );
  XNOR U35342 ( .A(n34034), .B(n34035), .Z(n32517) );
  ANDN U35343 ( .B(\modmult_1/xin[1023] ), .A(n34036), .Z(n34034) );
  IV U35344 ( .A(n34035), .Z(n34036) );
  XNOR U35345 ( .A(m[885]), .B(n34037), .Z(n34035) );
  NAND U35346 ( .A(n34038), .B(mul_pow), .Z(n34037) );
  XOR U35347 ( .A(m[885]), .B(c[885]), .Z(n34038) );
  XOR U35348 ( .A(n34039), .B(n34040), .Z(n34031) );
  ANDN U35349 ( .B(n34041), .A(n32514), .Z(n34039) );
  XNOR U35350 ( .A(\modmult_1/zin[0][883] ), .B(n34042), .Z(n32514) );
  IV U35351 ( .A(n34040), .Z(n34042) );
  XOR U35352 ( .A(n34040), .B(n32515), .Z(n34041) );
  XNOR U35353 ( .A(n34043), .B(n34044), .Z(n32515) );
  ANDN U35354 ( .B(\modmult_1/xin[1023] ), .A(n34045), .Z(n34043) );
  IV U35355 ( .A(n34044), .Z(n34045) );
  XNOR U35356 ( .A(m[884]), .B(n34046), .Z(n34044) );
  NAND U35357 ( .A(n34047), .B(mul_pow), .Z(n34046) );
  XOR U35358 ( .A(m[884]), .B(c[884]), .Z(n34047) );
  XOR U35359 ( .A(n34048), .B(n34049), .Z(n34040) );
  ANDN U35360 ( .B(n34050), .A(n32512), .Z(n34048) );
  XNOR U35361 ( .A(\modmult_1/zin[0][882] ), .B(n34051), .Z(n32512) );
  IV U35362 ( .A(n34049), .Z(n34051) );
  XOR U35363 ( .A(n34049), .B(n32513), .Z(n34050) );
  XNOR U35364 ( .A(n34052), .B(n34053), .Z(n32513) );
  ANDN U35365 ( .B(\modmult_1/xin[1023] ), .A(n34054), .Z(n34052) );
  IV U35366 ( .A(n34053), .Z(n34054) );
  XNOR U35367 ( .A(m[883]), .B(n34055), .Z(n34053) );
  NAND U35368 ( .A(n34056), .B(mul_pow), .Z(n34055) );
  XOR U35369 ( .A(m[883]), .B(c[883]), .Z(n34056) );
  XOR U35370 ( .A(n34057), .B(n34058), .Z(n34049) );
  ANDN U35371 ( .B(n34059), .A(n32510), .Z(n34057) );
  XNOR U35372 ( .A(\modmult_1/zin[0][881] ), .B(n34060), .Z(n32510) );
  IV U35373 ( .A(n34058), .Z(n34060) );
  XOR U35374 ( .A(n34058), .B(n32511), .Z(n34059) );
  XNOR U35375 ( .A(n34061), .B(n34062), .Z(n32511) );
  ANDN U35376 ( .B(\modmult_1/xin[1023] ), .A(n34063), .Z(n34061) );
  IV U35377 ( .A(n34062), .Z(n34063) );
  XNOR U35378 ( .A(m[882]), .B(n34064), .Z(n34062) );
  NAND U35379 ( .A(n34065), .B(mul_pow), .Z(n34064) );
  XOR U35380 ( .A(m[882]), .B(c[882]), .Z(n34065) );
  XOR U35381 ( .A(n34066), .B(n34067), .Z(n34058) );
  ANDN U35382 ( .B(n34068), .A(n32508), .Z(n34066) );
  XNOR U35383 ( .A(\modmult_1/zin[0][880] ), .B(n34069), .Z(n32508) );
  IV U35384 ( .A(n34067), .Z(n34069) );
  XOR U35385 ( .A(n34067), .B(n32509), .Z(n34068) );
  XNOR U35386 ( .A(n34070), .B(n34071), .Z(n32509) );
  ANDN U35387 ( .B(\modmult_1/xin[1023] ), .A(n34072), .Z(n34070) );
  IV U35388 ( .A(n34071), .Z(n34072) );
  XNOR U35389 ( .A(m[881]), .B(n34073), .Z(n34071) );
  NAND U35390 ( .A(n34074), .B(mul_pow), .Z(n34073) );
  XOR U35391 ( .A(m[881]), .B(c[881]), .Z(n34074) );
  XOR U35392 ( .A(n34075), .B(n34076), .Z(n34067) );
  ANDN U35393 ( .B(n34077), .A(n32506), .Z(n34075) );
  XNOR U35394 ( .A(\modmult_1/zin[0][879] ), .B(n34078), .Z(n32506) );
  IV U35395 ( .A(n34076), .Z(n34078) );
  XOR U35396 ( .A(n34076), .B(n32507), .Z(n34077) );
  XNOR U35397 ( .A(n34079), .B(n34080), .Z(n32507) );
  ANDN U35398 ( .B(\modmult_1/xin[1023] ), .A(n34081), .Z(n34079) );
  IV U35399 ( .A(n34080), .Z(n34081) );
  XNOR U35400 ( .A(m[880]), .B(n34082), .Z(n34080) );
  NAND U35401 ( .A(n34083), .B(mul_pow), .Z(n34082) );
  XOR U35402 ( .A(m[880]), .B(c[880]), .Z(n34083) );
  XOR U35403 ( .A(n34084), .B(n34085), .Z(n34076) );
  ANDN U35404 ( .B(n34086), .A(n32504), .Z(n34084) );
  XNOR U35405 ( .A(\modmult_1/zin[0][878] ), .B(n34087), .Z(n32504) );
  IV U35406 ( .A(n34085), .Z(n34087) );
  XOR U35407 ( .A(n34085), .B(n32505), .Z(n34086) );
  XNOR U35408 ( .A(n34088), .B(n34089), .Z(n32505) );
  ANDN U35409 ( .B(\modmult_1/xin[1023] ), .A(n34090), .Z(n34088) );
  IV U35410 ( .A(n34089), .Z(n34090) );
  XNOR U35411 ( .A(m[879]), .B(n34091), .Z(n34089) );
  NAND U35412 ( .A(n34092), .B(mul_pow), .Z(n34091) );
  XOR U35413 ( .A(m[879]), .B(c[879]), .Z(n34092) );
  XOR U35414 ( .A(n34093), .B(n34094), .Z(n34085) );
  ANDN U35415 ( .B(n34095), .A(n32502), .Z(n34093) );
  XNOR U35416 ( .A(\modmult_1/zin[0][877] ), .B(n34096), .Z(n32502) );
  IV U35417 ( .A(n34094), .Z(n34096) );
  XOR U35418 ( .A(n34094), .B(n32503), .Z(n34095) );
  XNOR U35419 ( .A(n34097), .B(n34098), .Z(n32503) );
  ANDN U35420 ( .B(\modmult_1/xin[1023] ), .A(n34099), .Z(n34097) );
  IV U35421 ( .A(n34098), .Z(n34099) );
  XNOR U35422 ( .A(m[878]), .B(n34100), .Z(n34098) );
  NAND U35423 ( .A(n34101), .B(mul_pow), .Z(n34100) );
  XOR U35424 ( .A(m[878]), .B(c[878]), .Z(n34101) );
  XOR U35425 ( .A(n34102), .B(n34103), .Z(n34094) );
  ANDN U35426 ( .B(n34104), .A(n32500), .Z(n34102) );
  XNOR U35427 ( .A(\modmult_1/zin[0][876] ), .B(n34105), .Z(n32500) );
  IV U35428 ( .A(n34103), .Z(n34105) );
  XOR U35429 ( .A(n34103), .B(n32501), .Z(n34104) );
  XNOR U35430 ( .A(n34106), .B(n34107), .Z(n32501) );
  ANDN U35431 ( .B(\modmult_1/xin[1023] ), .A(n34108), .Z(n34106) );
  IV U35432 ( .A(n34107), .Z(n34108) );
  XNOR U35433 ( .A(m[877]), .B(n34109), .Z(n34107) );
  NAND U35434 ( .A(n34110), .B(mul_pow), .Z(n34109) );
  XOR U35435 ( .A(m[877]), .B(c[877]), .Z(n34110) );
  XOR U35436 ( .A(n34111), .B(n34112), .Z(n34103) );
  ANDN U35437 ( .B(n34113), .A(n32498), .Z(n34111) );
  XNOR U35438 ( .A(\modmult_1/zin[0][875] ), .B(n34114), .Z(n32498) );
  IV U35439 ( .A(n34112), .Z(n34114) );
  XOR U35440 ( .A(n34112), .B(n32499), .Z(n34113) );
  XNOR U35441 ( .A(n34115), .B(n34116), .Z(n32499) );
  ANDN U35442 ( .B(\modmult_1/xin[1023] ), .A(n34117), .Z(n34115) );
  IV U35443 ( .A(n34116), .Z(n34117) );
  XNOR U35444 ( .A(m[876]), .B(n34118), .Z(n34116) );
  NAND U35445 ( .A(n34119), .B(mul_pow), .Z(n34118) );
  XOR U35446 ( .A(m[876]), .B(c[876]), .Z(n34119) );
  XOR U35447 ( .A(n34120), .B(n34121), .Z(n34112) );
  ANDN U35448 ( .B(n34122), .A(n32496), .Z(n34120) );
  XNOR U35449 ( .A(\modmult_1/zin[0][874] ), .B(n34123), .Z(n32496) );
  IV U35450 ( .A(n34121), .Z(n34123) );
  XOR U35451 ( .A(n34121), .B(n32497), .Z(n34122) );
  XNOR U35452 ( .A(n34124), .B(n34125), .Z(n32497) );
  ANDN U35453 ( .B(\modmult_1/xin[1023] ), .A(n34126), .Z(n34124) );
  IV U35454 ( .A(n34125), .Z(n34126) );
  XNOR U35455 ( .A(m[875]), .B(n34127), .Z(n34125) );
  NAND U35456 ( .A(n34128), .B(mul_pow), .Z(n34127) );
  XOR U35457 ( .A(m[875]), .B(c[875]), .Z(n34128) );
  XOR U35458 ( .A(n34129), .B(n34130), .Z(n34121) );
  ANDN U35459 ( .B(n34131), .A(n32494), .Z(n34129) );
  XNOR U35460 ( .A(\modmult_1/zin[0][873] ), .B(n34132), .Z(n32494) );
  IV U35461 ( .A(n34130), .Z(n34132) );
  XOR U35462 ( .A(n34130), .B(n32495), .Z(n34131) );
  XNOR U35463 ( .A(n34133), .B(n34134), .Z(n32495) );
  ANDN U35464 ( .B(\modmult_1/xin[1023] ), .A(n34135), .Z(n34133) );
  IV U35465 ( .A(n34134), .Z(n34135) );
  XNOR U35466 ( .A(m[874]), .B(n34136), .Z(n34134) );
  NAND U35467 ( .A(n34137), .B(mul_pow), .Z(n34136) );
  XOR U35468 ( .A(m[874]), .B(c[874]), .Z(n34137) );
  XOR U35469 ( .A(n34138), .B(n34139), .Z(n34130) );
  ANDN U35470 ( .B(n34140), .A(n32492), .Z(n34138) );
  XNOR U35471 ( .A(\modmult_1/zin[0][872] ), .B(n34141), .Z(n32492) );
  IV U35472 ( .A(n34139), .Z(n34141) );
  XOR U35473 ( .A(n34139), .B(n32493), .Z(n34140) );
  XNOR U35474 ( .A(n34142), .B(n34143), .Z(n32493) );
  ANDN U35475 ( .B(\modmult_1/xin[1023] ), .A(n34144), .Z(n34142) );
  IV U35476 ( .A(n34143), .Z(n34144) );
  XNOR U35477 ( .A(m[873]), .B(n34145), .Z(n34143) );
  NAND U35478 ( .A(n34146), .B(mul_pow), .Z(n34145) );
  XOR U35479 ( .A(m[873]), .B(c[873]), .Z(n34146) );
  XOR U35480 ( .A(n34147), .B(n34148), .Z(n34139) );
  ANDN U35481 ( .B(n34149), .A(n32490), .Z(n34147) );
  XNOR U35482 ( .A(\modmult_1/zin[0][871] ), .B(n34150), .Z(n32490) );
  IV U35483 ( .A(n34148), .Z(n34150) );
  XOR U35484 ( .A(n34148), .B(n32491), .Z(n34149) );
  XNOR U35485 ( .A(n34151), .B(n34152), .Z(n32491) );
  ANDN U35486 ( .B(\modmult_1/xin[1023] ), .A(n34153), .Z(n34151) );
  IV U35487 ( .A(n34152), .Z(n34153) );
  XNOR U35488 ( .A(m[872]), .B(n34154), .Z(n34152) );
  NAND U35489 ( .A(n34155), .B(mul_pow), .Z(n34154) );
  XOR U35490 ( .A(m[872]), .B(c[872]), .Z(n34155) );
  XOR U35491 ( .A(n34156), .B(n34157), .Z(n34148) );
  ANDN U35492 ( .B(n34158), .A(n32488), .Z(n34156) );
  XNOR U35493 ( .A(\modmult_1/zin[0][870] ), .B(n34159), .Z(n32488) );
  IV U35494 ( .A(n34157), .Z(n34159) );
  XOR U35495 ( .A(n34157), .B(n32489), .Z(n34158) );
  XNOR U35496 ( .A(n34160), .B(n34161), .Z(n32489) );
  ANDN U35497 ( .B(\modmult_1/xin[1023] ), .A(n34162), .Z(n34160) );
  IV U35498 ( .A(n34161), .Z(n34162) );
  XNOR U35499 ( .A(m[871]), .B(n34163), .Z(n34161) );
  NAND U35500 ( .A(n34164), .B(mul_pow), .Z(n34163) );
  XOR U35501 ( .A(m[871]), .B(c[871]), .Z(n34164) );
  XOR U35502 ( .A(n34165), .B(n34166), .Z(n34157) );
  ANDN U35503 ( .B(n34167), .A(n32486), .Z(n34165) );
  XNOR U35504 ( .A(\modmult_1/zin[0][869] ), .B(n34168), .Z(n32486) );
  IV U35505 ( .A(n34166), .Z(n34168) );
  XOR U35506 ( .A(n34166), .B(n32487), .Z(n34167) );
  XNOR U35507 ( .A(n34169), .B(n34170), .Z(n32487) );
  ANDN U35508 ( .B(\modmult_1/xin[1023] ), .A(n34171), .Z(n34169) );
  IV U35509 ( .A(n34170), .Z(n34171) );
  XNOR U35510 ( .A(m[870]), .B(n34172), .Z(n34170) );
  NAND U35511 ( .A(n34173), .B(mul_pow), .Z(n34172) );
  XOR U35512 ( .A(m[870]), .B(c[870]), .Z(n34173) );
  XOR U35513 ( .A(n34174), .B(n34175), .Z(n34166) );
  ANDN U35514 ( .B(n34176), .A(n32484), .Z(n34174) );
  XNOR U35515 ( .A(\modmult_1/zin[0][868] ), .B(n34177), .Z(n32484) );
  IV U35516 ( .A(n34175), .Z(n34177) );
  XOR U35517 ( .A(n34175), .B(n32485), .Z(n34176) );
  XNOR U35518 ( .A(n34178), .B(n34179), .Z(n32485) );
  ANDN U35519 ( .B(\modmult_1/xin[1023] ), .A(n34180), .Z(n34178) );
  IV U35520 ( .A(n34179), .Z(n34180) );
  XNOR U35521 ( .A(m[869]), .B(n34181), .Z(n34179) );
  NAND U35522 ( .A(n34182), .B(mul_pow), .Z(n34181) );
  XOR U35523 ( .A(m[869]), .B(c[869]), .Z(n34182) );
  XOR U35524 ( .A(n34183), .B(n34184), .Z(n34175) );
  ANDN U35525 ( .B(n34185), .A(n32482), .Z(n34183) );
  XNOR U35526 ( .A(\modmult_1/zin[0][867] ), .B(n34186), .Z(n32482) );
  IV U35527 ( .A(n34184), .Z(n34186) );
  XOR U35528 ( .A(n34184), .B(n32483), .Z(n34185) );
  XNOR U35529 ( .A(n34187), .B(n34188), .Z(n32483) );
  ANDN U35530 ( .B(\modmult_1/xin[1023] ), .A(n34189), .Z(n34187) );
  IV U35531 ( .A(n34188), .Z(n34189) );
  XNOR U35532 ( .A(m[868]), .B(n34190), .Z(n34188) );
  NAND U35533 ( .A(n34191), .B(mul_pow), .Z(n34190) );
  XOR U35534 ( .A(m[868]), .B(c[868]), .Z(n34191) );
  XOR U35535 ( .A(n34192), .B(n34193), .Z(n34184) );
  ANDN U35536 ( .B(n34194), .A(n32480), .Z(n34192) );
  XNOR U35537 ( .A(\modmult_1/zin[0][866] ), .B(n34195), .Z(n32480) );
  IV U35538 ( .A(n34193), .Z(n34195) );
  XOR U35539 ( .A(n34193), .B(n32481), .Z(n34194) );
  XNOR U35540 ( .A(n34196), .B(n34197), .Z(n32481) );
  ANDN U35541 ( .B(\modmult_1/xin[1023] ), .A(n34198), .Z(n34196) );
  IV U35542 ( .A(n34197), .Z(n34198) );
  XNOR U35543 ( .A(m[867]), .B(n34199), .Z(n34197) );
  NAND U35544 ( .A(n34200), .B(mul_pow), .Z(n34199) );
  XOR U35545 ( .A(m[867]), .B(c[867]), .Z(n34200) );
  XOR U35546 ( .A(n34201), .B(n34202), .Z(n34193) );
  ANDN U35547 ( .B(n34203), .A(n32478), .Z(n34201) );
  XNOR U35548 ( .A(\modmult_1/zin[0][865] ), .B(n34204), .Z(n32478) );
  IV U35549 ( .A(n34202), .Z(n34204) );
  XOR U35550 ( .A(n34202), .B(n32479), .Z(n34203) );
  XNOR U35551 ( .A(n34205), .B(n34206), .Z(n32479) );
  ANDN U35552 ( .B(\modmult_1/xin[1023] ), .A(n34207), .Z(n34205) );
  IV U35553 ( .A(n34206), .Z(n34207) );
  XNOR U35554 ( .A(m[866]), .B(n34208), .Z(n34206) );
  NAND U35555 ( .A(n34209), .B(mul_pow), .Z(n34208) );
  XOR U35556 ( .A(m[866]), .B(c[866]), .Z(n34209) );
  XOR U35557 ( .A(n34210), .B(n34211), .Z(n34202) );
  ANDN U35558 ( .B(n34212), .A(n32476), .Z(n34210) );
  XNOR U35559 ( .A(\modmult_1/zin[0][864] ), .B(n34213), .Z(n32476) );
  IV U35560 ( .A(n34211), .Z(n34213) );
  XOR U35561 ( .A(n34211), .B(n32477), .Z(n34212) );
  XNOR U35562 ( .A(n34214), .B(n34215), .Z(n32477) );
  ANDN U35563 ( .B(\modmult_1/xin[1023] ), .A(n34216), .Z(n34214) );
  IV U35564 ( .A(n34215), .Z(n34216) );
  XNOR U35565 ( .A(m[865]), .B(n34217), .Z(n34215) );
  NAND U35566 ( .A(n34218), .B(mul_pow), .Z(n34217) );
  XOR U35567 ( .A(m[865]), .B(c[865]), .Z(n34218) );
  XOR U35568 ( .A(n34219), .B(n34220), .Z(n34211) );
  ANDN U35569 ( .B(n34221), .A(n32474), .Z(n34219) );
  XNOR U35570 ( .A(\modmult_1/zin[0][863] ), .B(n34222), .Z(n32474) );
  IV U35571 ( .A(n34220), .Z(n34222) );
  XOR U35572 ( .A(n34220), .B(n32475), .Z(n34221) );
  XNOR U35573 ( .A(n34223), .B(n34224), .Z(n32475) );
  ANDN U35574 ( .B(\modmult_1/xin[1023] ), .A(n34225), .Z(n34223) );
  IV U35575 ( .A(n34224), .Z(n34225) );
  XNOR U35576 ( .A(m[864]), .B(n34226), .Z(n34224) );
  NAND U35577 ( .A(n34227), .B(mul_pow), .Z(n34226) );
  XOR U35578 ( .A(m[864]), .B(c[864]), .Z(n34227) );
  XOR U35579 ( .A(n34228), .B(n34229), .Z(n34220) );
  ANDN U35580 ( .B(n34230), .A(n32472), .Z(n34228) );
  XNOR U35581 ( .A(\modmult_1/zin[0][862] ), .B(n34231), .Z(n32472) );
  IV U35582 ( .A(n34229), .Z(n34231) );
  XOR U35583 ( .A(n34229), .B(n32473), .Z(n34230) );
  XNOR U35584 ( .A(n34232), .B(n34233), .Z(n32473) );
  ANDN U35585 ( .B(\modmult_1/xin[1023] ), .A(n34234), .Z(n34232) );
  IV U35586 ( .A(n34233), .Z(n34234) );
  XNOR U35587 ( .A(m[863]), .B(n34235), .Z(n34233) );
  NAND U35588 ( .A(n34236), .B(mul_pow), .Z(n34235) );
  XOR U35589 ( .A(m[863]), .B(c[863]), .Z(n34236) );
  XOR U35590 ( .A(n34237), .B(n34238), .Z(n34229) );
  ANDN U35591 ( .B(n34239), .A(n32470), .Z(n34237) );
  XNOR U35592 ( .A(\modmult_1/zin[0][861] ), .B(n34240), .Z(n32470) );
  IV U35593 ( .A(n34238), .Z(n34240) );
  XOR U35594 ( .A(n34238), .B(n32471), .Z(n34239) );
  XNOR U35595 ( .A(n34241), .B(n34242), .Z(n32471) );
  ANDN U35596 ( .B(\modmult_1/xin[1023] ), .A(n34243), .Z(n34241) );
  IV U35597 ( .A(n34242), .Z(n34243) );
  XNOR U35598 ( .A(m[862]), .B(n34244), .Z(n34242) );
  NAND U35599 ( .A(n34245), .B(mul_pow), .Z(n34244) );
  XOR U35600 ( .A(m[862]), .B(c[862]), .Z(n34245) );
  XOR U35601 ( .A(n34246), .B(n34247), .Z(n34238) );
  ANDN U35602 ( .B(n34248), .A(n32468), .Z(n34246) );
  XNOR U35603 ( .A(\modmult_1/zin[0][860] ), .B(n34249), .Z(n32468) );
  IV U35604 ( .A(n34247), .Z(n34249) );
  XOR U35605 ( .A(n34247), .B(n32469), .Z(n34248) );
  XNOR U35606 ( .A(n34250), .B(n34251), .Z(n32469) );
  ANDN U35607 ( .B(\modmult_1/xin[1023] ), .A(n34252), .Z(n34250) );
  IV U35608 ( .A(n34251), .Z(n34252) );
  XNOR U35609 ( .A(m[861]), .B(n34253), .Z(n34251) );
  NAND U35610 ( .A(n34254), .B(mul_pow), .Z(n34253) );
  XOR U35611 ( .A(m[861]), .B(c[861]), .Z(n34254) );
  XOR U35612 ( .A(n34255), .B(n34256), .Z(n34247) );
  ANDN U35613 ( .B(n34257), .A(n32466), .Z(n34255) );
  XNOR U35614 ( .A(\modmult_1/zin[0][859] ), .B(n34258), .Z(n32466) );
  IV U35615 ( .A(n34256), .Z(n34258) );
  XOR U35616 ( .A(n34256), .B(n32467), .Z(n34257) );
  XNOR U35617 ( .A(n34259), .B(n34260), .Z(n32467) );
  ANDN U35618 ( .B(\modmult_1/xin[1023] ), .A(n34261), .Z(n34259) );
  IV U35619 ( .A(n34260), .Z(n34261) );
  XNOR U35620 ( .A(m[860]), .B(n34262), .Z(n34260) );
  NAND U35621 ( .A(n34263), .B(mul_pow), .Z(n34262) );
  XOR U35622 ( .A(m[860]), .B(c[860]), .Z(n34263) );
  XOR U35623 ( .A(n34264), .B(n34265), .Z(n34256) );
  ANDN U35624 ( .B(n34266), .A(n32464), .Z(n34264) );
  XNOR U35625 ( .A(\modmult_1/zin[0][858] ), .B(n34267), .Z(n32464) );
  IV U35626 ( .A(n34265), .Z(n34267) );
  XOR U35627 ( .A(n34265), .B(n32465), .Z(n34266) );
  XNOR U35628 ( .A(n34268), .B(n34269), .Z(n32465) );
  ANDN U35629 ( .B(\modmult_1/xin[1023] ), .A(n34270), .Z(n34268) );
  IV U35630 ( .A(n34269), .Z(n34270) );
  XNOR U35631 ( .A(m[859]), .B(n34271), .Z(n34269) );
  NAND U35632 ( .A(n34272), .B(mul_pow), .Z(n34271) );
  XOR U35633 ( .A(m[859]), .B(c[859]), .Z(n34272) );
  XOR U35634 ( .A(n34273), .B(n34274), .Z(n34265) );
  ANDN U35635 ( .B(n34275), .A(n32462), .Z(n34273) );
  XNOR U35636 ( .A(\modmult_1/zin[0][857] ), .B(n34276), .Z(n32462) );
  IV U35637 ( .A(n34274), .Z(n34276) );
  XOR U35638 ( .A(n34274), .B(n32463), .Z(n34275) );
  XNOR U35639 ( .A(n34277), .B(n34278), .Z(n32463) );
  ANDN U35640 ( .B(\modmult_1/xin[1023] ), .A(n34279), .Z(n34277) );
  IV U35641 ( .A(n34278), .Z(n34279) );
  XNOR U35642 ( .A(m[858]), .B(n34280), .Z(n34278) );
  NAND U35643 ( .A(n34281), .B(mul_pow), .Z(n34280) );
  XOR U35644 ( .A(m[858]), .B(c[858]), .Z(n34281) );
  XOR U35645 ( .A(n34282), .B(n34283), .Z(n34274) );
  ANDN U35646 ( .B(n34284), .A(n32460), .Z(n34282) );
  XNOR U35647 ( .A(\modmult_1/zin[0][856] ), .B(n34285), .Z(n32460) );
  IV U35648 ( .A(n34283), .Z(n34285) );
  XOR U35649 ( .A(n34283), .B(n32461), .Z(n34284) );
  XNOR U35650 ( .A(n34286), .B(n34287), .Z(n32461) );
  ANDN U35651 ( .B(\modmult_1/xin[1023] ), .A(n34288), .Z(n34286) );
  IV U35652 ( .A(n34287), .Z(n34288) );
  XNOR U35653 ( .A(m[857]), .B(n34289), .Z(n34287) );
  NAND U35654 ( .A(n34290), .B(mul_pow), .Z(n34289) );
  XOR U35655 ( .A(m[857]), .B(c[857]), .Z(n34290) );
  XOR U35656 ( .A(n34291), .B(n34292), .Z(n34283) );
  ANDN U35657 ( .B(n34293), .A(n32458), .Z(n34291) );
  XNOR U35658 ( .A(\modmult_1/zin[0][855] ), .B(n34294), .Z(n32458) );
  IV U35659 ( .A(n34292), .Z(n34294) );
  XOR U35660 ( .A(n34292), .B(n32459), .Z(n34293) );
  XNOR U35661 ( .A(n34295), .B(n34296), .Z(n32459) );
  ANDN U35662 ( .B(\modmult_1/xin[1023] ), .A(n34297), .Z(n34295) );
  IV U35663 ( .A(n34296), .Z(n34297) );
  XNOR U35664 ( .A(m[856]), .B(n34298), .Z(n34296) );
  NAND U35665 ( .A(n34299), .B(mul_pow), .Z(n34298) );
  XOR U35666 ( .A(m[856]), .B(c[856]), .Z(n34299) );
  XOR U35667 ( .A(n34300), .B(n34301), .Z(n34292) );
  ANDN U35668 ( .B(n34302), .A(n32456), .Z(n34300) );
  XNOR U35669 ( .A(\modmult_1/zin[0][854] ), .B(n34303), .Z(n32456) );
  IV U35670 ( .A(n34301), .Z(n34303) );
  XOR U35671 ( .A(n34301), .B(n32457), .Z(n34302) );
  XNOR U35672 ( .A(n34304), .B(n34305), .Z(n32457) );
  ANDN U35673 ( .B(\modmult_1/xin[1023] ), .A(n34306), .Z(n34304) );
  IV U35674 ( .A(n34305), .Z(n34306) );
  XNOR U35675 ( .A(m[855]), .B(n34307), .Z(n34305) );
  NAND U35676 ( .A(n34308), .B(mul_pow), .Z(n34307) );
  XOR U35677 ( .A(m[855]), .B(c[855]), .Z(n34308) );
  XOR U35678 ( .A(n34309), .B(n34310), .Z(n34301) );
  ANDN U35679 ( .B(n34311), .A(n32454), .Z(n34309) );
  XNOR U35680 ( .A(\modmult_1/zin[0][853] ), .B(n34312), .Z(n32454) );
  IV U35681 ( .A(n34310), .Z(n34312) );
  XOR U35682 ( .A(n34310), .B(n32455), .Z(n34311) );
  XNOR U35683 ( .A(n34313), .B(n34314), .Z(n32455) );
  ANDN U35684 ( .B(\modmult_1/xin[1023] ), .A(n34315), .Z(n34313) );
  IV U35685 ( .A(n34314), .Z(n34315) );
  XNOR U35686 ( .A(m[854]), .B(n34316), .Z(n34314) );
  NAND U35687 ( .A(n34317), .B(mul_pow), .Z(n34316) );
  XOR U35688 ( .A(m[854]), .B(c[854]), .Z(n34317) );
  XOR U35689 ( .A(n34318), .B(n34319), .Z(n34310) );
  ANDN U35690 ( .B(n34320), .A(n32452), .Z(n34318) );
  XNOR U35691 ( .A(\modmult_1/zin[0][852] ), .B(n34321), .Z(n32452) );
  IV U35692 ( .A(n34319), .Z(n34321) );
  XOR U35693 ( .A(n34319), .B(n32453), .Z(n34320) );
  XNOR U35694 ( .A(n34322), .B(n34323), .Z(n32453) );
  ANDN U35695 ( .B(\modmult_1/xin[1023] ), .A(n34324), .Z(n34322) );
  IV U35696 ( .A(n34323), .Z(n34324) );
  XNOR U35697 ( .A(m[853]), .B(n34325), .Z(n34323) );
  NAND U35698 ( .A(n34326), .B(mul_pow), .Z(n34325) );
  XOR U35699 ( .A(m[853]), .B(c[853]), .Z(n34326) );
  XOR U35700 ( .A(n34327), .B(n34328), .Z(n34319) );
  ANDN U35701 ( .B(n34329), .A(n32450), .Z(n34327) );
  XNOR U35702 ( .A(\modmult_1/zin[0][851] ), .B(n34330), .Z(n32450) );
  IV U35703 ( .A(n34328), .Z(n34330) );
  XOR U35704 ( .A(n34328), .B(n32451), .Z(n34329) );
  XNOR U35705 ( .A(n34331), .B(n34332), .Z(n32451) );
  ANDN U35706 ( .B(\modmult_1/xin[1023] ), .A(n34333), .Z(n34331) );
  IV U35707 ( .A(n34332), .Z(n34333) );
  XNOR U35708 ( .A(m[852]), .B(n34334), .Z(n34332) );
  NAND U35709 ( .A(n34335), .B(mul_pow), .Z(n34334) );
  XOR U35710 ( .A(m[852]), .B(c[852]), .Z(n34335) );
  XOR U35711 ( .A(n34336), .B(n34337), .Z(n34328) );
  ANDN U35712 ( .B(n34338), .A(n32448), .Z(n34336) );
  XNOR U35713 ( .A(\modmult_1/zin[0][850] ), .B(n34339), .Z(n32448) );
  IV U35714 ( .A(n34337), .Z(n34339) );
  XOR U35715 ( .A(n34337), .B(n32449), .Z(n34338) );
  XNOR U35716 ( .A(n34340), .B(n34341), .Z(n32449) );
  ANDN U35717 ( .B(\modmult_1/xin[1023] ), .A(n34342), .Z(n34340) );
  IV U35718 ( .A(n34341), .Z(n34342) );
  XNOR U35719 ( .A(m[851]), .B(n34343), .Z(n34341) );
  NAND U35720 ( .A(n34344), .B(mul_pow), .Z(n34343) );
  XOR U35721 ( .A(m[851]), .B(c[851]), .Z(n34344) );
  XOR U35722 ( .A(n34345), .B(n34346), .Z(n34337) );
  ANDN U35723 ( .B(n34347), .A(n32446), .Z(n34345) );
  XNOR U35724 ( .A(\modmult_1/zin[0][849] ), .B(n34348), .Z(n32446) );
  IV U35725 ( .A(n34346), .Z(n34348) );
  XOR U35726 ( .A(n34346), .B(n32447), .Z(n34347) );
  XNOR U35727 ( .A(n34349), .B(n34350), .Z(n32447) );
  ANDN U35728 ( .B(\modmult_1/xin[1023] ), .A(n34351), .Z(n34349) );
  IV U35729 ( .A(n34350), .Z(n34351) );
  XNOR U35730 ( .A(m[850]), .B(n34352), .Z(n34350) );
  NAND U35731 ( .A(n34353), .B(mul_pow), .Z(n34352) );
  XOR U35732 ( .A(m[850]), .B(c[850]), .Z(n34353) );
  XOR U35733 ( .A(n34354), .B(n34355), .Z(n34346) );
  ANDN U35734 ( .B(n34356), .A(n32444), .Z(n34354) );
  XNOR U35735 ( .A(\modmult_1/zin[0][848] ), .B(n34357), .Z(n32444) );
  IV U35736 ( .A(n34355), .Z(n34357) );
  XOR U35737 ( .A(n34355), .B(n32445), .Z(n34356) );
  XNOR U35738 ( .A(n34358), .B(n34359), .Z(n32445) );
  ANDN U35739 ( .B(\modmult_1/xin[1023] ), .A(n34360), .Z(n34358) );
  IV U35740 ( .A(n34359), .Z(n34360) );
  XNOR U35741 ( .A(m[849]), .B(n34361), .Z(n34359) );
  NAND U35742 ( .A(n34362), .B(mul_pow), .Z(n34361) );
  XOR U35743 ( .A(m[849]), .B(c[849]), .Z(n34362) );
  XOR U35744 ( .A(n34363), .B(n34364), .Z(n34355) );
  ANDN U35745 ( .B(n34365), .A(n32442), .Z(n34363) );
  XNOR U35746 ( .A(\modmult_1/zin[0][847] ), .B(n34366), .Z(n32442) );
  IV U35747 ( .A(n34364), .Z(n34366) );
  XOR U35748 ( .A(n34364), .B(n32443), .Z(n34365) );
  XNOR U35749 ( .A(n34367), .B(n34368), .Z(n32443) );
  ANDN U35750 ( .B(\modmult_1/xin[1023] ), .A(n34369), .Z(n34367) );
  IV U35751 ( .A(n34368), .Z(n34369) );
  XNOR U35752 ( .A(m[848]), .B(n34370), .Z(n34368) );
  NAND U35753 ( .A(n34371), .B(mul_pow), .Z(n34370) );
  XOR U35754 ( .A(m[848]), .B(c[848]), .Z(n34371) );
  XOR U35755 ( .A(n34372), .B(n34373), .Z(n34364) );
  ANDN U35756 ( .B(n34374), .A(n32440), .Z(n34372) );
  XNOR U35757 ( .A(\modmult_1/zin[0][846] ), .B(n34375), .Z(n32440) );
  IV U35758 ( .A(n34373), .Z(n34375) );
  XOR U35759 ( .A(n34373), .B(n32441), .Z(n34374) );
  XNOR U35760 ( .A(n34376), .B(n34377), .Z(n32441) );
  ANDN U35761 ( .B(\modmult_1/xin[1023] ), .A(n34378), .Z(n34376) );
  IV U35762 ( .A(n34377), .Z(n34378) );
  XNOR U35763 ( .A(m[847]), .B(n34379), .Z(n34377) );
  NAND U35764 ( .A(n34380), .B(mul_pow), .Z(n34379) );
  XOR U35765 ( .A(m[847]), .B(c[847]), .Z(n34380) );
  XOR U35766 ( .A(n34381), .B(n34382), .Z(n34373) );
  ANDN U35767 ( .B(n34383), .A(n32438), .Z(n34381) );
  XNOR U35768 ( .A(\modmult_1/zin[0][845] ), .B(n34384), .Z(n32438) );
  IV U35769 ( .A(n34382), .Z(n34384) );
  XOR U35770 ( .A(n34382), .B(n32439), .Z(n34383) );
  XNOR U35771 ( .A(n34385), .B(n34386), .Z(n32439) );
  ANDN U35772 ( .B(\modmult_1/xin[1023] ), .A(n34387), .Z(n34385) );
  IV U35773 ( .A(n34386), .Z(n34387) );
  XNOR U35774 ( .A(m[846]), .B(n34388), .Z(n34386) );
  NAND U35775 ( .A(n34389), .B(mul_pow), .Z(n34388) );
  XOR U35776 ( .A(m[846]), .B(c[846]), .Z(n34389) );
  XOR U35777 ( .A(n34390), .B(n34391), .Z(n34382) );
  ANDN U35778 ( .B(n34392), .A(n32436), .Z(n34390) );
  XNOR U35779 ( .A(\modmult_1/zin[0][844] ), .B(n34393), .Z(n32436) );
  IV U35780 ( .A(n34391), .Z(n34393) );
  XOR U35781 ( .A(n34391), .B(n32437), .Z(n34392) );
  XNOR U35782 ( .A(n34394), .B(n34395), .Z(n32437) );
  ANDN U35783 ( .B(\modmult_1/xin[1023] ), .A(n34396), .Z(n34394) );
  IV U35784 ( .A(n34395), .Z(n34396) );
  XNOR U35785 ( .A(m[845]), .B(n34397), .Z(n34395) );
  NAND U35786 ( .A(n34398), .B(mul_pow), .Z(n34397) );
  XOR U35787 ( .A(m[845]), .B(c[845]), .Z(n34398) );
  XOR U35788 ( .A(n34399), .B(n34400), .Z(n34391) );
  ANDN U35789 ( .B(n34401), .A(n32434), .Z(n34399) );
  XNOR U35790 ( .A(\modmult_1/zin[0][843] ), .B(n34402), .Z(n32434) );
  IV U35791 ( .A(n34400), .Z(n34402) );
  XOR U35792 ( .A(n34400), .B(n32435), .Z(n34401) );
  XNOR U35793 ( .A(n34403), .B(n34404), .Z(n32435) );
  ANDN U35794 ( .B(\modmult_1/xin[1023] ), .A(n34405), .Z(n34403) );
  IV U35795 ( .A(n34404), .Z(n34405) );
  XNOR U35796 ( .A(m[844]), .B(n34406), .Z(n34404) );
  NAND U35797 ( .A(n34407), .B(mul_pow), .Z(n34406) );
  XOR U35798 ( .A(m[844]), .B(c[844]), .Z(n34407) );
  XOR U35799 ( .A(n34408), .B(n34409), .Z(n34400) );
  ANDN U35800 ( .B(n34410), .A(n32432), .Z(n34408) );
  XNOR U35801 ( .A(\modmult_1/zin[0][842] ), .B(n34411), .Z(n32432) );
  IV U35802 ( .A(n34409), .Z(n34411) );
  XOR U35803 ( .A(n34409), .B(n32433), .Z(n34410) );
  XNOR U35804 ( .A(n34412), .B(n34413), .Z(n32433) );
  ANDN U35805 ( .B(\modmult_1/xin[1023] ), .A(n34414), .Z(n34412) );
  IV U35806 ( .A(n34413), .Z(n34414) );
  XNOR U35807 ( .A(m[843]), .B(n34415), .Z(n34413) );
  NAND U35808 ( .A(n34416), .B(mul_pow), .Z(n34415) );
  XOR U35809 ( .A(m[843]), .B(c[843]), .Z(n34416) );
  XOR U35810 ( .A(n34417), .B(n34418), .Z(n34409) );
  ANDN U35811 ( .B(n34419), .A(n32430), .Z(n34417) );
  XNOR U35812 ( .A(\modmult_1/zin[0][841] ), .B(n34420), .Z(n32430) );
  IV U35813 ( .A(n34418), .Z(n34420) );
  XOR U35814 ( .A(n34418), .B(n32431), .Z(n34419) );
  XNOR U35815 ( .A(n34421), .B(n34422), .Z(n32431) );
  ANDN U35816 ( .B(\modmult_1/xin[1023] ), .A(n34423), .Z(n34421) );
  IV U35817 ( .A(n34422), .Z(n34423) );
  XNOR U35818 ( .A(m[842]), .B(n34424), .Z(n34422) );
  NAND U35819 ( .A(n34425), .B(mul_pow), .Z(n34424) );
  XOR U35820 ( .A(m[842]), .B(c[842]), .Z(n34425) );
  XOR U35821 ( .A(n34426), .B(n34427), .Z(n34418) );
  ANDN U35822 ( .B(n34428), .A(n32428), .Z(n34426) );
  XNOR U35823 ( .A(\modmult_1/zin[0][840] ), .B(n34429), .Z(n32428) );
  IV U35824 ( .A(n34427), .Z(n34429) );
  XOR U35825 ( .A(n34427), .B(n32429), .Z(n34428) );
  XNOR U35826 ( .A(n34430), .B(n34431), .Z(n32429) );
  ANDN U35827 ( .B(\modmult_1/xin[1023] ), .A(n34432), .Z(n34430) );
  IV U35828 ( .A(n34431), .Z(n34432) );
  XNOR U35829 ( .A(m[841]), .B(n34433), .Z(n34431) );
  NAND U35830 ( .A(n34434), .B(mul_pow), .Z(n34433) );
  XOR U35831 ( .A(m[841]), .B(c[841]), .Z(n34434) );
  XOR U35832 ( .A(n34435), .B(n34436), .Z(n34427) );
  ANDN U35833 ( .B(n34437), .A(n32426), .Z(n34435) );
  XNOR U35834 ( .A(\modmult_1/zin[0][839] ), .B(n34438), .Z(n32426) );
  IV U35835 ( .A(n34436), .Z(n34438) );
  XOR U35836 ( .A(n34436), .B(n32427), .Z(n34437) );
  XNOR U35837 ( .A(n34439), .B(n34440), .Z(n32427) );
  ANDN U35838 ( .B(\modmult_1/xin[1023] ), .A(n34441), .Z(n34439) );
  IV U35839 ( .A(n34440), .Z(n34441) );
  XNOR U35840 ( .A(m[840]), .B(n34442), .Z(n34440) );
  NAND U35841 ( .A(n34443), .B(mul_pow), .Z(n34442) );
  XOR U35842 ( .A(m[840]), .B(c[840]), .Z(n34443) );
  XOR U35843 ( .A(n34444), .B(n34445), .Z(n34436) );
  ANDN U35844 ( .B(n34446), .A(n32424), .Z(n34444) );
  XNOR U35845 ( .A(\modmult_1/zin[0][838] ), .B(n34447), .Z(n32424) );
  IV U35846 ( .A(n34445), .Z(n34447) );
  XOR U35847 ( .A(n34445), .B(n32425), .Z(n34446) );
  XNOR U35848 ( .A(n34448), .B(n34449), .Z(n32425) );
  ANDN U35849 ( .B(\modmult_1/xin[1023] ), .A(n34450), .Z(n34448) );
  IV U35850 ( .A(n34449), .Z(n34450) );
  XNOR U35851 ( .A(m[839]), .B(n34451), .Z(n34449) );
  NAND U35852 ( .A(n34452), .B(mul_pow), .Z(n34451) );
  XOR U35853 ( .A(m[839]), .B(c[839]), .Z(n34452) );
  XOR U35854 ( .A(n34453), .B(n34454), .Z(n34445) );
  ANDN U35855 ( .B(n34455), .A(n32422), .Z(n34453) );
  XNOR U35856 ( .A(\modmult_1/zin[0][837] ), .B(n34456), .Z(n32422) );
  IV U35857 ( .A(n34454), .Z(n34456) );
  XOR U35858 ( .A(n34454), .B(n32423), .Z(n34455) );
  XNOR U35859 ( .A(n34457), .B(n34458), .Z(n32423) );
  ANDN U35860 ( .B(\modmult_1/xin[1023] ), .A(n34459), .Z(n34457) );
  IV U35861 ( .A(n34458), .Z(n34459) );
  XNOR U35862 ( .A(m[838]), .B(n34460), .Z(n34458) );
  NAND U35863 ( .A(n34461), .B(mul_pow), .Z(n34460) );
  XOR U35864 ( .A(m[838]), .B(c[838]), .Z(n34461) );
  XOR U35865 ( .A(n34462), .B(n34463), .Z(n34454) );
  ANDN U35866 ( .B(n34464), .A(n32420), .Z(n34462) );
  XNOR U35867 ( .A(\modmult_1/zin[0][836] ), .B(n34465), .Z(n32420) );
  IV U35868 ( .A(n34463), .Z(n34465) );
  XOR U35869 ( .A(n34463), .B(n32421), .Z(n34464) );
  XNOR U35870 ( .A(n34466), .B(n34467), .Z(n32421) );
  ANDN U35871 ( .B(\modmult_1/xin[1023] ), .A(n34468), .Z(n34466) );
  IV U35872 ( .A(n34467), .Z(n34468) );
  XNOR U35873 ( .A(m[837]), .B(n34469), .Z(n34467) );
  NAND U35874 ( .A(n34470), .B(mul_pow), .Z(n34469) );
  XOR U35875 ( .A(m[837]), .B(c[837]), .Z(n34470) );
  XOR U35876 ( .A(n34471), .B(n34472), .Z(n34463) );
  ANDN U35877 ( .B(n34473), .A(n32418), .Z(n34471) );
  XNOR U35878 ( .A(\modmult_1/zin[0][835] ), .B(n34474), .Z(n32418) );
  IV U35879 ( .A(n34472), .Z(n34474) );
  XOR U35880 ( .A(n34472), .B(n32419), .Z(n34473) );
  XNOR U35881 ( .A(n34475), .B(n34476), .Z(n32419) );
  ANDN U35882 ( .B(\modmult_1/xin[1023] ), .A(n34477), .Z(n34475) );
  IV U35883 ( .A(n34476), .Z(n34477) );
  XNOR U35884 ( .A(m[836]), .B(n34478), .Z(n34476) );
  NAND U35885 ( .A(n34479), .B(mul_pow), .Z(n34478) );
  XOR U35886 ( .A(m[836]), .B(c[836]), .Z(n34479) );
  XOR U35887 ( .A(n34480), .B(n34481), .Z(n34472) );
  ANDN U35888 ( .B(n34482), .A(n32416), .Z(n34480) );
  XNOR U35889 ( .A(\modmult_1/zin[0][834] ), .B(n34483), .Z(n32416) );
  IV U35890 ( .A(n34481), .Z(n34483) );
  XOR U35891 ( .A(n34481), .B(n32417), .Z(n34482) );
  XNOR U35892 ( .A(n34484), .B(n34485), .Z(n32417) );
  ANDN U35893 ( .B(\modmult_1/xin[1023] ), .A(n34486), .Z(n34484) );
  IV U35894 ( .A(n34485), .Z(n34486) );
  XNOR U35895 ( .A(m[835]), .B(n34487), .Z(n34485) );
  NAND U35896 ( .A(n34488), .B(mul_pow), .Z(n34487) );
  XOR U35897 ( .A(m[835]), .B(c[835]), .Z(n34488) );
  XOR U35898 ( .A(n34489), .B(n34490), .Z(n34481) );
  ANDN U35899 ( .B(n34491), .A(n32414), .Z(n34489) );
  XNOR U35900 ( .A(\modmult_1/zin[0][833] ), .B(n34492), .Z(n32414) );
  IV U35901 ( .A(n34490), .Z(n34492) );
  XOR U35902 ( .A(n34490), .B(n32415), .Z(n34491) );
  XNOR U35903 ( .A(n34493), .B(n34494), .Z(n32415) );
  ANDN U35904 ( .B(\modmult_1/xin[1023] ), .A(n34495), .Z(n34493) );
  IV U35905 ( .A(n34494), .Z(n34495) );
  XNOR U35906 ( .A(m[834]), .B(n34496), .Z(n34494) );
  NAND U35907 ( .A(n34497), .B(mul_pow), .Z(n34496) );
  XOR U35908 ( .A(m[834]), .B(c[834]), .Z(n34497) );
  XOR U35909 ( .A(n34498), .B(n34499), .Z(n34490) );
  ANDN U35910 ( .B(n34500), .A(n32412), .Z(n34498) );
  XNOR U35911 ( .A(\modmult_1/zin[0][832] ), .B(n34501), .Z(n32412) );
  IV U35912 ( .A(n34499), .Z(n34501) );
  XOR U35913 ( .A(n34499), .B(n32413), .Z(n34500) );
  XNOR U35914 ( .A(n34502), .B(n34503), .Z(n32413) );
  ANDN U35915 ( .B(\modmult_1/xin[1023] ), .A(n34504), .Z(n34502) );
  IV U35916 ( .A(n34503), .Z(n34504) );
  XNOR U35917 ( .A(m[833]), .B(n34505), .Z(n34503) );
  NAND U35918 ( .A(n34506), .B(mul_pow), .Z(n34505) );
  XOR U35919 ( .A(m[833]), .B(c[833]), .Z(n34506) );
  XOR U35920 ( .A(n34507), .B(n34508), .Z(n34499) );
  ANDN U35921 ( .B(n34509), .A(n32410), .Z(n34507) );
  XNOR U35922 ( .A(\modmult_1/zin[0][831] ), .B(n34510), .Z(n32410) );
  IV U35923 ( .A(n34508), .Z(n34510) );
  XOR U35924 ( .A(n34508), .B(n32411), .Z(n34509) );
  XNOR U35925 ( .A(n34511), .B(n34512), .Z(n32411) );
  ANDN U35926 ( .B(\modmult_1/xin[1023] ), .A(n34513), .Z(n34511) );
  IV U35927 ( .A(n34512), .Z(n34513) );
  XNOR U35928 ( .A(m[832]), .B(n34514), .Z(n34512) );
  NAND U35929 ( .A(n34515), .B(mul_pow), .Z(n34514) );
  XOR U35930 ( .A(m[832]), .B(c[832]), .Z(n34515) );
  XOR U35931 ( .A(n34516), .B(n34517), .Z(n34508) );
  ANDN U35932 ( .B(n34518), .A(n32408), .Z(n34516) );
  XNOR U35933 ( .A(\modmult_1/zin[0][830] ), .B(n34519), .Z(n32408) );
  IV U35934 ( .A(n34517), .Z(n34519) );
  XOR U35935 ( .A(n34517), .B(n32409), .Z(n34518) );
  XNOR U35936 ( .A(n34520), .B(n34521), .Z(n32409) );
  ANDN U35937 ( .B(\modmult_1/xin[1023] ), .A(n34522), .Z(n34520) );
  IV U35938 ( .A(n34521), .Z(n34522) );
  XNOR U35939 ( .A(m[831]), .B(n34523), .Z(n34521) );
  NAND U35940 ( .A(n34524), .B(mul_pow), .Z(n34523) );
  XOR U35941 ( .A(m[831]), .B(c[831]), .Z(n34524) );
  XOR U35942 ( .A(n34525), .B(n34526), .Z(n34517) );
  ANDN U35943 ( .B(n34527), .A(n32406), .Z(n34525) );
  XNOR U35944 ( .A(\modmult_1/zin[0][829] ), .B(n34528), .Z(n32406) );
  IV U35945 ( .A(n34526), .Z(n34528) );
  XOR U35946 ( .A(n34526), .B(n32407), .Z(n34527) );
  XNOR U35947 ( .A(n34529), .B(n34530), .Z(n32407) );
  ANDN U35948 ( .B(\modmult_1/xin[1023] ), .A(n34531), .Z(n34529) );
  IV U35949 ( .A(n34530), .Z(n34531) );
  XNOR U35950 ( .A(m[830]), .B(n34532), .Z(n34530) );
  NAND U35951 ( .A(n34533), .B(mul_pow), .Z(n34532) );
  XOR U35952 ( .A(m[830]), .B(c[830]), .Z(n34533) );
  XOR U35953 ( .A(n34534), .B(n34535), .Z(n34526) );
  ANDN U35954 ( .B(n34536), .A(n32404), .Z(n34534) );
  XNOR U35955 ( .A(\modmult_1/zin[0][828] ), .B(n34537), .Z(n32404) );
  IV U35956 ( .A(n34535), .Z(n34537) );
  XOR U35957 ( .A(n34535), .B(n32405), .Z(n34536) );
  XNOR U35958 ( .A(n34538), .B(n34539), .Z(n32405) );
  ANDN U35959 ( .B(\modmult_1/xin[1023] ), .A(n34540), .Z(n34538) );
  IV U35960 ( .A(n34539), .Z(n34540) );
  XNOR U35961 ( .A(m[829]), .B(n34541), .Z(n34539) );
  NAND U35962 ( .A(n34542), .B(mul_pow), .Z(n34541) );
  XOR U35963 ( .A(m[829]), .B(c[829]), .Z(n34542) );
  XOR U35964 ( .A(n34543), .B(n34544), .Z(n34535) );
  ANDN U35965 ( .B(n34545), .A(n32402), .Z(n34543) );
  XNOR U35966 ( .A(\modmult_1/zin[0][827] ), .B(n34546), .Z(n32402) );
  IV U35967 ( .A(n34544), .Z(n34546) );
  XOR U35968 ( .A(n34544), .B(n32403), .Z(n34545) );
  XNOR U35969 ( .A(n34547), .B(n34548), .Z(n32403) );
  ANDN U35970 ( .B(\modmult_1/xin[1023] ), .A(n34549), .Z(n34547) );
  IV U35971 ( .A(n34548), .Z(n34549) );
  XNOR U35972 ( .A(m[828]), .B(n34550), .Z(n34548) );
  NAND U35973 ( .A(n34551), .B(mul_pow), .Z(n34550) );
  XOR U35974 ( .A(m[828]), .B(c[828]), .Z(n34551) );
  XOR U35975 ( .A(n34552), .B(n34553), .Z(n34544) );
  ANDN U35976 ( .B(n34554), .A(n32400), .Z(n34552) );
  XNOR U35977 ( .A(\modmult_1/zin[0][826] ), .B(n34555), .Z(n32400) );
  IV U35978 ( .A(n34553), .Z(n34555) );
  XOR U35979 ( .A(n34553), .B(n32401), .Z(n34554) );
  XNOR U35980 ( .A(n34556), .B(n34557), .Z(n32401) );
  ANDN U35981 ( .B(\modmult_1/xin[1023] ), .A(n34558), .Z(n34556) );
  IV U35982 ( .A(n34557), .Z(n34558) );
  XNOR U35983 ( .A(m[827]), .B(n34559), .Z(n34557) );
  NAND U35984 ( .A(n34560), .B(mul_pow), .Z(n34559) );
  XOR U35985 ( .A(m[827]), .B(c[827]), .Z(n34560) );
  XOR U35986 ( .A(n34561), .B(n34562), .Z(n34553) );
  ANDN U35987 ( .B(n34563), .A(n32398), .Z(n34561) );
  XNOR U35988 ( .A(\modmult_1/zin[0][825] ), .B(n34564), .Z(n32398) );
  IV U35989 ( .A(n34562), .Z(n34564) );
  XOR U35990 ( .A(n34562), .B(n32399), .Z(n34563) );
  XNOR U35991 ( .A(n34565), .B(n34566), .Z(n32399) );
  ANDN U35992 ( .B(\modmult_1/xin[1023] ), .A(n34567), .Z(n34565) );
  IV U35993 ( .A(n34566), .Z(n34567) );
  XNOR U35994 ( .A(m[826]), .B(n34568), .Z(n34566) );
  NAND U35995 ( .A(n34569), .B(mul_pow), .Z(n34568) );
  XOR U35996 ( .A(m[826]), .B(c[826]), .Z(n34569) );
  XOR U35997 ( .A(n34570), .B(n34571), .Z(n34562) );
  ANDN U35998 ( .B(n34572), .A(n32396), .Z(n34570) );
  XNOR U35999 ( .A(\modmult_1/zin[0][824] ), .B(n34573), .Z(n32396) );
  IV U36000 ( .A(n34571), .Z(n34573) );
  XOR U36001 ( .A(n34571), .B(n32397), .Z(n34572) );
  XNOR U36002 ( .A(n34574), .B(n34575), .Z(n32397) );
  ANDN U36003 ( .B(\modmult_1/xin[1023] ), .A(n34576), .Z(n34574) );
  IV U36004 ( .A(n34575), .Z(n34576) );
  XNOR U36005 ( .A(m[825]), .B(n34577), .Z(n34575) );
  NAND U36006 ( .A(n34578), .B(mul_pow), .Z(n34577) );
  XOR U36007 ( .A(m[825]), .B(c[825]), .Z(n34578) );
  XOR U36008 ( .A(n34579), .B(n34580), .Z(n34571) );
  ANDN U36009 ( .B(n34581), .A(n32394), .Z(n34579) );
  XNOR U36010 ( .A(\modmult_1/zin[0][823] ), .B(n34582), .Z(n32394) );
  IV U36011 ( .A(n34580), .Z(n34582) );
  XOR U36012 ( .A(n34580), .B(n32395), .Z(n34581) );
  XNOR U36013 ( .A(n34583), .B(n34584), .Z(n32395) );
  ANDN U36014 ( .B(\modmult_1/xin[1023] ), .A(n34585), .Z(n34583) );
  IV U36015 ( .A(n34584), .Z(n34585) );
  XNOR U36016 ( .A(m[824]), .B(n34586), .Z(n34584) );
  NAND U36017 ( .A(n34587), .B(mul_pow), .Z(n34586) );
  XOR U36018 ( .A(m[824]), .B(c[824]), .Z(n34587) );
  XOR U36019 ( .A(n34588), .B(n34589), .Z(n34580) );
  ANDN U36020 ( .B(n34590), .A(n32392), .Z(n34588) );
  XNOR U36021 ( .A(\modmult_1/zin[0][822] ), .B(n34591), .Z(n32392) );
  IV U36022 ( .A(n34589), .Z(n34591) );
  XOR U36023 ( .A(n34589), .B(n32393), .Z(n34590) );
  XNOR U36024 ( .A(n34592), .B(n34593), .Z(n32393) );
  ANDN U36025 ( .B(\modmult_1/xin[1023] ), .A(n34594), .Z(n34592) );
  IV U36026 ( .A(n34593), .Z(n34594) );
  XNOR U36027 ( .A(m[823]), .B(n34595), .Z(n34593) );
  NAND U36028 ( .A(n34596), .B(mul_pow), .Z(n34595) );
  XOR U36029 ( .A(m[823]), .B(c[823]), .Z(n34596) );
  XOR U36030 ( .A(n34597), .B(n34598), .Z(n34589) );
  ANDN U36031 ( .B(n34599), .A(n32390), .Z(n34597) );
  XNOR U36032 ( .A(\modmult_1/zin[0][821] ), .B(n34600), .Z(n32390) );
  IV U36033 ( .A(n34598), .Z(n34600) );
  XOR U36034 ( .A(n34598), .B(n32391), .Z(n34599) );
  XNOR U36035 ( .A(n34601), .B(n34602), .Z(n32391) );
  ANDN U36036 ( .B(\modmult_1/xin[1023] ), .A(n34603), .Z(n34601) );
  IV U36037 ( .A(n34602), .Z(n34603) );
  XNOR U36038 ( .A(m[822]), .B(n34604), .Z(n34602) );
  NAND U36039 ( .A(n34605), .B(mul_pow), .Z(n34604) );
  XOR U36040 ( .A(m[822]), .B(c[822]), .Z(n34605) );
  XOR U36041 ( .A(n34606), .B(n34607), .Z(n34598) );
  ANDN U36042 ( .B(n34608), .A(n32388), .Z(n34606) );
  XNOR U36043 ( .A(\modmult_1/zin[0][820] ), .B(n34609), .Z(n32388) );
  IV U36044 ( .A(n34607), .Z(n34609) );
  XOR U36045 ( .A(n34607), .B(n32389), .Z(n34608) );
  XNOR U36046 ( .A(n34610), .B(n34611), .Z(n32389) );
  ANDN U36047 ( .B(\modmult_1/xin[1023] ), .A(n34612), .Z(n34610) );
  IV U36048 ( .A(n34611), .Z(n34612) );
  XNOR U36049 ( .A(m[821]), .B(n34613), .Z(n34611) );
  NAND U36050 ( .A(n34614), .B(mul_pow), .Z(n34613) );
  XOR U36051 ( .A(m[821]), .B(c[821]), .Z(n34614) );
  XOR U36052 ( .A(n34615), .B(n34616), .Z(n34607) );
  ANDN U36053 ( .B(n34617), .A(n32386), .Z(n34615) );
  XNOR U36054 ( .A(\modmult_1/zin[0][819] ), .B(n34618), .Z(n32386) );
  IV U36055 ( .A(n34616), .Z(n34618) );
  XOR U36056 ( .A(n34616), .B(n32387), .Z(n34617) );
  XNOR U36057 ( .A(n34619), .B(n34620), .Z(n32387) );
  ANDN U36058 ( .B(\modmult_1/xin[1023] ), .A(n34621), .Z(n34619) );
  IV U36059 ( .A(n34620), .Z(n34621) );
  XNOR U36060 ( .A(m[820]), .B(n34622), .Z(n34620) );
  NAND U36061 ( .A(n34623), .B(mul_pow), .Z(n34622) );
  XOR U36062 ( .A(m[820]), .B(c[820]), .Z(n34623) );
  XOR U36063 ( .A(n34624), .B(n34625), .Z(n34616) );
  ANDN U36064 ( .B(n34626), .A(n32384), .Z(n34624) );
  XNOR U36065 ( .A(\modmult_1/zin[0][818] ), .B(n34627), .Z(n32384) );
  IV U36066 ( .A(n34625), .Z(n34627) );
  XOR U36067 ( .A(n34625), .B(n32385), .Z(n34626) );
  XNOR U36068 ( .A(n34628), .B(n34629), .Z(n32385) );
  ANDN U36069 ( .B(\modmult_1/xin[1023] ), .A(n34630), .Z(n34628) );
  IV U36070 ( .A(n34629), .Z(n34630) );
  XNOR U36071 ( .A(m[819]), .B(n34631), .Z(n34629) );
  NAND U36072 ( .A(n34632), .B(mul_pow), .Z(n34631) );
  XOR U36073 ( .A(m[819]), .B(c[819]), .Z(n34632) );
  XOR U36074 ( .A(n34633), .B(n34634), .Z(n34625) );
  ANDN U36075 ( .B(n34635), .A(n32382), .Z(n34633) );
  XNOR U36076 ( .A(\modmult_1/zin[0][817] ), .B(n34636), .Z(n32382) );
  IV U36077 ( .A(n34634), .Z(n34636) );
  XOR U36078 ( .A(n34634), .B(n32383), .Z(n34635) );
  XNOR U36079 ( .A(n34637), .B(n34638), .Z(n32383) );
  ANDN U36080 ( .B(\modmult_1/xin[1023] ), .A(n34639), .Z(n34637) );
  IV U36081 ( .A(n34638), .Z(n34639) );
  XNOR U36082 ( .A(m[818]), .B(n34640), .Z(n34638) );
  NAND U36083 ( .A(n34641), .B(mul_pow), .Z(n34640) );
  XOR U36084 ( .A(m[818]), .B(c[818]), .Z(n34641) );
  XOR U36085 ( .A(n34642), .B(n34643), .Z(n34634) );
  ANDN U36086 ( .B(n34644), .A(n32380), .Z(n34642) );
  XNOR U36087 ( .A(\modmult_1/zin[0][816] ), .B(n34645), .Z(n32380) );
  IV U36088 ( .A(n34643), .Z(n34645) );
  XOR U36089 ( .A(n34643), .B(n32381), .Z(n34644) );
  XNOR U36090 ( .A(n34646), .B(n34647), .Z(n32381) );
  ANDN U36091 ( .B(\modmult_1/xin[1023] ), .A(n34648), .Z(n34646) );
  IV U36092 ( .A(n34647), .Z(n34648) );
  XNOR U36093 ( .A(m[817]), .B(n34649), .Z(n34647) );
  NAND U36094 ( .A(n34650), .B(mul_pow), .Z(n34649) );
  XOR U36095 ( .A(m[817]), .B(c[817]), .Z(n34650) );
  XOR U36096 ( .A(n34651), .B(n34652), .Z(n34643) );
  ANDN U36097 ( .B(n34653), .A(n32378), .Z(n34651) );
  XNOR U36098 ( .A(\modmult_1/zin[0][815] ), .B(n34654), .Z(n32378) );
  IV U36099 ( .A(n34652), .Z(n34654) );
  XOR U36100 ( .A(n34652), .B(n32379), .Z(n34653) );
  XNOR U36101 ( .A(n34655), .B(n34656), .Z(n32379) );
  ANDN U36102 ( .B(\modmult_1/xin[1023] ), .A(n34657), .Z(n34655) );
  IV U36103 ( .A(n34656), .Z(n34657) );
  XNOR U36104 ( .A(m[816]), .B(n34658), .Z(n34656) );
  NAND U36105 ( .A(n34659), .B(mul_pow), .Z(n34658) );
  XOR U36106 ( .A(m[816]), .B(c[816]), .Z(n34659) );
  XOR U36107 ( .A(n34660), .B(n34661), .Z(n34652) );
  ANDN U36108 ( .B(n34662), .A(n32376), .Z(n34660) );
  XNOR U36109 ( .A(\modmult_1/zin[0][814] ), .B(n34663), .Z(n32376) );
  IV U36110 ( .A(n34661), .Z(n34663) );
  XOR U36111 ( .A(n34661), .B(n32377), .Z(n34662) );
  XNOR U36112 ( .A(n34664), .B(n34665), .Z(n32377) );
  ANDN U36113 ( .B(\modmult_1/xin[1023] ), .A(n34666), .Z(n34664) );
  IV U36114 ( .A(n34665), .Z(n34666) );
  XNOR U36115 ( .A(m[815]), .B(n34667), .Z(n34665) );
  NAND U36116 ( .A(n34668), .B(mul_pow), .Z(n34667) );
  XOR U36117 ( .A(m[815]), .B(c[815]), .Z(n34668) );
  XOR U36118 ( .A(n34669), .B(n34670), .Z(n34661) );
  ANDN U36119 ( .B(n34671), .A(n32374), .Z(n34669) );
  XNOR U36120 ( .A(\modmult_1/zin[0][813] ), .B(n34672), .Z(n32374) );
  IV U36121 ( .A(n34670), .Z(n34672) );
  XOR U36122 ( .A(n34670), .B(n32375), .Z(n34671) );
  XNOR U36123 ( .A(n34673), .B(n34674), .Z(n32375) );
  ANDN U36124 ( .B(\modmult_1/xin[1023] ), .A(n34675), .Z(n34673) );
  IV U36125 ( .A(n34674), .Z(n34675) );
  XNOR U36126 ( .A(m[814]), .B(n34676), .Z(n34674) );
  NAND U36127 ( .A(n34677), .B(mul_pow), .Z(n34676) );
  XOR U36128 ( .A(m[814]), .B(c[814]), .Z(n34677) );
  XOR U36129 ( .A(n34678), .B(n34679), .Z(n34670) );
  ANDN U36130 ( .B(n34680), .A(n32372), .Z(n34678) );
  XNOR U36131 ( .A(\modmult_1/zin[0][812] ), .B(n34681), .Z(n32372) );
  IV U36132 ( .A(n34679), .Z(n34681) );
  XOR U36133 ( .A(n34679), .B(n32373), .Z(n34680) );
  XNOR U36134 ( .A(n34682), .B(n34683), .Z(n32373) );
  ANDN U36135 ( .B(\modmult_1/xin[1023] ), .A(n34684), .Z(n34682) );
  IV U36136 ( .A(n34683), .Z(n34684) );
  XNOR U36137 ( .A(m[813]), .B(n34685), .Z(n34683) );
  NAND U36138 ( .A(n34686), .B(mul_pow), .Z(n34685) );
  XOR U36139 ( .A(m[813]), .B(c[813]), .Z(n34686) );
  XOR U36140 ( .A(n34687), .B(n34688), .Z(n34679) );
  ANDN U36141 ( .B(n34689), .A(n32370), .Z(n34687) );
  XNOR U36142 ( .A(\modmult_1/zin[0][811] ), .B(n34690), .Z(n32370) );
  IV U36143 ( .A(n34688), .Z(n34690) );
  XOR U36144 ( .A(n34688), .B(n32371), .Z(n34689) );
  XNOR U36145 ( .A(n34691), .B(n34692), .Z(n32371) );
  ANDN U36146 ( .B(\modmult_1/xin[1023] ), .A(n34693), .Z(n34691) );
  IV U36147 ( .A(n34692), .Z(n34693) );
  XNOR U36148 ( .A(m[812]), .B(n34694), .Z(n34692) );
  NAND U36149 ( .A(n34695), .B(mul_pow), .Z(n34694) );
  XOR U36150 ( .A(m[812]), .B(c[812]), .Z(n34695) );
  XOR U36151 ( .A(n34696), .B(n34697), .Z(n34688) );
  ANDN U36152 ( .B(n34698), .A(n32368), .Z(n34696) );
  XNOR U36153 ( .A(\modmult_1/zin[0][810] ), .B(n34699), .Z(n32368) );
  IV U36154 ( .A(n34697), .Z(n34699) );
  XOR U36155 ( .A(n34697), .B(n32369), .Z(n34698) );
  XNOR U36156 ( .A(n34700), .B(n34701), .Z(n32369) );
  ANDN U36157 ( .B(\modmult_1/xin[1023] ), .A(n34702), .Z(n34700) );
  IV U36158 ( .A(n34701), .Z(n34702) );
  XNOR U36159 ( .A(m[811]), .B(n34703), .Z(n34701) );
  NAND U36160 ( .A(n34704), .B(mul_pow), .Z(n34703) );
  XOR U36161 ( .A(m[811]), .B(c[811]), .Z(n34704) );
  XOR U36162 ( .A(n34705), .B(n34706), .Z(n34697) );
  ANDN U36163 ( .B(n34707), .A(n32366), .Z(n34705) );
  XNOR U36164 ( .A(\modmult_1/zin[0][809] ), .B(n34708), .Z(n32366) );
  IV U36165 ( .A(n34706), .Z(n34708) );
  XOR U36166 ( .A(n34706), .B(n32367), .Z(n34707) );
  XNOR U36167 ( .A(n34709), .B(n34710), .Z(n32367) );
  ANDN U36168 ( .B(\modmult_1/xin[1023] ), .A(n34711), .Z(n34709) );
  IV U36169 ( .A(n34710), .Z(n34711) );
  XNOR U36170 ( .A(m[810]), .B(n34712), .Z(n34710) );
  NAND U36171 ( .A(n34713), .B(mul_pow), .Z(n34712) );
  XOR U36172 ( .A(m[810]), .B(c[810]), .Z(n34713) );
  XOR U36173 ( .A(n34714), .B(n34715), .Z(n34706) );
  ANDN U36174 ( .B(n34716), .A(n32364), .Z(n34714) );
  XNOR U36175 ( .A(\modmult_1/zin[0][808] ), .B(n34717), .Z(n32364) );
  IV U36176 ( .A(n34715), .Z(n34717) );
  XOR U36177 ( .A(n34715), .B(n32365), .Z(n34716) );
  XNOR U36178 ( .A(n34718), .B(n34719), .Z(n32365) );
  ANDN U36179 ( .B(\modmult_1/xin[1023] ), .A(n34720), .Z(n34718) );
  IV U36180 ( .A(n34719), .Z(n34720) );
  XNOR U36181 ( .A(m[809]), .B(n34721), .Z(n34719) );
  NAND U36182 ( .A(n34722), .B(mul_pow), .Z(n34721) );
  XOR U36183 ( .A(m[809]), .B(c[809]), .Z(n34722) );
  XOR U36184 ( .A(n34723), .B(n34724), .Z(n34715) );
  ANDN U36185 ( .B(n34725), .A(n32362), .Z(n34723) );
  XNOR U36186 ( .A(\modmult_1/zin[0][807] ), .B(n34726), .Z(n32362) );
  IV U36187 ( .A(n34724), .Z(n34726) );
  XOR U36188 ( .A(n34724), .B(n32363), .Z(n34725) );
  XNOR U36189 ( .A(n34727), .B(n34728), .Z(n32363) );
  ANDN U36190 ( .B(\modmult_1/xin[1023] ), .A(n34729), .Z(n34727) );
  IV U36191 ( .A(n34728), .Z(n34729) );
  XNOR U36192 ( .A(m[808]), .B(n34730), .Z(n34728) );
  NAND U36193 ( .A(n34731), .B(mul_pow), .Z(n34730) );
  XOR U36194 ( .A(m[808]), .B(c[808]), .Z(n34731) );
  XOR U36195 ( .A(n34732), .B(n34733), .Z(n34724) );
  ANDN U36196 ( .B(n34734), .A(n32360), .Z(n34732) );
  XNOR U36197 ( .A(\modmult_1/zin[0][806] ), .B(n34735), .Z(n32360) );
  IV U36198 ( .A(n34733), .Z(n34735) );
  XOR U36199 ( .A(n34733), .B(n32361), .Z(n34734) );
  XNOR U36200 ( .A(n34736), .B(n34737), .Z(n32361) );
  ANDN U36201 ( .B(\modmult_1/xin[1023] ), .A(n34738), .Z(n34736) );
  IV U36202 ( .A(n34737), .Z(n34738) );
  XNOR U36203 ( .A(m[807]), .B(n34739), .Z(n34737) );
  NAND U36204 ( .A(n34740), .B(mul_pow), .Z(n34739) );
  XOR U36205 ( .A(m[807]), .B(c[807]), .Z(n34740) );
  XOR U36206 ( .A(n34741), .B(n34742), .Z(n34733) );
  ANDN U36207 ( .B(n34743), .A(n32358), .Z(n34741) );
  XNOR U36208 ( .A(\modmult_1/zin[0][805] ), .B(n34744), .Z(n32358) );
  IV U36209 ( .A(n34742), .Z(n34744) );
  XOR U36210 ( .A(n34742), .B(n32359), .Z(n34743) );
  XNOR U36211 ( .A(n34745), .B(n34746), .Z(n32359) );
  ANDN U36212 ( .B(\modmult_1/xin[1023] ), .A(n34747), .Z(n34745) );
  IV U36213 ( .A(n34746), .Z(n34747) );
  XNOR U36214 ( .A(m[806]), .B(n34748), .Z(n34746) );
  NAND U36215 ( .A(n34749), .B(mul_pow), .Z(n34748) );
  XOR U36216 ( .A(m[806]), .B(c[806]), .Z(n34749) );
  XOR U36217 ( .A(n34750), .B(n34751), .Z(n34742) );
  ANDN U36218 ( .B(n34752), .A(n32356), .Z(n34750) );
  XNOR U36219 ( .A(\modmult_1/zin[0][804] ), .B(n34753), .Z(n32356) );
  IV U36220 ( .A(n34751), .Z(n34753) );
  XOR U36221 ( .A(n34751), .B(n32357), .Z(n34752) );
  XNOR U36222 ( .A(n34754), .B(n34755), .Z(n32357) );
  ANDN U36223 ( .B(\modmult_1/xin[1023] ), .A(n34756), .Z(n34754) );
  IV U36224 ( .A(n34755), .Z(n34756) );
  XNOR U36225 ( .A(m[805]), .B(n34757), .Z(n34755) );
  NAND U36226 ( .A(n34758), .B(mul_pow), .Z(n34757) );
  XOR U36227 ( .A(m[805]), .B(c[805]), .Z(n34758) );
  XOR U36228 ( .A(n34759), .B(n34760), .Z(n34751) );
  ANDN U36229 ( .B(n34761), .A(n32354), .Z(n34759) );
  XNOR U36230 ( .A(\modmult_1/zin[0][803] ), .B(n34762), .Z(n32354) );
  IV U36231 ( .A(n34760), .Z(n34762) );
  XOR U36232 ( .A(n34760), .B(n32355), .Z(n34761) );
  XNOR U36233 ( .A(n34763), .B(n34764), .Z(n32355) );
  ANDN U36234 ( .B(\modmult_1/xin[1023] ), .A(n34765), .Z(n34763) );
  IV U36235 ( .A(n34764), .Z(n34765) );
  XNOR U36236 ( .A(m[804]), .B(n34766), .Z(n34764) );
  NAND U36237 ( .A(n34767), .B(mul_pow), .Z(n34766) );
  XOR U36238 ( .A(m[804]), .B(c[804]), .Z(n34767) );
  XOR U36239 ( .A(n34768), .B(n34769), .Z(n34760) );
  ANDN U36240 ( .B(n34770), .A(n32352), .Z(n34768) );
  XNOR U36241 ( .A(\modmult_1/zin[0][802] ), .B(n34771), .Z(n32352) );
  IV U36242 ( .A(n34769), .Z(n34771) );
  XOR U36243 ( .A(n34769), .B(n32353), .Z(n34770) );
  XNOR U36244 ( .A(n34772), .B(n34773), .Z(n32353) );
  ANDN U36245 ( .B(\modmult_1/xin[1023] ), .A(n34774), .Z(n34772) );
  IV U36246 ( .A(n34773), .Z(n34774) );
  XNOR U36247 ( .A(m[803]), .B(n34775), .Z(n34773) );
  NAND U36248 ( .A(n34776), .B(mul_pow), .Z(n34775) );
  XOR U36249 ( .A(m[803]), .B(c[803]), .Z(n34776) );
  XOR U36250 ( .A(n34777), .B(n34778), .Z(n34769) );
  ANDN U36251 ( .B(n34779), .A(n32350), .Z(n34777) );
  XNOR U36252 ( .A(\modmult_1/zin[0][801] ), .B(n34780), .Z(n32350) );
  IV U36253 ( .A(n34778), .Z(n34780) );
  XOR U36254 ( .A(n34778), .B(n32351), .Z(n34779) );
  XNOR U36255 ( .A(n34781), .B(n34782), .Z(n32351) );
  ANDN U36256 ( .B(\modmult_1/xin[1023] ), .A(n34783), .Z(n34781) );
  IV U36257 ( .A(n34782), .Z(n34783) );
  XNOR U36258 ( .A(m[802]), .B(n34784), .Z(n34782) );
  NAND U36259 ( .A(n34785), .B(mul_pow), .Z(n34784) );
  XOR U36260 ( .A(m[802]), .B(c[802]), .Z(n34785) );
  XOR U36261 ( .A(n34786), .B(n34787), .Z(n34778) );
  ANDN U36262 ( .B(n34788), .A(n32348), .Z(n34786) );
  XNOR U36263 ( .A(\modmult_1/zin[0][800] ), .B(n34789), .Z(n32348) );
  IV U36264 ( .A(n34787), .Z(n34789) );
  XOR U36265 ( .A(n34787), .B(n32349), .Z(n34788) );
  XNOR U36266 ( .A(n34790), .B(n34791), .Z(n32349) );
  ANDN U36267 ( .B(\modmult_1/xin[1023] ), .A(n34792), .Z(n34790) );
  IV U36268 ( .A(n34791), .Z(n34792) );
  XNOR U36269 ( .A(m[801]), .B(n34793), .Z(n34791) );
  NAND U36270 ( .A(n34794), .B(mul_pow), .Z(n34793) );
  XOR U36271 ( .A(m[801]), .B(c[801]), .Z(n34794) );
  XOR U36272 ( .A(n34795), .B(n34796), .Z(n34787) );
  ANDN U36273 ( .B(n34797), .A(n32346), .Z(n34795) );
  XNOR U36274 ( .A(\modmult_1/zin[0][799] ), .B(n34798), .Z(n32346) );
  IV U36275 ( .A(n34796), .Z(n34798) );
  XOR U36276 ( .A(n34796), .B(n32347), .Z(n34797) );
  XNOR U36277 ( .A(n34799), .B(n34800), .Z(n32347) );
  ANDN U36278 ( .B(\modmult_1/xin[1023] ), .A(n34801), .Z(n34799) );
  IV U36279 ( .A(n34800), .Z(n34801) );
  XNOR U36280 ( .A(m[800]), .B(n34802), .Z(n34800) );
  NAND U36281 ( .A(n34803), .B(mul_pow), .Z(n34802) );
  XOR U36282 ( .A(m[800]), .B(c[800]), .Z(n34803) );
  XOR U36283 ( .A(n34804), .B(n34805), .Z(n34796) );
  ANDN U36284 ( .B(n34806), .A(n32344), .Z(n34804) );
  XNOR U36285 ( .A(\modmult_1/zin[0][798] ), .B(n34807), .Z(n32344) );
  IV U36286 ( .A(n34805), .Z(n34807) );
  XOR U36287 ( .A(n34805), .B(n32345), .Z(n34806) );
  XNOR U36288 ( .A(n34808), .B(n34809), .Z(n32345) );
  ANDN U36289 ( .B(\modmult_1/xin[1023] ), .A(n34810), .Z(n34808) );
  IV U36290 ( .A(n34809), .Z(n34810) );
  XNOR U36291 ( .A(m[799]), .B(n34811), .Z(n34809) );
  NAND U36292 ( .A(n34812), .B(mul_pow), .Z(n34811) );
  XOR U36293 ( .A(m[799]), .B(c[799]), .Z(n34812) );
  XOR U36294 ( .A(n34813), .B(n34814), .Z(n34805) );
  ANDN U36295 ( .B(n34815), .A(n32342), .Z(n34813) );
  XNOR U36296 ( .A(\modmult_1/zin[0][797] ), .B(n34816), .Z(n32342) );
  IV U36297 ( .A(n34814), .Z(n34816) );
  XOR U36298 ( .A(n34814), .B(n32343), .Z(n34815) );
  XNOR U36299 ( .A(n34817), .B(n34818), .Z(n32343) );
  ANDN U36300 ( .B(\modmult_1/xin[1023] ), .A(n34819), .Z(n34817) );
  IV U36301 ( .A(n34818), .Z(n34819) );
  XNOR U36302 ( .A(m[798]), .B(n34820), .Z(n34818) );
  NAND U36303 ( .A(n34821), .B(mul_pow), .Z(n34820) );
  XOR U36304 ( .A(m[798]), .B(c[798]), .Z(n34821) );
  XOR U36305 ( .A(n34822), .B(n34823), .Z(n34814) );
  ANDN U36306 ( .B(n34824), .A(n32340), .Z(n34822) );
  XNOR U36307 ( .A(\modmult_1/zin[0][796] ), .B(n34825), .Z(n32340) );
  IV U36308 ( .A(n34823), .Z(n34825) );
  XOR U36309 ( .A(n34823), .B(n32341), .Z(n34824) );
  XNOR U36310 ( .A(n34826), .B(n34827), .Z(n32341) );
  ANDN U36311 ( .B(\modmult_1/xin[1023] ), .A(n34828), .Z(n34826) );
  IV U36312 ( .A(n34827), .Z(n34828) );
  XNOR U36313 ( .A(m[797]), .B(n34829), .Z(n34827) );
  NAND U36314 ( .A(n34830), .B(mul_pow), .Z(n34829) );
  XOR U36315 ( .A(m[797]), .B(c[797]), .Z(n34830) );
  XOR U36316 ( .A(n34831), .B(n34832), .Z(n34823) );
  ANDN U36317 ( .B(n34833), .A(n32338), .Z(n34831) );
  XNOR U36318 ( .A(\modmult_1/zin[0][795] ), .B(n34834), .Z(n32338) );
  IV U36319 ( .A(n34832), .Z(n34834) );
  XOR U36320 ( .A(n34832), .B(n32339), .Z(n34833) );
  XNOR U36321 ( .A(n34835), .B(n34836), .Z(n32339) );
  ANDN U36322 ( .B(\modmult_1/xin[1023] ), .A(n34837), .Z(n34835) );
  IV U36323 ( .A(n34836), .Z(n34837) );
  XNOR U36324 ( .A(m[796]), .B(n34838), .Z(n34836) );
  NAND U36325 ( .A(n34839), .B(mul_pow), .Z(n34838) );
  XOR U36326 ( .A(m[796]), .B(c[796]), .Z(n34839) );
  XOR U36327 ( .A(n34840), .B(n34841), .Z(n34832) );
  ANDN U36328 ( .B(n34842), .A(n32336), .Z(n34840) );
  XNOR U36329 ( .A(\modmult_1/zin[0][794] ), .B(n34843), .Z(n32336) );
  IV U36330 ( .A(n34841), .Z(n34843) );
  XOR U36331 ( .A(n34841), .B(n32337), .Z(n34842) );
  XNOR U36332 ( .A(n34844), .B(n34845), .Z(n32337) );
  ANDN U36333 ( .B(\modmult_1/xin[1023] ), .A(n34846), .Z(n34844) );
  IV U36334 ( .A(n34845), .Z(n34846) );
  XNOR U36335 ( .A(m[795]), .B(n34847), .Z(n34845) );
  NAND U36336 ( .A(n34848), .B(mul_pow), .Z(n34847) );
  XOR U36337 ( .A(m[795]), .B(c[795]), .Z(n34848) );
  XOR U36338 ( .A(n34849), .B(n34850), .Z(n34841) );
  ANDN U36339 ( .B(n34851), .A(n32334), .Z(n34849) );
  XNOR U36340 ( .A(\modmult_1/zin[0][793] ), .B(n34852), .Z(n32334) );
  IV U36341 ( .A(n34850), .Z(n34852) );
  XOR U36342 ( .A(n34850), .B(n32335), .Z(n34851) );
  XNOR U36343 ( .A(n34853), .B(n34854), .Z(n32335) );
  ANDN U36344 ( .B(\modmult_1/xin[1023] ), .A(n34855), .Z(n34853) );
  IV U36345 ( .A(n34854), .Z(n34855) );
  XNOR U36346 ( .A(m[794]), .B(n34856), .Z(n34854) );
  NAND U36347 ( .A(n34857), .B(mul_pow), .Z(n34856) );
  XOR U36348 ( .A(m[794]), .B(c[794]), .Z(n34857) );
  XOR U36349 ( .A(n34858), .B(n34859), .Z(n34850) );
  ANDN U36350 ( .B(n34860), .A(n32332), .Z(n34858) );
  XNOR U36351 ( .A(\modmult_1/zin[0][792] ), .B(n34861), .Z(n32332) );
  IV U36352 ( .A(n34859), .Z(n34861) );
  XOR U36353 ( .A(n34859), .B(n32333), .Z(n34860) );
  XNOR U36354 ( .A(n34862), .B(n34863), .Z(n32333) );
  ANDN U36355 ( .B(\modmult_1/xin[1023] ), .A(n34864), .Z(n34862) );
  IV U36356 ( .A(n34863), .Z(n34864) );
  XNOR U36357 ( .A(m[793]), .B(n34865), .Z(n34863) );
  NAND U36358 ( .A(n34866), .B(mul_pow), .Z(n34865) );
  XOR U36359 ( .A(m[793]), .B(c[793]), .Z(n34866) );
  XOR U36360 ( .A(n34867), .B(n34868), .Z(n34859) );
  ANDN U36361 ( .B(n34869), .A(n32330), .Z(n34867) );
  XNOR U36362 ( .A(\modmult_1/zin[0][791] ), .B(n34870), .Z(n32330) );
  IV U36363 ( .A(n34868), .Z(n34870) );
  XOR U36364 ( .A(n34868), .B(n32331), .Z(n34869) );
  XNOR U36365 ( .A(n34871), .B(n34872), .Z(n32331) );
  ANDN U36366 ( .B(\modmult_1/xin[1023] ), .A(n34873), .Z(n34871) );
  IV U36367 ( .A(n34872), .Z(n34873) );
  XNOR U36368 ( .A(m[792]), .B(n34874), .Z(n34872) );
  NAND U36369 ( .A(n34875), .B(mul_pow), .Z(n34874) );
  XOR U36370 ( .A(m[792]), .B(c[792]), .Z(n34875) );
  XOR U36371 ( .A(n34876), .B(n34877), .Z(n34868) );
  ANDN U36372 ( .B(n34878), .A(n32328), .Z(n34876) );
  XNOR U36373 ( .A(\modmult_1/zin[0][790] ), .B(n34879), .Z(n32328) );
  IV U36374 ( .A(n34877), .Z(n34879) );
  XOR U36375 ( .A(n34877), .B(n32329), .Z(n34878) );
  XNOR U36376 ( .A(n34880), .B(n34881), .Z(n32329) );
  ANDN U36377 ( .B(\modmult_1/xin[1023] ), .A(n34882), .Z(n34880) );
  IV U36378 ( .A(n34881), .Z(n34882) );
  XNOR U36379 ( .A(m[791]), .B(n34883), .Z(n34881) );
  NAND U36380 ( .A(n34884), .B(mul_pow), .Z(n34883) );
  XOR U36381 ( .A(m[791]), .B(c[791]), .Z(n34884) );
  XOR U36382 ( .A(n34885), .B(n34886), .Z(n34877) );
  ANDN U36383 ( .B(n34887), .A(n32326), .Z(n34885) );
  XNOR U36384 ( .A(\modmult_1/zin[0][789] ), .B(n34888), .Z(n32326) );
  IV U36385 ( .A(n34886), .Z(n34888) );
  XOR U36386 ( .A(n34886), .B(n32327), .Z(n34887) );
  XNOR U36387 ( .A(n34889), .B(n34890), .Z(n32327) );
  ANDN U36388 ( .B(\modmult_1/xin[1023] ), .A(n34891), .Z(n34889) );
  IV U36389 ( .A(n34890), .Z(n34891) );
  XNOR U36390 ( .A(m[790]), .B(n34892), .Z(n34890) );
  NAND U36391 ( .A(n34893), .B(mul_pow), .Z(n34892) );
  XOR U36392 ( .A(m[790]), .B(c[790]), .Z(n34893) );
  XOR U36393 ( .A(n34894), .B(n34895), .Z(n34886) );
  ANDN U36394 ( .B(n34896), .A(n32324), .Z(n34894) );
  XNOR U36395 ( .A(\modmult_1/zin[0][788] ), .B(n34897), .Z(n32324) );
  IV U36396 ( .A(n34895), .Z(n34897) );
  XOR U36397 ( .A(n34895), .B(n32325), .Z(n34896) );
  XNOR U36398 ( .A(n34898), .B(n34899), .Z(n32325) );
  ANDN U36399 ( .B(\modmult_1/xin[1023] ), .A(n34900), .Z(n34898) );
  IV U36400 ( .A(n34899), .Z(n34900) );
  XNOR U36401 ( .A(m[789]), .B(n34901), .Z(n34899) );
  NAND U36402 ( .A(n34902), .B(mul_pow), .Z(n34901) );
  XOR U36403 ( .A(m[789]), .B(c[789]), .Z(n34902) );
  XOR U36404 ( .A(n34903), .B(n34904), .Z(n34895) );
  ANDN U36405 ( .B(n34905), .A(n32322), .Z(n34903) );
  XNOR U36406 ( .A(\modmult_1/zin[0][787] ), .B(n34906), .Z(n32322) );
  IV U36407 ( .A(n34904), .Z(n34906) );
  XOR U36408 ( .A(n34904), .B(n32323), .Z(n34905) );
  XNOR U36409 ( .A(n34907), .B(n34908), .Z(n32323) );
  ANDN U36410 ( .B(\modmult_1/xin[1023] ), .A(n34909), .Z(n34907) );
  IV U36411 ( .A(n34908), .Z(n34909) );
  XNOR U36412 ( .A(m[788]), .B(n34910), .Z(n34908) );
  NAND U36413 ( .A(n34911), .B(mul_pow), .Z(n34910) );
  XOR U36414 ( .A(m[788]), .B(c[788]), .Z(n34911) );
  XOR U36415 ( .A(n34912), .B(n34913), .Z(n34904) );
  ANDN U36416 ( .B(n34914), .A(n32320), .Z(n34912) );
  XNOR U36417 ( .A(\modmult_1/zin[0][786] ), .B(n34915), .Z(n32320) );
  IV U36418 ( .A(n34913), .Z(n34915) );
  XOR U36419 ( .A(n34913), .B(n32321), .Z(n34914) );
  XNOR U36420 ( .A(n34916), .B(n34917), .Z(n32321) );
  ANDN U36421 ( .B(\modmult_1/xin[1023] ), .A(n34918), .Z(n34916) );
  IV U36422 ( .A(n34917), .Z(n34918) );
  XNOR U36423 ( .A(m[787]), .B(n34919), .Z(n34917) );
  NAND U36424 ( .A(n34920), .B(mul_pow), .Z(n34919) );
  XOR U36425 ( .A(m[787]), .B(c[787]), .Z(n34920) );
  XOR U36426 ( .A(n34921), .B(n34922), .Z(n34913) );
  ANDN U36427 ( .B(n34923), .A(n32318), .Z(n34921) );
  XNOR U36428 ( .A(\modmult_1/zin[0][785] ), .B(n34924), .Z(n32318) );
  IV U36429 ( .A(n34922), .Z(n34924) );
  XOR U36430 ( .A(n34922), .B(n32319), .Z(n34923) );
  XNOR U36431 ( .A(n34925), .B(n34926), .Z(n32319) );
  ANDN U36432 ( .B(\modmult_1/xin[1023] ), .A(n34927), .Z(n34925) );
  IV U36433 ( .A(n34926), .Z(n34927) );
  XNOR U36434 ( .A(m[786]), .B(n34928), .Z(n34926) );
  NAND U36435 ( .A(n34929), .B(mul_pow), .Z(n34928) );
  XOR U36436 ( .A(m[786]), .B(c[786]), .Z(n34929) );
  XOR U36437 ( .A(n34930), .B(n34931), .Z(n34922) );
  ANDN U36438 ( .B(n34932), .A(n32316), .Z(n34930) );
  XNOR U36439 ( .A(\modmult_1/zin[0][784] ), .B(n34933), .Z(n32316) );
  IV U36440 ( .A(n34931), .Z(n34933) );
  XOR U36441 ( .A(n34931), .B(n32317), .Z(n34932) );
  XNOR U36442 ( .A(n34934), .B(n34935), .Z(n32317) );
  ANDN U36443 ( .B(\modmult_1/xin[1023] ), .A(n34936), .Z(n34934) );
  IV U36444 ( .A(n34935), .Z(n34936) );
  XNOR U36445 ( .A(m[785]), .B(n34937), .Z(n34935) );
  NAND U36446 ( .A(n34938), .B(mul_pow), .Z(n34937) );
  XOR U36447 ( .A(m[785]), .B(c[785]), .Z(n34938) );
  XOR U36448 ( .A(n34939), .B(n34940), .Z(n34931) );
  ANDN U36449 ( .B(n34941), .A(n32314), .Z(n34939) );
  XNOR U36450 ( .A(\modmult_1/zin[0][783] ), .B(n34942), .Z(n32314) );
  IV U36451 ( .A(n34940), .Z(n34942) );
  XOR U36452 ( .A(n34940), .B(n32315), .Z(n34941) );
  XNOR U36453 ( .A(n34943), .B(n34944), .Z(n32315) );
  ANDN U36454 ( .B(\modmult_1/xin[1023] ), .A(n34945), .Z(n34943) );
  IV U36455 ( .A(n34944), .Z(n34945) );
  XNOR U36456 ( .A(m[784]), .B(n34946), .Z(n34944) );
  NAND U36457 ( .A(n34947), .B(mul_pow), .Z(n34946) );
  XOR U36458 ( .A(m[784]), .B(c[784]), .Z(n34947) );
  XOR U36459 ( .A(n34948), .B(n34949), .Z(n34940) );
  ANDN U36460 ( .B(n34950), .A(n32312), .Z(n34948) );
  XNOR U36461 ( .A(\modmult_1/zin[0][782] ), .B(n34951), .Z(n32312) );
  IV U36462 ( .A(n34949), .Z(n34951) );
  XOR U36463 ( .A(n34949), .B(n32313), .Z(n34950) );
  XNOR U36464 ( .A(n34952), .B(n34953), .Z(n32313) );
  ANDN U36465 ( .B(\modmult_1/xin[1023] ), .A(n34954), .Z(n34952) );
  IV U36466 ( .A(n34953), .Z(n34954) );
  XNOR U36467 ( .A(m[783]), .B(n34955), .Z(n34953) );
  NAND U36468 ( .A(n34956), .B(mul_pow), .Z(n34955) );
  XOR U36469 ( .A(m[783]), .B(c[783]), .Z(n34956) );
  XOR U36470 ( .A(n34957), .B(n34958), .Z(n34949) );
  ANDN U36471 ( .B(n34959), .A(n32310), .Z(n34957) );
  XNOR U36472 ( .A(\modmult_1/zin[0][781] ), .B(n34960), .Z(n32310) );
  IV U36473 ( .A(n34958), .Z(n34960) );
  XOR U36474 ( .A(n34958), .B(n32311), .Z(n34959) );
  XNOR U36475 ( .A(n34961), .B(n34962), .Z(n32311) );
  ANDN U36476 ( .B(\modmult_1/xin[1023] ), .A(n34963), .Z(n34961) );
  IV U36477 ( .A(n34962), .Z(n34963) );
  XNOR U36478 ( .A(m[782]), .B(n34964), .Z(n34962) );
  NAND U36479 ( .A(n34965), .B(mul_pow), .Z(n34964) );
  XOR U36480 ( .A(m[782]), .B(c[782]), .Z(n34965) );
  XOR U36481 ( .A(n34966), .B(n34967), .Z(n34958) );
  ANDN U36482 ( .B(n34968), .A(n32308), .Z(n34966) );
  XNOR U36483 ( .A(\modmult_1/zin[0][780] ), .B(n34969), .Z(n32308) );
  IV U36484 ( .A(n34967), .Z(n34969) );
  XOR U36485 ( .A(n34967), .B(n32309), .Z(n34968) );
  XNOR U36486 ( .A(n34970), .B(n34971), .Z(n32309) );
  ANDN U36487 ( .B(\modmult_1/xin[1023] ), .A(n34972), .Z(n34970) );
  IV U36488 ( .A(n34971), .Z(n34972) );
  XNOR U36489 ( .A(m[781]), .B(n34973), .Z(n34971) );
  NAND U36490 ( .A(n34974), .B(mul_pow), .Z(n34973) );
  XOR U36491 ( .A(m[781]), .B(c[781]), .Z(n34974) );
  XOR U36492 ( .A(n34975), .B(n34976), .Z(n34967) );
  ANDN U36493 ( .B(n34977), .A(n32306), .Z(n34975) );
  XNOR U36494 ( .A(\modmult_1/zin[0][779] ), .B(n34978), .Z(n32306) );
  IV U36495 ( .A(n34976), .Z(n34978) );
  XOR U36496 ( .A(n34976), .B(n32307), .Z(n34977) );
  XNOR U36497 ( .A(n34979), .B(n34980), .Z(n32307) );
  ANDN U36498 ( .B(\modmult_1/xin[1023] ), .A(n34981), .Z(n34979) );
  IV U36499 ( .A(n34980), .Z(n34981) );
  XNOR U36500 ( .A(m[780]), .B(n34982), .Z(n34980) );
  NAND U36501 ( .A(n34983), .B(mul_pow), .Z(n34982) );
  XOR U36502 ( .A(m[780]), .B(c[780]), .Z(n34983) );
  XOR U36503 ( .A(n34984), .B(n34985), .Z(n34976) );
  ANDN U36504 ( .B(n34986), .A(n32304), .Z(n34984) );
  XNOR U36505 ( .A(\modmult_1/zin[0][778] ), .B(n34987), .Z(n32304) );
  IV U36506 ( .A(n34985), .Z(n34987) );
  XOR U36507 ( .A(n34985), .B(n32305), .Z(n34986) );
  XNOR U36508 ( .A(n34988), .B(n34989), .Z(n32305) );
  ANDN U36509 ( .B(\modmult_1/xin[1023] ), .A(n34990), .Z(n34988) );
  IV U36510 ( .A(n34989), .Z(n34990) );
  XNOR U36511 ( .A(m[779]), .B(n34991), .Z(n34989) );
  NAND U36512 ( .A(n34992), .B(mul_pow), .Z(n34991) );
  XOR U36513 ( .A(m[779]), .B(c[779]), .Z(n34992) );
  XOR U36514 ( .A(n34993), .B(n34994), .Z(n34985) );
  ANDN U36515 ( .B(n34995), .A(n32302), .Z(n34993) );
  XNOR U36516 ( .A(\modmult_1/zin[0][777] ), .B(n34996), .Z(n32302) );
  IV U36517 ( .A(n34994), .Z(n34996) );
  XOR U36518 ( .A(n34994), .B(n32303), .Z(n34995) );
  XNOR U36519 ( .A(n34997), .B(n34998), .Z(n32303) );
  ANDN U36520 ( .B(\modmult_1/xin[1023] ), .A(n34999), .Z(n34997) );
  IV U36521 ( .A(n34998), .Z(n34999) );
  XNOR U36522 ( .A(m[778]), .B(n35000), .Z(n34998) );
  NAND U36523 ( .A(n35001), .B(mul_pow), .Z(n35000) );
  XOR U36524 ( .A(m[778]), .B(c[778]), .Z(n35001) );
  XOR U36525 ( .A(n35002), .B(n35003), .Z(n34994) );
  ANDN U36526 ( .B(n35004), .A(n32300), .Z(n35002) );
  XNOR U36527 ( .A(\modmult_1/zin[0][776] ), .B(n35005), .Z(n32300) );
  IV U36528 ( .A(n35003), .Z(n35005) );
  XOR U36529 ( .A(n35003), .B(n32301), .Z(n35004) );
  XNOR U36530 ( .A(n35006), .B(n35007), .Z(n32301) );
  ANDN U36531 ( .B(\modmult_1/xin[1023] ), .A(n35008), .Z(n35006) );
  IV U36532 ( .A(n35007), .Z(n35008) );
  XNOR U36533 ( .A(m[777]), .B(n35009), .Z(n35007) );
  NAND U36534 ( .A(n35010), .B(mul_pow), .Z(n35009) );
  XOR U36535 ( .A(m[777]), .B(c[777]), .Z(n35010) );
  XOR U36536 ( .A(n35011), .B(n35012), .Z(n35003) );
  ANDN U36537 ( .B(n35013), .A(n32298), .Z(n35011) );
  XNOR U36538 ( .A(\modmult_1/zin[0][775] ), .B(n35014), .Z(n32298) );
  IV U36539 ( .A(n35012), .Z(n35014) );
  XOR U36540 ( .A(n35012), .B(n32299), .Z(n35013) );
  XNOR U36541 ( .A(n35015), .B(n35016), .Z(n32299) );
  ANDN U36542 ( .B(\modmult_1/xin[1023] ), .A(n35017), .Z(n35015) );
  IV U36543 ( .A(n35016), .Z(n35017) );
  XNOR U36544 ( .A(m[776]), .B(n35018), .Z(n35016) );
  NAND U36545 ( .A(n35019), .B(mul_pow), .Z(n35018) );
  XOR U36546 ( .A(m[776]), .B(c[776]), .Z(n35019) );
  XOR U36547 ( .A(n35020), .B(n35021), .Z(n35012) );
  ANDN U36548 ( .B(n35022), .A(n32296), .Z(n35020) );
  XNOR U36549 ( .A(\modmult_1/zin[0][774] ), .B(n35023), .Z(n32296) );
  IV U36550 ( .A(n35021), .Z(n35023) );
  XOR U36551 ( .A(n35021), .B(n32297), .Z(n35022) );
  XNOR U36552 ( .A(n35024), .B(n35025), .Z(n32297) );
  ANDN U36553 ( .B(\modmult_1/xin[1023] ), .A(n35026), .Z(n35024) );
  IV U36554 ( .A(n35025), .Z(n35026) );
  XNOR U36555 ( .A(m[775]), .B(n35027), .Z(n35025) );
  NAND U36556 ( .A(n35028), .B(mul_pow), .Z(n35027) );
  XOR U36557 ( .A(m[775]), .B(c[775]), .Z(n35028) );
  XOR U36558 ( .A(n35029), .B(n35030), .Z(n35021) );
  ANDN U36559 ( .B(n35031), .A(n32294), .Z(n35029) );
  XNOR U36560 ( .A(\modmult_1/zin[0][773] ), .B(n35032), .Z(n32294) );
  IV U36561 ( .A(n35030), .Z(n35032) );
  XOR U36562 ( .A(n35030), .B(n32295), .Z(n35031) );
  XNOR U36563 ( .A(n35033), .B(n35034), .Z(n32295) );
  ANDN U36564 ( .B(\modmult_1/xin[1023] ), .A(n35035), .Z(n35033) );
  IV U36565 ( .A(n35034), .Z(n35035) );
  XNOR U36566 ( .A(m[774]), .B(n35036), .Z(n35034) );
  NAND U36567 ( .A(n35037), .B(mul_pow), .Z(n35036) );
  XOR U36568 ( .A(m[774]), .B(c[774]), .Z(n35037) );
  XOR U36569 ( .A(n35038), .B(n35039), .Z(n35030) );
  ANDN U36570 ( .B(n35040), .A(n32292), .Z(n35038) );
  XNOR U36571 ( .A(\modmult_1/zin[0][772] ), .B(n35041), .Z(n32292) );
  IV U36572 ( .A(n35039), .Z(n35041) );
  XOR U36573 ( .A(n35039), .B(n32293), .Z(n35040) );
  XNOR U36574 ( .A(n35042), .B(n35043), .Z(n32293) );
  ANDN U36575 ( .B(\modmult_1/xin[1023] ), .A(n35044), .Z(n35042) );
  IV U36576 ( .A(n35043), .Z(n35044) );
  XNOR U36577 ( .A(m[773]), .B(n35045), .Z(n35043) );
  NAND U36578 ( .A(n35046), .B(mul_pow), .Z(n35045) );
  XOR U36579 ( .A(m[773]), .B(c[773]), .Z(n35046) );
  XOR U36580 ( .A(n35047), .B(n35048), .Z(n35039) );
  ANDN U36581 ( .B(n35049), .A(n32290), .Z(n35047) );
  XNOR U36582 ( .A(\modmult_1/zin[0][771] ), .B(n35050), .Z(n32290) );
  IV U36583 ( .A(n35048), .Z(n35050) );
  XOR U36584 ( .A(n35048), .B(n32291), .Z(n35049) );
  XNOR U36585 ( .A(n35051), .B(n35052), .Z(n32291) );
  ANDN U36586 ( .B(\modmult_1/xin[1023] ), .A(n35053), .Z(n35051) );
  IV U36587 ( .A(n35052), .Z(n35053) );
  XNOR U36588 ( .A(m[772]), .B(n35054), .Z(n35052) );
  NAND U36589 ( .A(n35055), .B(mul_pow), .Z(n35054) );
  XOR U36590 ( .A(m[772]), .B(c[772]), .Z(n35055) );
  XOR U36591 ( .A(n35056), .B(n35057), .Z(n35048) );
  ANDN U36592 ( .B(n35058), .A(n32288), .Z(n35056) );
  XNOR U36593 ( .A(\modmult_1/zin[0][770] ), .B(n35059), .Z(n32288) );
  IV U36594 ( .A(n35057), .Z(n35059) );
  XOR U36595 ( .A(n35057), .B(n32289), .Z(n35058) );
  XNOR U36596 ( .A(n35060), .B(n35061), .Z(n32289) );
  ANDN U36597 ( .B(\modmult_1/xin[1023] ), .A(n35062), .Z(n35060) );
  IV U36598 ( .A(n35061), .Z(n35062) );
  XNOR U36599 ( .A(m[771]), .B(n35063), .Z(n35061) );
  NAND U36600 ( .A(n35064), .B(mul_pow), .Z(n35063) );
  XOR U36601 ( .A(m[771]), .B(c[771]), .Z(n35064) );
  XOR U36602 ( .A(n35065), .B(n35066), .Z(n35057) );
  ANDN U36603 ( .B(n35067), .A(n32286), .Z(n35065) );
  XNOR U36604 ( .A(\modmult_1/zin[0][769] ), .B(n35068), .Z(n32286) );
  IV U36605 ( .A(n35066), .Z(n35068) );
  XOR U36606 ( .A(n35066), .B(n32287), .Z(n35067) );
  XNOR U36607 ( .A(n35069), .B(n35070), .Z(n32287) );
  ANDN U36608 ( .B(\modmult_1/xin[1023] ), .A(n35071), .Z(n35069) );
  IV U36609 ( .A(n35070), .Z(n35071) );
  XNOR U36610 ( .A(m[770]), .B(n35072), .Z(n35070) );
  NAND U36611 ( .A(n35073), .B(mul_pow), .Z(n35072) );
  XOR U36612 ( .A(m[770]), .B(c[770]), .Z(n35073) );
  XOR U36613 ( .A(n35074), .B(n35075), .Z(n35066) );
  ANDN U36614 ( .B(n35076), .A(n32284), .Z(n35074) );
  XNOR U36615 ( .A(\modmult_1/zin[0][768] ), .B(n35077), .Z(n32284) );
  IV U36616 ( .A(n35075), .Z(n35077) );
  XOR U36617 ( .A(n35075), .B(n32285), .Z(n35076) );
  XNOR U36618 ( .A(n35078), .B(n35079), .Z(n32285) );
  ANDN U36619 ( .B(\modmult_1/xin[1023] ), .A(n35080), .Z(n35078) );
  IV U36620 ( .A(n35079), .Z(n35080) );
  XNOR U36621 ( .A(m[769]), .B(n35081), .Z(n35079) );
  NAND U36622 ( .A(n35082), .B(mul_pow), .Z(n35081) );
  XOR U36623 ( .A(m[769]), .B(c[769]), .Z(n35082) );
  XOR U36624 ( .A(n35083), .B(n35084), .Z(n35075) );
  ANDN U36625 ( .B(n35085), .A(n32282), .Z(n35083) );
  XNOR U36626 ( .A(\modmult_1/zin[0][767] ), .B(n35086), .Z(n32282) );
  IV U36627 ( .A(n35084), .Z(n35086) );
  XOR U36628 ( .A(n35084), .B(n32283), .Z(n35085) );
  XNOR U36629 ( .A(n35087), .B(n35088), .Z(n32283) );
  ANDN U36630 ( .B(\modmult_1/xin[1023] ), .A(n35089), .Z(n35087) );
  IV U36631 ( .A(n35088), .Z(n35089) );
  XNOR U36632 ( .A(m[768]), .B(n35090), .Z(n35088) );
  NAND U36633 ( .A(n35091), .B(mul_pow), .Z(n35090) );
  XOR U36634 ( .A(m[768]), .B(c[768]), .Z(n35091) );
  XOR U36635 ( .A(n35092), .B(n35093), .Z(n35084) );
  ANDN U36636 ( .B(n35094), .A(n32280), .Z(n35092) );
  XNOR U36637 ( .A(\modmult_1/zin[0][766] ), .B(n35095), .Z(n32280) );
  IV U36638 ( .A(n35093), .Z(n35095) );
  XOR U36639 ( .A(n35093), .B(n32281), .Z(n35094) );
  XNOR U36640 ( .A(n35096), .B(n35097), .Z(n32281) );
  ANDN U36641 ( .B(\modmult_1/xin[1023] ), .A(n35098), .Z(n35096) );
  IV U36642 ( .A(n35097), .Z(n35098) );
  XNOR U36643 ( .A(m[767]), .B(n35099), .Z(n35097) );
  NAND U36644 ( .A(n35100), .B(mul_pow), .Z(n35099) );
  XOR U36645 ( .A(m[767]), .B(c[767]), .Z(n35100) );
  XOR U36646 ( .A(n35101), .B(n35102), .Z(n35093) );
  ANDN U36647 ( .B(n35103), .A(n32278), .Z(n35101) );
  XNOR U36648 ( .A(\modmult_1/zin[0][765] ), .B(n35104), .Z(n32278) );
  IV U36649 ( .A(n35102), .Z(n35104) );
  XOR U36650 ( .A(n35102), .B(n32279), .Z(n35103) );
  XNOR U36651 ( .A(n35105), .B(n35106), .Z(n32279) );
  ANDN U36652 ( .B(\modmult_1/xin[1023] ), .A(n35107), .Z(n35105) );
  IV U36653 ( .A(n35106), .Z(n35107) );
  XNOR U36654 ( .A(m[766]), .B(n35108), .Z(n35106) );
  NAND U36655 ( .A(n35109), .B(mul_pow), .Z(n35108) );
  XOR U36656 ( .A(m[766]), .B(c[766]), .Z(n35109) );
  XOR U36657 ( .A(n35110), .B(n35111), .Z(n35102) );
  ANDN U36658 ( .B(n35112), .A(n32276), .Z(n35110) );
  XNOR U36659 ( .A(\modmult_1/zin[0][764] ), .B(n35113), .Z(n32276) );
  IV U36660 ( .A(n35111), .Z(n35113) );
  XOR U36661 ( .A(n35111), .B(n32277), .Z(n35112) );
  XNOR U36662 ( .A(n35114), .B(n35115), .Z(n32277) );
  ANDN U36663 ( .B(\modmult_1/xin[1023] ), .A(n35116), .Z(n35114) );
  IV U36664 ( .A(n35115), .Z(n35116) );
  XNOR U36665 ( .A(m[765]), .B(n35117), .Z(n35115) );
  NAND U36666 ( .A(n35118), .B(mul_pow), .Z(n35117) );
  XOR U36667 ( .A(m[765]), .B(c[765]), .Z(n35118) );
  XOR U36668 ( .A(n35119), .B(n35120), .Z(n35111) );
  ANDN U36669 ( .B(n35121), .A(n32274), .Z(n35119) );
  XNOR U36670 ( .A(\modmult_1/zin[0][763] ), .B(n35122), .Z(n32274) );
  IV U36671 ( .A(n35120), .Z(n35122) );
  XOR U36672 ( .A(n35120), .B(n32275), .Z(n35121) );
  XNOR U36673 ( .A(n35123), .B(n35124), .Z(n32275) );
  ANDN U36674 ( .B(\modmult_1/xin[1023] ), .A(n35125), .Z(n35123) );
  IV U36675 ( .A(n35124), .Z(n35125) );
  XNOR U36676 ( .A(m[764]), .B(n35126), .Z(n35124) );
  NAND U36677 ( .A(n35127), .B(mul_pow), .Z(n35126) );
  XOR U36678 ( .A(m[764]), .B(c[764]), .Z(n35127) );
  XOR U36679 ( .A(n35128), .B(n35129), .Z(n35120) );
  ANDN U36680 ( .B(n35130), .A(n32272), .Z(n35128) );
  XNOR U36681 ( .A(\modmult_1/zin[0][762] ), .B(n35131), .Z(n32272) );
  IV U36682 ( .A(n35129), .Z(n35131) );
  XOR U36683 ( .A(n35129), .B(n32273), .Z(n35130) );
  XNOR U36684 ( .A(n35132), .B(n35133), .Z(n32273) );
  ANDN U36685 ( .B(\modmult_1/xin[1023] ), .A(n35134), .Z(n35132) );
  IV U36686 ( .A(n35133), .Z(n35134) );
  XNOR U36687 ( .A(m[763]), .B(n35135), .Z(n35133) );
  NAND U36688 ( .A(n35136), .B(mul_pow), .Z(n35135) );
  XOR U36689 ( .A(m[763]), .B(c[763]), .Z(n35136) );
  XOR U36690 ( .A(n35137), .B(n35138), .Z(n35129) );
  ANDN U36691 ( .B(n35139), .A(n32270), .Z(n35137) );
  XNOR U36692 ( .A(\modmult_1/zin[0][761] ), .B(n35140), .Z(n32270) );
  IV U36693 ( .A(n35138), .Z(n35140) );
  XOR U36694 ( .A(n35138), .B(n32271), .Z(n35139) );
  XNOR U36695 ( .A(n35141), .B(n35142), .Z(n32271) );
  ANDN U36696 ( .B(\modmult_1/xin[1023] ), .A(n35143), .Z(n35141) );
  IV U36697 ( .A(n35142), .Z(n35143) );
  XNOR U36698 ( .A(m[762]), .B(n35144), .Z(n35142) );
  NAND U36699 ( .A(n35145), .B(mul_pow), .Z(n35144) );
  XOR U36700 ( .A(m[762]), .B(c[762]), .Z(n35145) );
  XOR U36701 ( .A(n35146), .B(n35147), .Z(n35138) );
  ANDN U36702 ( .B(n35148), .A(n32268), .Z(n35146) );
  XNOR U36703 ( .A(\modmult_1/zin[0][760] ), .B(n35149), .Z(n32268) );
  IV U36704 ( .A(n35147), .Z(n35149) );
  XOR U36705 ( .A(n35147), .B(n32269), .Z(n35148) );
  XNOR U36706 ( .A(n35150), .B(n35151), .Z(n32269) );
  ANDN U36707 ( .B(\modmult_1/xin[1023] ), .A(n35152), .Z(n35150) );
  IV U36708 ( .A(n35151), .Z(n35152) );
  XNOR U36709 ( .A(m[761]), .B(n35153), .Z(n35151) );
  NAND U36710 ( .A(n35154), .B(mul_pow), .Z(n35153) );
  XOR U36711 ( .A(m[761]), .B(c[761]), .Z(n35154) );
  XOR U36712 ( .A(n35155), .B(n35156), .Z(n35147) );
  ANDN U36713 ( .B(n35157), .A(n32266), .Z(n35155) );
  XNOR U36714 ( .A(\modmult_1/zin[0][759] ), .B(n35158), .Z(n32266) );
  IV U36715 ( .A(n35156), .Z(n35158) );
  XOR U36716 ( .A(n35156), .B(n32267), .Z(n35157) );
  XNOR U36717 ( .A(n35159), .B(n35160), .Z(n32267) );
  ANDN U36718 ( .B(\modmult_1/xin[1023] ), .A(n35161), .Z(n35159) );
  IV U36719 ( .A(n35160), .Z(n35161) );
  XNOR U36720 ( .A(m[760]), .B(n35162), .Z(n35160) );
  NAND U36721 ( .A(n35163), .B(mul_pow), .Z(n35162) );
  XOR U36722 ( .A(m[760]), .B(c[760]), .Z(n35163) );
  XOR U36723 ( .A(n35164), .B(n35165), .Z(n35156) );
  ANDN U36724 ( .B(n35166), .A(n32264), .Z(n35164) );
  XNOR U36725 ( .A(\modmult_1/zin[0][758] ), .B(n35167), .Z(n32264) );
  IV U36726 ( .A(n35165), .Z(n35167) );
  XOR U36727 ( .A(n35165), .B(n32265), .Z(n35166) );
  XNOR U36728 ( .A(n35168), .B(n35169), .Z(n32265) );
  ANDN U36729 ( .B(\modmult_1/xin[1023] ), .A(n35170), .Z(n35168) );
  IV U36730 ( .A(n35169), .Z(n35170) );
  XNOR U36731 ( .A(m[759]), .B(n35171), .Z(n35169) );
  NAND U36732 ( .A(n35172), .B(mul_pow), .Z(n35171) );
  XOR U36733 ( .A(m[759]), .B(c[759]), .Z(n35172) );
  XOR U36734 ( .A(n35173), .B(n35174), .Z(n35165) );
  ANDN U36735 ( .B(n35175), .A(n32262), .Z(n35173) );
  XNOR U36736 ( .A(\modmult_1/zin[0][757] ), .B(n35176), .Z(n32262) );
  IV U36737 ( .A(n35174), .Z(n35176) );
  XOR U36738 ( .A(n35174), .B(n32263), .Z(n35175) );
  XNOR U36739 ( .A(n35177), .B(n35178), .Z(n32263) );
  ANDN U36740 ( .B(\modmult_1/xin[1023] ), .A(n35179), .Z(n35177) );
  IV U36741 ( .A(n35178), .Z(n35179) );
  XNOR U36742 ( .A(m[758]), .B(n35180), .Z(n35178) );
  NAND U36743 ( .A(n35181), .B(mul_pow), .Z(n35180) );
  XOR U36744 ( .A(m[758]), .B(c[758]), .Z(n35181) );
  XOR U36745 ( .A(n35182), .B(n35183), .Z(n35174) );
  ANDN U36746 ( .B(n35184), .A(n32260), .Z(n35182) );
  XNOR U36747 ( .A(\modmult_1/zin[0][756] ), .B(n35185), .Z(n32260) );
  IV U36748 ( .A(n35183), .Z(n35185) );
  XOR U36749 ( .A(n35183), .B(n32261), .Z(n35184) );
  XNOR U36750 ( .A(n35186), .B(n35187), .Z(n32261) );
  ANDN U36751 ( .B(\modmult_1/xin[1023] ), .A(n35188), .Z(n35186) );
  IV U36752 ( .A(n35187), .Z(n35188) );
  XNOR U36753 ( .A(m[757]), .B(n35189), .Z(n35187) );
  NAND U36754 ( .A(n35190), .B(mul_pow), .Z(n35189) );
  XOR U36755 ( .A(m[757]), .B(c[757]), .Z(n35190) );
  XOR U36756 ( .A(n35191), .B(n35192), .Z(n35183) );
  ANDN U36757 ( .B(n35193), .A(n32258), .Z(n35191) );
  XNOR U36758 ( .A(\modmult_1/zin[0][755] ), .B(n35194), .Z(n32258) );
  IV U36759 ( .A(n35192), .Z(n35194) );
  XOR U36760 ( .A(n35192), .B(n32259), .Z(n35193) );
  XNOR U36761 ( .A(n35195), .B(n35196), .Z(n32259) );
  ANDN U36762 ( .B(\modmult_1/xin[1023] ), .A(n35197), .Z(n35195) );
  IV U36763 ( .A(n35196), .Z(n35197) );
  XNOR U36764 ( .A(m[756]), .B(n35198), .Z(n35196) );
  NAND U36765 ( .A(n35199), .B(mul_pow), .Z(n35198) );
  XOR U36766 ( .A(m[756]), .B(c[756]), .Z(n35199) );
  XOR U36767 ( .A(n35200), .B(n35201), .Z(n35192) );
  ANDN U36768 ( .B(n35202), .A(n32256), .Z(n35200) );
  XNOR U36769 ( .A(\modmult_1/zin[0][754] ), .B(n35203), .Z(n32256) );
  IV U36770 ( .A(n35201), .Z(n35203) );
  XOR U36771 ( .A(n35201), .B(n32257), .Z(n35202) );
  XNOR U36772 ( .A(n35204), .B(n35205), .Z(n32257) );
  ANDN U36773 ( .B(\modmult_1/xin[1023] ), .A(n35206), .Z(n35204) );
  IV U36774 ( .A(n35205), .Z(n35206) );
  XNOR U36775 ( .A(m[755]), .B(n35207), .Z(n35205) );
  NAND U36776 ( .A(n35208), .B(mul_pow), .Z(n35207) );
  XOR U36777 ( .A(m[755]), .B(c[755]), .Z(n35208) );
  XOR U36778 ( .A(n35209), .B(n35210), .Z(n35201) );
  ANDN U36779 ( .B(n35211), .A(n32254), .Z(n35209) );
  XNOR U36780 ( .A(\modmult_1/zin[0][753] ), .B(n35212), .Z(n32254) );
  IV U36781 ( .A(n35210), .Z(n35212) );
  XOR U36782 ( .A(n35210), .B(n32255), .Z(n35211) );
  XNOR U36783 ( .A(n35213), .B(n35214), .Z(n32255) );
  ANDN U36784 ( .B(\modmult_1/xin[1023] ), .A(n35215), .Z(n35213) );
  IV U36785 ( .A(n35214), .Z(n35215) );
  XNOR U36786 ( .A(m[754]), .B(n35216), .Z(n35214) );
  NAND U36787 ( .A(n35217), .B(mul_pow), .Z(n35216) );
  XOR U36788 ( .A(m[754]), .B(c[754]), .Z(n35217) );
  XOR U36789 ( .A(n35218), .B(n35219), .Z(n35210) );
  ANDN U36790 ( .B(n35220), .A(n32252), .Z(n35218) );
  XNOR U36791 ( .A(\modmult_1/zin[0][752] ), .B(n35221), .Z(n32252) );
  IV U36792 ( .A(n35219), .Z(n35221) );
  XOR U36793 ( .A(n35219), .B(n32253), .Z(n35220) );
  XNOR U36794 ( .A(n35222), .B(n35223), .Z(n32253) );
  ANDN U36795 ( .B(\modmult_1/xin[1023] ), .A(n35224), .Z(n35222) );
  IV U36796 ( .A(n35223), .Z(n35224) );
  XNOR U36797 ( .A(m[753]), .B(n35225), .Z(n35223) );
  NAND U36798 ( .A(n35226), .B(mul_pow), .Z(n35225) );
  XOR U36799 ( .A(m[753]), .B(c[753]), .Z(n35226) );
  XOR U36800 ( .A(n35227), .B(n35228), .Z(n35219) );
  ANDN U36801 ( .B(n35229), .A(n32250), .Z(n35227) );
  XNOR U36802 ( .A(\modmult_1/zin[0][751] ), .B(n35230), .Z(n32250) );
  IV U36803 ( .A(n35228), .Z(n35230) );
  XOR U36804 ( .A(n35228), .B(n32251), .Z(n35229) );
  XNOR U36805 ( .A(n35231), .B(n35232), .Z(n32251) );
  ANDN U36806 ( .B(\modmult_1/xin[1023] ), .A(n35233), .Z(n35231) );
  IV U36807 ( .A(n35232), .Z(n35233) );
  XNOR U36808 ( .A(m[752]), .B(n35234), .Z(n35232) );
  NAND U36809 ( .A(n35235), .B(mul_pow), .Z(n35234) );
  XOR U36810 ( .A(m[752]), .B(c[752]), .Z(n35235) );
  XOR U36811 ( .A(n35236), .B(n35237), .Z(n35228) );
  ANDN U36812 ( .B(n35238), .A(n32248), .Z(n35236) );
  XNOR U36813 ( .A(\modmult_1/zin[0][750] ), .B(n35239), .Z(n32248) );
  IV U36814 ( .A(n35237), .Z(n35239) );
  XOR U36815 ( .A(n35237), .B(n32249), .Z(n35238) );
  XNOR U36816 ( .A(n35240), .B(n35241), .Z(n32249) );
  ANDN U36817 ( .B(\modmult_1/xin[1023] ), .A(n35242), .Z(n35240) );
  IV U36818 ( .A(n35241), .Z(n35242) );
  XNOR U36819 ( .A(m[751]), .B(n35243), .Z(n35241) );
  NAND U36820 ( .A(n35244), .B(mul_pow), .Z(n35243) );
  XOR U36821 ( .A(m[751]), .B(c[751]), .Z(n35244) );
  XOR U36822 ( .A(n35245), .B(n35246), .Z(n35237) );
  ANDN U36823 ( .B(n35247), .A(n32246), .Z(n35245) );
  XNOR U36824 ( .A(\modmult_1/zin[0][749] ), .B(n35248), .Z(n32246) );
  IV U36825 ( .A(n35246), .Z(n35248) );
  XOR U36826 ( .A(n35246), .B(n32247), .Z(n35247) );
  XNOR U36827 ( .A(n35249), .B(n35250), .Z(n32247) );
  ANDN U36828 ( .B(\modmult_1/xin[1023] ), .A(n35251), .Z(n35249) );
  IV U36829 ( .A(n35250), .Z(n35251) );
  XNOR U36830 ( .A(m[750]), .B(n35252), .Z(n35250) );
  NAND U36831 ( .A(n35253), .B(mul_pow), .Z(n35252) );
  XOR U36832 ( .A(m[750]), .B(c[750]), .Z(n35253) );
  XOR U36833 ( .A(n35254), .B(n35255), .Z(n35246) );
  ANDN U36834 ( .B(n35256), .A(n32244), .Z(n35254) );
  XNOR U36835 ( .A(\modmult_1/zin[0][748] ), .B(n35257), .Z(n32244) );
  IV U36836 ( .A(n35255), .Z(n35257) );
  XOR U36837 ( .A(n35255), .B(n32245), .Z(n35256) );
  XNOR U36838 ( .A(n35258), .B(n35259), .Z(n32245) );
  ANDN U36839 ( .B(\modmult_1/xin[1023] ), .A(n35260), .Z(n35258) );
  IV U36840 ( .A(n35259), .Z(n35260) );
  XNOR U36841 ( .A(m[749]), .B(n35261), .Z(n35259) );
  NAND U36842 ( .A(n35262), .B(mul_pow), .Z(n35261) );
  XOR U36843 ( .A(m[749]), .B(c[749]), .Z(n35262) );
  XOR U36844 ( .A(n35263), .B(n35264), .Z(n35255) );
  ANDN U36845 ( .B(n35265), .A(n32242), .Z(n35263) );
  XNOR U36846 ( .A(\modmult_1/zin[0][747] ), .B(n35266), .Z(n32242) );
  IV U36847 ( .A(n35264), .Z(n35266) );
  XOR U36848 ( .A(n35264), .B(n32243), .Z(n35265) );
  XNOR U36849 ( .A(n35267), .B(n35268), .Z(n32243) );
  ANDN U36850 ( .B(\modmult_1/xin[1023] ), .A(n35269), .Z(n35267) );
  IV U36851 ( .A(n35268), .Z(n35269) );
  XNOR U36852 ( .A(m[748]), .B(n35270), .Z(n35268) );
  NAND U36853 ( .A(n35271), .B(mul_pow), .Z(n35270) );
  XOR U36854 ( .A(m[748]), .B(c[748]), .Z(n35271) );
  XOR U36855 ( .A(n35272), .B(n35273), .Z(n35264) );
  ANDN U36856 ( .B(n35274), .A(n32240), .Z(n35272) );
  XNOR U36857 ( .A(\modmult_1/zin[0][746] ), .B(n35275), .Z(n32240) );
  IV U36858 ( .A(n35273), .Z(n35275) );
  XOR U36859 ( .A(n35273), .B(n32241), .Z(n35274) );
  XNOR U36860 ( .A(n35276), .B(n35277), .Z(n32241) );
  ANDN U36861 ( .B(\modmult_1/xin[1023] ), .A(n35278), .Z(n35276) );
  IV U36862 ( .A(n35277), .Z(n35278) );
  XNOR U36863 ( .A(m[747]), .B(n35279), .Z(n35277) );
  NAND U36864 ( .A(n35280), .B(mul_pow), .Z(n35279) );
  XOR U36865 ( .A(m[747]), .B(c[747]), .Z(n35280) );
  XOR U36866 ( .A(n35281), .B(n35282), .Z(n35273) );
  ANDN U36867 ( .B(n35283), .A(n32238), .Z(n35281) );
  XNOR U36868 ( .A(\modmult_1/zin[0][745] ), .B(n35284), .Z(n32238) );
  IV U36869 ( .A(n35282), .Z(n35284) );
  XOR U36870 ( .A(n35282), .B(n32239), .Z(n35283) );
  XNOR U36871 ( .A(n35285), .B(n35286), .Z(n32239) );
  ANDN U36872 ( .B(\modmult_1/xin[1023] ), .A(n35287), .Z(n35285) );
  IV U36873 ( .A(n35286), .Z(n35287) );
  XNOR U36874 ( .A(m[746]), .B(n35288), .Z(n35286) );
  NAND U36875 ( .A(n35289), .B(mul_pow), .Z(n35288) );
  XOR U36876 ( .A(m[746]), .B(c[746]), .Z(n35289) );
  XOR U36877 ( .A(n35290), .B(n35291), .Z(n35282) );
  ANDN U36878 ( .B(n35292), .A(n32236), .Z(n35290) );
  XNOR U36879 ( .A(\modmult_1/zin[0][744] ), .B(n35293), .Z(n32236) );
  IV U36880 ( .A(n35291), .Z(n35293) );
  XOR U36881 ( .A(n35291), .B(n32237), .Z(n35292) );
  XNOR U36882 ( .A(n35294), .B(n35295), .Z(n32237) );
  ANDN U36883 ( .B(\modmult_1/xin[1023] ), .A(n35296), .Z(n35294) );
  IV U36884 ( .A(n35295), .Z(n35296) );
  XNOR U36885 ( .A(m[745]), .B(n35297), .Z(n35295) );
  NAND U36886 ( .A(n35298), .B(mul_pow), .Z(n35297) );
  XOR U36887 ( .A(m[745]), .B(c[745]), .Z(n35298) );
  XOR U36888 ( .A(n35299), .B(n35300), .Z(n35291) );
  ANDN U36889 ( .B(n35301), .A(n32234), .Z(n35299) );
  XNOR U36890 ( .A(\modmult_1/zin[0][743] ), .B(n35302), .Z(n32234) );
  IV U36891 ( .A(n35300), .Z(n35302) );
  XOR U36892 ( .A(n35300), .B(n32235), .Z(n35301) );
  XNOR U36893 ( .A(n35303), .B(n35304), .Z(n32235) );
  ANDN U36894 ( .B(\modmult_1/xin[1023] ), .A(n35305), .Z(n35303) );
  IV U36895 ( .A(n35304), .Z(n35305) );
  XNOR U36896 ( .A(m[744]), .B(n35306), .Z(n35304) );
  NAND U36897 ( .A(n35307), .B(mul_pow), .Z(n35306) );
  XOR U36898 ( .A(m[744]), .B(c[744]), .Z(n35307) );
  XOR U36899 ( .A(n35308), .B(n35309), .Z(n35300) );
  ANDN U36900 ( .B(n35310), .A(n32232), .Z(n35308) );
  XNOR U36901 ( .A(\modmult_1/zin[0][742] ), .B(n35311), .Z(n32232) );
  IV U36902 ( .A(n35309), .Z(n35311) );
  XOR U36903 ( .A(n35309), .B(n32233), .Z(n35310) );
  XNOR U36904 ( .A(n35312), .B(n35313), .Z(n32233) );
  ANDN U36905 ( .B(\modmult_1/xin[1023] ), .A(n35314), .Z(n35312) );
  IV U36906 ( .A(n35313), .Z(n35314) );
  XNOR U36907 ( .A(m[743]), .B(n35315), .Z(n35313) );
  NAND U36908 ( .A(n35316), .B(mul_pow), .Z(n35315) );
  XOR U36909 ( .A(m[743]), .B(c[743]), .Z(n35316) );
  XOR U36910 ( .A(n35317), .B(n35318), .Z(n35309) );
  ANDN U36911 ( .B(n35319), .A(n32230), .Z(n35317) );
  XNOR U36912 ( .A(\modmult_1/zin[0][741] ), .B(n35320), .Z(n32230) );
  IV U36913 ( .A(n35318), .Z(n35320) );
  XOR U36914 ( .A(n35318), .B(n32231), .Z(n35319) );
  XNOR U36915 ( .A(n35321), .B(n35322), .Z(n32231) );
  ANDN U36916 ( .B(\modmult_1/xin[1023] ), .A(n35323), .Z(n35321) );
  IV U36917 ( .A(n35322), .Z(n35323) );
  XNOR U36918 ( .A(m[742]), .B(n35324), .Z(n35322) );
  NAND U36919 ( .A(n35325), .B(mul_pow), .Z(n35324) );
  XOR U36920 ( .A(m[742]), .B(c[742]), .Z(n35325) );
  XOR U36921 ( .A(n35326), .B(n35327), .Z(n35318) );
  ANDN U36922 ( .B(n35328), .A(n32228), .Z(n35326) );
  XNOR U36923 ( .A(\modmult_1/zin[0][740] ), .B(n35329), .Z(n32228) );
  IV U36924 ( .A(n35327), .Z(n35329) );
  XOR U36925 ( .A(n35327), .B(n32229), .Z(n35328) );
  XNOR U36926 ( .A(n35330), .B(n35331), .Z(n32229) );
  ANDN U36927 ( .B(\modmult_1/xin[1023] ), .A(n35332), .Z(n35330) );
  IV U36928 ( .A(n35331), .Z(n35332) );
  XNOR U36929 ( .A(m[741]), .B(n35333), .Z(n35331) );
  NAND U36930 ( .A(n35334), .B(mul_pow), .Z(n35333) );
  XOR U36931 ( .A(m[741]), .B(c[741]), .Z(n35334) );
  XOR U36932 ( .A(n35335), .B(n35336), .Z(n35327) );
  ANDN U36933 ( .B(n35337), .A(n32226), .Z(n35335) );
  XNOR U36934 ( .A(\modmult_1/zin[0][739] ), .B(n35338), .Z(n32226) );
  IV U36935 ( .A(n35336), .Z(n35338) );
  XOR U36936 ( .A(n35336), .B(n32227), .Z(n35337) );
  XNOR U36937 ( .A(n35339), .B(n35340), .Z(n32227) );
  ANDN U36938 ( .B(\modmult_1/xin[1023] ), .A(n35341), .Z(n35339) );
  IV U36939 ( .A(n35340), .Z(n35341) );
  XNOR U36940 ( .A(m[740]), .B(n35342), .Z(n35340) );
  NAND U36941 ( .A(n35343), .B(mul_pow), .Z(n35342) );
  XOR U36942 ( .A(m[740]), .B(c[740]), .Z(n35343) );
  XOR U36943 ( .A(n35344), .B(n35345), .Z(n35336) );
  ANDN U36944 ( .B(n35346), .A(n32224), .Z(n35344) );
  XNOR U36945 ( .A(\modmult_1/zin[0][738] ), .B(n35347), .Z(n32224) );
  IV U36946 ( .A(n35345), .Z(n35347) );
  XOR U36947 ( .A(n35345), .B(n32225), .Z(n35346) );
  XNOR U36948 ( .A(n35348), .B(n35349), .Z(n32225) );
  ANDN U36949 ( .B(\modmult_1/xin[1023] ), .A(n35350), .Z(n35348) );
  IV U36950 ( .A(n35349), .Z(n35350) );
  XNOR U36951 ( .A(m[739]), .B(n35351), .Z(n35349) );
  NAND U36952 ( .A(n35352), .B(mul_pow), .Z(n35351) );
  XOR U36953 ( .A(m[739]), .B(c[739]), .Z(n35352) );
  XOR U36954 ( .A(n35353), .B(n35354), .Z(n35345) );
  ANDN U36955 ( .B(n35355), .A(n32222), .Z(n35353) );
  XNOR U36956 ( .A(\modmult_1/zin[0][737] ), .B(n35356), .Z(n32222) );
  IV U36957 ( .A(n35354), .Z(n35356) );
  XOR U36958 ( .A(n35354), .B(n32223), .Z(n35355) );
  XNOR U36959 ( .A(n35357), .B(n35358), .Z(n32223) );
  ANDN U36960 ( .B(\modmult_1/xin[1023] ), .A(n35359), .Z(n35357) );
  IV U36961 ( .A(n35358), .Z(n35359) );
  XNOR U36962 ( .A(m[738]), .B(n35360), .Z(n35358) );
  NAND U36963 ( .A(n35361), .B(mul_pow), .Z(n35360) );
  XOR U36964 ( .A(m[738]), .B(c[738]), .Z(n35361) );
  XOR U36965 ( .A(n35362), .B(n35363), .Z(n35354) );
  ANDN U36966 ( .B(n35364), .A(n32220), .Z(n35362) );
  XNOR U36967 ( .A(\modmult_1/zin[0][736] ), .B(n35365), .Z(n32220) );
  IV U36968 ( .A(n35363), .Z(n35365) );
  XOR U36969 ( .A(n35363), .B(n32221), .Z(n35364) );
  XNOR U36970 ( .A(n35366), .B(n35367), .Z(n32221) );
  ANDN U36971 ( .B(\modmult_1/xin[1023] ), .A(n35368), .Z(n35366) );
  IV U36972 ( .A(n35367), .Z(n35368) );
  XNOR U36973 ( .A(m[737]), .B(n35369), .Z(n35367) );
  NAND U36974 ( .A(n35370), .B(mul_pow), .Z(n35369) );
  XOR U36975 ( .A(m[737]), .B(c[737]), .Z(n35370) );
  XOR U36976 ( .A(n35371), .B(n35372), .Z(n35363) );
  ANDN U36977 ( .B(n35373), .A(n32218), .Z(n35371) );
  XNOR U36978 ( .A(\modmult_1/zin[0][735] ), .B(n35374), .Z(n32218) );
  IV U36979 ( .A(n35372), .Z(n35374) );
  XOR U36980 ( .A(n35372), .B(n32219), .Z(n35373) );
  XNOR U36981 ( .A(n35375), .B(n35376), .Z(n32219) );
  ANDN U36982 ( .B(\modmult_1/xin[1023] ), .A(n35377), .Z(n35375) );
  IV U36983 ( .A(n35376), .Z(n35377) );
  XNOR U36984 ( .A(m[736]), .B(n35378), .Z(n35376) );
  NAND U36985 ( .A(n35379), .B(mul_pow), .Z(n35378) );
  XOR U36986 ( .A(m[736]), .B(c[736]), .Z(n35379) );
  XOR U36987 ( .A(n35380), .B(n35381), .Z(n35372) );
  ANDN U36988 ( .B(n35382), .A(n32216), .Z(n35380) );
  XNOR U36989 ( .A(\modmult_1/zin[0][734] ), .B(n35383), .Z(n32216) );
  IV U36990 ( .A(n35381), .Z(n35383) );
  XOR U36991 ( .A(n35381), .B(n32217), .Z(n35382) );
  XNOR U36992 ( .A(n35384), .B(n35385), .Z(n32217) );
  ANDN U36993 ( .B(\modmult_1/xin[1023] ), .A(n35386), .Z(n35384) );
  IV U36994 ( .A(n35385), .Z(n35386) );
  XNOR U36995 ( .A(m[735]), .B(n35387), .Z(n35385) );
  NAND U36996 ( .A(n35388), .B(mul_pow), .Z(n35387) );
  XOR U36997 ( .A(m[735]), .B(c[735]), .Z(n35388) );
  XOR U36998 ( .A(n35389), .B(n35390), .Z(n35381) );
  ANDN U36999 ( .B(n35391), .A(n32214), .Z(n35389) );
  XNOR U37000 ( .A(\modmult_1/zin[0][733] ), .B(n35392), .Z(n32214) );
  IV U37001 ( .A(n35390), .Z(n35392) );
  XOR U37002 ( .A(n35390), .B(n32215), .Z(n35391) );
  XNOR U37003 ( .A(n35393), .B(n35394), .Z(n32215) );
  ANDN U37004 ( .B(\modmult_1/xin[1023] ), .A(n35395), .Z(n35393) );
  IV U37005 ( .A(n35394), .Z(n35395) );
  XNOR U37006 ( .A(m[734]), .B(n35396), .Z(n35394) );
  NAND U37007 ( .A(n35397), .B(mul_pow), .Z(n35396) );
  XOR U37008 ( .A(m[734]), .B(c[734]), .Z(n35397) );
  XOR U37009 ( .A(n35398), .B(n35399), .Z(n35390) );
  ANDN U37010 ( .B(n35400), .A(n32212), .Z(n35398) );
  XNOR U37011 ( .A(\modmult_1/zin[0][732] ), .B(n35401), .Z(n32212) );
  IV U37012 ( .A(n35399), .Z(n35401) );
  XOR U37013 ( .A(n35399), .B(n32213), .Z(n35400) );
  XNOR U37014 ( .A(n35402), .B(n35403), .Z(n32213) );
  ANDN U37015 ( .B(\modmult_1/xin[1023] ), .A(n35404), .Z(n35402) );
  IV U37016 ( .A(n35403), .Z(n35404) );
  XNOR U37017 ( .A(m[733]), .B(n35405), .Z(n35403) );
  NAND U37018 ( .A(n35406), .B(mul_pow), .Z(n35405) );
  XOR U37019 ( .A(m[733]), .B(c[733]), .Z(n35406) );
  XOR U37020 ( .A(n35407), .B(n35408), .Z(n35399) );
  ANDN U37021 ( .B(n35409), .A(n32210), .Z(n35407) );
  XNOR U37022 ( .A(\modmult_1/zin[0][731] ), .B(n35410), .Z(n32210) );
  IV U37023 ( .A(n35408), .Z(n35410) );
  XOR U37024 ( .A(n35408), .B(n32211), .Z(n35409) );
  XNOR U37025 ( .A(n35411), .B(n35412), .Z(n32211) );
  ANDN U37026 ( .B(\modmult_1/xin[1023] ), .A(n35413), .Z(n35411) );
  IV U37027 ( .A(n35412), .Z(n35413) );
  XNOR U37028 ( .A(m[732]), .B(n35414), .Z(n35412) );
  NAND U37029 ( .A(n35415), .B(mul_pow), .Z(n35414) );
  XOR U37030 ( .A(m[732]), .B(c[732]), .Z(n35415) );
  XOR U37031 ( .A(n35416), .B(n35417), .Z(n35408) );
  ANDN U37032 ( .B(n35418), .A(n32208), .Z(n35416) );
  XNOR U37033 ( .A(\modmult_1/zin[0][730] ), .B(n35419), .Z(n32208) );
  IV U37034 ( .A(n35417), .Z(n35419) );
  XOR U37035 ( .A(n35417), .B(n32209), .Z(n35418) );
  XNOR U37036 ( .A(n35420), .B(n35421), .Z(n32209) );
  ANDN U37037 ( .B(\modmult_1/xin[1023] ), .A(n35422), .Z(n35420) );
  IV U37038 ( .A(n35421), .Z(n35422) );
  XNOR U37039 ( .A(m[731]), .B(n35423), .Z(n35421) );
  NAND U37040 ( .A(n35424), .B(mul_pow), .Z(n35423) );
  XOR U37041 ( .A(m[731]), .B(c[731]), .Z(n35424) );
  XOR U37042 ( .A(n35425), .B(n35426), .Z(n35417) );
  ANDN U37043 ( .B(n35427), .A(n32206), .Z(n35425) );
  XNOR U37044 ( .A(\modmult_1/zin[0][729] ), .B(n35428), .Z(n32206) );
  IV U37045 ( .A(n35426), .Z(n35428) );
  XOR U37046 ( .A(n35426), .B(n32207), .Z(n35427) );
  XNOR U37047 ( .A(n35429), .B(n35430), .Z(n32207) );
  ANDN U37048 ( .B(\modmult_1/xin[1023] ), .A(n35431), .Z(n35429) );
  IV U37049 ( .A(n35430), .Z(n35431) );
  XNOR U37050 ( .A(m[730]), .B(n35432), .Z(n35430) );
  NAND U37051 ( .A(n35433), .B(mul_pow), .Z(n35432) );
  XOR U37052 ( .A(m[730]), .B(c[730]), .Z(n35433) );
  XOR U37053 ( .A(n35434), .B(n35435), .Z(n35426) );
  ANDN U37054 ( .B(n35436), .A(n32204), .Z(n35434) );
  XNOR U37055 ( .A(\modmult_1/zin[0][728] ), .B(n35437), .Z(n32204) );
  IV U37056 ( .A(n35435), .Z(n35437) );
  XOR U37057 ( .A(n35435), .B(n32205), .Z(n35436) );
  XNOR U37058 ( .A(n35438), .B(n35439), .Z(n32205) );
  ANDN U37059 ( .B(\modmult_1/xin[1023] ), .A(n35440), .Z(n35438) );
  IV U37060 ( .A(n35439), .Z(n35440) );
  XNOR U37061 ( .A(m[729]), .B(n35441), .Z(n35439) );
  NAND U37062 ( .A(n35442), .B(mul_pow), .Z(n35441) );
  XOR U37063 ( .A(m[729]), .B(c[729]), .Z(n35442) );
  XOR U37064 ( .A(n35443), .B(n35444), .Z(n35435) );
  ANDN U37065 ( .B(n35445), .A(n32202), .Z(n35443) );
  XNOR U37066 ( .A(\modmult_1/zin[0][727] ), .B(n35446), .Z(n32202) );
  IV U37067 ( .A(n35444), .Z(n35446) );
  XOR U37068 ( .A(n35444), .B(n32203), .Z(n35445) );
  XNOR U37069 ( .A(n35447), .B(n35448), .Z(n32203) );
  ANDN U37070 ( .B(\modmult_1/xin[1023] ), .A(n35449), .Z(n35447) );
  IV U37071 ( .A(n35448), .Z(n35449) );
  XNOR U37072 ( .A(m[728]), .B(n35450), .Z(n35448) );
  NAND U37073 ( .A(n35451), .B(mul_pow), .Z(n35450) );
  XOR U37074 ( .A(m[728]), .B(c[728]), .Z(n35451) );
  XOR U37075 ( .A(n35452), .B(n35453), .Z(n35444) );
  ANDN U37076 ( .B(n35454), .A(n32200), .Z(n35452) );
  XNOR U37077 ( .A(\modmult_1/zin[0][726] ), .B(n35455), .Z(n32200) );
  IV U37078 ( .A(n35453), .Z(n35455) );
  XOR U37079 ( .A(n35453), .B(n32201), .Z(n35454) );
  XNOR U37080 ( .A(n35456), .B(n35457), .Z(n32201) );
  ANDN U37081 ( .B(\modmult_1/xin[1023] ), .A(n35458), .Z(n35456) );
  IV U37082 ( .A(n35457), .Z(n35458) );
  XNOR U37083 ( .A(m[727]), .B(n35459), .Z(n35457) );
  NAND U37084 ( .A(n35460), .B(mul_pow), .Z(n35459) );
  XOR U37085 ( .A(m[727]), .B(c[727]), .Z(n35460) );
  XOR U37086 ( .A(n35461), .B(n35462), .Z(n35453) );
  ANDN U37087 ( .B(n35463), .A(n32198), .Z(n35461) );
  XNOR U37088 ( .A(\modmult_1/zin[0][725] ), .B(n35464), .Z(n32198) );
  IV U37089 ( .A(n35462), .Z(n35464) );
  XOR U37090 ( .A(n35462), .B(n32199), .Z(n35463) );
  XNOR U37091 ( .A(n35465), .B(n35466), .Z(n32199) );
  ANDN U37092 ( .B(\modmult_1/xin[1023] ), .A(n35467), .Z(n35465) );
  IV U37093 ( .A(n35466), .Z(n35467) );
  XNOR U37094 ( .A(m[726]), .B(n35468), .Z(n35466) );
  NAND U37095 ( .A(n35469), .B(mul_pow), .Z(n35468) );
  XOR U37096 ( .A(m[726]), .B(c[726]), .Z(n35469) );
  XOR U37097 ( .A(n35470), .B(n35471), .Z(n35462) );
  ANDN U37098 ( .B(n35472), .A(n32196), .Z(n35470) );
  XNOR U37099 ( .A(\modmult_1/zin[0][724] ), .B(n35473), .Z(n32196) );
  IV U37100 ( .A(n35471), .Z(n35473) );
  XOR U37101 ( .A(n35471), .B(n32197), .Z(n35472) );
  XNOR U37102 ( .A(n35474), .B(n35475), .Z(n32197) );
  ANDN U37103 ( .B(\modmult_1/xin[1023] ), .A(n35476), .Z(n35474) );
  IV U37104 ( .A(n35475), .Z(n35476) );
  XNOR U37105 ( .A(m[725]), .B(n35477), .Z(n35475) );
  NAND U37106 ( .A(n35478), .B(mul_pow), .Z(n35477) );
  XOR U37107 ( .A(m[725]), .B(c[725]), .Z(n35478) );
  XOR U37108 ( .A(n35479), .B(n35480), .Z(n35471) );
  ANDN U37109 ( .B(n35481), .A(n32194), .Z(n35479) );
  XNOR U37110 ( .A(\modmult_1/zin[0][723] ), .B(n35482), .Z(n32194) );
  IV U37111 ( .A(n35480), .Z(n35482) );
  XOR U37112 ( .A(n35480), .B(n32195), .Z(n35481) );
  XNOR U37113 ( .A(n35483), .B(n35484), .Z(n32195) );
  ANDN U37114 ( .B(\modmult_1/xin[1023] ), .A(n35485), .Z(n35483) );
  IV U37115 ( .A(n35484), .Z(n35485) );
  XNOR U37116 ( .A(m[724]), .B(n35486), .Z(n35484) );
  NAND U37117 ( .A(n35487), .B(mul_pow), .Z(n35486) );
  XOR U37118 ( .A(m[724]), .B(c[724]), .Z(n35487) );
  XOR U37119 ( .A(n35488), .B(n35489), .Z(n35480) );
  ANDN U37120 ( .B(n35490), .A(n32192), .Z(n35488) );
  XNOR U37121 ( .A(\modmult_1/zin[0][722] ), .B(n35491), .Z(n32192) );
  IV U37122 ( .A(n35489), .Z(n35491) );
  XOR U37123 ( .A(n35489), .B(n32193), .Z(n35490) );
  XNOR U37124 ( .A(n35492), .B(n35493), .Z(n32193) );
  ANDN U37125 ( .B(\modmult_1/xin[1023] ), .A(n35494), .Z(n35492) );
  IV U37126 ( .A(n35493), .Z(n35494) );
  XNOR U37127 ( .A(m[723]), .B(n35495), .Z(n35493) );
  NAND U37128 ( .A(n35496), .B(mul_pow), .Z(n35495) );
  XOR U37129 ( .A(m[723]), .B(c[723]), .Z(n35496) );
  XOR U37130 ( .A(n35497), .B(n35498), .Z(n35489) );
  ANDN U37131 ( .B(n35499), .A(n32190), .Z(n35497) );
  XNOR U37132 ( .A(\modmult_1/zin[0][721] ), .B(n35500), .Z(n32190) );
  IV U37133 ( .A(n35498), .Z(n35500) );
  XOR U37134 ( .A(n35498), .B(n32191), .Z(n35499) );
  XNOR U37135 ( .A(n35501), .B(n35502), .Z(n32191) );
  ANDN U37136 ( .B(\modmult_1/xin[1023] ), .A(n35503), .Z(n35501) );
  IV U37137 ( .A(n35502), .Z(n35503) );
  XNOR U37138 ( .A(m[722]), .B(n35504), .Z(n35502) );
  NAND U37139 ( .A(n35505), .B(mul_pow), .Z(n35504) );
  XOR U37140 ( .A(m[722]), .B(c[722]), .Z(n35505) );
  XOR U37141 ( .A(n35506), .B(n35507), .Z(n35498) );
  ANDN U37142 ( .B(n35508), .A(n32188), .Z(n35506) );
  XNOR U37143 ( .A(\modmult_1/zin[0][720] ), .B(n35509), .Z(n32188) );
  IV U37144 ( .A(n35507), .Z(n35509) );
  XOR U37145 ( .A(n35507), .B(n32189), .Z(n35508) );
  XNOR U37146 ( .A(n35510), .B(n35511), .Z(n32189) );
  ANDN U37147 ( .B(\modmult_1/xin[1023] ), .A(n35512), .Z(n35510) );
  IV U37148 ( .A(n35511), .Z(n35512) );
  XNOR U37149 ( .A(m[721]), .B(n35513), .Z(n35511) );
  NAND U37150 ( .A(n35514), .B(mul_pow), .Z(n35513) );
  XOR U37151 ( .A(m[721]), .B(c[721]), .Z(n35514) );
  XOR U37152 ( .A(n35515), .B(n35516), .Z(n35507) );
  ANDN U37153 ( .B(n35517), .A(n32186), .Z(n35515) );
  XNOR U37154 ( .A(\modmult_1/zin[0][719] ), .B(n35518), .Z(n32186) );
  IV U37155 ( .A(n35516), .Z(n35518) );
  XOR U37156 ( .A(n35516), .B(n32187), .Z(n35517) );
  XNOR U37157 ( .A(n35519), .B(n35520), .Z(n32187) );
  ANDN U37158 ( .B(\modmult_1/xin[1023] ), .A(n35521), .Z(n35519) );
  IV U37159 ( .A(n35520), .Z(n35521) );
  XNOR U37160 ( .A(m[720]), .B(n35522), .Z(n35520) );
  NAND U37161 ( .A(n35523), .B(mul_pow), .Z(n35522) );
  XOR U37162 ( .A(m[720]), .B(c[720]), .Z(n35523) );
  XOR U37163 ( .A(n35524), .B(n35525), .Z(n35516) );
  ANDN U37164 ( .B(n35526), .A(n32184), .Z(n35524) );
  XNOR U37165 ( .A(\modmult_1/zin[0][718] ), .B(n35527), .Z(n32184) );
  IV U37166 ( .A(n35525), .Z(n35527) );
  XOR U37167 ( .A(n35525), .B(n32185), .Z(n35526) );
  XNOR U37168 ( .A(n35528), .B(n35529), .Z(n32185) );
  ANDN U37169 ( .B(\modmult_1/xin[1023] ), .A(n35530), .Z(n35528) );
  IV U37170 ( .A(n35529), .Z(n35530) );
  XNOR U37171 ( .A(m[719]), .B(n35531), .Z(n35529) );
  NAND U37172 ( .A(n35532), .B(mul_pow), .Z(n35531) );
  XOR U37173 ( .A(m[719]), .B(c[719]), .Z(n35532) );
  XOR U37174 ( .A(n35533), .B(n35534), .Z(n35525) );
  ANDN U37175 ( .B(n35535), .A(n32182), .Z(n35533) );
  XNOR U37176 ( .A(\modmult_1/zin[0][717] ), .B(n35536), .Z(n32182) );
  IV U37177 ( .A(n35534), .Z(n35536) );
  XOR U37178 ( .A(n35534), .B(n32183), .Z(n35535) );
  XNOR U37179 ( .A(n35537), .B(n35538), .Z(n32183) );
  ANDN U37180 ( .B(\modmult_1/xin[1023] ), .A(n35539), .Z(n35537) );
  IV U37181 ( .A(n35538), .Z(n35539) );
  XNOR U37182 ( .A(m[718]), .B(n35540), .Z(n35538) );
  NAND U37183 ( .A(n35541), .B(mul_pow), .Z(n35540) );
  XOR U37184 ( .A(m[718]), .B(c[718]), .Z(n35541) );
  XOR U37185 ( .A(n35542), .B(n35543), .Z(n35534) );
  ANDN U37186 ( .B(n35544), .A(n32180), .Z(n35542) );
  XNOR U37187 ( .A(\modmult_1/zin[0][716] ), .B(n35545), .Z(n32180) );
  IV U37188 ( .A(n35543), .Z(n35545) );
  XOR U37189 ( .A(n35543), .B(n32181), .Z(n35544) );
  XNOR U37190 ( .A(n35546), .B(n35547), .Z(n32181) );
  ANDN U37191 ( .B(\modmult_1/xin[1023] ), .A(n35548), .Z(n35546) );
  IV U37192 ( .A(n35547), .Z(n35548) );
  XNOR U37193 ( .A(m[717]), .B(n35549), .Z(n35547) );
  NAND U37194 ( .A(n35550), .B(mul_pow), .Z(n35549) );
  XOR U37195 ( .A(m[717]), .B(c[717]), .Z(n35550) );
  XOR U37196 ( .A(n35551), .B(n35552), .Z(n35543) );
  ANDN U37197 ( .B(n35553), .A(n32178), .Z(n35551) );
  XNOR U37198 ( .A(\modmult_1/zin[0][715] ), .B(n35554), .Z(n32178) );
  IV U37199 ( .A(n35552), .Z(n35554) );
  XOR U37200 ( .A(n35552), .B(n32179), .Z(n35553) );
  XNOR U37201 ( .A(n35555), .B(n35556), .Z(n32179) );
  ANDN U37202 ( .B(\modmult_1/xin[1023] ), .A(n35557), .Z(n35555) );
  IV U37203 ( .A(n35556), .Z(n35557) );
  XNOR U37204 ( .A(m[716]), .B(n35558), .Z(n35556) );
  NAND U37205 ( .A(n35559), .B(mul_pow), .Z(n35558) );
  XOR U37206 ( .A(m[716]), .B(c[716]), .Z(n35559) );
  XOR U37207 ( .A(n35560), .B(n35561), .Z(n35552) );
  ANDN U37208 ( .B(n35562), .A(n32176), .Z(n35560) );
  XNOR U37209 ( .A(\modmult_1/zin[0][714] ), .B(n35563), .Z(n32176) );
  IV U37210 ( .A(n35561), .Z(n35563) );
  XOR U37211 ( .A(n35561), .B(n32177), .Z(n35562) );
  XNOR U37212 ( .A(n35564), .B(n35565), .Z(n32177) );
  ANDN U37213 ( .B(\modmult_1/xin[1023] ), .A(n35566), .Z(n35564) );
  IV U37214 ( .A(n35565), .Z(n35566) );
  XNOR U37215 ( .A(m[715]), .B(n35567), .Z(n35565) );
  NAND U37216 ( .A(n35568), .B(mul_pow), .Z(n35567) );
  XOR U37217 ( .A(m[715]), .B(c[715]), .Z(n35568) );
  XOR U37218 ( .A(n35569), .B(n35570), .Z(n35561) );
  ANDN U37219 ( .B(n35571), .A(n32174), .Z(n35569) );
  XNOR U37220 ( .A(\modmult_1/zin[0][713] ), .B(n35572), .Z(n32174) );
  IV U37221 ( .A(n35570), .Z(n35572) );
  XOR U37222 ( .A(n35570), .B(n32175), .Z(n35571) );
  XNOR U37223 ( .A(n35573), .B(n35574), .Z(n32175) );
  ANDN U37224 ( .B(\modmult_1/xin[1023] ), .A(n35575), .Z(n35573) );
  IV U37225 ( .A(n35574), .Z(n35575) );
  XNOR U37226 ( .A(m[714]), .B(n35576), .Z(n35574) );
  NAND U37227 ( .A(n35577), .B(mul_pow), .Z(n35576) );
  XOR U37228 ( .A(m[714]), .B(c[714]), .Z(n35577) );
  XOR U37229 ( .A(n35578), .B(n35579), .Z(n35570) );
  ANDN U37230 ( .B(n35580), .A(n32172), .Z(n35578) );
  XNOR U37231 ( .A(\modmult_1/zin[0][712] ), .B(n35581), .Z(n32172) );
  IV U37232 ( .A(n35579), .Z(n35581) );
  XOR U37233 ( .A(n35579), .B(n32173), .Z(n35580) );
  XNOR U37234 ( .A(n35582), .B(n35583), .Z(n32173) );
  ANDN U37235 ( .B(\modmult_1/xin[1023] ), .A(n35584), .Z(n35582) );
  IV U37236 ( .A(n35583), .Z(n35584) );
  XNOR U37237 ( .A(m[713]), .B(n35585), .Z(n35583) );
  NAND U37238 ( .A(n35586), .B(mul_pow), .Z(n35585) );
  XOR U37239 ( .A(m[713]), .B(c[713]), .Z(n35586) );
  XOR U37240 ( .A(n35587), .B(n35588), .Z(n35579) );
  ANDN U37241 ( .B(n35589), .A(n32170), .Z(n35587) );
  XNOR U37242 ( .A(\modmult_1/zin[0][711] ), .B(n35590), .Z(n32170) );
  IV U37243 ( .A(n35588), .Z(n35590) );
  XOR U37244 ( .A(n35588), .B(n32171), .Z(n35589) );
  XNOR U37245 ( .A(n35591), .B(n35592), .Z(n32171) );
  ANDN U37246 ( .B(\modmult_1/xin[1023] ), .A(n35593), .Z(n35591) );
  IV U37247 ( .A(n35592), .Z(n35593) );
  XNOR U37248 ( .A(m[712]), .B(n35594), .Z(n35592) );
  NAND U37249 ( .A(n35595), .B(mul_pow), .Z(n35594) );
  XOR U37250 ( .A(m[712]), .B(c[712]), .Z(n35595) );
  XOR U37251 ( .A(n35596), .B(n35597), .Z(n35588) );
  ANDN U37252 ( .B(n35598), .A(n32168), .Z(n35596) );
  XNOR U37253 ( .A(\modmult_1/zin[0][710] ), .B(n35599), .Z(n32168) );
  IV U37254 ( .A(n35597), .Z(n35599) );
  XOR U37255 ( .A(n35597), .B(n32169), .Z(n35598) );
  XNOR U37256 ( .A(n35600), .B(n35601), .Z(n32169) );
  ANDN U37257 ( .B(\modmult_1/xin[1023] ), .A(n35602), .Z(n35600) );
  IV U37258 ( .A(n35601), .Z(n35602) );
  XNOR U37259 ( .A(m[711]), .B(n35603), .Z(n35601) );
  NAND U37260 ( .A(n35604), .B(mul_pow), .Z(n35603) );
  XOR U37261 ( .A(m[711]), .B(c[711]), .Z(n35604) );
  XOR U37262 ( .A(n35605), .B(n35606), .Z(n35597) );
  ANDN U37263 ( .B(n35607), .A(n32166), .Z(n35605) );
  XNOR U37264 ( .A(\modmult_1/zin[0][709] ), .B(n35608), .Z(n32166) );
  IV U37265 ( .A(n35606), .Z(n35608) );
  XOR U37266 ( .A(n35606), .B(n32167), .Z(n35607) );
  XNOR U37267 ( .A(n35609), .B(n35610), .Z(n32167) );
  ANDN U37268 ( .B(\modmult_1/xin[1023] ), .A(n35611), .Z(n35609) );
  IV U37269 ( .A(n35610), .Z(n35611) );
  XNOR U37270 ( .A(m[710]), .B(n35612), .Z(n35610) );
  NAND U37271 ( .A(n35613), .B(mul_pow), .Z(n35612) );
  XOR U37272 ( .A(m[710]), .B(c[710]), .Z(n35613) );
  XOR U37273 ( .A(n35614), .B(n35615), .Z(n35606) );
  ANDN U37274 ( .B(n35616), .A(n32164), .Z(n35614) );
  XNOR U37275 ( .A(\modmult_1/zin[0][708] ), .B(n35617), .Z(n32164) );
  IV U37276 ( .A(n35615), .Z(n35617) );
  XOR U37277 ( .A(n35615), .B(n32165), .Z(n35616) );
  XNOR U37278 ( .A(n35618), .B(n35619), .Z(n32165) );
  ANDN U37279 ( .B(\modmult_1/xin[1023] ), .A(n35620), .Z(n35618) );
  IV U37280 ( .A(n35619), .Z(n35620) );
  XNOR U37281 ( .A(m[709]), .B(n35621), .Z(n35619) );
  NAND U37282 ( .A(n35622), .B(mul_pow), .Z(n35621) );
  XOR U37283 ( .A(m[709]), .B(c[709]), .Z(n35622) );
  XOR U37284 ( .A(n35623), .B(n35624), .Z(n35615) );
  ANDN U37285 ( .B(n35625), .A(n32162), .Z(n35623) );
  XNOR U37286 ( .A(\modmult_1/zin[0][707] ), .B(n35626), .Z(n32162) );
  IV U37287 ( .A(n35624), .Z(n35626) );
  XOR U37288 ( .A(n35624), .B(n32163), .Z(n35625) );
  XNOR U37289 ( .A(n35627), .B(n35628), .Z(n32163) );
  ANDN U37290 ( .B(\modmult_1/xin[1023] ), .A(n35629), .Z(n35627) );
  IV U37291 ( .A(n35628), .Z(n35629) );
  XNOR U37292 ( .A(m[708]), .B(n35630), .Z(n35628) );
  NAND U37293 ( .A(n35631), .B(mul_pow), .Z(n35630) );
  XOR U37294 ( .A(m[708]), .B(c[708]), .Z(n35631) );
  XOR U37295 ( .A(n35632), .B(n35633), .Z(n35624) );
  ANDN U37296 ( .B(n35634), .A(n32160), .Z(n35632) );
  XNOR U37297 ( .A(\modmult_1/zin[0][706] ), .B(n35635), .Z(n32160) );
  IV U37298 ( .A(n35633), .Z(n35635) );
  XOR U37299 ( .A(n35633), .B(n32161), .Z(n35634) );
  XNOR U37300 ( .A(n35636), .B(n35637), .Z(n32161) );
  ANDN U37301 ( .B(\modmult_1/xin[1023] ), .A(n35638), .Z(n35636) );
  IV U37302 ( .A(n35637), .Z(n35638) );
  XNOR U37303 ( .A(m[707]), .B(n35639), .Z(n35637) );
  NAND U37304 ( .A(n35640), .B(mul_pow), .Z(n35639) );
  XOR U37305 ( .A(m[707]), .B(c[707]), .Z(n35640) );
  XOR U37306 ( .A(n35641), .B(n35642), .Z(n35633) );
  ANDN U37307 ( .B(n35643), .A(n32158), .Z(n35641) );
  XNOR U37308 ( .A(\modmult_1/zin[0][705] ), .B(n35644), .Z(n32158) );
  IV U37309 ( .A(n35642), .Z(n35644) );
  XOR U37310 ( .A(n35642), .B(n32159), .Z(n35643) );
  XNOR U37311 ( .A(n35645), .B(n35646), .Z(n32159) );
  ANDN U37312 ( .B(\modmult_1/xin[1023] ), .A(n35647), .Z(n35645) );
  IV U37313 ( .A(n35646), .Z(n35647) );
  XNOR U37314 ( .A(m[706]), .B(n35648), .Z(n35646) );
  NAND U37315 ( .A(n35649), .B(mul_pow), .Z(n35648) );
  XOR U37316 ( .A(m[706]), .B(c[706]), .Z(n35649) );
  XOR U37317 ( .A(n35650), .B(n35651), .Z(n35642) );
  ANDN U37318 ( .B(n35652), .A(n32156), .Z(n35650) );
  XNOR U37319 ( .A(\modmult_1/zin[0][704] ), .B(n35653), .Z(n32156) );
  IV U37320 ( .A(n35651), .Z(n35653) );
  XOR U37321 ( .A(n35651), .B(n32157), .Z(n35652) );
  XNOR U37322 ( .A(n35654), .B(n35655), .Z(n32157) );
  ANDN U37323 ( .B(\modmult_1/xin[1023] ), .A(n35656), .Z(n35654) );
  IV U37324 ( .A(n35655), .Z(n35656) );
  XNOR U37325 ( .A(m[705]), .B(n35657), .Z(n35655) );
  NAND U37326 ( .A(n35658), .B(mul_pow), .Z(n35657) );
  XOR U37327 ( .A(m[705]), .B(c[705]), .Z(n35658) );
  XOR U37328 ( .A(n35659), .B(n35660), .Z(n35651) );
  ANDN U37329 ( .B(n35661), .A(n32154), .Z(n35659) );
  XNOR U37330 ( .A(\modmult_1/zin[0][703] ), .B(n35662), .Z(n32154) );
  IV U37331 ( .A(n35660), .Z(n35662) );
  XOR U37332 ( .A(n35660), .B(n32155), .Z(n35661) );
  XNOR U37333 ( .A(n35663), .B(n35664), .Z(n32155) );
  ANDN U37334 ( .B(\modmult_1/xin[1023] ), .A(n35665), .Z(n35663) );
  IV U37335 ( .A(n35664), .Z(n35665) );
  XNOR U37336 ( .A(m[704]), .B(n35666), .Z(n35664) );
  NAND U37337 ( .A(n35667), .B(mul_pow), .Z(n35666) );
  XOR U37338 ( .A(m[704]), .B(c[704]), .Z(n35667) );
  XOR U37339 ( .A(n35668), .B(n35669), .Z(n35660) );
  ANDN U37340 ( .B(n35670), .A(n32152), .Z(n35668) );
  XNOR U37341 ( .A(\modmult_1/zin[0][702] ), .B(n35671), .Z(n32152) );
  IV U37342 ( .A(n35669), .Z(n35671) );
  XOR U37343 ( .A(n35669), .B(n32153), .Z(n35670) );
  XNOR U37344 ( .A(n35672), .B(n35673), .Z(n32153) );
  ANDN U37345 ( .B(\modmult_1/xin[1023] ), .A(n35674), .Z(n35672) );
  IV U37346 ( .A(n35673), .Z(n35674) );
  XNOR U37347 ( .A(m[703]), .B(n35675), .Z(n35673) );
  NAND U37348 ( .A(n35676), .B(mul_pow), .Z(n35675) );
  XOR U37349 ( .A(m[703]), .B(c[703]), .Z(n35676) );
  XOR U37350 ( .A(n35677), .B(n35678), .Z(n35669) );
  ANDN U37351 ( .B(n35679), .A(n32150), .Z(n35677) );
  XNOR U37352 ( .A(\modmult_1/zin[0][701] ), .B(n35680), .Z(n32150) );
  IV U37353 ( .A(n35678), .Z(n35680) );
  XOR U37354 ( .A(n35678), .B(n32151), .Z(n35679) );
  XNOR U37355 ( .A(n35681), .B(n35682), .Z(n32151) );
  ANDN U37356 ( .B(\modmult_1/xin[1023] ), .A(n35683), .Z(n35681) );
  IV U37357 ( .A(n35682), .Z(n35683) );
  XNOR U37358 ( .A(m[702]), .B(n35684), .Z(n35682) );
  NAND U37359 ( .A(n35685), .B(mul_pow), .Z(n35684) );
  XOR U37360 ( .A(m[702]), .B(c[702]), .Z(n35685) );
  XOR U37361 ( .A(n35686), .B(n35687), .Z(n35678) );
  ANDN U37362 ( .B(n35688), .A(n32148), .Z(n35686) );
  XNOR U37363 ( .A(\modmult_1/zin[0][700] ), .B(n35689), .Z(n32148) );
  IV U37364 ( .A(n35687), .Z(n35689) );
  XOR U37365 ( .A(n35687), .B(n32149), .Z(n35688) );
  XNOR U37366 ( .A(n35690), .B(n35691), .Z(n32149) );
  ANDN U37367 ( .B(\modmult_1/xin[1023] ), .A(n35692), .Z(n35690) );
  IV U37368 ( .A(n35691), .Z(n35692) );
  XNOR U37369 ( .A(m[701]), .B(n35693), .Z(n35691) );
  NAND U37370 ( .A(n35694), .B(mul_pow), .Z(n35693) );
  XOR U37371 ( .A(m[701]), .B(c[701]), .Z(n35694) );
  XOR U37372 ( .A(n35695), .B(n35696), .Z(n35687) );
  ANDN U37373 ( .B(n35697), .A(n32146), .Z(n35695) );
  XNOR U37374 ( .A(\modmult_1/zin[0][699] ), .B(n35698), .Z(n32146) );
  IV U37375 ( .A(n35696), .Z(n35698) );
  XOR U37376 ( .A(n35696), .B(n32147), .Z(n35697) );
  XNOR U37377 ( .A(n35699), .B(n35700), .Z(n32147) );
  ANDN U37378 ( .B(\modmult_1/xin[1023] ), .A(n35701), .Z(n35699) );
  IV U37379 ( .A(n35700), .Z(n35701) );
  XNOR U37380 ( .A(m[700]), .B(n35702), .Z(n35700) );
  NAND U37381 ( .A(n35703), .B(mul_pow), .Z(n35702) );
  XOR U37382 ( .A(m[700]), .B(c[700]), .Z(n35703) );
  XOR U37383 ( .A(n35704), .B(n35705), .Z(n35696) );
  ANDN U37384 ( .B(n35706), .A(n32144), .Z(n35704) );
  XNOR U37385 ( .A(\modmult_1/zin[0][698] ), .B(n35707), .Z(n32144) );
  IV U37386 ( .A(n35705), .Z(n35707) );
  XOR U37387 ( .A(n35705), .B(n32145), .Z(n35706) );
  XNOR U37388 ( .A(n35708), .B(n35709), .Z(n32145) );
  ANDN U37389 ( .B(\modmult_1/xin[1023] ), .A(n35710), .Z(n35708) );
  IV U37390 ( .A(n35709), .Z(n35710) );
  XNOR U37391 ( .A(m[699]), .B(n35711), .Z(n35709) );
  NAND U37392 ( .A(n35712), .B(mul_pow), .Z(n35711) );
  XOR U37393 ( .A(m[699]), .B(c[699]), .Z(n35712) );
  XOR U37394 ( .A(n35713), .B(n35714), .Z(n35705) );
  ANDN U37395 ( .B(n35715), .A(n32142), .Z(n35713) );
  XNOR U37396 ( .A(\modmult_1/zin[0][697] ), .B(n35716), .Z(n32142) );
  IV U37397 ( .A(n35714), .Z(n35716) );
  XOR U37398 ( .A(n35714), .B(n32143), .Z(n35715) );
  XNOR U37399 ( .A(n35717), .B(n35718), .Z(n32143) );
  ANDN U37400 ( .B(\modmult_1/xin[1023] ), .A(n35719), .Z(n35717) );
  IV U37401 ( .A(n35718), .Z(n35719) );
  XNOR U37402 ( .A(m[698]), .B(n35720), .Z(n35718) );
  NAND U37403 ( .A(n35721), .B(mul_pow), .Z(n35720) );
  XOR U37404 ( .A(m[698]), .B(c[698]), .Z(n35721) );
  XOR U37405 ( .A(n35722), .B(n35723), .Z(n35714) );
  ANDN U37406 ( .B(n35724), .A(n32140), .Z(n35722) );
  XNOR U37407 ( .A(\modmult_1/zin[0][696] ), .B(n35725), .Z(n32140) );
  IV U37408 ( .A(n35723), .Z(n35725) );
  XOR U37409 ( .A(n35723), .B(n32141), .Z(n35724) );
  XNOR U37410 ( .A(n35726), .B(n35727), .Z(n32141) );
  ANDN U37411 ( .B(\modmult_1/xin[1023] ), .A(n35728), .Z(n35726) );
  IV U37412 ( .A(n35727), .Z(n35728) );
  XNOR U37413 ( .A(m[697]), .B(n35729), .Z(n35727) );
  NAND U37414 ( .A(n35730), .B(mul_pow), .Z(n35729) );
  XOR U37415 ( .A(m[697]), .B(c[697]), .Z(n35730) );
  XOR U37416 ( .A(n35731), .B(n35732), .Z(n35723) );
  ANDN U37417 ( .B(n35733), .A(n32138), .Z(n35731) );
  XNOR U37418 ( .A(\modmult_1/zin[0][695] ), .B(n35734), .Z(n32138) );
  IV U37419 ( .A(n35732), .Z(n35734) );
  XOR U37420 ( .A(n35732), .B(n32139), .Z(n35733) );
  XNOR U37421 ( .A(n35735), .B(n35736), .Z(n32139) );
  ANDN U37422 ( .B(\modmult_1/xin[1023] ), .A(n35737), .Z(n35735) );
  IV U37423 ( .A(n35736), .Z(n35737) );
  XNOR U37424 ( .A(m[696]), .B(n35738), .Z(n35736) );
  NAND U37425 ( .A(n35739), .B(mul_pow), .Z(n35738) );
  XOR U37426 ( .A(m[696]), .B(c[696]), .Z(n35739) );
  XOR U37427 ( .A(n35740), .B(n35741), .Z(n35732) );
  ANDN U37428 ( .B(n35742), .A(n32136), .Z(n35740) );
  XNOR U37429 ( .A(\modmult_1/zin[0][694] ), .B(n35743), .Z(n32136) );
  IV U37430 ( .A(n35741), .Z(n35743) );
  XOR U37431 ( .A(n35741), .B(n32137), .Z(n35742) );
  XNOR U37432 ( .A(n35744), .B(n35745), .Z(n32137) );
  ANDN U37433 ( .B(\modmult_1/xin[1023] ), .A(n35746), .Z(n35744) );
  IV U37434 ( .A(n35745), .Z(n35746) );
  XNOR U37435 ( .A(m[695]), .B(n35747), .Z(n35745) );
  NAND U37436 ( .A(n35748), .B(mul_pow), .Z(n35747) );
  XOR U37437 ( .A(m[695]), .B(c[695]), .Z(n35748) );
  XOR U37438 ( .A(n35749), .B(n35750), .Z(n35741) );
  ANDN U37439 ( .B(n35751), .A(n32134), .Z(n35749) );
  XNOR U37440 ( .A(\modmult_1/zin[0][693] ), .B(n35752), .Z(n32134) );
  IV U37441 ( .A(n35750), .Z(n35752) );
  XOR U37442 ( .A(n35750), .B(n32135), .Z(n35751) );
  XNOR U37443 ( .A(n35753), .B(n35754), .Z(n32135) );
  ANDN U37444 ( .B(\modmult_1/xin[1023] ), .A(n35755), .Z(n35753) );
  IV U37445 ( .A(n35754), .Z(n35755) );
  XNOR U37446 ( .A(m[694]), .B(n35756), .Z(n35754) );
  NAND U37447 ( .A(n35757), .B(mul_pow), .Z(n35756) );
  XOR U37448 ( .A(m[694]), .B(c[694]), .Z(n35757) );
  XOR U37449 ( .A(n35758), .B(n35759), .Z(n35750) );
  ANDN U37450 ( .B(n35760), .A(n32132), .Z(n35758) );
  XNOR U37451 ( .A(\modmult_1/zin[0][692] ), .B(n35761), .Z(n32132) );
  IV U37452 ( .A(n35759), .Z(n35761) );
  XOR U37453 ( .A(n35759), .B(n32133), .Z(n35760) );
  XNOR U37454 ( .A(n35762), .B(n35763), .Z(n32133) );
  ANDN U37455 ( .B(\modmult_1/xin[1023] ), .A(n35764), .Z(n35762) );
  IV U37456 ( .A(n35763), .Z(n35764) );
  XNOR U37457 ( .A(m[693]), .B(n35765), .Z(n35763) );
  NAND U37458 ( .A(n35766), .B(mul_pow), .Z(n35765) );
  XOR U37459 ( .A(m[693]), .B(c[693]), .Z(n35766) );
  XOR U37460 ( .A(n35767), .B(n35768), .Z(n35759) );
  ANDN U37461 ( .B(n35769), .A(n32130), .Z(n35767) );
  XNOR U37462 ( .A(\modmult_1/zin[0][691] ), .B(n35770), .Z(n32130) );
  IV U37463 ( .A(n35768), .Z(n35770) );
  XOR U37464 ( .A(n35768), .B(n32131), .Z(n35769) );
  XNOR U37465 ( .A(n35771), .B(n35772), .Z(n32131) );
  ANDN U37466 ( .B(\modmult_1/xin[1023] ), .A(n35773), .Z(n35771) );
  IV U37467 ( .A(n35772), .Z(n35773) );
  XNOR U37468 ( .A(m[692]), .B(n35774), .Z(n35772) );
  NAND U37469 ( .A(n35775), .B(mul_pow), .Z(n35774) );
  XOR U37470 ( .A(m[692]), .B(c[692]), .Z(n35775) );
  XOR U37471 ( .A(n35776), .B(n35777), .Z(n35768) );
  ANDN U37472 ( .B(n35778), .A(n32128), .Z(n35776) );
  XNOR U37473 ( .A(\modmult_1/zin[0][690] ), .B(n35779), .Z(n32128) );
  IV U37474 ( .A(n35777), .Z(n35779) );
  XOR U37475 ( .A(n35777), .B(n32129), .Z(n35778) );
  XNOR U37476 ( .A(n35780), .B(n35781), .Z(n32129) );
  ANDN U37477 ( .B(\modmult_1/xin[1023] ), .A(n35782), .Z(n35780) );
  IV U37478 ( .A(n35781), .Z(n35782) );
  XNOR U37479 ( .A(m[691]), .B(n35783), .Z(n35781) );
  NAND U37480 ( .A(n35784), .B(mul_pow), .Z(n35783) );
  XOR U37481 ( .A(m[691]), .B(c[691]), .Z(n35784) );
  XOR U37482 ( .A(n35785), .B(n35786), .Z(n35777) );
  ANDN U37483 ( .B(n35787), .A(n32126), .Z(n35785) );
  XNOR U37484 ( .A(\modmult_1/zin[0][689] ), .B(n35788), .Z(n32126) );
  IV U37485 ( .A(n35786), .Z(n35788) );
  XOR U37486 ( .A(n35786), .B(n32127), .Z(n35787) );
  XNOR U37487 ( .A(n35789), .B(n35790), .Z(n32127) );
  ANDN U37488 ( .B(\modmult_1/xin[1023] ), .A(n35791), .Z(n35789) );
  IV U37489 ( .A(n35790), .Z(n35791) );
  XNOR U37490 ( .A(m[690]), .B(n35792), .Z(n35790) );
  NAND U37491 ( .A(n35793), .B(mul_pow), .Z(n35792) );
  XOR U37492 ( .A(m[690]), .B(c[690]), .Z(n35793) );
  XOR U37493 ( .A(n35794), .B(n35795), .Z(n35786) );
  ANDN U37494 ( .B(n35796), .A(n32124), .Z(n35794) );
  XNOR U37495 ( .A(\modmult_1/zin[0][688] ), .B(n35797), .Z(n32124) );
  IV U37496 ( .A(n35795), .Z(n35797) );
  XOR U37497 ( .A(n35795), .B(n32125), .Z(n35796) );
  XNOR U37498 ( .A(n35798), .B(n35799), .Z(n32125) );
  ANDN U37499 ( .B(\modmult_1/xin[1023] ), .A(n35800), .Z(n35798) );
  IV U37500 ( .A(n35799), .Z(n35800) );
  XNOR U37501 ( .A(m[689]), .B(n35801), .Z(n35799) );
  NAND U37502 ( .A(n35802), .B(mul_pow), .Z(n35801) );
  XOR U37503 ( .A(m[689]), .B(c[689]), .Z(n35802) );
  XOR U37504 ( .A(n35803), .B(n35804), .Z(n35795) );
  ANDN U37505 ( .B(n35805), .A(n32122), .Z(n35803) );
  XNOR U37506 ( .A(\modmult_1/zin[0][687] ), .B(n35806), .Z(n32122) );
  IV U37507 ( .A(n35804), .Z(n35806) );
  XOR U37508 ( .A(n35804), .B(n32123), .Z(n35805) );
  XNOR U37509 ( .A(n35807), .B(n35808), .Z(n32123) );
  ANDN U37510 ( .B(\modmult_1/xin[1023] ), .A(n35809), .Z(n35807) );
  IV U37511 ( .A(n35808), .Z(n35809) );
  XNOR U37512 ( .A(m[688]), .B(n35810), .Z(n35808) );
  NAND U37513 ( .A(n35811), .B(mul_pow), .Z(n35810) );
  XOR U37514 ( .A(m[688]), .B(c[688]), .Z(n35811) );
  XOR U37515 ( .A(n35812), .B(n35813), .Z(n35804) );
  ANDN U37516 ( .B(n35814), .A(n32120), .Z(n35812) );
  XNOR U37517 ( .A(\modmult_1/zin[0][686] ), .B(n35815), .Z(n32120) );
  IV U37518 ( .A(n35813), .Z(n35815) );
  XOR U37519 ( .A(n35813), .B(n32121), .Z(n35814) );
  XNOR U37520 ( .A(n35816), .B(n35817), .Z(n32121) );
  ANDN U37521 ( .B(\modmult_1/xin[1023] ), .A(n35818), .Z(n35816) );
  IV U37522 ( .A(n35817), .Z(n35818) );
  XNOR U37523 ( .A(m[687]), .B(n35819), .Z(n35817) );
  NAND U37524 ( .A(n35820), .B(mul_pow), .Z(n35819) );
  XOR U37525 ( .A(m[687]), .B(c[687]), .Z(n35820) );
  XOR U37526 ( .A(n35821), .B(n35822), .Z(n35813) );
  ANDN U37527 ( .B(n35823), .A(n32118), .Z(n35821) );
  XNOR U37528 ( .A(\modmult_1/zin[0][685] ), .B(n35824), .Z(n32118) );
  IV U37529 ( .A(n35822), .Z(n35824) );
  XOR U37530 ( .A(n35822), .B(n32119), .Z(n35823) );
  XNOR U37531 ( .A(n35825), .B(n35826), .Z(n32119) );
  ANDN U37532 ( .B(\modmult_1/xin[1023] ), .A(n35827), .Z(n35825) );
  IV U37533 ( .A(n35826), .Z(n35827) );
  XNOR U37534 ( .A(m[686]), .B(n35828), .Z(n35826) );
  NAND U37535 ( .A(n35829), .B(mul_pow), .Z(n35828) );
  XOR U37536 ( .A(m[686]), .B(c[686]), .Z(n35829) );
  XOR U37537 ( .A(n35830), .B(n35831), .Z(n35822) );
  ANDN U37538 ( .B(n35832), .A(n32116), .Z(n35830) );
  XNOR U37539 ( .A(\modmult_1/zin[0][684] ), .B(n35833), .Z(n32116) );
  IV U37540 ( .A(n35831), .Z(n35833) );
  XOR U37541 ( .A(n35831), .B(n32117), .Z(n35832) );
  XNOR U37542 ( .A(n35834), .B(n35835), .Z(n32117) );
  ANDN U37543 ( .B(\modmult_1/xin[1023] ), .A(n35836), .Z(n35834) );
  IV U37544 ( .A(n35835), .Z(n35836) );
  XNOR U37545 ( .A(m[685]), .B(n35837), .Z(n35835) );
  NAND U37546 ( .A(n35838), .B(mul_pow), .Z(n35837) );
  XOR U37547 ( .A(m[685]), .B(c[685]), .Z(n35838) );
  XOR U37548 ( .A(n35839), .B(n35840), .Z(n35831) );
  ANDN U37549 ( .B(n35841), .A(n32114), .Z(n35839) );
  XNOR U37550 ( .A(\modmult_1/zin[0][683] ), .B(n35842), .Z(n32114) );
  IV U37551 ( .A(n35840), .Z(n35842) );
  XOR U37552 ( .A(n35840), .B(n32115), .Z(n35841) );
  XNOR U37553 ( .A(n35843), .B(n35844), .Z(n32115) );
  ANDN U37554 ( .B(\modmult_1/xin[1023] ), .A(n35845), .Z(n35843) );
  IV U37555 ( .A(n35844), .Z(n35845) );
  XNOR U37556 ( .A(m[684]), .B(n35846), .Z(n35844) );
  NAND U37557 ( .A(n35847), .B(mul_pow), .Z(n35846) );
  XOR U37558 ( .A(m[684]), .B(c[684]), .Z(n35847) );
  XOR U37559 ( .A(n35848), .B(n35849), .Z(n35840) );
  ANDN U37560 ( .B(n35850), .A(n32112), .Z(n35848) );
  XNOR U37561 ( .A(\modmult_1/zin[0][682] ), .B(n35851), .Z(n32112) );
  IV U37562 ( .A(n35849), .Z(n35851) );
  XOR U37563 ( .A(n35849), .B(n32113), .Z(n35850) );
  XNOR U37564 ( .A(n35852), .B(n35853), .Z(n32113) );
  ANDN U37565 ( .B(\modmult_1/xin[1023] ), .A(n35854), .Z(n35852) );
  IV U37566 ( .A(n35853), .Z(n35854) );
  XNOR U37567 ( .A(m[683]), .B(n35855), .Z(n35853) );
  NAND U37568 ( .A(n35856), .B(mul_pow), .Z(n35855) );
  XOR U37569 ( .A(m[683]), .B(c[683]), .Z(n35856) );
  XOR U37570 ( .A(n35857), .B(n35858), .Z(n35849) );
  ANDN U37571 ( .B(n35859), .A(n32110), .Z(n35857) );
  XNOR U37572 ( .A(\modmult_1/zin[0][681] ), .B(n35860), .Z(n32110) );
  IV U37573 ( .A(n35858), .Z(n35860) );
  XOR U37574 ( .A(n35858), .B(n32111), .Z(n35859) );
  XNOR U37575 ( .A(n35861), .B(n35862), .Z(n32111) );
  ANDN U37576 ( .B(\modmult_1/xin[1023] ), .A(n35863), .Z(n35861) );
  IV U37577 ( .A(n35862), .Z(n35863) );
  XNOR U37578 ( .A(m[682]), .B(n35864), .Z(n35862) );
  NAND U37579 ( .A(n35865), .B(mul_pow), .Z(n35864) );
  XOR U37580 ( .A(m[682]), .B(c[682]), .Z(n35865) );
  XOR U37581 ( .A(n35866), .B(n35867), .Z(n35858) );
  ANDN U37582 ( .B(n35868), .A(n32108), .Z(n35866) );
  XNOR U37583 ( .A(\modmult_1/zin[0][680] ), .B(n35869), .Z(n32108) );
  IV U37584 ( .A(n35867), .Z(n35869) );
  XOR U37585 ( .A(n35867), .B(n32109), .Z(n35868) );
  XNOR U37586 ( .A(n35870), .B(n35871), .Z(n32109) );
  ANDN U37587 ( .B(\modmult_1/xin[1023] ), .A(n35872), .Z(n35870) );
  IV U37588 ( .A(n35871), .Z(n35872) );
  XNOR U37589 ( .A(m[681]), .B(n35873), .Z(n35871) );
  NAND U37590 ( .A(n35874), .B(mul_pow), .Z(n35873) );
  XOR U37591 ( .A(m[681]), .B(c[681]), .Z(n35874) );
  XOR U37592 ( .A(n35875), .B(n35876), .Z(n35867) );
  ANDN U37593 ( .B(n35877), .A(n32106), .Z(n35875) );
  XNOR U37594 ( .A(\modmult_1/zin[0][679] ), .B(n35878), .Z(n32106) );
  IV U37595 ( .A(n35876), .Z(n35878) );
  XOR U37596 ( .A(n35876), .B(n32107), .Z(n35877) );
  XNOR U37597 ( .A(n35879), .B(n35880), .Z(n32107) );
  ANDN U37598 ( .B(\modmult_1/xin[1023] ), .A(n35881), .Z(n35879) );
  IV U37599 ( .A(n35880), .Z(n35881) );
  XNOR U37600 ( .A(m[680]), .B(n35882), .Z(n35880) );
  NAND U37601 ( .A(n35883), .B(mul_pow), .Z(n35882) );
  XOR U37602 ( .A(m[680]), .B(c[680]), .Z(n35883) );
  XOR U37603 ( .A(n35884), .B(n35885), .Z(n35876) );
  ANDN U37604 ( .B(n35886), .A(n32104), .Z(n35884) );
  XNOR U37605 ( .A(\modmult_1/zin[0][678] ), .B(n35887), .Z(n32104) );
  IV U37606 ( .A(n35885), .Z(n35887) );
  XOR U37607 ( .A(n35885), .B(n32105), .Z(n35886) );
  XNOR U37608 ( .A(n35888), .B(n35889), .Z(n32105) );
  ANDN U37609 ( .B(\modmult_1/xin[1023] ), .A(n35890), .Z(n35888) );
  IV U37610 ( .A(n35889), .Z(n35890) );
  XNOR U37611 ( .A(m[679]), .B(n35891), .Z(n35889) );
  NAND U37612 ( .A(n35892), .B(mul_pow), .Z(n35891) );
  XOR U37613 ( .A(m[679]), .B(c[679]), .Z(n35892) );
  XOR U37614 ( .A(n35893), .B(n35894), .Z(n35885) );
  ANDN U37615 ( .B(n35895), .A(n32102), .Z(n35893) );
  XNOR U37616 ( .A(\modmult_1/zin[0][677] ), .B(n35896), .Z(n32102) );
  IV U37617 ( .A(n35894), .Z(n35896) );
  XOR U37618 ( .A(n35894), .B(n32103), .Z(n35895) );
  XNOR U37619 ( .A(n35897), .B(n35898), .Z(n32103) );
  ANDN U37620 ( .B(\modmult_1/xin[1023] ), .A(n35899), .Z(n35897) );
  IV U37621 ( .A(n35898), .Z(n35899) );
  XNOR U37622 ( .A(m[678]), .B(n35900), .Z(n35898) );
  NAND U37623 ( .A(n35901), .B(mul_pow), .Z(n35900) );
  XOR U37624 ( .A(m[678]), .B(c[678]), .Z(n35901) );
  XOR U37625 ( .A(n35902), .B(n35903), .Z(n35894) );
  ANDN U37626 ( .B(n35904), .A(n32100), .Z(n35902) );
  XNOR U37627 ( .A(\modmult_1/zin[0][676] ), .B(n35905), .Z(n32100) );
  IV U37628 ( .A(n35903), .Z(n35905) );
  XOR U37629 ( .A(n35903), .B(n32101), .Z(n35904) );
  XNOR U37630 ( .A(n35906), .B(n35907), .Z(n32101) );
  ANDN U37631 ( .B(\modmult_1/xin[1023] ), .A(n35908), .Z(n35906) );
  IV U37632 ( .A(n35907), .Z(n35908) );
  XNOR U37633 ( .A(m[677]), .B(n35909), .Z(n35907) );
  NAND U37634 ( .A(n35910), .B(mul_pow), .Z(n35909) );
  XOR U37635 ( .A(m[677]), .B(c[677]), .Z(n35910) );
  XOR U37636 ( .A(n35911), .B(n35912), .Z(n35903) );
  ANDN U37637 ( .B(n35913), .A(n32098), .Z(n35911) );
  XNOR U37638 ( .A(\modmult_1/zin[0][675] ), .B(n35914), .Z(n32098) );
  IV U37639 ( .A(n35912), .Z(n35914) );
  XOR U37640 ( .A(n35912), .B(n32099), .Z(n35913) );
  XNOR U37641 ( .A(n35915), .B(n35916), .Z(n32099) );
  ANDN U37642 ( .B(\modmult_1/xin[1023] ), .A(n35917), .Z(n35915) );
  IV U37643 ( .A(n35916), .Z(n35917) );
  XNOR U37644 ( .A(m[676]), .B(n35918), .Z(n35916) );
  NAND U37645 ( .A(n35919), .B(mul_pow), .Z(n35918) );
  XOR U37646 ( .A(m[676]), .B(c[676]), .Z(n35919) );
  XOR U37647 ( .A(n35920), .B(n35921), .Z(n35912) );
  ANDN U37648 ( .B(n35922), .A(n32096), .Z(n35920) );
  XNOR U37649 ( .A(\modmult_1/zin[0][674] ), .B(n35923), .Z(n32096) );
  IV U37650 ( .A(n35921), .Z(n35923) );
  XOR U37651 ( .A(n35921), .B(n32097), .Z(n35922) );
  XNOR U37652 ( .A(n35924), .B(n35925), .Z(n32097) );
  ANDN U37653 ( .B(\modmult_1/xin[1023] ), .A(n35926), .Z(n35924) );
  IV U37654 ( .A(n35925), .Z(n35926) );
  XNOR U37655 ( .A(m[675]), .B(n35927), .Z(n35925) );
  NAND U37656 ( .A(n35928), .B(mul_pow), .Z(n35927) );
  XOR U37657 ( .A(m[675]), .B(c[675]), .Z(n35928) );
  XOR U37658 ( .A(n35929), .B(n35930), .Z(n35921) );
  ANDN U37659 ( .B(n35931), .A(n32094), .Z(n35929) );
  XNOR U37660 ( .A(\modmult_1/zin[0][673] ), .B(n35932), .Z(n32094) );
  IV U37661 ( .A(n35930), .Z(n35932) );
  XOR U37662 ( .A(n35930), .B(n32095), .Z(n35931) );
  XNOR U37663 ( .A(n35933), .B(n35934), .Z(n32095) );
  ANDN U37664 ( .B(\modmult_1/xin[1023] ), .A(n35935), .Z(n35933) );
  IV U37665 ( .A(n35934), .Z(n35935) );
  XNOR U37666 ( .A(m[674]), .B(n35936), .Z(n35934) );
  NAND U37667 ( .A(n35937), .B(mul_pow), .Z(n35936) );
  XOR U37668 ( .A(m[674]), .B(c[674]), .Z(n35937) );
  XOR U37669 ( .A(n35938), .B(n35939), .Z(n35930) );
  ANDN U37670 ( .B(n35940), .A(n32092), .Z(n35938) );
  XNOR U37671 ( .A(\modmult_1/zin[0][672] ), .B(n35941), .Z(n32092) );
  IV U37672 ( .A(n35939), .Z(n35941) );
  XOR U37673 ( .A(n35939), .B(n32093), .Z(n35940) );
  XNOR U37674 ( .A(n35942), .B(n35943), .Z(n32093) );
  ANDN U37675 ( .B(\modmult_1/xin[1023] ), .A(n35944), .Z(n35942) );
  IV U37676 ( .A(n35943), .Z(n35944) );
  XNOR U37677 ( .A(m[673]), .B(n35945), .Z(n35943) );
  NAND U37678 ( .A(n35946), .B(mul_pow), .Z(n35945) );
  XOR U37679 ( .A(m[673]), .B(c[673]), .Z(n35946) );
  XOR U37680 ( .A(n35947), .B(n35948), .Z(n35939) );
  ANDN U37681 ( .B(n35949), .A(n32090), .Z(n35947) );
  XNOR U37682 ( .A(\modmult_1/zin[0][671] ), .B(n35950), .Z(n32090) );
  IV U37683 ( .A(n35948), .Z(n35950) );
  XOR U37684 ( .A(n35948), .B(n32091), .Z(n35949) );
  XNOR U37685 ( .A(n35951), .B(n35952), .Z(n32091) );
  ANDN U37686 ( .B(\modmult_1/xin[1023] ), .A(n35953), .Z(n35951) );
  IV U37687 ( .A(n35952), .Z(n35953) );
  XNOR U37688 ( .A(m[672]), .B(n35954), .Z(n35952) );
  NAND U37689 ( .A(n35955), .B(mul_pow), .Z(n35954) );
  XOR U37690 ( .A(m[672]), .B(c[672]), .Z(n35955) );
  XOR U37691 ( .A(n35956), .B(n35957), .Z(n35948) );
  ANDN U37692 ( .B(n35958), .A(n32088), .Z(n35956) );
  XNOR U37693 ( .A(\modmult_1/zin[0][670] ), .B(n35959), .Z(n32088) );
  IV U37694 ( .A(n35957), .Z(n35959) );
  XOR U37695 ( .A(n35957), .B(n32089), .Z(n35958) );
  XNOR U37696 ( .A(n35960), .B(n35961), .Z(n32089) );
  ANDN U37697 ( .B(\modmult_1/xin[1023] ), .A(n35962), .Z(n35960) );
  IV U37698 ( .A(n35961), .Z(n35962) );
  XNOR U37699 ( .A(m[671]), .B(n35963), .Z(n35961) );
  NAND U37700 ( .A(n35964), .B(mul_pow), .Z(n35963) );
  XOR U37701 ( .A(m[671]), .B(c[671]), .Z(n35964) );
  XOR U37702 ( .A(n35965), .B(n35966), .Z(n35957) );
  ANDN U37703 ( .B(n35967), .A(n32086), .Z(n35965) );
  XNOR U37704 ( .A(\modmult_1/zin[0][669] ), .B(n35968), .Z(n32086) );
  IV U37705 ( .A(n35966), .Z(n35968) );
  XOR U37706 ( .A(n35966), .B(n32087), .Z(n35967) );
  XNOR U37707 ( .A(n35969), .B(n35970), .Z(n32087) );
  ANDN U37708 ( .B(\modmult_1/xin[1023] ), .A(n35971), .Z(n35969) );
  IV U37709 ( .A(n35970), .Z(n35971) );
  XNOR U37710 ( .A(m[670]), .B(n35972), .Z(n35970) );
  NAND U37711 ( .A(n35973), .B(mul_pow), .Z(n35972) );
  XOR U37712 ( .A(m[670]), .B(c[670]), .Z(n35973) );
  XOR U37713 ( .A(n35974), .B(n35975), .Z(n35966) );
  ANDN U37714 ( .B(n35976), .A(n32084), .Z(n35974) );
  XNOR U37715 ( .A(\modmult_1/zin[0][668] ), .B(n35977), .Z(n32084) );
  IV U37716 ( .A(n35975), .Z(n35977) );
  XOR U37717 ( .A(n35975), .B(n32085), .Z(n35976) );
  XNOR U37718 ( .A(n35978), .B(n35979), .Z(n32085) );
  ANDN U37719 ( .B(\modmult_1/xin[1023] ), .A(n35980), .Z(n35978) );
  IV U37720 ( .A(n35979), .Z(n35980) );
  XNOR U37721 ( .A(m[669]), .B(n35981), .Z(n35979) );
  NAND U37722 ( .A(n35982), .B(mul_pow), .Z(n35981) );
  XOR U37723 ( .A(m[669]), .B(c[669]), .Z(n35982) );
  XOR U37724 ( .A(n35983), .B(n35984), .Z(n35975) );
  ANDN U37725 ( .B(n35985), .A(n32082), .Z(n35983) );
  XNOR U37726 ( .A(\modmult_1/zin[0][667] ), .B(n35986), .Z(n32082) );
  IV U37727 ( .A(n35984), .Z(n35986) );
  XOR U37728 ( .A(n35984), .B(n32083), .Z(n35985) );
  XNOR U37729 ( .A(n35987), .B(n35988), .Z(n32083) );
  ANDN U37730 ( .B(\modmult_1/xin[1023] ), .A(n35989), .Z(n35987) );
  IV U37731 ( .A(n35988), .Z(n35989) );
  XNOR U37732 ( .A(m[668]), .B(n35990), .Z(n35988) );
  NAND U37733 ( .A(n35991), .B(mul_pow), .Z(n35990) );
  XOR U37734 ( .A(m[668]), .B(c[668]), .Z(n35991) );
  XOR U37735 ( .A(n35992), .B(n35993), .Z(n35984) );
  ANDN U37736 ( .B(n35994), .A(n32080), .Z(n35992) );
  XNOR U37737 ( .A(\modmult_1/zin[0][666] ), .B(n35995), .Z(n32080) );
  IV U37738 ( .A(n35993), .Z(n35995) );
  XOR U37739 ( .A(n35993), .B(n32081), .Z(n35994) );
  XNOR U37740 ( .A(n35996), .B(n35997), .Z(n32081) );
  ANDN U37741 ( .B(\modmult_1/xin[1023] ), .A(n35998), .Z(n35996) );
  IV U37742 ( .A(n35997), .Z(n35998) );
  XNOR U37743 ( .A(m[667]), .B(n35999), .Z(n35997) );
  NAND U37744 ( .A(n36000), .B(mul_pow), .Z(n35999) );
  XOR U37745 ( .A(m[667]), .B(c[667]), .Z(n36000) );
  XOR U37746 ( .A(n36001), .B(n36002), .Z(n35993) );
  ANDN U37747 ( .B(n36003), .A(n32078), .Z(n36001) );
  XNOR U37748 ( .A(\modmult_1/zin[0][665] ), .B(n36004), .Z(n32078) );
  IV U37749 ( .A(n36002), .Z(n36004) );
  XOR U37750 ( .A(n36002), .B(n32079), .Z(n36003) );
  XNOR U37751 ( .A(n36005), .B(n36006), .Z(n32079) );
  ANDN U37752 ( .B(\modmult_1/xin[1023] ), .A(n36007), .Z(n36005) );
  IV U37753 ( .A(n36006), .Z(n36007) );
  XNOR U37754 ( .A(m[666]), .B(n36008), .Z(n36006) );
  NAND U37755 ( .A(n36009), .B(mul_pow), .Z(n36008) );
  XOR U37756 ( .A(m[666]), .B(c[666]), .Z(n36009) );
  XOR U37757 ( .A(n36010), .B(n36011), .Z(n36002) );
  ANDN U37758 ( .B(n36012), .A(n32076), .Z(n36010) );
  XNOR U37759 ( .A(\modmult_1/zin[0][664] ), .B(n36013), .Z(n32076) );
  IV U37760 ( .A(n36011), .Z(n36013) );
  XOR U37761 ( .A(n36011), .B(n32077), .Z(n36012) );
  XNOR U37762 ( .A(n36014), .B(n36015), .Z(n32077) );
  ANDN U37763 ( .B(\modmult_1/xin[1023] ), .A(n36016), .Z(n36014) );
  IV U37764 ( .A(n36015), .Z(n36016) );
  XNOR U37765 ( .A(m[665]), .B(n36017), .Z(n36015) );
  NAND U37766 ( .A(n36018), .B(mul_pow), .Z(n36017) );
  XOR U37767 ( .A(m[665]), .B(c[665]), .Z(n36018) );
  XOR U37768 ( .A(n36019), .B(n36020), .Z(n36011) );
  ANDN U37769 ( .B(n36021), .A(n32074), .Z(n36019) );
  XNOR U37770 ( .A(\modmult_1/zin[0][663] ), .B(n36022), .Z(n32074) );
  IV U37771 ( .A(n36020), .Z(n36022) );
  XOR U37772 ( .A(n36020), .B(n32075), .Z(n36021) );
  XNOR U37773 ( .A(n36023), .B(n36024), .Z(n32075) );
  ANDN U37774 ( .B(\modmult_1/xin[1023] ), .A(n36025), .Z(n36023) );
  IV U37775 ( .A(n36024), .Z(n36025) );
  XNOR U37776 ( .A(m[664]), .B(n36026), .Z(n36024) );
  NAND U37777 ( .A(n36027), .B(mul_pow), .Z(n36026) );
  XOR U37778 ( .A(m[664]), .B(c[664]), .Z(n36027) );
  XOR U37779 ( .A(n36028), .B(n36029), .Z(n36020) );
  ANDN U37780 ( .B(n36030), .A(n32072), .Z(n36028) );
  XNOR U37781 ( .A(\modmult_1/zin[0][662] ), .B(n36031), .Z(n32072) );
  IV U37782 ( .A(n36029), .Z(n36031) );
  XOR U37783 ( .A(n36029), .B(n32073), .Z(n36030) );
  XNOR U37784 ( .A(n36032), .B(n36033), .Z(n32073) );
  ANDN U37785 ( .B(\modmult_1/xin[1023] ), .A(n36034), .Z(n36032) );
  IV U37786 ( .A(n36033), .Z(n36034) );
  XNOR U37787 ( .A(m[663]), .B(n36035), .Z(n36033) );
  NAND U37788 ( .A(n36036), .B(mul_pow), .Z(n36035) );
  XOR U37789 ( .A(m[663]), .B(c[663]), .Z(n36036) );
  XOR U37790 ( .A(n36037), .B(n36038), .Z(n36029) );
  ANDN U37791 ( .B(n36039), .A(n32070), .Z(n36037) );
  XNOR U37792 ( .A(\modmult_1/zin[0][661] ), .B(n36040), .Z(n32070) );
  IV U37793 ( .A(n36038), .Z(n36040) );
  XOR U37794 ( .A(n36038), .B(n32071), .Z(n36039) );
  XNOR U37795 ( .A(n36041), .B(n36042), .Z(n32071) );
  ANDN U37796 ( .B(\modmult_1/xin[1023] ), .A(n36043), .Z(n36041) );
  IV U37797 ( .A(n36042), .Z(n36043) );
  XNOR U37798 ( .A(m[662]), .B(n36044), .Z(n36042) );
  NAND U37799 ( .A(n36045), .B(mul_pow), .Z(n36044) );
  XOR U37800 ( .A(m[662]), .B(c[662]), .Z(n36045) );
  XOR U37801 ( .A(n36046), .B(n36047), .Z(n36038) );
  ANDN U37802 ( .B(n36048), .A(n32068), .Z(n36046) );
  XNOR U37803 ( .A(\modmult_1/zin[0][660] ), .B(n36049), .Z(n32068) );
  IV U37804 ( .A(n36047), .Z(n36049) );
  XOR U37805 ( .A(n36047), .B(n32069), .Z(n36048) );
  XNOR U37806 ( .A(n36050), .B(n36051), .Z(n32069) );
  ANDN U37807 ( .B(\modmult_1/xin[1023] ), .A(n36052), .Z(n36050) );
  IV U37808 ( .A(n36051), .Z(n36052) );
  XNOR U37809 ( .A(m[661]), .B(n36053), .Z(n36051) );
  NAND U37810 ( .A(n36054), .B(mul_pow), .Z(n36053) );
  XOR U37811 ( .A(m[661]), .B(c[661]), .Z(n36054) );
  XOR U37812 ( .A(n36055), .B(n36056), .Z(n36047) );
  ANDN U37813 ( .B(n36057), .A(n32066), .Z(n36055) );
  XNOR U37814 ( .A(\modmult_1/zin[0][659] ), .B(n36058), .Z(n32066) );
  IV U37815 ( .A(n36056), .Z(n36058) );
  XOR U37816 ( .A(n36056), .B(n32067), .Z(n36057) );
  XNOR U37817 ( .A(n36059), .B(n36060), .Z(n32067) );
  ANDN U37818 ( .B(\modmult_1/xin[1023] ), .A(n36061), .Z(n36059) );
  IV U37819 ( .A(n36060), .Z(n36061) );
  XNOR U37820 ( .A(m[660]), .B(n36062), .Z(n36060) );
  NAND U37821 ( .A(n36063), .B(mul_pow), .Z(n36062) );
  XOR U37822 ( .A(m[660]), .B(c[660]), .Z(n36063) );
  XOR U37823 ( .A(n36064), .B(n36065), .Z(n36056) );
  ANDN U37824 ( .B(n36066), .A(n32064), .Z(n36064) );
  XNOR U37825 ( .A(\modmult_1/zin[0][658] ), .B(n36067), .Z(n32064) );
  IV U37826 ( .A(n36065), .Z(n36067) );
  XOR U37827 ( .A(n36065), .B(n32065), .Z(n36066) );
  XNOR U37828 ( .A(n36068), .B(n36069), .Z(n32065) );
  ANDN U37829 ( .B(\modmult_1/xin[1023] ), .A(n36070), .Z(n36068) );
  IV U37830 ( .A(n36069), .Z(n36070) );
  XNOR U37831 ( .A(m[659]), .B(n36071), .Z(n36069) );
  NAND U37832 ( .A(n36072), .B(mul_pow), .Z(n36071) );
  XOR U37833 ( .A(m[659]), .B(c[659]), .Z(n36072) );
  XOR U37834 ( .A(n36073), .B(n36074), .Z(n36065) );
  ANDN U37835 ( .B(n36075), .A(n32062), .Z(n36073) );
  XNOR U37836 ( .A(\modmult_1/zin[0][657] ), .B(n36076), .Z(n32062) );
  IV U37837 ( .A(n36074), .Z(n36076) );
  XOR U37838 ( .A(n36074), .B(n32063), .Z(n36075) );
  XNOR U37839 ( .A(n36077), .B(n36078), .Z(n32063) );
  ANDN U37840 ( .B(\modmult_1/xin[1023] ), .A(n36079), .Z(n36077) );
  IV U37841 ( .A(n36078), .Z(n36079) );
  XNOR U37842 ( .A(m[658]), .B(n36080), .Z(n36078) );
  NAND U37843 ( .A(n36081), .B(mul_pow), .Z(n36080) );
  XOR U37844 ( .A(m[658]), .B(c[658]), .Z(n36081) );
  XOR U37845 ( .A(n36082), .B(n36083), .Z(n36074) );
  ANDN U37846 ( .B(n36084), .A(n32060), .Z(n36082) );
  XNOR U37847 ( .A(\modmult_1/zin[0][656] ), .B(n36085), .Z(n32060) );
  IV U37848 ( .A(n36083), .Z(n36085) );
  XOR U37849 ( .A(n36083), .B(n32061), .Z(n36084) );
  XNOR U37850 ( .A(n36086), .B(n36087), .Z(n32061) );
  ANDN U37851 ( .B(\modmult_1/xin[1023] ), .A(n36088), .Z(n36086) );
  IV U37852 ( .A(n36087), .Z(n36088) );
  XNOR U37853 ( .A(m[657]), .B(n36089), .Z(n36087) );
  NAND U37854 ( .A(n36090), .B(mul_pow), .Z(n36089) );
  XOR U37855 ( .A(m[657]), .B(c[657]), .Z(n36090) );
  XOR U37856 ( .A(n36091), .B(n36092), .Z(n36083) );
  ANDN U37857 ( .B(n36093), .A(n32058), .Z(n36091) );
  XNOR U37858 ( .A(\modmult_1/zin[0][655] ), .B(n36094), .Z(n32058) );
  IV U37859 ( .A(n36092), .Z(n36094) );
  XOR U37860 ( .A(n36092), .B(n32059), .Z(n36093) );
  XNOR U37861 ( .A(n36095), .B(n36096), .Z(n32059) );
  ANDN U37862 ( .B(\modmult_1/xin[1023] ), .A(n36097), .Z(n36095) );
  IV U37863 ( .A(n36096), .Z(n36097) );
  XNOR U37864 ( .A(m[656]), .B(n36098), .Z(n36096) );
  NAND U37865 ( .A(n36099), .B(mul_pow), .Z(n36098) );
  XOR U37866 ( .A(m[656]), .B(c[656]), .Z(n36099) );
  XOR U37867 ( .A(n36100), .B(n36101), .Z(n36092) );
  ANDN U37868 ( .B(n36102), .A(n32056), .Z(n36100) );
  XNOR U37869 ( .A(\modmult_1/zin[0][654] ), .B(n36103), .Z(n32056) );
  IV U37870 ( .A(n36101), .Z(n36103) );
  XOR U37871 ( .A(n36101), .B(n32057), .Z(n36102) );
  XNOR U37872 ( .A(n36104), .B(n36105), .Z(n32057) );
  ANDN U37873 ( .B(\modmult_1/xin[1023] ), .A(n36106), .Z(n36104) );
  IV U37874 ( .A(n36105), .Z(n36106) );
  XNOR U37875 ( .A(m[655]), .B(n36107), .Z(n36105) );
  NAND U37876 ( .A(n36108), .B(mul_pow), .Z(n36107) );
  XOR U37877 ( .A(m[655]), .B(c[655]), .Z(n36108) );
  XOR U37878 ( .A(n36109), .B(n36110), .Z(n36101) );
  ANDN U37879 ( .B(n36111), .A(n32054), .Z(n36109) );
  XNOR U37880 ( .A(\modmult_1/zin[0][653] ), .B(n36112), .Z(n32054) );
  IV U37881 ( .A(n36110), .Z(n36112) );
  XOR U37882 ( .A(n36110), .B(n32055), .Z(n36111) );
  XNOR U37883 ( .A(n36113), .B(n36114), .Z(n32055) );
  ANDN U37884 ( .B(\modmult_1/xin[1023] ), .A(n36115), .Z(n36113) );
  IV U37885 ( .A(n36114), .Z(n36115) );
  XNOR U37886 ( .A(m[654]), .B(n36116), .Z(n36114) );
  NAND U37887 ( .A(n36117), .B(mul_pow), .Z(n36116) );
  XOR U37888 ( .A(m[654]), .B(c[654]), .Z(n36117) );
  XOR U37889 ( .A(n36118), .B(n36119), .Z(n36110) );
  ANDN U37890 ( .B(n36120), .A(n32052), .Z(n36118) );
  XNOR U37891 ( .A(\modmult_1/zin[0][652] ), .B(n36121), .Z(n32052) );
  IV U37892 ( .A(n36119), .Z(n36121) );
  XOR U37893 ( .A(n36119), .B(n32053), .Z(n36120) );
  XNOR U37894 ( .A(n36122), .B(n36123), .Z(n32053) );
  ANDN U37895 ( .B(\modmult_1/xin[1023] ), .A(n36124), .Z(n36122) );
  IV U37896 ( .A(n36123), .Z(n36124) );
  XNOR U37897 ( .A(m[653]), .B(n36125), .Z(n36123) );
  NAND U37898 ( .A(n36126), .B(mul_pow), .Z(n36125) );
  XOR U37899 ( .A(m[653]), .B(c[653]), .Z(n36126) );
  XOR U37900 ( .A(n36127), .B(n36128), .Z(n36119) );
  ANDN U37901 ( .B(n36129), .A(n32050), .Z(n36127) );
  XNOR U37902 ( .A(\modmult_1/zin[0][651] ), .B(n36130), .Z(n32050) );
  IV U37903 ( .A(n36128), .Z(n36130) );
  XOR U37904 ( .A(n36128), .B(n32051), .Z(n36129) );
  XNOR U37905 ( .A(n36131), .B(n36132), .Z(n32051) );
  ANDN U37906 ( .B(\modmult_1/xin[1023] ), .A(n36133), .Z(n36131) );
  IV U37907 ( .A(n36132), .Z(n36133) );
  XNOR U37908 ( .A(m[652]), .B(n36134), .Z(n36132) );
  NAND U37909 ( .A(n36135), .B(mul_pow), .Z(n36134) );
  XOR U37910 ( .A(m[652]), .B(c[652]), .Z(n36135) );
  XOR U37911 ( .A(n36136), .B(n36137), .Z(n36128) );
  ANDN U37912 ( .B(n36138), .A(n32048), .Z(n36136) );
  XNOR U37913 ( .A(\modmult_1/zin[0][650] ), .B(n36139), .Z(n32048) );
  IV U37914 ( .A(n36137), .Z(n36139) );
  XOR U37915 ( .A(n36137), .B(n32049), .Z(n36138) );
  XNOR U37916 ( .A(n36140), .B(n36141), .Z(n32049) );
  ANDN U37917 ( .B(\modmult_1/xin[1023] ), .A(n36142), .Z(n36140) );
  IV U37918 ( .A(n36141), .Z(n36142) );
  XNOR U37919 ( .A(m[651]), .B(n36143), .Z(n36141) );
  NAND U37920 ( .A(n36144), .B(mul_pow), .Z(n36143) );
  XOR U37921 ( .A(m[651]), .B(c[651]), .Z(n36144) );
  XOR U37922 ( .A(n36145), .B(n36146), .Z(n36137) );
  ANDN U37923 ( .B(n36147), .A(n32046), .Z(n36145) );
  XNOR U37924 ( .A(\modmult_1/zin[0][649] ), .B(n36148), .Z(n32046) );
  IV U37925 ( .A(n36146), .Z(n36148) );
  XOR U37926 ( .A(n36146), .B(n32047), .Z(n36147) );
  XNOR U37927 ( .A(n36149), .B(n36150), .Z(n32047) );
  ANDN U37928 ( .B(\modmult_1/xin[1023] ), .A(n36151), .Z(n36149) );
  IV U37929 ( .A(n36150), .Z(n36151) );
  XNOR U37930 ( .A(m[650]), .B(n36152), .Z(n36150) );
  NAND U37931 ( .A(n36153), .B(mul_pow), .Z(n36152) );
  XOR U37932 ( .A(m[650]), .B(c[650]), .Z(n36153) );
  XOR U37933 ( .A(n36154), .B(n36155), .Z(n36146) );
  ANDN U37934 ( .B(n36156), .A(n32044), .Z(n36154) );
  XNOR U37935 ( .A(\modmult_1/zin[0][648] ), .B(n36157), .Z(n32044) );
  IV U37936 ( .A(n36155), .Z(n36157) );
  XOR U37937 ( .A(n36155), .B(n32045), .Z(n36156) );
  XNOR U37938 ( .A(n36158), .B(n36159), .Z(n32045) );
  ANDN U37939 ( .B(\modmult_1/xin[1023] ), .A(n36160), .Z(n36158) );
  IV U37940 ( .A(n36159), .Z(n36160) );
  XNOR U37941 ( .A(m[649]), .B(n36161), .Z(n36159) );
  NAND U37942 ( .A(n36162), .B(mul_pow), .Z(n36161) );
  XOR U37943 ( .A(m[649]), .B(c[649]), .Z(n36162) );
  XOR U37944 ( .A(n36163), .B(n36164), .Z(n36155) );
  ANDN U37945 ( .B(n36165), .A(n32042), .Z(n36163) );
  XNOR U37946 ( .A(\modmult_1/zin[0][647] ), .B(n36166), .Z(n32042) );
  IV U37947 ( .A(n36164), .Z(n36166) );
  XOR U37948 ( .A(n36164), .B(n32043), .Z(n36165) );
  XNOR U37949 ( .A(n36167), .B(n36168), .Z(n32043) );
  ANDN U37950 ( .B(\modmult_1/xin[1023] ), .A(n36169), .Z(n36167) );
  IV U37951 ( .A(n36168), .Z(n36169) );
  XNOR U37952 ( .A(m[648]), .B(n36170), .Z(n36168) );
  NAND U37953 ( .A(n36171), .B(mul_pow), .Z(n36170) );
  XOR U37954 ( .A(m[648]), .B(c[648]), .Z(n36171) );
  XOR U37955 ( .A(n36172), .B(n36173), .Z(n36164) );
  ANDN U37956 ( .B(n36174), .A(n32040), .Z(n36172) );
  XNOR U37957 ( .A(\modmult_1/zin[0][646] ), .B(n36175), .Z(n32040) );
  IV U37958 ( .A(n36173), .Z(n36175) );
  XOR U37959 ( .A(n36173), .B(n32041), .Z(n36174) );
  XNOR U37960 ( .A(n36176), .B(n36177), .Z(n32041) );
  ANDN U37961 ( .B(\modmult_1/xin[1023] ), .A(n36178), .Z(n36176) );
  IV U37962 ( .A(n36177), .Z(n36178) );
  XNOR U37963 ( .A(m[647]), .B(n36179), .Z(n36177) );
  NAND U37964 ( .A(n36180), .B(mul_pow), .Z(n36179) );
  XOR U37965 ( .A(m[647]), .B(c[647]), .Z(n36180) );
  XOR U37966 ( .A(n36181), .B(n36182), .Z(n36173) );
  ANDN U37967 ( .B(n36183), .A(n32038), .Z(n36181) );
  XNOR U37968 ( .A(\modmult_1/zin[0][645] ), .B(n36184), .Z(n32038) );
  IV U37969 ( .A(n36182), .Z(n36184) );
  XOR U37970 ( .A(n36182), .B(n32039), .Z(n36183) );
  XNOR U37971 ( .A(n36185), .B(n36186), .Z(n32039) );
  ANDN U37972 ( .B(\modmult_1/xin[1023] ), .A(n36187), .Z(n36185) );
  IV U37973 ( .A(n36186), .Z(n36187) );
  XNOR U37974 ( .A(m[646]), .B(n36188), .Z(n36186) );
  NAND U37975 ( .A(n36189), .B(mul_pow), .Z(n36188) );
  XOR U37976 ( .A(m[646]), .B(c[646]), .Z(n36189) );
  XOR U37977 ( .A(n36190), .B(n36191), .Z(n36182) );
  ANDN U37978 ( .B(n36192), .A(n32036), .Z(n36190) );
  XNOR U37979 ( .A(\modmult_1/zin[0][644] ), .B(n36193), .Z(n32036) );
  IV U37980 ( .A(n36191), .Z(n36193) );
  XOR U37981 ( .A(n36191), .B(n32037), .Z(n36192) );
  XNOR U37982 ( .A(n36194), .B(n36195), .Z(n32037) );
  ANDN U37983 ( .B(\modmult_1/xin[1023] ), .A(n36196), .Z(n36194) );
  IV U37984 ( .A(n36195), .Z(n36196) );
  XNOR U37985 ( .A(m[645]), .B(n36197), .Z(n36195) );
  NAND U37986 ( .A(n36198), .B(mul_pow), .Z(n36197) );
  XOR U37987 ( .A(m[645]), .B(c[645]), .Z(n36198) );
  XOR U37988 ( .A(n36199), .B(n36200), .Z(n36191) );
  ANDN U37989 ( .B(n36201), .A(n32034), .Z(n36199) );
  XNOR U37990 ( .A(\modmult_1/zin[0][643] ), .B(n36202), .Z(n32034) );
  IV U37991 ( .A(n36200), .Z(n36202) );
  XOR U37992 ( .A(n36200), .B(n32035), .Z(n36201) );
  XNOR U37993 ( .A(n36203), .B(n36204), .Z(n32035) );
  ANDN U37994 ( .B(\modmult_1/xin[1023] ), .A(n36205), .Z(n36203) );
  IV U37995 ( .A(n36204), .Z(n36205) );
  XNOR U37996 ( .A(m[644]), .B(n36206), .Z(n36204) );
  NAND U37997 ( .A(n36207), .B(mul_pow), .Z(n36206) );
  XOR U37998 ( .A(m[644]), .B(c[644]), .Z(n36207) );
  XOR U37999 ( .A(n36208), .B(n36209), .Z(n36200) );
  ANDN U38000 ( .B(n36210), .A(n32032), .Z(n36208) );
  XNOR U38001 ( .A(\modmult_1/zin[0][642] ), .B(n36211), .Z(n32032) );
  IV U38002 ( .A(n36209), .Z(n36211) );
  XOR U38003 ( .A(n36209), .B(n32033), .Z(n36210) );
  XNOR U38004 ( .A(n36212), .B(n36213), .Z(n32033) );
  ANDN U38005 ( .B(\modmult_1/xin[1023] ), .A(n36214), .Z(n36212) );
  IV U38006 ( .A(n36213), .Z(n36214) );
  XNOR U38007 ( .A(m[643]), .B(n36215), .Z(n36213) );
  NAND U38008 ( .A(n36216), .B(mul_pow), .Z(n36215) );
  XOR U38009 ( .A(m[643]), .B(c[643]), .Z(n36216) );
  XOR U38010 ( .A(n36217), .B(n36218), .Z(n36209) );
  ANDN U38011 ( .B(n36219), .A(n32030), .Z(n36217) );
  XNOR U38012 ( .A(\modmult_1/zin[0][641] ), .B(n36220), .Z(n32030) );
  IV U38013 ( .A(n36218), .Z(n36220) );
  XOR U38014 ( .A(n36218), .B(n32031), .Z(n36219) );
  XNOR U38015 ( .A(n36221), .B(n36222), .Z(n32031) );
  ANDN U38016 ( .B(\modmult_1/xin[1023] ), .A(n36223), .Z(n36221) );
  IV U38017 ( .A(n36222), .Z(n36223) );
  XNOR U38018 ( .A(m[642]), .B(n36224), .Z(n36222) );
  NAND U38019 ( .A(n36225), .B(mul_pow), .Z(n36224) );
  XOR U38020 ( .A(m[642]), .B(c[642]), .Z(n36225) );
  XOR U38021 ( .A(n36226), .B(n36227), .Z(n36218) );
  ANDN U38022 ( .B(n36228), .A(n32028), .Z(n36226) );
  XNOR U38023 ( .A(\modmult_1/zin[0][640] ), .B(n36229), .Z(n32028) );
  IV U38024 ( .A(n36227), .Z(n36229) );
  XOR U38025 ( .A(n36227), .B(n32029), .Z(n36228) );
  XNOR U38026 ( .A(n36230), .B(n36231), .Z(n32029) );
  ANDN U38027 ( .B(\modmult_1/xin[1023] ), .A(n36232), .Z(n36230) );
  IV U38028 ( .A(n36231), .Z(n36232) );
  XNOR U38029 ( .A(m[641]), .B(n36233), .Z(n36231) );
  NAND U38030 ( .A(n36234), .B(mul_pow), .Z(n36233) );
  XOR U38031 ( .A(m[641]), .B(c[641]), .Z(n36234) );
  XOR U38032 ( .A(n36235), .B(n36236), .Z(n36227) );
  ANDN U38033 ( .B(n36237), .A(n32026), .Z(n36235) );
  XNOR U38034 ( .A(\modmult_1/zin[0][639] ), .B(n36238), .Z(n32026) );
  IV U38035 ( .A(n36236), .Z(n36238) );
  XOR U38036 ( .A(n36236), .B(n32027), .Z(n36237) );
  XNOR U38037 ( .A(n36239), .B(n36240), .Z(n32027) );
  ANDN U38038 ( .B(\modmult_1/xin[1023] ), .A(n36241), .Z(n36239) );
  IV U38039 ( .A(n36240), .Z(n36241) );
  XNOR U38040 ( .A(m[640]), .B(n36242), .Z(n36240) );
  NAND U38041 ( .A(n36243), .B(mul_pow), .Z(n36242) );
  XOR U38042 ( .A(m[640]), .B(c[640]), .Z(n36243) );
  XOR U38043 ( .A(n36244), .B(n36245), .Z(n36236) );
  ANDN U38044 ( .B(n36246), .A(n32024), .Z(n36244) );
  XNOR U38045 ( .A(\modmult_1/zin[0][638] ), .B(n36247), .Z(n32024) );
  IV U38046 ( .A(n36245), .Z(n36247) );
  XOR U38047 ( .A(n36245), .B(n32025), .Z(n36246) );
  XNOR U38048 ( .A(n36248), .B(n36249), .Z(n32025) );
  ANDN U38049 ( .B(\modmult_1/xin[1023] ), .A(n36250), .Z(n36248) );
  IV U38050 ( .A(n36249), .Z(n36250) );
  XNOR U38051 ( .A(m[639]), .B(n36251), .Z(n36249) );
  NAND U38052 ( .A(n36252), .B(mul_pow), .Z(n36251) );
  XOR U38053 ( .A(m[639]), .B(c[639]), .Z(n36252) );
  XOR U38054 ( .A(n36253), .B(n36254), .Z(n36245) );
  ANDN U38055 ( .B(n36255), .A(n32022), .Z(n36253) );
  XNOR U38056 ( .A(\modmult_1/zin[0][637] ), .B(n36256), .Z(n32022) );
  IV U38057 ( .A(n36254), .Z(n36256) );
  XOR U38058 ( .A(n36254), .B(n32023), .Z(n36255) );
  XNOR U38059 ( .A(n36257), .B(n36258), .Z(n32023) );
  ANDN U38060 ( .B(\modmult_1/xin[1023] ), .A(n36259), .Z(n36257) );
  IV U38061 ( .A(n36258), .Z(n36259) );
  XNOR U38062 ( .A(m[638]), .B(n36260), .Z(n36258) );
  NAND U38063 ( .A(n36261), .B(mul_pow), .Z(n36260) );
  XOR U38064 ( .A(m[638]), .B(c[638]), .Z(n36261) );
  XOR U38065 ( .A(n36262), .B(n36263), .Z(n36254) );
  ANDN U38066 ( .B(n36264), .A(n32020), .Z(n36262) );
  XNOR U38067 ( .A(\modmult_1/zin[0][636] ), .B(n36265), .Z(n32020) );
  IV U38068 ( .A(n36263), .Z(n36265) );
  XOR U38069 ( .A(n36263), .B(n32021), .Z(n36264) );
  XNOR U38070 ( .A(n36266), .B(n36267), .Z(n32021) );
  ANDN U38071 ( .B(\modmult_1/xin[1023] ), .A(n36268), .Z(n36266) );
  IV U38072 ( .A(n36267), .Z(n36268) );
  XNOR U38073 ( .A(m[637]), .B(n36269), .Z(n36267) );
  NAND U38074 ( .A(n36270), .B(mul_pow), .Z(n36269) );
  XOR U38075 ( .A(m[637]), .B(c[637]), .Z(n36270) );
  XOR U38076 ( .A(n36271), .B(n36272), .Z(n36263) );
  ANDN U38077 ( .B(n36273), .A(n32018), .Z(n36271) );
  XNOR U38078 ( .A(\modmult_1/zin[0][635] ), .B(n36274), .Z(n32018) );
  IV U38079 ( .A(n36272), .Z(n36274) );
  XOR U38080 ( .A(n36272), .B(n32019), .Z(n36273) );
  XNOR U38081 ( .A(n36275), .B(n36276), .Z(n32019) );
  ANDN U38082 ( .B(\modmult_1/xin[1023] ), .A(n36277), .Z(n36275) );
  IV U38083 ( .A(n36276), .Z(n36277) );
  XNOR U38084 ( .A(m[636]), .B(n36278), .Z(n36276) );
  NAND U38085 ( .A(n36279), .B(mul_pow), .Z(n36278) );
  XOR U38086 ( .A(m[636]), .B(c[636]), .Z(n36279) );
  XOR U38087 ( .A(n36280), .B(n36281), .Z(n36272) );
  ANDN U38088 ( .B(n36282), .A(n32016), .Z(n36280) );
  XNOR U38089 ( .A(\modmult_1/zin[0][634] ), .B(n36283), .Z(n32016) );
  IV U38090 ( .A(n36281), .Z(n36283) );
  XOR U38091 ( .A(n36281), .B(n32017), .Z(n36282) );
  XNOR U38092 ( .A(n36284), .B(n36285), .Z(n32017) );
  ANDN U38093 ( .B(\modmult_1/xin[1023] ), .A(n36286), .Z(n36284) );
  IV U38094 ( .A(n36285), .Z(n36286) );
  XNOR U38095 ( .A(m[635]), .B(n36287), .Z(n36285) );
  NAND U38096 ( .A(n36288), .B(mul_pow), .Z(n36287) );
  XOR U38097 ( .A(m[635]), .B(c[635]), .Z(n36288) );
  XOR U38098 ( .A(n36289), .B(n36290), .Z(n36281) );
  ANDN U38099 ( .B(n36291), .A(n32014), .Z(n36289) );
  XNOR U38100 ( .A(\modmult_1/zin[0][633] ), .B(n36292), .Z(n32014) );
  IV U38101 ( .A(n36290), .Z(n36292) );
  XOR U38102 ( .A(n36290), .B(n32015), .Z(n36291) );
  XNOR U38103 ( .A(n36293), .B(n36294), .Z(n32015) );
  ANDN U38104 ( .B(\modmult_1/xin[1023] ), .A(n36295), .Z(n36293) );
  IV U38105 ( .A(n36294), .Z(n36295) );
  XNOR U38106 ( .A(m[634]), .B(n36296), .Z(n36294) );
  NAND U38107 ( .A(n36297), .B(mul_pow), .Z(n36296) );
  XOR U38108 ( .A(m[634]), .B(c[634]), .Z(n36297) );
  XOR U38109 ( .A(n36298), .B(n36299), .Z(n36290) );
  ANDN U38110 ( .B(n36300), .A(n32012), .Z(n36298) );
  XNOR U38111 ( .A(\modmult_1/zin[0][632] ), .B(n36301), .Z(n32012) );
  IV U38112 ( .A(n36299), .Z(n36301) );
  XOR U38113 ( .A(n36299), .B(n32013), .Z(n36300) );
  XNOR U38114 ( .A(n36302), .B(n36303), .Z(n32013) );
  ANDN U38115 ( .B(\modmult_1/xin[1023] ), .A(n36304), .Z(n36302) );
  IV U38116 ( .A(n36303), .Z(n36304) );
  XNOR U38117 ( .A(m[633]), .B(n36305), .Z(n36303) );
  NAND U38118 ( .A(n36306), .B(mul_pow), .Z(n36305) );
  XOR U38119 ( .A(m[633]), .B(c[633]), .Z(n36306) );
  XOR U38120 ( .A(n36307), .B(n36308), .Z(n36299) );
  ANDN U38121 ( .B(n36309), .A(n32010), .Z(n36307) );
  XNOR U38122 ( .A(\modmult_1/zin[0][631] ), .B(n36310), .Z(n32010) );
  IV U38123 ( .A(n36308), .Z(n36310) );
  XOR U38124 ( .A(n36308), .B(n32011), .Z(n36309) );
  XNOR U38125 ( .A(n36311), .B(n36312), .Z(n32011) );
  ANDN U38126 ( .B(\modmult_1/xin[1023] ), .A(n36313), .Z(n36311) );
  IV U38127 ( .A(n36312), .Z(n36313) );
  XNOR U38128 ( .A(m[632]), .B(n36314), .Z(n36312) );
  NAND U38129 ( .A(n36315), .B(mul_pow), .Z(n36314) );
  XOR U38130 ( .A(m[632]), .B(c[632]), .Z(n36315) );
  XOR U38131 ( .A(n36316), .B(n36317), .Z(n36308) );
  ANDN U38132 ( .B(n36318), .A(n32008), .Z(n36316) );
  XNOR U38133 ( .A(\modmult_1/zin[0][630] ), .B(n36319), .Z(n32008) );
  IV U38134 ( .A(n36317), .Z(n36319) );
  XOR U38135 ( .A(n36317), .B(n32009), .Z(n36318) );
  XNOR U38136 ( .A(n36320), .B(n36321), .Z(n32009) );
  ANDN U38137 ( .B(\modmult_1/xin[1023] ), .A(n36322), .Z(n36320) );
  IV U38138 ( .A(n36321), .Z(n36322) );
  XNOR U38139 ( .A(m[631]), .B(n36323), .Z(n36321) );
  NAND U38140 ( .A(n36324), .B(mul_pow), .Z(n36323) );
  XOR U38141 ( .A(m[631]), .B(c[631]), .Z(n36324) );
  XOR U38142 ( .A(n36325), .B(n36326), .Z(n36317) );
  ANDN U38143 ( .B(n36327), .A(n32006), .Z(n36325) );
  XNOR U38144 ( .A(\modmult_1/zin[0][629] ), .B(n36328), .Z(n32006) );
  IV U38145 ( .A(n36326), .Z(n36328) );
  XOR U38146 ( .A(n36326), .B(n32007), .Z(n36327) );
  XNOR U38147 ( .A(n36329), .B(n36330), .Z(n32007) );
  ANDN U38148 ( .B(\modmult_1/xin[1023] ), .A(n36331), .Z(n36329) );
  IV U38149 ( .A(n36330), .Z(n36331) );
  XNOR U38150 ( .A(m[630]), .B(n36332), .Z(n36330) );
  NAND U38151 ( .A(n36333), .B(mul_pow), .Z(n36332) );
  XOR U38152 ( .A(m[630]), .B(c[630]), .Z(n36333) );
  XOR U38153 ( .A(n36334), .B(n36335), .Z(n36326) );
  ANDN U38154 ( .B(n36336), .A(n32004), .Z(n36334) );
  XNOR U38155 ( .A(\modmult_1/zin[0][628] ), .B(n36337), .Z(n32004) );
  IV U38156 ( .A(n36335), .Z(n36337) );
  XOR U38157 ( .A(n36335), .B(n32005), .Z(n36336) );
  XNOR U38158 ( .A(n36338), .B(n36339), .Z(n32005) );
  ANDN U38159 ( .B(\modmult_1/xin[1023] ), .A(n36340), .Z(n36338) );
  IV U38160 ( .A(n36339), .Z(n36340) );
  XNOR U38161 ( .A(m[629]), .B(n36341), .Z(n36339) );
  NAND U38162 ( .A(n36342), .B(mul_pow), .Z(n36341) );
  XOR U38163 ( .A(m[629]), .B(c[629]), .Z(n36342) );
  XOR U38164 ( .A(n36343), .B(n36344), .Z(n36335) );
  ANDN U38165 ( .B(n36345), .A(n32002), .Z(n36343) );
  XNOR U38166 ( .A(\modmult_1/zin[0][627] ), .B(n36346), .Z(n32002) );
  IV U38167 ( .A(n36344), .Z(n36346) );
  XOR U38168 ( .A(n36344), .B(n32003), .Z(n36345) );
  XNOR U38169 ( .A(n36347), .B(n36348), .Z(n32003) );
  ANDN U38170 ( .B(\modmult_1/xin[1023] ), .A(n36349), .Z(n36347) );
  IV U38171 ( .A(n36348), .Z(n36349) );
  XNOR U38172 ( .A(m[628]), .B(n36350), .Z(n36348) );
  NAND U38173 ( .A(n36351), .B(mul_pow), .Z(n36350) );
  XOR U38174 ( .A(m[628]), .B(c[628]), .Z(n36351) );
  XOR U38175 ( .A(n36352), .B(n36353), .Z(n36344) );
  ANDN U38176 ( .B(n36354), .A(n32000), .Z(n36352) );
  XNOR U38177 ( .A(\modmult_1/zin[0][626] ), .B(n36355), .Z(n32000) );
  IV U38178 ( .A(n36353), .Z(n36355) );
  XOR U38179 ( .A(n36353), .B(n32001), .Z(n36354) );
  XNOR U38180 ( .A(n36356), .B(n36357), .Z(n32001) );
  ANDN U38181 ( .B(\modmult_1/xin[1023] ), .A(n36358), .Z(n36356) );
  IV U38182 ( .A(n36357), .Z(n36358) );
  XNOR U38183 ( .A(m[627]), .B(n36359), .Z(n36357) );
  NAND U38184 ( .A(n36360), .B(mul_pow), .Z(n36359) );
  XOR U38185 ( .A(m[627]), .B(c[627]), .Z(n36360) );
  XOR U38186 ( .A(n36361), .B(n36362), .Z(n36353) );
  ANDN U38187 ( .B(n36363), .A(n31998), .Z(n36361) );
  XNOR U38188 ( .A(\modmult_1/zin[0][625] ), .B(n36364), .Z(n31998) );
  IV U38189 ( .A(n36362), .Z(n36364) );
  XOR U38190 ( .A(n36362), .B(n31999), .Z(n36363) );
  XNOR U38191 ( .A(n36365), .B(n36366), .Z(n31999) );
  ANDN U38192 ( .B(\modmult_1/xin[1023] ), .A(n36367), .Z(n36365) );
  IV U38193 ( .A(n36366), .Z(n36367) );
  XNOR U38194 ( .A(m[626]), .B(n36368), .Z(n36366) );
  NAND U38195 ( .A(n36369), .B(mul_pow), .Z(n36368) );
  XOR U38196 ( .A(m[626]), .B(c[626]), .Z(n36369) );
  XOR U38197 ( .A(n36370), .B(n36371), .Z(n36362) );
  ANDN U38198 ( .B(n36372), .A(n31996), .Z(n36370) );
  XNOR U38199 ( .A(\modmult_1/zin[0][624] ), .B(n36373), .Z(n31996) );
  IV U38200 ( .A(n36371), .Z(n36373) );
  XOR U38201 ( .A(n36371), .B(n31997), .Z(n36372) );
  XNOR U38202 ( .A(n36374), .B(n36375), .Z(n31997) );
  ANDN U38203 ( .B(\modmult_1/xin[1023] ), .A(n36376), .Z(n36374) );
  IV U38204 ( .A(n36375), .Z(n36376) );
  XNOR U38205 ( .A(m[625]), .B(n36377), .Z(n36375) );
  NAND U38206 ( .A(n36378), .B(mul_pow), .Z(n36377) );
  XOR U38207 ( .A(m[625]), .B(c[625]), .Z(n36378) );
  XOR U38208 ( .A(n36379), .B(n36380), .Z(n36371) );
  ANDN U38209 ( .B(n36381), .A(n31994), .Z(n36379) );
  XNOR U38210 ( .A(\modmult_1/zin[0][623] ), .B(n36382), .Z(n31994) );
  IV U38211 ( .A(n36380), .Z(n36382) );
  XOR U38212 ( .A(n36380), .B(n31995), .Z(n36381) );
  XNOR U38213 ( .A(n36383), .B(n36384), .Z(n31995) );
  ANDN U38214 ( .B(\modmult_1/xin[1023] ), .A(n36385), .Z(n36383) );
  IV U38215 ( .A(n36384), .Z(n36385) );
  XNOR U38216 ( .A(m[624]), .B(n36386), .Z(n36384) );
  NAND U38217 ( .A(n36387), .B(mul_pow), .Z(n36386) );
  XOR U38218 ( .A(m[624]), .B(c[624]), .Z(n36387) );
  XOR U38219 ( .A(n36388), .B(n36389), .Z(n36380) );
  ANDN U38220 ( .B(n36390), .A(n31992), .Z(n36388) );
  XNOR U38221 ( .A(\modmult_1/zin[0][622] ), .B(n36391), .Z(n31992) );
  IV U38222 ( .A(n36389), .Z(n36391) );
  XOR U38223 ( .A(n36389), .B(n31993), .Z(n36390) );
  XNOR U38224 ( .A(n36392), .B(n36393), .Z(n31993) );
  ANDN U38225 ( .B(\modmult_1/xin[1023] ), .A(n36394), .Z(n36392) );
  IV U38226 ( .A(n36393), .Z(n36394) );
  XNOR U38227 ( .A(m[623]), .B(n36395), .Z(n36393) );
  NAND U38228 ( .A(n36396), .B(mul_pow), .Z(n36395) );
  XOR U38229 ( .A(m[623]), .B(c[623]), .Z(n36396) );
  XOR U38230 ( .A(n36397), .B(n36398), .Z(n36389) );
  ANDN U38231 ( .B(n36399), .A(n31990), .Z(n36397) );
  XNOR U38232 ( .A(\modmult_1/zin[0][621] ), .B(n36400), .Z(n31990) );
  IV U38233 ( .A(n36398), .Z(n36400) );
  XOR U38234 ( .A(n36398), .B(n31991), .Z(n36399) );
  XNOR U38235 ( .A(n36401), .B(n36402), .Z(n31991) );
  ANDN U38236 ( .B(\modmult_1/xin[1023] ), .A(n36403), .Z(n36401) );
  IV U38237 ( .A(n36402), .Z(n36403) );
  XNOR U38238 ( .A(m[622]), .B(n36404), .Z(n36402) );
  NAND U38239 ( .A(n36405), .B(mul_pow), .Z(n36404) );
  XOR U38240 ( .A(m[622]), .B(c[622]), .Z(n36405) );
  XOR U38241 ( .A(n36406), .B(n36407), .Z(n36398) );
  ANDN U38242 ( .B(n36408), .A(n31988), .Z(n36406) );
  XNOR U38243 ( .A(\modmult_1/zin[0][620] ), .B(n36409), .Z(n31988) );
  IV U38244 ( .A(n36407), .Z(n36409) );
  XOR U38245 ( .A(n36407), .B(n31989), .Z(n36408) );
  XNOR U38246 ( .A(n36410), .B(n36411), .Z(n31989) );
  ANDN U38247 ( .B(\modmult_1/xin[1023] ), .A(n36412), .Z(n36410) );
  IV U38248 ( .A(n36411), .Z(n36412) );
  XNOR U38249 ( .A(m[621]), .B(n36413), .Z(n36411) );
  NAND U38250 ( .A(n36414), .B(mul_pow), .Z(n36413) );
  XOR U38251 ( .A(m[621]), .B(c[621]), .Z(n36414) );
  XOR U38252 ( .A(n36415), .B(n36416), .Z(n36407) );
  ANDN U38253 ( .B(n36417), .A(n31986), .Z(n36415) );
  XNOR U38254 ( .A(\modmult_1/zin[0][619] ), .B(n36418), .Z(n31986) );
  IV U38255 ( .A(n36416), .Z(n36418) );
  XOR U38256 ( .A(n36416), .B(n31987), .Z(n36417) );
  XNOR U38257 ( .A(n36419), .B(n36420), .Z(n31987) );
  ANDN U38258 ( .B(\modmult_1/xin[1023] ), .A(n36421), .Z(n36419) );
  IV U38259 ( .A(n36420), .Z(n36421) );
  XNOR U38260 ( .A(m[620]), .B(n36422), .Z(n36420) );
  NAND U38261 ( .A(n36423), .B(mul_pow), .Z(n36422) );
  XOR U38262 ( .A(m[620]), .B(c[620]), .Z(n36423) );
  XOR U38263 ( .A(n36424), .B(n36425), .Z(n36416) );
  ANDN U38264 ( .B(n36426), .A(n31984), .Z(n36424) );
  XNOR U38265 ( .A(\modmult_1/zin[0][618] ), .B(n36427), .Z(n31984) );
  IV U38266 ( .A(n36425), .Z(n36427) );
  XOR U38267 ( .A(n36425), .B(n31985), .Z(n36426) );
  XNOR U38268 ( .A(n36428), .B(n36429), .Z(n31985) );
  ANDN U38269 ( .B(\modmult_1/xin[1023] ), .A(n36430), .Z(n36428) );
  IV U38270 ( .A(n36429), .Z(n36430) );
  XNOR U38271 ( .A(m[619]), .B(n36431), .Z(n36429) );
  NAND U38272 ( .A(n36432), .B(mul_pow), .Z(n36431) );
  XOR U38273 ( .A(m[619]), .B(c[619]), .Z(n36432) );
  XOR U38274 ( .A(n36433), .B(n36434), .Z(n36425) );
  ANDN U38275 ( .B(n36435), .A(n31982), .Z(n36433) );
  XNOR U38276 ( .A(\modmult_1/zin[0][617] ), .B(n36436), .Z(n31982) );
  IV U38277 ( .A(n36434), .Z(n36436) );
  XOR U38278 ( .A(n36434), .B(n31983), .Z(n36435) );
  XNOR U38279 ( .A(n36437), .B(n36438), .Z(n31983) );
  ANDN U38280 ( .B(\modmult_1/xin[1023] ), .A(n36439), .Z(n36437) );
  IV U38281 ( .A(n36438), .Z(n36439) );
  XNOR U38282 ( .A(m[618]), .B(n36440), .Z(n36438) );
  NAND U38283 ( .A(n36441), .B(mul_pow), .Z(n36440) );
  XOR U38284 ( .A(m[618]), .B(c[618]), .Z(n36441) );
  XOR U38285 ( .A(n36442), .B(n36443), .Z(n36434) );
  ANDN U38286 ( .B(n36444), .A(n31980), .Z(n36442) );
  XNOR U38287 ( .A(\modmult_1/zin[0][616] ), .B(n36445), .Z(n31980) );
  IV U38288 ( .A(n36443), .Z(n36445) );
  XOR U38289 ( .A(n36443), .B(n31981), .Z(n36444) );
  XNOR U38290 ( .A(n36446), .B(n36447), .Z(n31981) );
  ANDN U38291 ( .B(\modmult_1/xin[1023] ), .A(n36448), .Z(n36446) );
  IV U38292 ( .A(n36447), .Z(n36448) );
  XNOR U38293 ( .A(m[617]), .B(n36449), .Z(n36447) );
  NAND U38294 ( .A(n36450), .B(mul_pow), .Z(n36449) );
  XOR U38295 ( .A(m[617]), .B(c[617]), .Z(n36450) );
  XOR U38296 ( .A(n36451), .B(n36452), .Z(n36443) );
  ANDN U38297 ( .B(n36453), .A(n31978), .Z(n36451) );
  XNOR U38298 ( .A(\modmult_1/zin[0][615] ), .B(n36454), .Z(n31978) );
  IV U38299 ( .A(n36452), .Z(n36454) );
  XOR U38300 ( .A(n36452), .B(n31979), .Z(n36453) );
  XNOR U38301 ( .A(n36455), .B(n36456), .Z(n31979) );
  ANDN U38302 ( .B(\modmult_1/xin[1023] ), .A(n36457), .Z(n36455) );
  IV U38303 ( .A(n36456), .Z(n36457) );
  XNOR U38304 ( .A(m[616]), .B(n36458), .Z(n36456) );
  NAND U38305 ( .A(n36459), .B(mul_pow), .Z(n36458) );
  XOR U38306 ( .A(m[616]), .B(c[616]), .Z(n36459) );
  XOR U38307 ( .A(n36460), .B(n36461), .Z(n36452) );
  ANDN U38308 ( .B(n36462), .A(n31976), .Z(n36460) );
  XNOR U38309 ( .A(\modmult_1/zin[0][614] ), .B(n36463), .Z(n31976) );
  IV U38310 ( .A(n36461), .Z(n36463) );
  XOR U38311 ( .A(n36461), .B(n31977), .Z(n36462) );
  XNOR U38312 ( .A(n36464), .B(n36465), .Z(n31977) );
  ANDN U38313 ( .B(\modmult_1/xin[1023] ), .A(n36466), .Z(n36464) );
  IV U38314 ( .A(n36465), .Z(n36466) );
  XNOR U38315 ( .A(m[615]), .B(n36467), .Z(n36465) );
  NAND U38316 ( .A(n36468), .B(mul_pow), .Z(n36467) );
  XOR U38317 ( .A(m[615]), .B(c[615]), .Z(n36468) );
  XOR U38318 ( .A(n36469), .B(n36470), .Z(n36461) );
  ANDN U38319 ( .B(n36471), .A(n31974), .Z(n36469) );
  XNOR U38320 ( .A(\modmult_1/zin[0][613] ), .B(n36472), .Z(n31974) );
  IV U38321 ( .A(n36470), .Z(n36472) );
  XOR U38322 ( .A(n36470), .B(n31975), .Z(n36471) );
  XNOR U38323 ( .A(n36473), .B(n36474), .Z(n31975) );
  ANDN U38324 ( .B(\modmult_1/xin[1023] ), .A(n36475), .Z(n36473) );
  IV U38325 ( .A(n36474), .Z(n36475) );
  XNOR U38326 ( .A(m[614]), .B(n36476), .Z(n36474) );
  NAND U38327 ( .A(n36477), .B(mul_pow), .Z(n36476) );
  XOR U38328 ( .A(m[614]), .B(c[614]), .Z(n36477) );
  XOR U38329 ( .A(n36478), .B(n36479), .Z(n36470) );
  ANDN U38330 ( .B(n36480), .A(n31972), .Z(n36478) );
  XNOR U38331 ( .A(\modmult_1/zin[0][612] ), .B(n36481), .Z(n31972) );
  IV U38332 ( .A(n36479), .Z(n36481) );
  XOR U38333 ( .A(n36479), .B(n31973), .Z(n36480) );
  XNOR U38334 ( .A(n36482), .B(n36483), .Z(n31973) );
  ANDN U38335 ( .B(\modmult_1/xin[1023] ), .A(n36484), .Z(n36482) );
  IV U38336 ( .A(n36483), .Z(n36484) );
  XNOR U38337 ( .A(m[613]), .B(n36485), .Z(n36483) );
  NAND U38338 ( .A(n36486), .B(mul_pow), .Z(n36485) );
  XOR U38339 ( .A(m[613]), .B(c[613]), .Z(n36486) );
  XOR U38340 ( .A(n36487), .B(n36488), .Z(n36479) );
  ANDN U38341 ( .B(n36489), .A(n31970), .Z(n36487) );
  XNOR U38342 ( .A(\modmult_1/zin[0][611] ), .B(n36490), .Z(n31970) );
  IV U38343 ( .A(n36488), .Z(n36490) );
  XOR U38344 ( .A(n36488), .B(n31971), .Z(n36489) );
  XNOR U38345 ( .A(n36491), .B(n36492), .Z(n31971) );
  ANDN U38346 ( .B(\modmult_1/xin[1023] ), .A(n36493), .Z(n36491) );
  IV U38347 ( .A(n36492), .Z(n36493) );
  XNOR U38348 ( .A(m[612]), .B(n36494), .Z(n36492) );
  NAND U38349 ( .A(n36495), .B(mul_pow), .Z(n36494) );
  XOR U38350 ( .A(m[612]), .B(c[612]), .Z(n36495) );
  XOR U38351 ( .A(n36496), .B(n36497), .Z(n36488) );
  ANDN U38352 ( .B(n36498), .A(n31968), .Z(n36496) );
  XNOR U38353 ( .A(\modmult_1/zin[0][610] ), .B(n36499), .Z(n31968) );
  IV U38354 ( .A(n36497), .Z(n36499) );
  XOR U38355 ( .A(n36497), .B(n31969), .Z(n36498) );
  XNOR U38356 ( .A(n36500), .B(n36501), .Z(n31969) );
  ANDN U38357 ( .B(\modmult_1/xin[1023] ), .A(n36502), .Z(n36500) );
  IV U38358 ( .A(n36501), .Z(n36502) );
  XNOR U38359 ( .A(m[611]), .B(n36503), .Z(n36501) );
  NAND U38360 ( .A(n36504), .B(mul_pow), .Z(n36503) );
  XOR U38361 ( .A(m[611]), .B(c[611]), .Z(n36504) );
  XOR U38362 ( .A(n36505), .B(n36506), .Z(n36497) );
  ANDN U38363 ( .B(n36507), .A(n31966), .Z(n36505) );
  XNOR U38364 ( .A(\modmult_1/zin[0][609] ), .B(n36508), .Z(n31966) );
  IV U38365 ( .A(n36506), .Z(n36508) );
  XOR U38366 ( .A(n36506), .B(n31967), .Z(n36507) );
  XNOR U38367 ( .A(n36509), .B(n36510), .Z(n31967) );
  ANDN U38368 ( .B(\modmult_1/xin[1023] ), .A(n36511), .Z(n36509) );
  IV U38369 ( .A(n36510), .Z(n36511) );
  XNOR U38370 ( .A(m[610]), .B(n36512), .Z(n36510) );
  NAND U38371 ( .A(n36513), .B(mul_pow), .Z(n36512) );
  XOR U38372 ( .A(m[610]), .B(c[610]), .Z(n36513) );
  XOR U38373 ( .A(n36514), .B(n36515), .Z(n36506) );
  ANDN U38374 ( .B(n36516), .A(n31964), .Z(n36514) );
  XNOR U38375 ( .A(\modmult_1/zin[0][608] ), .B(n36517), .Z(n31964) );
  IV U38376 ( .A(n36515), .Z(n36517) );
  XOR U38377 ( .A(n36515), .B(n31965), .Z(n36516) );
  XNOR U38378 ( .A(n36518), .B(n36519), .Z(n31965) );
  ANDN U38379 ( .B(\modmult_1/xin[1023] ), .A(n36520), .Z(n36518) );
  IV U38380 ( .A(n36519), .Z(n36520) );
  XNOR U38381 ( .A(m[609]), .B(n36521), .Z(n36519) );
  NAND U38382 ( .A(n36522), .B(mul_pow), .Z(n36521) );
  XOR U38383 ( .A(m[609]), .B(c[609]), .Z(n36522) );
  XOR U38384 ( .A(n36523), .B(n36524), .Z(n36515) );
  ANDN U38385 ( .B(n36525), .A(n31962), .Z(n36523) );
  XNOR U38386 ( .A(\modmult_1/zin[0][607] ), .B(n36526), .Z(n31962) );
  IV U38387 ( .A(n36524), .Z(n36526) );
  XOR U38388 ( .A(n36524), .B(n31963), .Z(n36525) );
  XNOR U38389 ( .A(n36527), .B(n36528), .Z(n31963) );
  ANDN U38390 ( .B(\modmult_1/xin[1023] ), .A(n36529), .Z(n36527) );
  IV U38391 ( .A(n36528), .Z(n36529) );
  XNOR U38392 ( .A(m[608]), .B(n36530), .Z(n36528) );
  NAND U38393 ( .A(n36531), .B(mul_pow), .Z(n36530) );
  XOR U38394 ( .A(m[608]), .B(c[608]), .Z(n36531) );
  XOR U38395 ( .A(n36532), .B(n36533), .Z(n36524) );
  ANDN U38396 ( .B(n36534), .A(n31960), .Z(n36532) );
  XNOR U38397 ( .A(\modmult_1/zin[0][606] ), .B(n36535), .Z(n31960) );
  IV U38398 ( .A(n36533), .Z(n36535) );
  XOR U38399 ( .A(n36533), .B(n31961), .Z(n36534) );
  XNOR U38400 ( .A(n36536), .B(n36537), .Z(n31961) );
  ANDN U38401 ( .B(\modmult_1/xin[1023] ), .A(n36538), .Z(n36536) );
  IV U38402 ( .A(n36537), .Z(n36538) );
  XNOR U38403 ( .A(m[607]), .B(n36539), .Z(n36537) );
  NAND U38404 ( .A(n36540), .B(mul_pow), .Z(n36539) );
  XOR U38405 ( .A(m[607]), .B(c[607]), .Z(n36540) );
  XOR U38406 ( .A(n36541), .B(n36542), .Z(n36533) );
  ANDN U38407 ( .B(n36543), .A(n31958), .Z(n36541) );
  XNOR U38408 ( .A(\modmult_1/zin[0][605] ), .B(n36544), .Z(n31958) );
  IV U38409 ( .A(n36542), .Z(n36544) );
  XOR U38410 ( .A(n36542), .B(n31959), .Z(n36543) );
  XNOR U38411 ( .A(n36545), .B(n36546), .Z(n31959) );
  ANDN U38412 ( .B(\modmult_1/xin[1023] ), .A(n36547), .Z(n36545) );
  IV U38413 ( .A(n36546), .Z(n36547) );
  XNOR U38414 ( .A(m[606]), .B(n36548), .Z(n36546) );
  NAND U38415 ( .A(n36549), .B(mul_pow), .Z(n36548) );
  XOR U38416 ( .A(m[606]), .B(c[606]), .Z(n36549) );
  XOR U38417 ( .A(n36550), .B(n36551), .Z(n36542) );
  ANDN U38418 ( .B(n36552), .A(n31956), .Z(n36550) );
  XNOR U38419 ( .A(\modmult_1/zin[0][604] ), .B(n36553), .Z(n31956) );
  IV U38420 ( .A(n36551), .Z(n36553) );
  XOR U38421 ( .A(n36551), .B(n31957), .Z(n36552) );
  XNOR U38422 ( .A(n36554), .B(n36555), .Z(n31957) );
  ANDN U38423 ( .B(\modmult_1/xin[1023] ), .A(n36556), .Z(n36554) );
  IV U38424 ( .A(n36555), .Z(n36556) );
  XNOR U38425 ( .A(m[605]), .B(n36557), .Z(n36555) );
  NAND U38426 ( .A(n36558), .B(mul_pow), .Z(n36557) );
  XOR U38427 ( .A(m[605]), .B(c[605]), .Z(n36558) );
  XOR U38428 ( .A(n36559), .B(n36560), .Z(n36551) );
  ANDN U38429 ( .B(n36561), .A(n31954), .Z(n36559) );
  XNOR U38430 ( .A(\modmult_1/zin[0][603] ), .B(n36562), .Z(n31954) );
  IV U38431 ( .A(n36560), .Z(n36562) );
  XOR U38432 ( .A(n36560), .B(n31955), .Z(n36561) );
  XNOR U38433 ( .A(n36563), .B(n36564), .Z(n31955) );
  ANDN U38434 ( .B(\modmult_1/xin[1023] ), .A(n36565), .Z(n36563) );
  IV U38435 ( .A(n36564), .Z(n36565) );
  XNOR U38436 ( .A(m[604]), .B(n36566), .Z(n36564) );
  NAND U38437 ( .A(n36567), .B(mul_pow), .Z(n36566) );
  XOR U38438 ( .A(m[604]), .B(c[604]), .Z(n36567) );
  XOR U38439 ( .A(n36568), .B(n36569), .Z(n36560) );
  ANDN U38440 ( .B(n36570), .A(n31952), .Z(n36568) );
  XNOR U38441 ( .A(\modmult_1/zin[0][602] ), .B(n36571), .Z(n31952) );
  IV U38442 ( .A(n36569), .Z(n36571) );
  XOR U38443 ( .A(n36569), .B(n31953), .Z(n36570) );
  XNOR U38444 ( .A(n36572), .B(n36573), .Z(n31953) );
  ANDN U38445 ( .B(\modmult_1/xin[1023] ), .A(n36574), .Z(n36572) );
  IV U38446 ( .A(n36573), .Z(n36574) );
  XNOR U38447 ( .A(m[603]), .B(n36575), .Z(n36573) );
  NAND U38448 ( .A(n36576), .B(mul_pow), .Z(n36575) );
  XOR U38449 ( .A(m[603]), .B(c[603]), .Z(n36576) );
  XOR U38450 ( .A(n36577), .B(n36578), .Z(n36569) );
  ANDN U38451 ( .B(n36579), .A(n31950), .Z(n36577) );
  XNOR U38452 ( .A(\modmult_1/zin[0][601] ), .B(n36580), .Z(n31950) );
  IV U38453 ( .A(n36578), .Z(n36580) );
  XOR U38454 ( .A(n36578), .B(n31951), .Z(n36579) );
  XNOR U38455 ( .A(n36581), .B(n36582), .Z(n31951) );
  ANDN U38456 ( .B(\modmult_1/xin[1023] ), .A(n36583), .Z(n36581) );
  IV U38457 ( .A(n36582), .Z(n36583) );
  XNOR U38458 ( .A(m[602]), .B(n36584), .Z(n36582) );
  NAND U38459 ( .A(n36585), .B(mul_pow), .Z(n36584) );
  XOR U38460 ( .A(m[602]), .B(c[602]), .Z(n36585) );
  XOR U38461 ( .A(n36586), .B(n36587), .Z(n36578) );
  ANDN U38462 ( .B(n36588), .A(n31948), .Z(n36586) );
  XNOR U38463 ( .A(\modmult_1/zin[0][600] ), .B(n36589), .Z(n31948) );
  IV U38464 ( .A(n36587), .Z(n36589) );
  XOR U38465 ( .A(n36587), .B(n31949), .Z(n36588) );
  XNOR U38466 ( .A(n36590), .B(n36591), .Z(n31949) );
  ANDN U38467 ( .B(\modmult_1/xin[1023] ), .A(n36592), .Z(n36590) );
  IV U38468 ( .A(n36591), .Z(n36592) );
  XNOR U38469 ( .A(m[601]), .B(n36593), .Z(n36591) );
  NAND U38470 ( .A(n36594), .B(mul_pow), .Z(n36593) );
  XOR U38471 ( .A(m[601]), .B(c[601]), .Z(n36594) );
  XOR U38472 ( .A(n36595), .B(n36596), .Z(n36587) );
  ANDN U38473 ( .B(n36597), .A(n31946), .Z(n36595) );
  XNOR U38474 ( .A(\modmult_1/zin[0][599] ), .B(n36598), .Z(n31946) );
  IV U38475 ( .A(n36596), .Z(n36598) );
  XOR U38476 ( .A(n36596), .B(n31947), .Z(n36597) );
  XNOR U38477 ( .A(n36599), .B(n36600), .Z(n31947) );
  ANDN U38478 ( .B(\modmult_1/xin[1023] ), .A(n36601), .Z(n36599) );
  IV U38479 ( .A(n36600), .Z(n36601) );
  XNOR U38480 ( .A(m[600]), .B(n36602), .Z(n36600) );
  NAND U38481 ( .A(n36603), .B(mul_pow), .Z(n36602) );
  XOR U38482 ( .A(m[600]), .B(c[600]), .Z(n36603) );
  XOR U38483 ( .A(n36604), .B(n36605), .Z(n36596) );
  ANDN U38484 ( .B(n36606), .A(n31944), .Z(n36604) );
  XNOR U38485 ( .A(\modmult_1/zin[0][598] ), .B(n36607), .Z(n31944) );
  IV U38486 ( .A(n36605), .Z(n36607) );
  XOR U38487 ( .A(n36605), .B(n31945), .Z(n36606) );
  XNOR U38488 ( .A(n36608), .B(n36609), .Z(n31945) );
  ANDN U38489 ( .B(\modmult_1/xin[1023] ), .A(n36610), .Z(n36608) );
  IV U38490 ( .A(n36609), .Z(n36610) );
  XNOR U38491 ( .A(m[599]), .B(n36611), .Z(n36609) );
  NAND U38492 ( .A(n36612), .B(mul_pow), .Z(n36611) );
  XOR U38493 ( .A(m[599]), .B(c[599]), .Z(n36612) );
  XOR U38494 ( .A(n36613), .B(n36614), .Z(n36605) );
  ANDN U38495 ( .B(n36615), .A(n31942), .Z(n36613) );
  XNOR U38496 ( .A(\modmult_1/zin[0][597] ), .B(n36616), .Z(n31942) );
  IV U38497 ( .A(n36614), .Z(n36616) );
  XOR U38498 ( .A(n36614), .B(n31943), .Z(n36615) );
  XNOR U38499 ( .A(n36617), .B(n36618), .Z(n31943) );
  ANDN U38500 ( .B(\modmult_1/xin[1023] ), .A(n36619), .Z(n36617) );
  IV U38501 ( .A(n36618), .Z(n36619) );
  XNOR U38502 ( .A(m[598]), .B(n36620), .Z(n36618) );
  NAND U38503 ( .A(n36621), .B(mul_pow), .Z(n36620) );
  XOR U38504 ( .A(m[598]), .B(c[598]), .Z(n36621) );
  XOR U38505 ( .A(n36622), .B(n36623), .Z(n36614) );
  ANDN U38506 ( .B(n36624), .A(n31940), .Z(n36622) );
  XNOR U38507 ( .A(\modmult_1/zin[0][596] ), .B(n36625), .Z(n31940) );
  IV U38508 ( .A(n36623), .Z(n36625) );
  XOR U38509 ( .A(n36623), .B(n31941), .Z(n36624) );
  XNOR U38510 ( .A(n36626), .B(n36627), .Z(n31941) );
  ANDN U38511 ( .B(\modmult_1/xin[1023] ), .A(n36628), .Z(n36626) );
  IV U38512 ( .A(n36627), .Z(n36628) );
  XNOR U38513 ( .A(m[597]), .B(n36629), .Z(n36627) );
  NAND U38514 ( .A(n36630), .B(mul_pow), .Z(n36629) );
  XOR U38515 ( .A(m[597]), .B(c[597]), .Z(n36630) );
  XOR U38516 ( .A(n36631), .B(n36632), .Z(n36623) );
  ANDN U38517 ( .B(n36633), .A(n31938), .Z(n36631) );
  XNOR U38518 ( .A(\modmult_1/zin[0][595] ), .B(n36634), .Z(n31938) );
  IV U38519 ( .A(n36632), .Z(n36634) );
  XOR U38520 ( .A(n36632), .B(n31939), .Z(n36633) );
  XNOR U38521 ( .A(n36635), .B(n36636), .Z(n31939) );
  ANDN U38522 ( .B(\modmult_1/xin[1023] ), .A(n36637), .Z(n36635) );
  IV U38523 ( .A(n36636), .Z(n36637) );
  XNOR U38524 ( .A(m[596]), .B(n36638), .Z(n36636) );
  NAND U38525 ( .A(n36639), .B(mul_pow), .Z(n36638) );
  XOR U38526 ( .A(m[596]), .B(c[596]), .Z(n36639) );
  XOR U38527 ( .A(n36640), .B(n36641), .Z(n36632) );
  ANDN U38528 ( .B(n36642), .A(n31936), .Z(n36640) );
  XNOR U38529 ( .A(\modmult_1/zin[0][594] ), .B(n36643), .Z(n31936) );
  IV U38530 ( .A(n36641), .Z(n36643) );
  XOR U38531 ( .A(n36641), .B(n31937), .Z(n36642) );
  XNOR U38532 ( .A(n36644), .B(n36645), .Z(n31937) );
  ANDN U38533 ( .B(\modmult_1/xin[1023] ), .A(n36646), .Z(n36644) );
  IV U38534 ( .A(n36645), .Z(n36646) );
  XNOR U38535 ( .A(m[595]), .B(n36647), .Z(n36645) );
  NAND U38536 ( .A(n36648), .B(mul_pow), .Z(n36647) );
  XOR U38537 ( .A(m[595]), .B(c[595]), .Z(n36648) );
  XOR U38538 ( .A(n36649), .B(n36650), .Z(n36641) );
  ANDN U38539 ( .B(n36651), .A(n31934), .Z(n36649) );
  XNOR U38540 ( .A(\modmult_1/zin[0][593] ), .B(n36652), .Z(n31934) );
  IV U38541 ( .A(n36650), .Z(n36652) );
  XOR U38542 ( .A(n36650), .B(n31935), .Z(n36651) );
  XNOR U38543 ( .A(n36653), .B(n36654), .Z(n31935) );
  ANDN U38544 ( .B(\modmult_1/xin[1023] ), .A(n36655), .Z(n36653) );
  IV U38545 ( .A(n36654), .Z(n36655) );
  XNOR U38546 ( .A(m[594]), .B(n36656), .Z(n36654) );
  NAND U38547 ( .A(n36657), .B(mul_pow), .Z(n36656) );
  XOR U38548 ( .A(m[594]), .B(c[594]), .Z(n36657) );
  XOR U38549 ( .A(n36658), .B(n36659), .Z(n36650) );
  ANDN U38550 ( .B(n36660), .A(n31932), .Z(n36658) );
  XNOR U38551 ( .A(\modmult_1/zin[0][592] ), .B(n36661), .Z(n31932) );
  IV U38552 ( .A(n36659), .Z(n36661) );
  XOR U38553 ( .A(n36659), .B(n31933), .Z(n36660) );
  XNOR U38554 ( .A(n36662), .B(n36663), .Z(n31933) );
  ANDN U38555 ( .B(\modmult_1/xin[1023] ), .A(n36664), .Z(n36662) );
  IV U38556 ( .A(n36663), .Z(n36664) );
  XNOR U38557 ( .A(m[593]), .B(n36665), .Z(n36663) );
  NAND U38558 ( .A(n36666), .B(mul_pow), .Z(n36665) );
  XOR U38559 ( .A(m[593]), .B(c[593]), .Z(n36666) );
  XOR U38560 ( .A(n36667), .B(n36668), .Z(n36659) );
  ANDN U38561 ( .B(n36669), .A(n31930), .Z(n36667) );
  XNOR U38562 ( .A(\modmult_1/zin[0][591] ), .B(n36670), .Z(n31930) );
  IV U38563 ( .A(n36668), .Z(n36670) );
  XOR U38564 ( .A(n36668), .B(n31931), .Z(n36669) );
  XNOR U38565 ( .A(n36671), .B(n36672), .Z(n31931) );
  ANDN U38566 ( .B(\modmult_1/xin[1023] ), .A(n36673), .Z(n36671) );
  IV U38567 ( .A(n36672), .Z(n36673) );
  XNOR U38568 ( .A(m[592]), .B(n36674), .Z(n36672) );
  NAND U38569 ( .A(n36675), .B(mul_pow), .Z(n36674) );
  XOR U38570 ( .A(m[592]), .B(c[592]), .Z(n36675) );
  XOR U38571 ( .A(n36676), .B(n36677), .Z(n36668) );
  ANDN U38572 ( .B(n36678), .A(n31928), .Z(n36676) );
  XNOR U38573 ( .A(\modmult_1/zin[0][590] ), .B(n36679), .Z(n31928) );
  IV U38574 ( .A(n36677), .Z(n36679) );
  XOR U38575 ( .A(n36677), .B(n31929), .Z(n36678) );
  XNOR U38576 ( .A(n36680), .B(n36681), .Z(n31929) );
  ANDN U38577 ( .B(\modmult_1/xin[1023] ), .A(n36682), .Z(n36680) );
  IV U38578 ( .A(n36681), .Z(n36682) );
  XNOR U38579 ( .A(m[591]), .B(n36683), .Z(n36681) );
  NAND U38580 ( .A(n36684), .B(mul_pow), .Z(n36683) );
  XOR U38581 ( .A(m[591]), .B(c[591]), .Z(n36684) );
  XOR U38582 ( .A(n36685), .B(n36686), .Z(n36677) );
  ANDN U38583 ( .B(n36687), .A(n31926), .Z(n36685) );
  XNOR U38584 ( .A(\modmult_1/zin[0][589] ), .B(n36688), .Z(n31926) );
  IV U38585 ( .A(n36686), .Z(n36688) );
  XOR U38586 ( .A(n36686), .B(n31927), .Z(n36687) );
  XNOR U38587 ( .A(n36689), .B(n36690), .Z(n31927) );
  ANDN U38588 ( .B(\modmult_1/xin[1023] ), .A(n36691), .Z(n36689) );
  IV U38589 ( .A(n36690), .Z(n36691) );
  XNOR U38590 ( .A(m[590]), .B(n36692), .Z(n36690) );
  NAND U38591 ( .A(n36693), .B(mul_pow), .Z(n36692) );
  XOR U38592 ( .A(m[590]), .B(c[590]), .Z(n36693) );
  XOR U38593 ( .A(n36694), .B(n36695), .Z(n36686) );
  ANDN U38594 ( .B(n36696), .A(n31924), .Z(n36694) );
  XNOR U38595 ( .A(\modmult_1/zin[0][588] ), .B(n36697), .Z(n31924) );
  IV U38596 ( .A(n36695), .Z(n36697) );
  XOR U38597 ( .A(n36695), .B(n31925), .Z(n36696) );
  XNOR U38598 ( .A(n36698), .B(n36699), .Z(n31925) );
  ANDN U38599 ( .B(\modmult_1/xin[1023] ), .A(n36700), .Z(n36698) );
  IV U38600 ( .A(n36699), .Z(n36700) );
  XNOR U38601 ( .A(m[589]), .B(n36701), .Z(n36699) );
  NAND U38602 ( .A(n36702), .B(mul_pow), .Z(n36701) );
  XOR U38603 ( .A(m[589]), .B(c[589]), .Z(n36702) );
  XOR U38604 ( .A(n36703), .B(n36704), .Z(n36695) );
  ANDN U38605 ( .B(n36705), .A(n31922), .Z(n36703) );
  XNOR U38606 ( .A(\modmult_1/zin[0][587] ), .B(n36706), .Z(n31922) );
  IV U38607 ( .A(n36704), .Z(n36706) );
  XOR U38608 ( .A(n36704), .B(n31923), .Z(n36705) );
  XNOR U38609 ( .A(n36707), .B(n36708), .Z(n31923) );
  ANDN U38610 ( .B(\modmult_1/xin[1023] ), .A(n36709), .Z(n36707) );
  IV U38611 ( .A(n36708), .Z(n36709) );
  XNOR U38612 ( .A(m[588]), .B(n36710), .Z(n36708) );
  NAND U38613 ( .A(n36711), .B(mul_pow), .Z(n36710) );
  XOR U38614 ( .A(m[588]), .B(c[588]), .Z(n36711) );
  XOR U38615 ( .A(n36712), .B(n36713), .Z(n36704) );
  ANDN U38616 ( .B(n36714), .A(n31920), .Z(n36712) );
  XNOR U38617 ( .A(\modmult_1/zin[0][586] ), .B(n36715), .Z(n31920) );
  IV U38618 ( .A(n36713), .Z(n36715) );
  XOR U38619 ( .A(n36713), .B(n31921), .Z(n36714) );
  XNOR U38620 ( .A(n36716), .B(n36717), .Z(n31921) );
  ANDN U38621 ( .B(\modmult_1/xin[1023] ), .A(n36718), .Z(n36716) );
  IV U38622 ( .A(n36717), .Z(n36718) );
  XNOR U38623 ( .A(m[587]), .B(n36719), .Z(n36717) );
  NAND U38624 ( .A(n36720), .B(mul_pow), .Z(n36719) );
  XOR U38625 ( .A(m[587]), .B(c[587]), .Z(n36720) );
  XOR U38626 ( .A(n36721), .B(n36722), .Z(n36713) );
  ANDN U38627 ( .B(n36723), .A(n31918), .Z(n36721) );
  XNOR U38628 ( .A(\modmult_1/zin[0][585] ), .B(n36724), .Z(n31918) );
  IV U38629 ( .A(n36722), .Z(n36724) );
  XOR U38630 ( .A(n36722), .B(n31919), .Z(n36723) );
  XNOR U38631 ( .A(n36725), .B(n36726), .Z(n31919) );
  ANDN U38632 ( .B(\modmult_1/xin[1023] ), .A(n36727), .Z(n36725) );
  IV U38633 ( .A(n36726), .Z(n36727) );
  XNOR U38634 ( .A(m[586]), .B(n36728), .Z(n36726) );
  NAND U38635 ( .A(n36729), .B(mul_pow), .Z(n36728) );
  XOR U38636 ( .A(m[586]), .B(c[586]), .Z(n36729) );
  XOR U38637 ( .A(n36730), .B(n36731), .Z(n36722) );
  ANDN U38638 ( .B(n36732), .A(n31916), .Z(n36730) );
  XNOR U38639 ( .A(\modmult_1/zin[0][584] ), .B(n36733), .Z(n31916) );
  IV U38640 ( .A(n36731), .Z(n36733) );
  XOR U38641 ( .A(n36731), .B(n31917), .Z(n36732) );
  XNOR U38642 ( .A(n36734), .B(n36735), .Z(n31917) );
  ANDN U38643 ( .B(\modmult_1/xin[1023] ), .A(n36736), .Z(n36734) );
  IV U38644 ( .A(n36735), .Z(n36736) );
  XNOR U38645 ( .A(m[585]), .B(n36737), .Z(n36735) );
  NAND U38646 ( .A(n36738), .B(mul_pow), .Z(n36737) );
  XOR U38647 ( .A(m[585]), .B(c[585]), .Z(n36738) );
  XOR U38648 ( .A(n36739), .B(n36740), .Z(n36731) );
  ANDN U38649 ( .B(n36741), .A(n31914), .Z(n36739) );
  XNOR U38650 ( .A(\modmult_1/zin[0][583] ), .B(n36742), .Z(n31914) );
  IV U38651 ( .A(n36740), .Z(n36742) );
  XOR U38652 ( .A(n36740), .B(n31915), .Z(n36741) );
  XNOR U38653 ( .A(n36743), .B(n36744), .Z(n31915) );
  ANDN U38654 ( .B(\modmult_1/xin[1023] ), .A(n36745), .Z(n36743) );
  IV U38655 ( .A(n36744), .Z(n36745) );
  XNOR U38656 ( .A(m[584]), .B(n36746), .Z(n36744) );
  NAND U38657 ( .A(n36747), .B(mul_pow), .Z(n36746) );
  XOR U38658 ( .A(m[584]), .B(c[584]), .Z(n36747) );
  XOR U38659 ( .A(n36748), .B(n36749), .Z(n36740) );
  ANDN U38660 ( .B(n36750), .A(n31912), .Z(n36748) );
  XNOR U38661 ( .A(\modmult_1/zin[0][582] ), .B(n36751), .Z(n31912) );
  IV U38662 ( .A(n36749), .Z(n36751) );
  XOR U38663 ( .A(n36749), .B(n31913), .Z(n36750) );
  XNOR U38664 ( .A(n36752), .B(n36753), .Z(n31913) );
  ANDN U38665 ( .B(\modmult_1/xin[1023] ), .A(n36754), .Z(n36752) );
  IV U38666 ( .A(n36753), .Z(n36754) );
  XNOR U38667 ( .A(m[583]), .B(n36755), .Z(n36753) );
  NAND U38668 ( .A(n36756), .B(mul_pow), .Z(n36755) );
  XOR U38669 ( .A(m[583]), .B(c[583]), .Z(n36756) );
  XOR U38670 ( .A(n36757), .B(n36758), .Z(n36749) );
  ANDN U38671 ( .B(n36759), .A(n31910), .Z(n36757) );
  XNOR U38672 ( .A(\modmult_1/zin[0][581] ), .B(n36760), .Z(n31910) );
  IV U38673 ( .A(n36758), .Z(n36760) );
  XOR U38674 ( .A(n36758), .B(n31911), .Z(n36759) );
  XNOR U38675 ( .A(n36761), .B(n36762), .Z(n31911) );
  ANDN U38676 ( .B(\modmult_1/xin[1023] ), .A(n36763), .Z(n36761) );
  IV U38677 ( .A(n36762), .Z(n36763) );
  XNOR U38678 ( .A(m[582]), .B(n36764), .Z(n36762) );
  NAND U38679 ( .A(n36765), .B(mul_pow), .Z(n36764) );
  XOR U38680 ( .A(m[582]), .B(c[582]), .Z(n36765) );
  XOR U38681 ( .A(n36766), .B(n36767), .Z(n36758) );
  ANDN U38682 ( .B(n36768), .A(n31908), .Z(n36766) );
  XNOR U38683 ( .A(\modmult_1/zin[0][580] ), .B(n36769), .Z(n31908) );
  IV U38684 ( .A(n36767), .Z(n36769) );
  XOR U38685 ( .A(n36767), .B(n31909), .Z(n36768) );
  XNOR U38686 ( .A(n36770), .B(n36771), .Z(n31909) );
  ANDN U38687 ( .B(\modmult_1/xin[1023] ), .A(n36772), .Z(n36770) );
  IV U38688 ( .A(n36771), .Z(n36772) );
  XNOR U38689 ( .A(m[581]), .B(n36773), .Z(n36771) );
  NAND U38690 ( .A(n36774), .B(mul_pow), .Z(n36773) );
  XOR U38691 ( .A(m[581]), .B(c[581]), .Z(n36774) );
  XOR U38692 ( .A(n36775), .B(n36776), .Z(n36767) );
  ANDN U38693 ( .B(n36777), .A(n31906), .Z(n36775) );
  XNOR U38694 ( .A(\modmult_1/zin[0][579] ), .B(n36778), .Z(n31906) );
  IV U38695 ( .A(n36776), .Z(n36778) );
  XOR U38696 ( .A(n36776), .B(n31907), .Z(n36777) );
  XNOR U38697 ( .A(n36779), .B(n36780), .Z(n31907) );
  ANDN U38698 ( .B(\modmult_1/xin[1023] ), .A(n36781), .Z(n36779) );
  IV U38699 ( .A(n36780), .Z(n36781) );
  XNOR U38700 ( .A(m[580]), .B(n36782), .Z(n36780) );
  NAND U38701 ( .A(n36783), .B(mul_pow), .Z(n36782) );
  XOR U38702 ( .A(m[580]), .B(c[580]), .Z(n36783) );
  XOR U38703 ( .A(n36784), .B(n36785), .Z(n36776) );
  ANDN U38704 ( .B(n36786), .A(n31904), .Z(n36784) );
  XNOR U38705 ( .A(\modmult_1/zin[0][578] ), .B(n36787), .Z(n31904) );
  IV U38706 ( .A(n36785), .Z(n36787) );
  XOR U38707 ( .A(n36785), .B(n31905), .Z(n36786) );
  XNOR U38708 ( .A(n36788), .B(n36789), .Z(n31905) );
  ANDN U38709 ( .B(\modmult_1/xin[1023] ), .A(n36790), .Z(n36788) );
  IV U38710 ( .A(n36789), .Z(n36790) );
  XNOR U38711 ( .A(m[579]), .B(n36791), .Z(n36789) );
  NAND U38712 ( .A(n36792), .B(mul_pow), .Z(n36791) );
  XOR U38713 ( .A(m[579]), .B(c[579]), .Z(n36792) );
  XOR U38714 ( .A(n36793), .B(n36794), .Z(n36785) );
  ANDN U38715 ( .B(n36795), .A(n31902), .Z(n36793) );
  XNOR U38716 ( .A(\modmult_1/zin[0][577] ), .B(n36796), .Z(n31902) );
  IV U38717 ( .A(n36794), .Z(n36796) );
  XOR U38718 ( .A(n36794), .B(n31903), .Z(n36795) );
  XNOR U38719 ( .A(n36797), .B(n36798), .Z(n31903) );
  ANDN U38720 ( .B(\modmult_1/xin[1023] ), .A(n36799), .Z(n36797) );
  IV U38721 ( .A(n36798), .Z(n36799) );
  XNOR U38722 ( .A(m[578]), .B(n36800), .Z(n36798) );
  NAND U38723 ( .A(n36801), .B(mul_pow), .Z(n36800) );
  XOR U38724 ( .A(m[578]), .B(c[578]), .Z(n36801) );
  XOR U38725 ( .A(n36802), .B(n36803), .Z(n36794) );
  ANDN U38726 ( .B(n36804), .A(n31900), .Z(n36802) );
  XNOR U38727 ( .A(\modmult_1/zin[0][576] ), .B(n36805), .Z(n31900) );
  IV U38728 ( .A(n36803), .Z(n36805) );
  XOR U38729 ( .A(n36803), .B(n31901), .Z(n36804) );
  XNOR U38730 ( .A(n36806), .B(n36807), .Z(n31901) );
  ANDN U38731 ( .B(\modmult_1/xin[1023] ), .A(n36808), .Z(n36806) );
  IV U38732 ( .A(n36807), .Z(n36808) );
  XNOR U38733 ( .A(m[577]), .B(n36809), .Z(n36807) );
  NAND U38734 ( .A(n36810), .B(mul_pow), .Z(n36809) );
  XOR U38735 ( .A(m[577]), .B(c[577]), .Z(n36810) );
  XOR U38736 ( .A(n36811), .B(n36812), .Z(n36803) );
  ANDN U38737 ( .B(n36813), .A(n31898), .Z(n36811) );
  XNOR U38738 ( .A(\modmult_1/zin[0][575] ), .B(n36814), .Z(n31898) );
  IV U38739 ( .A(n36812), .Z(n36814) );
  XOR U38740 ( .A(n36812), .B(n31899), .Z(n36813) );
  XNOR U38741 ( .A(n36815), .B(n36816), .Z(n31899) );
  ANDN U38742 ( .B(\modmult_1/xin[1023] ), .A(n36817), .Z(n36815) );
  IV U38743 ( .A(n36816), .Z(n36817) );
  XNOR U38744 ( .A(m[576]), .B(n36818), .Z(n36816) );
  NAND U38745 ( .A(n36819), .B(mul_pow), .Z(n36818) );
  XOR U38746 ( .A(m[576]), .B(c[576]), .Z(n36819) );
  XOR U38747 ( .A(n36820), .B(n36821), .Z(n36812) );
  ANDN U38748 ( .B(n36822), .A(n31896), .Z(n36820) );
  XNOR U38749 ( .A(\modmult_1/zin[0][574] ), .B(n36823), .Z(n31896) );
  IV U38750 ( .A(n36821), .Z(n36823) );
  XOR U38751 ( .A(n36821), .B(n31897), .Z(n36822) );
  XNOR U38752 ( .A(n36824), .B(n36825), .Z(n31897) );
  ANDN U38753 ( .B(\modmult_1/xin[1023] ), .A(n36826), .Z(n36824) );
  IV U38754 ( .A(n36825), .Z(n36826) );
  XNOR U38755 ( .A(m[575]), .B(n36827), .Z(n36825) );
  NAND U38756 ( .A(n36828), .B(mul_pow), .Z(n36827) );
  XOR U38757 ( .A(m[575]), .B(c[575]), .Z(n36828) );
  XOR U38758 ( .A(n36829), .B(n36830), .Z(n36821) );
  ANDN U38759 ( .B(n36831), .A(n31894), .Z(n36829) );
  XNOR U38760 ( .A(\modmult_1/zin[0][573] ), .B(n36832), .Z(n31894) );
  IV U38761 ( .A(n36830), .Z(n36832) );
  XOR U38762 ( .A(n36830), .B(n31895), .Z(n36831) );
  XNOR U38763 ( .A(n36833), .B(n36834), .Z(n31895) );
  ANDN U38764 ( .B(\modmult_1/xin[1023] ), .A(n36835), .Z(n36833) );
  IV U38765 ( .A(n36834), .Z(n36835) );
  XNOR U38766 ( .A(m[574]), .B(n36836), .Z(n36834) );
  NAND U38767 ( .A(n36837), .B(mul_pow), .Z(n36836) );
  XOR U38768 ( .A(m[574]), .B(c[574]), .Z(n36837) );
  XOR U38769 ( .A(n36838), .B(n36839), .Z(n36830) );
  ANDN U38770 ( .B(n36840), .A(n31892), .Z(n36838) );
  XNOR U38771 ( .A(\modmult_1/zin[0][572] ), .B(n36841), .Z(n31892) );
  IV U38772 ( .A(n36839), .Z(n36841) );
  XOR U38773 ( .A(n36839), .B(n31893), .Z(n36840) );
  XNOR U38774 ( .A(n36842), .B(n36843), .Z(n31893) );
  ANDN U38775 ( .B(\modmult_1/xin[1023] ), .A(n36844), .Z(n36842) );
  IV U38776 ( .A(n36843), .Z(n36844) );
  XNOR U38777 ( .A(m[573]), .B(n36845), .Z(n36843) );
  NAND U38778 ( .A(n36846), .B(mul_pow), .Z(n36845) );
  XOR U38779 ( .A(m[573]), .B(c[573]), .Z(n36846) );
  XOR U38780 ( .A(n36847), .B(n36848), .Z(n36839) );
  ANDN U38781 ( .B(n36849), .A(n31890), .Z(n36847) );
  XNOR U38782 ( .A(\modmult_1/zin[0][571] ), .B(n36850), .Z(n31890) );
  IV U38783 ( .A(n36848), .Z(n36850) );
  XOR U38784 ( .A(n36848), .B(n31891), .Z(n36849) );
  XNOR U38785 ( .A(n36851), .B(n36852), .Z(n31891) );
  ANDN U38786 ( .B(\modmult_1/xin[1023] ), .A(n36853), .Z(n36851) );
  IV U38787 ( .A(n36852), .Z(n36853) );
  XNOR U38788 ( .A(m[572]), .B(n36854), .Z(n36852) );
  NAND U38789 ( .A(n36855), .B(mul_pow), .Z(n36854) );
  XOR U38790 ( .A(m[572]), .B(c[572]), .Z(n36855) );
  XOR U38791 ( .A(n36856), .B(n36857), .Z(n36848) );
  ANDN U38792 ( .B(n36858), .A(n31888), .Z(n36856) );
  XNOR U38793 ( .A(\modmult_1/zin[0][570] ), .B(n36859), .Z(n31888) );
  IV U38794 ( .A(n36857), .Z(n36859) );
  XOR U38795 ( .A(n36857), .B(n31889), .Z(n36858) );
  XNOR U38796 ( .A(n36860), .B(n36861), .Z(n31889) );
  ANDN U38797 ( .B(\modmult_1/xin[1023] ), .A(n36862), .Z(n36860) );
  IV U38798 ( .A(n36861), .Z(n36862) );
  XNOR U38799 ( .A(m[571]), .B(n36863), .Z(n36861) );
  NAND U38800 ( .A(n36864), .B(mul_pow), .Z(n36863) );
  XOR U38801 ( .A(m[571]), .B(c[571]), .Z(n36864) );
  XOR U38802 ( .A(n36865), .B(n36866), .Z(n36857) );
  ANDN U38803 ( .B(n36867), .A(n31886), .Z(n36865) );
  XNOR U38804 ( .A(\modmult_1/zin[0][569] ), .B(n36868), .Z(n31886) );
  IV U38805 ( .A(n36866), .Z(n36868) );
  XOR U38806 ( .A(n36866), .B(n31887), .Z(n36867) );
  XNOR U38807 ( .A(n36869), .B(n36870), .Z(n31887) );
  ANDN U38808 ( .B(\modmult_1/xin[1023] ), .A(n36871), .Z(n36869) );
  IV U38809 ( .A(n36870), .Z(n36871) );
  XNOR U38810 ( .A(m[570]), .B(n36872), .Z(n36870) );
  NAND U38811 ( .A(n36873), .B(mul_pow), .Z(n36872) );
  XOR U38812 ( .A(m[570]), .B(c[570]), .Z(n36873) );
  XOR U38813 ( .A(n36874), .B(n36875), .Z(n36866) );
  ANDN U38814 ( .B(n36876), .A(n31884), .Z(n36874) );
  XNOR U38815 ( .A(\modmult_1/zin[0][568] ), .B(n36877), .Z(n31884) );
  IV U38816 ( .A(n36875), .Z(n36877) );
  XOR U38817 ( .A(n36875), .B(n31885), .Z(n36876) );
  XNOR U38818 ( .A(n36878), .B(n36879), .Z(n31885) );
  ANDN U38819 ( .B(\modmult_1/xin[1023] ), .A(n36880), .Z(n36878) );
  IV U38820 ( .A(n36879), .Z(n36880) );
  XNOR U38821 ( .A(m[569]), .B(n36881), .Z(n36879) );
  NAND U38822 ( .A(n36882), .B(mul_pow), .Z(n36881) );
  XOR U38823 ( .A(m[569]), .B(c[569]), .Z(n36882) );
  XOR U38824 ( .A(n36883), .B(n36884), .Z(n36875) );
  ANDN U38825 ( .B(n36885), .A(n31882), .Z(n36883) );
  XNOR U38826 ( .A(\modmult_1/zin[0][567] ), .B(n36886), .Z(n31882) );
  IV U38827 ( .A(n36884), .Z(n36886) );
  XOR U38828 ( .A(n36884), .B(n31883), .Z(n36885) );
  XNOR U38829 ( .A(n36887), .B(n36888), .Z(n31883) );
  ANDN U38830 ( .B(\modmult_1/xin[1023] ), .A(n36889), .Z(n36887) );
  IV U38831 ( .A(n36888), .Z(n36889) );
  XNOR U38832 ( .A(m[568]), .B(n36890), .Z(n36888) );
  NAND U38833 ( .A(n36891), .B(mul_pow), .Z(n36890) );
  XOR U38834 ( .A(m[568]), .B(c[568]), .Z(n36891) );
  XOR U38835 ( .A(n36892), .B(n36893), .Z(n36884) );
  ANDN U38836 ( .B(n36894), .A(n31880), .Z(n36892) );
  XNOR U38837 ( .A(\modmult_1/zin[0][566] ), .B(n36895), .Z(n31880) );
  IV U38838 ( .A(n36893), .Z(n36895) );
  XOR U38839 ( .A(n36893), .B(n31881), .Z(n36894) );
  XNOR U38840 ( .A(n36896), .B(n36897), .Z(n31881) );
  ANDN U38841 ( .B(\modmult_1/xin[1023] ), .A(n36898), .Z(n36896) );
  IV U38842 ( .A(n36897), .Z(n36898) );
  XNOR U38843 ( .A(m[567]), .B(n36899), .Z(n36897) );
  NAND U38844 ( .A(n36900), .B(mul_pow), .Z(n36899) );
  XOR U38845 ( .A(m[567]), .B(c[567]), .Z(n36900) );
  XOR U38846 ( .A(n36901), .B(n36902), .Z(n36893) );
  ANDN U38847 ( .B(n36903), .A(n31878), .Z(n36901) );
  XNOR U38848 ( .A(\modmult_1/zin[0][565] ), .B(n36904), .Z(n31878) );
  IV U38849 ( .A(n36902), .Z(n36904) );
  XOR U38850 ( .A(n36902), .B(n31879), .Z(n36903) );
  XNOR U38851 ( .A(n36905), .B(n36906), .Z(n31879) );
  ANDN U38852 ( .B(\modmult_1/xin[1023] ), .A(n36907), .Z(n36905) );
  IV U38853 ( .A(n36906), .Z(n36907) );
  XNOR U38854 ( .A(m[566]), .B(n36908), .Z(n36906) );
  NAND U38855 ( .A(n36909), .B(mul_pow), .Z(n36908) );
  XOR U38856 ( .A(m[566]), .B(c[566]), .Z(n36909) );
  XOR U38857 ( .A(n36910), .B(n36911), .Z(n36902) );
  ANDN U38858 ( .B(n36912), .A(n31876), .Z(n36910) );
  XNOR U38859 ( .A(\modmult_1/zin[0][564] ), .B(n36913), .Z(n31876) );
  IV U38860 ( .A(n36911), .Z(n36913) );
  XOR U38861 ( .A(n36911), .B(n31877), .Z(n36912) );
  XNOR U38862 ( .A(n36914), .B(n36915), .Z(n31877) );
  ANDN U38863 ( .B(\modmult_1/xin[1023] ), .A(n36916), .Z(n36914) );
  IV U38864 ( .A(n36915), .Z(n36916) );
  XNOR U38865 ( .A(m[565]), .B(n36917), .Z(n36915) );
  NAND U38866 ( .A(n36918), .B(mul_pow), .Z(n36917) );
  XOR U38867 ( .A(m[565]), .B(c[565]), .Z(n36918) );
  XOR U38868 ( .A(n36919), .B(n36920), .Z(n36911) );
  ANDN U38869 ( .B(n36921), .A(n31874), .Z(n36919) );
  XNOR U38870 ( .A(\modmult_1/zin[0][563] ), .B(n36922), .Z(n31874) );
  IV U38871 ( .A(n36920), .Z(n36922) );
  XOR U38872 ( .A(n36920), .B(n31875), .Z(n36921) );
  XNOR U38873 ( .A(n36923), .B(n36924), .Z(n31875) );
  ANDN U38874 ( .B(\modmult_1/xin[1023] ), .A(n36925), .Z(n36923) );
  IV U38875 ( .A(n36924), .Z(n36925) );
  XNOR U38876 ( .A(m[564]), .B(n36926), .Z(n36924) );
  NAND U38877 ( .A(n36927), .B(mul_pow), .Z(n36926) );
  XOR U38878 ( .A(m[564]), .B(c[564]), .Z(n36927) );
  XOR U38879 ( .A(n36928), .B(n36929), .Z(n36920) );
  ANDN U38880 ( .B(n36930), .A(n31872), .Z(n36928) );
  XNOR U38881 ( .A(\modmult_1/zin[0][562] ), .B(n36931), .Z(n31872) );
  IV U38882 ( .A(n36929), .Z(n36931) );
  XOR U38883 ( .A(n36929), .B(n31873), .Z(n36930) );
  XNOR U38884 ( .A(n36932), .B(n36933), .Z(n31873) );
  ANDN U38885 ( .B(\modmult_1/xin[1023] ), .A(n36934), .Z(n36932) );
  IV U38886 ( .A(n36933), .Z(n36934) );
  XNOR U38887 ( .A(m[563]), .B(n36935), .Z(n36933) );
  NAND U38888 ( .A(n36936), .B(mul_pow), .Z(n36935) );
  XOR U38889 ( .A(m[563]), .B(c[563]), .Z(n36936) );
  XOR U38890 ( .A(n36937), .B(n36938), .Z(n36929) );
  ANDN U38891 ( .B(n36939), .A(n31870), .Z(n36937) );
  XNOR U38892 ( .A(\modmult_1/zin[0][561] ), .B(n36940), .Z(n31870) );
  IV U38893 ( .A(n36938), .Z(n36940) );
  XOR U38894 ( .A(n36938), .B(n31871), .Z(n36939) );
  XNOR U38895 ( .A(n36941), .B(n36942), .Z(n31871) );
  ANDN U38896 ( .B(\modmult_1/xin[1023] ), .A(n36943), .Z(n36941) );
  IV U38897 ( .A(n36942), .Z(n36943) );
  XNOR U38898 ( .A(m[562]), .B(n36944), .Z(n36942) );
  NAND U38899 ( .A(n36945), .B(mul_pow), .Z(n36944) );
  XOR U38900 ( .A(m[562]), .B(c[562]), .Z(n36945) );
  XOR U38901 ( .A(n36946), .B(n36947), .Z(n36938) );
  ANDN U38902 ( .B(n36948), .A(n31868), .Z(n36946) );
  XNOR U38903 ( .A(\modmult_1/zin[0][560] ), .B(n36949), .Z(n31868) );
  IV U38904 ( .A(n36947), .Z(n36949) );
  XOR U38905 ( .A(n36947), .B(n31869), .Z(n36948) );
  XNOR U38906 ( .A(n36950), .B(n36951), .Z(n31869) );
  ANDN U38907 ( .B(\modmult_1/xin[1023] ), .A(n36952), .Z(n36950) );
  IV U38908 ( .A(n36951), .Z(n36952) );
  XNOR U38909 ( .A(m[561]), .B(n36953), .Z(n36951) );
  NAND U38910 ( .A(n36954), .B(mul_pow), .Z(n36953) );
  XOR U38911 ( .A(m[561]), .B(c[561]), .Z(n36954) );
  XOR U38912 ( .A(n36955), .B(n36956), .Z(n36947) );
  ANDN U38913 ( .B(n36957), .A(n31866), .Z(n36955) );
  XNOR U38914 ( .A(\modmult_1/zin[0][559] ), .B(n36958), .Z(n31866) );
  IV U38915 ( .A(n36956), .Z(n36958) );
  XOR U38916 ( .A(n36956), .B(n31867), .Z(n36957) );
  XNOR U38917 ( .A(n36959), .B(n36960), .Z(n31867) );
  ANDN U38918 ( .B(\modmult_1/xin[1023] ), .A(n36961), .Z(n36959) );
  IV U38919 ( .A(n36960), .Z(n36961) );
  XNOR U38920 ( .A(m[560]), .B(n36962), .Z(n36960) );
  NAND U38921 ( .A(n36963), .B(mul_pow), .Z(n36962) );
  XOR U38922 ( .A(m[560]), .B(c[560]), .Z(n36963) );
  XOR U38923 ( .A(n36964), .B(n36965), .Z(n36956) );
  ANDN U38924 ( .B(n36966), .A(n31864), .Z(n36964) );
  XNOR U38925 ( .A(\modmult_1/zin[0][558] ), .B(n36967), .Z(n31864) );
  IV U38926 ( .A(n36965), .Z(n36967) );
  XOR U38927 ( .A(n36965), .B(n31865), .Z(n36966) );
  XNOR U38928 ( .A(n36968), .B(n36969), .Z(n31865) );
  ANDN U38929 ( .B(\modmult_1/xin[1023] ), .A(n36970), .Z(n36968) );
  IV U38930 ( .A(n36969), .Z(n36970) );
  XNOR U38931 ( .A(m[559]), .B(n36971), .Z(n36969) );
  NAND U38932 ( .A(n36972), .B(mul_pow), .Z(n36971) );
  XOR U38933 ( .A(m[559]), .B(c[559]), .Z(n36972) );
  XOR U38934 ( .A(n36973), .B(n36974), .Z(n36965) );
  ANDN U38935 ( .B(n36975), .A(n31862), .Z(n36973) );
  XNOR U38936 ( .A(\modmult_1/zin[0][557] ), .B(n36976), .Z(n31862) );
  IV U38937 ( .A(n36974), .Z(n36976) );
  XOR U38938 ( .A(n36974), .B(n31863), .Z(n36975) );
  XNOR U38939 ( .A(n36977), .B(n36978), .Z(n31863) );
  ANDN U38940 ( .B(\modmult_1/xin[1023] ), .A(n36979), .Z(n36977) );
  IV U38941 ( .A(n36978), .Z(n36979) );
  XNOR U38942 ( .A(m[558]), .B(n36980), .Z(n36978) );
  NAND U38943 ( .A(n36981), .B(mul_pow), .Z(n36980) );
  XOR U38944 ( .A(m[558]), .B(c[558]), .Z(n36981) );
  XOR U38945 ( .A(n36982), .B(n36983), .Z(n36974) );
  ANDN U38946 ( .B(n36984), .A(n31860), .Z(n36982) );
  XNOR U38947 ( .A(\modmult_1/zin[0][556] ), .B(n36985), .Z(n31860) );
  IV U38948 ( .A(n36983), .Z(n36985) );
  XOR U38949 ( .A(n36983), .B(n31861), .Z(n36984) );
  XNOR U38950 ( .A(n36986), .B(n36987), .Z(n31861) );
  ANDN U38951 ( .B(\modmult_1/xin[1023] ), .A(n36988), .Z(n36986) );
  IV U38952 ( .A(n36987), .Z(n36988) );
  XNOR U38953 ( .A(m[557]), .B(n36989), .Z(n36987) );
  NAND U38954 ( .A(n36990), .B(mul_pow), .Z(n36989) );
  XOR U38955 ( .A(m[557]), .B(c[557]), .Z(n36990) );
  XOR U38956 ( .A(n36991), .B(n36992), .Z(n36983) );
  ANDN U38957 ( .B(n36993), .A(n31858), .Z(n36991) );
  XNOR U38958 ( .A(\modmult_1/zin[0][555] ), .B(n36994), .Z(n31858) );
  IV U38959 ( .A(n36992), .Z(n36994) );
  XOR U38960 ( .A(n36992), .B(n31859), .Z(n36993) );
  XNOR U38961 ( .A(n36995), .B(n36996), .Z(n31859) );
  ANDN U38962 ( .B(\modmult_1/xin[1023] ), .A(n36997), .Z(n36995) );
  IV U38963 ( .A(n36996), .Z(n36997) );
  XNOR U38964 ( .A(m[556]), .B(n36998), .Z(n36996) );
  NAND U38965 ( .A(n36999), .B(mul_pow), .Z(n36998) );
  XOR U38966 ( .A(m[556]), .B(c[556]), .Z(n36999) );
  XOR U38967 ( .A(n37000), .B(n37001), .Z(n36992) );
  ANDN U38968 ( .B(n37002), .A(n31856), .Z(n37000) );
  XNOR U38969 ( .A(\modmult_1/zin[0][554] ), .B(n37003), .Z(n31856) );
  IV U38970 ( .A(n37001), .Z(n37003) );
  XOR U38971 ( .A(n37001), .B(n31857), .Z(n37002) );
  XNOR U38972 ( .A(n37004), .B(n37005), .Z(n31857) );
  ANDN U38973 ( .B(\modmult_1/xin[1023] ), .A(n37006), .Z(n37004) );
  IV U38974 ( .A(n37005), .Z(n37006) );
  XNOR U38975 ( .A(m[555]), .B(n37007), .Z(n37005) );
  NAND U38976 ( .A(n37008), .B(mul_pow), .Z(n37007) );
  XOR U38977 ( .A(m[555]), .B(c[555]), .Z(n37008) );
  XOR U38978 ( .A(n37009), .B(n37010), .Z(n37001) );
  ANDN U38979 ( .B(n37011), .A(n31854), .Z(n37009) );
  XNOR U38980 ( .A(\modmult_1/zin[0][553] ), .B(n37012), .Z(n31854) );
  IV U38981 ( .A(n37010), .Z(n37012) );
  XOR U38982 ( .A(n37010), .B(n31855), .Z(n37011) );
  XNOR U38983 ( .A(n37013), .B(n37014), .Z(n31855) );
  ANDN U38984 ( .B(\modmult_1/xin[1023] ), .A(n37015), .Z(n37013) );
  IV U38985 ( .A(n37014), .Z(n37015) );
  XNOR U38986 ( .A(m[554]), .B(n37016), .Z(n37014) );
  NAND U38987 ( .A(n37017), .B(mul_pow), .Z(n37016) );
  XOR U38988 ( .A(m[554]), .B(c[554]), .Z(n37017) );
  XOR U38989 ( .A(n37018), .B(n37019), .Z(n37010) );
  ANDN U38990 ( .B(n37020), .A(n31852), .Z(n37018) );
  XNOR U38991 ( .A(\modmult_1/zin[0][552] ), .B(n37021), .Z(n31852) );
  IV U38992 ( .A(n37019), .Z(n37021) );
  XOR U38993 ( .A(n37019), .B(n31853), .Z(n37020) );
  XNOR U38994 ( .A(n37022), .B(n37023), .Z(n31853) );
  ANDN U38995 ( .B(\modmult_1/xin[1023] ), .A(n37024), .Z(n37022) );
  IV U38996 ( .A(n37023), .Z(n37024) );
  XNOR U38997 ( .A(m[553]), .B(n37025), .Z(n37023) );
  NAND U38998 ( .A(n37026), .B(mul_pow), .Z(n37025) );
  XOR U38999 ( .A(m[553]), .B(c[553]), .Z(n37026) );
  XOR U39000 ( .A(n37027), .B(n37028), .Z(n37019) );
  ANDN U39001 ( .B(n37029), .A(n31850), .Z(n37027) );
  XNOR U39002 ( .A(\modmult_1/zin[0][551] ), .B(n37030), .Z(n31850) );
  IV U39003 ( .A(n37028), .Z(n37030) );
  XOR U39004 ( .A(n37028), .B(n31851), .Z(n37029) );
  XNOR U39005 ( .A(n37031), .B(n37032), .Z(n31851) );
  ANDN U39006 ( .B(\modmult_1/xin[1023] ), .A(n37033), .Z(n37031) );
  IV U39007 ( .A(n37032), .Z(n37033) );
  XNOR U39008 ( .A(m[552]), .B(n37034), .Z(n37032) );
  NAND U39009 ( .A(n37035), .B(mul_pow), .Z(n37034) );
  XOR U39010 ( .A(m[552]), .B(c[552]), .Z(n37035) );
  XOR U39011 ( .A(n37036), .B(n37037), .Z(n37028) );
  ANDN U39012 ( .B(n37038), .A(n31848), .Z(n37036) );
  XNOR U39013 ( .A(\modmult_1/zin[0][550] ), .B(n37039), .Z(n31848) );
  IV U39014 ( .A(n37037), .Z(n37039) );
  XOR U39015 ( .A(n37037), .B(n31849), .Z(n37038) );
  XNOR U39016 ( .A(n37040), .B(n37041), .Z(n31849) );
  ANDN U39017 ( .B(\modmult_1/xin[1023] ), .A(n37042), .Z(n37040) );
  IV U39018 ( .A(n37041), .Z(n37042) );
  XNOR U39019 ( .A(m[551]), .B(n37043), .Z(n37041) );
  NAND U39020 ( .A(n37044), .B(mul_pow), .Z(n37043) );
  XOR U39021 ( .A(m[551]), .B(c[551]), .Z(n37044) );
  XOR U39022 ( .A(n37045), .B(n37046), .Z(n37037) );
  ANDN U39023 ( .B(n37047), .A(n31846), .Z(n37045) );
  XNOR U39024 ( .A(\modmult_1/zin[0][549] ), .B(n37048), .Z(n31846) );
  IV U39025 ( .A(n37046), .Z(n37048) );
  XOR U39026 ( .A(n37046), .B(n31847), .Z(n37047) );
  XNOR U39027 ( .A(n37049), .B(n37050), .Z(n31847) );
  ANDN U39028 ( .B(\modmult_1/xin[1023] ), .A(n37051), .Z(n37049) );
  IV U39029 ( .A(n37050), .Z(n37051) );
  XNOR U39030 ( .A(m[550]), .B(n37052), .Z(n37050) );
  NAND U39031 ( .A(n37053), .B(mul_pow), .Z(n37052) );
  XOR U39032 ( .A(m[550]), .B(c[550]), .Z(n37053) );
  XOR U39033 ( .A(n37054), .B(n37055), .Z(n37046) );
  ANDN U39034 ( .B(n37056), .A(n31844), .Z(n37054) );
  XNOR U39035 ( .A(\modmult_1/zin[0][548] ), .B(n37057), .Z(n31844) );
  IV U39036 ( .A(n37055), .Z(n37057) );
  XOR U39037 ( .A(n37055), .B(n31845), .Z(n37056) );
  XNOR U39038 ( .A(n37058), .B(n37059), .Z(n31845) );
  ANDN U39039 ( .B(\modmult_1/xin[1023] ), .A(n37060), .Z(n37058) );
  IV U39040 ( .A(n37059), .Z(n37060) );
  XNOR U39041 ( .A(m[549]), .B(n37061), .Z(n37059) );
  NAND U39042 ( .A(n37062), .B(mul_pow), .Z(n37061) );
  XOR U39043 ( .A(m[549]), .B(c[549]), .Z(n37062) );
  XOR U39044 ( .A(n37063), .B(n37064), .Z(n37055) );
  ANDN U39045 ( .B(n37065), .A(n31842), .Z(n37063) );
  XNOR U39046 ( .A(\modmult_1/zin[0][547] ), .B(n37066), .Z(n31842) );
  IV U39047 ( .A(n37064), .Z(n37066) );
  XOR U39048 ( .A(n37064), .B(n31843), .Z(n37065) );
  XNOR U39049 ( .A(n37067), .B(n37068), .Z(n31843) );
  ANDN U39050 ( .B(\modmult_1/xin[1023] ), .A(n37069), .Z(n37067) );
  IV U39051 ( .A(n37068), .Z(n37069) );
  XNOR U39052 ( .A(m[548]), .B(n37070), .Z(n37068) );
  NAND U39053 ( .A(n37071), .B(mul_pow), .Z(n37070) );
  XOR U39054 ( .A(m[548]), .B(c[548]), .Z(n37071) );
  XOR U39055 ( .A(n37072), .B(n37073), .Z(n37064) );
  ANDN U39056 ( .B(n37074), .A(n31840), .Z(n37072) );
  XNOR U39057 ( .A(\modmult_1/zin[0][546] ), .B(n37075), .Z(n31840) );
  IV U39058 ( .A(n37073), .Z(n37075) );
  XOR U39059 ( .A(n37073), .B(n31841), .Z(n37074) );
  XNOR U39060 ( .A(n37076), .B(n37077), .Z(n31841) );
  ANDN U39061 ( .B(\modmult_1/xin[1023] ), .A(n37078), .Z(n37076) );
  IV U39062 ( .A(n37077), .Z(n37078) );
  XNOR U39063 ( .A(m[547]), .B(n37079), .Z(n37077) );
  NAND U39064 ( .A(n37080), .B(mul_pow), .Z(n37079) );
  XOR U39065 ( .A(m[547]), .B(c[547]), .Z(n37080) );
  XOR U39066 ( .A(n37081), .B(n37082), .Z(n37073) );
  ANDN U39067 ( .B(n37083), .A(n31838), .Z(n37081) );
  XNOR U39068 ( .A(\modmult_1/zin[0][545] ), .B(n37084), .Z(n31838) );
  IV U39069 ( .A(n37082), .Z(n37084) );
  XOR U39070 ( .A(n37082), .B(n31839), .Z(n37083) );
  XNOR U39071 ( .A(n37085), .B(n37086), .Z(n31839) );
  ANDN U39072 ( .B(\modmult_1/xin[1023] ), .A(n37087), .Z(n37085) );
  IV U39073 ( .A(n37086), .Z(n37087) );
  XNOR U39074 ( .A(m[546]), .B(n37088), .Z(n37086) );
  NAND U39075 ( .A(n37089), .B(mul_pow), .Z(n37088) );
  XOR U39076 ( .A(m[546]), .B(c[546]), .Z(n37089) );
  XOR U39077 ( .A(n37090), .B(n37091), .Z(n37082) );
  ANDN U39078 ( .B(n37092), .A(n31836), .Z(n37090) );
  XNOR U39079 ( .A(\modmult_1/zin[0][544] ), .B(n37093), .Z(n31836) );
  IV U39080 ( .A(n37091), .Z(n37093) );
  XOR U39081 ( .A(n37091), .B(n31837), .Z(n37092) );
  XNOR U39082 ( .A(n37094), .B(n37095), .Z(n31837) );
  ANDN U39083 ( .B(\modmult_1/xin[1023] ), .A(n37096), .Z(n37094) );
  IV U39084 ( .A(n37095), .Z(n37096) );
  XNOR U39085 ( .A(m[545]), .B(n37097), .Z(n37095) );
  NAND U39086 ( .A(n37098), .B(mul_pow), .Z(n37097) );
  XOR U39087 ( .A(m[545]), .B(c[545]), .Z(n37098) );
  XOR U39088 ( .A(n37099), .B(n37100), .Z(n37091) );
  ANDN U39089 ( .B(n37101), .A(n31834), .Z(n37099) );
  XNOR U39090 ( .A(\modmult_1/zin[0][543] ), .B(n37102), .Z(n31834) );
  IV U39091 ( .A(n37100), .Z(n37102) );
  XOR U39092 ( .A(n37100), .B(n31835), .Z(n37101) );
  XNOR U39093 ( .A(n37103), .B(n37104), .Z(n31835) );
  ANDN U39094 ( .B(\modmult_1/xin[1023] ), .A(n37105), .Z(n37103) );
  IV U39095 ( .A(n37104), .Z(n37105) );
  XNOR U39096 ( .A(m[544]), .B(n37106), .Z(n37104) );
  NAND U39097 ( .A(n37107), .B(mul_pow), .Z(n37106) );
  XOR U39098 ( .A(m[544]), .B(c[544]), .Z(n37107) );
  XOR U39099 ( .A(n37108), .B(n37109), .Z(n37100) );
  ANDN U39100 ( .B(n37110), .A(n31832), .Z(n37108) );
  XNOR U39101 ( .A(\modmult_1/zin[0][542] ), .B(n37111), .Z(n31832) );
  IV U39102 ( .A(n37109), .Z(n37111) );
  XOR U39103 ( .A(n37109), .B(n31833), .Z(n37110) );
  XNOR U39104 ( .A(n37112), .B(n37113), .Z(n31833) );
  ANDN U39105 ( .B(\modmult_1/xin[1023] ), .A(n37114), .Z(n37112) );
  IV U39106 ( .A(n37113), .Z(n37114) );
  XNOR U39107 ( .A(m[543]), .B(n37115), .Z(n37113) );
  NAND U39108 ( .A(n37116), .B(mul_pow), .Z(n37115) );
  XOR U39109 ( .A(m[543]), .B(c[543]), .Z(n37116) );
  XOR U39110 ( .A(n37117), .B(n37118), .Z(n37109) );
  ANDN U39111 ( .B(n37119), .A(n31830), .Z(n37117) );
  XNOR U39112 ( .A(\modmult_1/zin[0][541] ), .B(n37120), .Z(n31830) );
  IV U39113 ( .A(n37118), .Z(n37120) );
  XOR U39114 ( .A(n37118), .B(n31831), .Z(n37119) );
  XNOR U39115 ( .A(n37121), .B(n37122), .Z(n31831) );
  ANDN U39116 ( .B(\modmult_1/xin[1023] ), .A(n37123), .Z(n37121) );
  IV U39117 ( .A(n37122), .Z(n37123) );
  XNOR U39118 ( .A(m[542]), .B(n37124), .Z(n37122) );
  NAND U39119 ( .A(n37125), .B(mul_pow), .Z(n37124) );
  XOR U39120 ( .A(m[542]), .B(c[542]), .Z(n37125) );
  XOR U39121 ( .A(n37126), .B(n37127), .Z(n37118) );
  ANDN U39122 ( .B(n37128), .A(n31828), .Z(n37126) );
  XNOR U39123 ( .A(\modmult_1/zin[0][540] ), .B(n37129), .Z(n31828) );
  IV U39124 ( .A(n37127), .Z(n37129) );
  XOR U39125 ( .A(n37127), .B(n31829), .Z(n37128) );
  XNOR U39126 ( .A(n37130), .B(n37131), .Z(n31829) );
  ANDN U39127 ( .B(\modmult_1/xin[1023] ), .A(n37132), .Z(n37130) );
  IV U39128 ( .A(n37131), .Z(n37132) );
  XNOR U39129 ( .A(m[541]), .B(n37133), .Z(n37131) );
  NAND U39130 ( .A(n37134), .B(mul_pow), .Z(n37133) );
  XOR U39131 ( .A(m[541]), .B(c[541]), .Z(n37134) );
  XOR U39132 ( .A(n37135), .B(n37136), .Z(n37127) );
  ANDN U39133 ( .B(n37137), .A(n31826), .Z(n37135) );
  XNOR U39134 ( .A(\modmult_1/zin[0][539] ), .B(n37138), .Z(n31826) );
  IV U39135 ( .A(n37136), .Z(n37138) );
  XOR U39136 ( .A(n37136), .B(n31827), .Z(n37137) );
  XNOR U39137 ( .A(n37139), .B(n37140), .Z(n31827) );
  ANDN U39138 ( .B(\modmult_1/xin[1023] ), .A(n37141), .Z(n37139) );
  IV U39139 ( .A(n37140), .Z(n37141) );
  XNOR U39140 ( .A(m[540]), .B(n37142), .Z(n37140) );
  NAND U39141 ( .A(n37143), .B(mul_pow), .Z(n37142) );
  XOR U39142 ( .A(m[540]), .B(c[540]), .Z(n37143) );
  XOR U39143 ( .A(n37144), .B(n37145), .Z(n37136) );
  ANDN U39144 ( .B(n37146), .A(n31824), .Z(n37144) );
  XNOR U39145 ( .A(\modmult_1/zin[0][538] ), .B(n37147), .Z(n31824) );
  IV U39146 ( .A(n37145), .Z(n37147) );
  XOR U39147 ( .A(n37145), .B(n31825), .Z(n37146) );
  XNOR U39148 ( .A(n37148), .B(n37149), .Z(n31825) );
  ANDN U39149 ( .B(\modmult_1/xin[1023] ), .A(n37150), .Z(n37148) );
  IV U39150 ( .A(n37149), .Z(n37150) );
  XNOR U39151 ( .A(m[539]), .B(n37151), .Z(n37149) );
  NAND U39152 ( .A(n37152), .B(mul_pow), .Z(n37151) );
  XOR U39153 ( .A(m[539]), .B(c[539]), .Z(n37152) );
  XOR U39154 ( .A(n37153), .B(n37154), .Z(n37145) );
  ANDN U39155 ( .B(n37155), .A(n31822), .Z(n37153) );
  XNOR U39156 ( .A(\modmult_1/zin[0][537] ), .B(n37156), .Z(n31822) );
  IV U39157 ( .A(n37154), .Z(n37156) );
  XOR U39158 ( .A(n37154), .B(n31823), .Z(n37155) );
  XNOR U39159 ( .A(n37157), .B(n37158), .Z(n31823) );
  ANDN U39160 ( .B(\modmult_1/xin[1023] ), .A(n37159), .Z(n37157) );
  IV U39161 ( .A(n37158), .Z(n37159) );
  XNOR U39162 ( .A(m[538]), .B(n37160), .Z(n37158) );
  NAND U39163 ( .A(n37161), .B(mul_pow), .Z(n37160) );
  XOR U39164 ( .A(m[538]), .B(c[538]), .Z(n37161) );
  XOR U39165 ( .A(n37162), .B(n37163), .Z(n37154) );
  ANDN U39166 ( .B(n37164), .A(n31820), .Z(n37162) );
  XNOR U39167 ( .A(\modmult_1/zin[0][536] ), .B(n37165), .Z(n31820) );
  IV U39168 ( .A(n37163), .Z(n37165) );
  XOR U39169 ( .A(n37163), .B(n31821), .Z(n37164) );
  XNOR U39170 ( .A(n37166), .B(n37167), .Z(n31821) );
  ANDN U39171 ( .B(\modmult_1/xin[1023] ), .A(n37168), .Z(n37166) );
  IV U39172 ( .A(n37167), .Z(n37168) );
  XNOR U39173 ( .A(m[537]), .B(n37169), .Z(n37167) );
  NAND U39174 ( .A(n37170), .B(mul_pow), .Z(n37169) );
  XOR U39175 ( .A(m[537]), .B(c[537]), .Z(n37170) );
  XOR U39176 ( .A(n37171), .B(n37172), .Z(n37163) );
  ANDN U39177 ( .B(n37173), .A(n31818), .Z(n37171) );
  XNOR U39178 ( .A(\modmult_1/zin[0][535] ), .B(n37174), .Z(n31818) );
  IV U39179 ( .A(n37172), .Z(n37174) );
  XOR U39180 ( .A(n37172), .B(n31819), .Z(n37173) );
  XNOR U39181 ( .A(n37175), .B(n37176), .Z(n31819) );
  ANDN U39182 ( .B(\modmult_1/xin[1023] ), .A(n37177), .Z(n37175) );
  IV U39183 ( .A(n37176), .Z(n37177) );
  XNOR U39184 ( .A(m[536]), .B(n37178), .Z(n37176) );
  NAND U39185 ( .A(n37179), .B(mul_pow), .Z(n37178) );
  XOR U39186 ( .A(m[536]), .B(c[536]), .Z(n37179) );
  XOR U39187 ( .A(n37180), .B(n37181), .Z(n37172) );
  ANDN U39188 ( .B(n37182), .A(n31816), .Z(n37180) );
  XNOR U39189 ( .A(\modmult_1/zin[0][534] ), .B(n37183), .Z(n31816) );
  IV U39190 ( .A(n37181), .Z(n37183) );
  XOR U39191 ( .A(n37181), .B(n31817), .Z(n37182) );
  XNOR U39192 ( .A(n37184), .B(n37185), .Z(n31817) );
  ANDN U39193 ( .B(\modmult_1/xin[1023] ), .A(n37186), .Z(n37184) );
  IV U39194 ( .A(n37185), .Z(n37186) );
  XNOR U39195 ( .A(m[535]), .B(n37187), .Z(n37185) );
  NAND U39196 ( .A(n37188), .B(mul_pow), .Z(n37187) );
  XOR U39197 ( .A(m[535]), .B(c[535]), .Z(n37188) );
  XOR U39198 ( .A(n37189), .B(n37190), .Z(n37181) );
  ANDN U39199 ( .B(n37191), .A(n31814), .Z(n37189) );
  XNOR U39200 ( .A(\modmult_1/zin[0][533] ), .B(n37192), .Z(n31814) );
  IV U39201 ( .A(n37190), .Z(n37192) );
  XOR U39202 ( .A(n37190), .B(n31815), .Z(n37191) );
  XNOR U39203 ( .A(n37193), .B(n37194), .Z(n31815) );
  ANDN U39204 ( .B(\modmult_1/xin[1023] ), .A(n37195), .Z(n37193) );
  IV U39205 ( .A(n37194), .Z(n37195) );
  XNOR U39206 ( .A(m[534]), .B(n37196), .Z(n37194) );
  NAND U39207 ( .A(n37197), .B(mul_pow), .Z(n37196) );
  XOR U39208 ( .A(m[534]), .B(c[534]), .Z(n37197) );
  XOR U39209 ( .A(n37198), .B(n37199), .Z(n37190) );
  ANDN U39210 ( .B(n37200), .A(n31812), .Z(n37198) );
  XNOR U39211 ( .A(\modmult_1/zin[0][532] ), .B(n37201), .Z(n31812) );
  IV U39212 ( .A(n37199), .Z(n37201) );
  XOR U39213 ( .A(n37199), .B(n31813), .Z(n37200) );
  XNOR U39214 ( .A(n37202), .B(n37203), .Z(n31813) );
  ANDN U39215 ( .B(\modmult_1/xin[1023] ), .A(n37204), .Z(n37202) );
  IV U39216 ( .A(n37203), .Z(n37204) );
  XNOR U39217 ( .A(m[533]), .B(n37205), .Z(n37203) );
  NAND U39218 ( .A(n37206), .B(mul_pow), .Z(n37205) );
  XOR U39219 ( .A(m[533]), .B(c[533]), .Z(n37206) );
  XOR U39220 ( .A(n37207), .B(n37208), .Z(n37199) );
  ANDN U39221 ( .B(n37209), .A(n31810), .Z(n37207) );
  XNOR U39222 ( .A(\modmult_1/zin[0][531] ), .B(n37210), .Z(n31810) );
  IV U39223 ( .A(n37208), .Z(n37210) );
  XOR U39224 ( .A(n37208), .B(n31811), .Z(n37209) );
  XNOR U39225 ( .A(n37211), .B(n37212), .Z(n31811) );
  ANDN U39226 ( .B(\modmult_1/xin[1023] ), .A(n37213), .Z(n37211) );
  IV U39227 ( .A(n37212), .Z(n37213) );
  XNOR U39228 ( .A(m[532]), .B(n37214), .Z(n37212) );
  NAND U39229 ( .A(n37215), .B(mul_pow), .Z(n37214) );
  XOR U39230 ( .A(m[532]), .B(c[532]), .Z(n37215) );
  XOR U39231 ( .A(n37216), .B(n37217), .Z(n37208) );
  ANDN U39232 ( .B(n37218), .A(n31808), .Z(n37216) );
  XNOR U39233 ( .A(\modmult_1/zin[0][530] ), .B(n37219), .Z(n31808) );
  IV U39234 ( .A(n37217), .Z(n37219) );
  XOR U39235 ( .A(n37217), .B(n31809), .Z(n37218) );
  XNOR U39236 ( .A(n37220), .B(n37221), .Z(n31809) );
  ANDN U39237 ( .B(\modmult_1/xin[1023] ), .A(n37222), .Z(n37220) );
  IV U39238 ( .A(n37221), .Z(n37222) );
  XNOR U39239 ( .A(m[531]), .B(n37223), .Z(n37221) );
  NAND U39240 ( .A(n37224), .B(mul_pow), .Z(n37223) );
  XOR U39241 ( .A(m[531]), .B(c[531]), .Z(n37224) );
  XOR U39242 ( .A(n37225), .B(n37226), .Z(n37217) );
  ANDN U39243 ( .B(n37227), .A(n31806), .Z(n37225) );
  XNOR U39244 ( .A(\modmult_1/zin[0][529] ), .B(n37228), .Z(n31806) );
  IV U39245 ( .A(n37226), .Z(n37228) );
  XOR U39246 ( .A(n37226), .B(n31807), .Z(n37227) );
  XNOR U39247 ( .A(n37229), .B(n37230), .Z(n31807) );
  ANDN U39248 ( .B(\modmult_1/xin[1023] ), .A(n37231), .Z(n37229) );
  IV U39249 ( .A(n37230), .Z(n37231) );
  XNOR U39250 ( .A(m[530]), .B(n37232), .Z(n37230) );
  NAND U39251 ( .A(n37233), .B(mul_pow), .Z(n37232) );
  XOR U39252 ( .A(m[530]), .B(c[530]), .Z(n37233) );
  XOR U39253 ( .A(n37234), .B(n37235), .Z(n37226) );
  ANDN U39254 ( .B(n37236), .A(n31804), .Z(n37234) );
  XNOR U39255 ( .A(\modmult_1/zin[0][528] ), .B(n37237), .Z(n31804) );
  IV U39256 ( .A(n37235), .Z(n37237) );
  XOR U39257 ( .A(n37235), .B(n31805), .Z(n37236) );
  XNOR U39258 ( .A(n37238), .B(n37239), .Z(n31805) );
  ANDN U39259 ( .B(\modmult_1/xin[1023] ), .A(n37240), .Z(n37238) );
  IV U39260 ( .A(n37239), .Z(n37240) );
  XNOR U39261 ( .A(m[529]), .B(n37241), .Z(n37239) );
  NAND U39262 ( .A(n37242), .B(mul_pow), .Z(n37241) );
  XOR U39263 ( .A(m[529]), .B(c[529]), .Z(n37242) );
  XOR U39264 ( .A(n37243), .B(n37244), .Z(n37235) );
  ANDN U39265 ( .B(n37245), .A(n31802), .Z(n37243) );
  XNOR U39266 ( .A(\modmult_1/zin[0][527] ), .B(n37246), .Z(n31802) );
  IV U39267 ( .A(n37244), .Z(n37246) );
  XOR U39268 ( .A(n37244), .B(n31803), .Z(n37245) );
  XNOR U39269 ( .A(n37247), .B(n37248), .Z(n31803) );
  ANDN U39270 ( .B(\modmult_1/xin[1023] ), .A(n37249), .Z(n37247) );
  IV U39271 ( .A(n37248), .Z(n37249) );
  XNOR U39272 ( .A(m[528]), .B(n37250), .Z(n37248) );
  NAND U39273 ( .A(n37251), .B(mul_pow), .Z(n37250) );
  XOR U39274 ( .A(m[528]), .B(c[528]), .Z(n37251) );
  XOR U39275 ( .A(n37252), .B(n37253), .Z(n37244) );
  ANDN U39276 ( .B(n37254), .A(n31800), .Z(n37252) );
  XNOR U39277 ( .A(\modmult_1/zin[0][526] ), .B(n37255), .Z(n31800) );
  IV U39278 ( .A(n37253), .Z(n37255) );
  XOR U39279 ( .A(n37253), .B(n31801), .Z(n37254) );
  XNOR U39280 ( .A(n37256), .B(n37257), .Z(n31801) );
  ANDN U39281 ( .B(\modmult_1/xin[1023] ), .A(n37258), .Z(n37256) );
  IV U39282 ( .A(n37257), .Z(n37258) );
  XNOR U39283 ( .A(m[527]), .B(n37259), .Z(n37257) );
  NAND U39284 ( .A(n37260), .B(mul_pow), .Z(n37259) );
  XOR U39285 ( .A(m[527]), .B(c[527]), .Z(n37260) );
  XOR U39286 ( .A(n37261), .B(n37262), .Z(n37253) );
  ANDN U39287 ( .B(n37263), .A(n31798), .Z(n37261) );
  XNOR U39288 ( .A(\modmult_1/zin[0][525] ), .B(n37264), .Z(n31798) );
  IV U39289 ( .A(n37262), .Z(n37264) );
  XOR U39290 ( .A(n37262), .B(n31799), .Z(n37263) );
  XNOR U39291 ( .A(n37265), .B(n37266), .Z(n31799) );
  ANDN U39292 ( .B(\modmult_1/xin[1023] ), .A(n37267), .Z(n37265) );
  IV U39293 ( .A(n37266), .Z(n37267) );
  XNOR U39294 ( .A(m[526]), .B(n37268), .Z(n37266) );
  NAND U39295 ( .A(n37269), .B(mul_pow), .Z(n37268) );
  XOR U39296 ( .A(m[526]), .B(c[526]), .Z(n37269) );
  XOR U39297 ( .A(n37270), .B(n37271), .Z(n37262) );
  ANDN U39298 ( .B(n37272), .A(n31796), .Z(n37270) );
  XNOR U39299 ( .A(\modmult_1/zin[0][524] ), .B(n37273), .Z(n31796) );
  IV U39300 ( .A(n37271), .Z(n37273) );
  XOR U39301 ( .A(n37271), .B(n31797), .Z(n37272) );
  XNOR U39302 ( .A(n37274), .B(n37275), .Z(n31797) );
  ANDN U39303 ( .B(\modmult_1/xin[1023] ), .A(n37276), .Z(n37274) );
  IV U39304 ( .A(n37275), .Z(n37276) );
  XNOR U39305 ( .A(m[525]), .B(n37277), .Z(n37275) );
  NAND U39306 ( .A(n37278), .B(mul_pow), .Z(n37277) );
  XOR U39307 ( .A(m[525]), .B(c[525]), .Z(n37278) );
  XOR U39308 ( .A(n37279), .B(n37280), .Z(n37271) );
  ANDN U39309 ( .B(n37281), .A(n31794), .Z(n37279) );
  XNOR U39310 ( .A(\modmult_1/zin[0][523] ), .B(n37282), .Z(n31794) );
  IV U39311 ( .A(n37280), .Z(n37282) );
  XOR U39312 ( .A(n37280), .B(n31795), .Z(n37281) );
  XNOR U39313 ( .A(n37283), .B(n37284), .Z(n31795) );
  ANDN U39314 ( .B(\modmult_1/xin[1023] ), .A(n37285), .Z(n37283) );
  IV U39315 ( .A(n37284), .Z(n37285) );
  XNOR U39316 ( .A(m[524]), .B(n37286), .Z(n37284) );
  NAND U39317 ( .A(n37287), .B(mul_pow), .Z(n37286) );
  XOR U39318 ( .A(m[524]), .B(c[524]), .Z(n37287) );
  XOR U39319 ( .A(n37288), .B(n37289), .Z(n37280) );
  ANDN U39320 ( .B(n37290), .A(n31792), .Z(n37288) );
  XNOR U39321 ( .A(\modmult_1/zin[0][522] ), .B(n37291), .Z(n31792) );
  IV U39322 ( .A(n37289), .Z(n37291) );
  XOR U39323 ( .A(n37289), .B(n31793), .Z(n37290) );
  XNOR U39324 ( .A(n37292), .B(n37293), .Z(n31793) );
  ANDN U39325 ( .B(\modmult_1/xin[1023] ), .A(n37294), .Z(n37292) );
  IV U39326 ( .A(n37293), .Z(n37294) );
  XNOR U39327 ( .A(m[523]), .B(n37295), .Z(n37293) );
  NAND U39328 ( .A(n37296), .B(mul_pow), .Z(n37295) );
  XOR U39329 ( .A(m[523]), .B(c[523]), .Z(n37296) );
  XOR U39330 ( .A(n37297), .B(n37298), .Z(n37289) );
  ANDN U39331 ( .B(n37299), .A(n31790), .Z(n37297) );
  XNOR U39332 ( .A(\modmult_1/zin[0][521] ), .B(n37300), .Z(n31790) );
  IV U39333 ( .A(n37298), .Z(n37300) );
  XOR U39334 ( .A(n37298), .B(n31791), .Z(n37299) );
  XNOR U39335 ( .A(n37301), .B(n37302), .Z(n31791) );
  ANDN U39336 ( .B(\modmult_1/xin[1023] ), .A(n37303), .Z(n37301) );
  IV U39337 ( .A(n37302), .Z(n37303) );
  XNOR U39338 ( .A(m[522]), .B(n37304), .Z(n37302) );
  NAND U39339 ( .A(n37305), .B(mul_pow), .Z(n37304) );
  XOR U39340 ( .A(m[522]), .B(c[522]), .Z(n37305) );
  XOR U39341 ( .A(n37306), .B(n37307), .Z(n37298) );
  ANDN U39342 ( .B(n37308), .A(n31788), .Z(n37306) );
  XNOR U39343 ( .A(\modmult_1/zin[0][520] ), .B(n37309), .Z(n31788) );
  IV U39344 ( .A(n37307), .Z(n37309) );
  XOR U39345 ( .A(n37307), .B(n31789), .Z(n37308) );
  XNOR U39346 ( .A(n37310), .B(n37311), .Z(n31789) );
  ANDN U39347 ( .B(\modmult_1/xin[1023] ), .A(n37312), .Z(n37310) );
  IV U39348 ( .A(n37311), .Z(n37312) );
  XNOR U39349 ( .A(m[521]), .B(n37313), .Z(n37311) );
  NAND U39350 ( .A(n37314), .B(mul_pow), .Z(n37313) );
  XOR U39351 ( .A(m[521]), .B(c[521]), .Z(n37314) );
  XOR U39352 ( .A(n37315), .B(n37316), .Z(n37307) );
  ANDN U39353 ( .B(n37317), .A(n31786), .Z(n37315) );
  XNOR U39354 ( .A(\modmult_1/zin[0][519] ), .B(n37318), .Z(n31786) );
  IV U39355 ( .A(n37316), .Z(n37318) );
  XOR U39356 ( .A(n37316), .B(n31787), .Z(n37317) );
  XNOR U39357 ( .A(n37319), .B(n37320), .Z(n31787) );
  ANDN U39358 ( .B(\modmult_1/xin[1023] ), .A(n37321), .Z(n37319) );
  IV U39359 ( .A(n37320), .Z(n37321) );
  XNOR U39360 ( .A(m[520]), .B(n37322), .Z(n37320) );
  NAND U39361 ( .A(n37323), .B(mul_pow), .Z(n37322) );
  XOR U39362 ( .A(m[520]), .B(c[520]), .Z(n37323) );
  XOR U39363 ( .A(n37324), .B(n37325), .Z(n37316) );
  ANDN U39364 ( .B(n37326), .A(n31784), .Z(n37324) );
  XNOR U39365 ( .A(\modmult_1/zin[0][518] ), .B(n37327), .Z(n31784) );
  IV U39366 ( .A(n37325), .Z(n37327) );
  XOR U39367 ( .A(n37325), .B(n31785), .Z(n37326) );
  XNOR U39368 ( .A(n37328), .B(n37329), .Z(n31785) );
  ANDN U39369 ( .B(\modmult_1/xin[1023] ), .A(n37330), .Z(n37328) );
  IV U39370 ( .A(n37329), .Z(n37330) );
  XNOR U39371 ( .A(m[519]), .B(n37331), .Z(n37329) );
  NAND U39372 ( .A(n37332), .B(mul_pow), .Z(n37331) );
  XOR U39373 ( .A(m[519]), .B(c[519]), .Z(n37332) );
  XOR U39374 ( .A(n37333), .B(n37334), .Z(n37325) );
  ANDN U39375 ( .B(n37335), .A(n31782), .Z(n37333) );
  XNOR U39376 ( .A(\modmult_1/zin[0][517] ), .B(n37336), .Z(n31782) );
  IV U39377 ( .A(n37334), .Z(n37336) );
  XOR U39378 ( .A(n37334), .B(n31783), .Z(n37335) );
  XNOR U39379 ( .A(n37337), .B(n37338), .Z(n31783) );
  ANDN U39380 ( .B(\modmult_1/xin[1023] ), .A(n37339), .Z(n37337) );
  IV U39381 ( .A(n37338), .Z(n37339) );
  XNOR U39382 ( .A(m[518]), .B(n37340), .Z(n37338) );
  NAND U39383 ( .A(n37341), .B(mul_pow), .Z(n37340) );
  XOR U39384 ( .A(m[518]), .B(c[518]), .Z(n37341) );
  XOR U39385 ( .A(n37342), .B(n37343), .Z(n37334) );
  ANDN U39386 ( .B(n37344), .A(n31780), .Z(n37342) );
  XNOR U39387 ( .A(\modmult_1/zin[0][516] ), .B(n37345), .Z(n31780) );
  IV U39388 ( .A(n37343), .Z(n37345) );
  XOR U39389 ( .A(n37343), .B(n31781), .Z(n37344) );
  XNOR U39390 ( .A(n37346), .B(n37347), .Z(n31781) );
  ANDN U39391 ( .B(\modmult_1/xin[1023] ), .A(n37348), .Z(n37346) );
  IV U39392 ( .A(n37347), .Z(n37348) );
  XNOR U39393 ( .A(m[517]), .B(n37349), .Z(n37347) );
  NAND U39394 ( .A(n37350), .B(mul_pow), .Z(n37349) );
  XOR U39395 ( .A(m[517]), .B(c[517]), .Z(n37350) );
  XOR U39396 ( .A(n37351), .B(n37352), .Z(n37343) );
  ANDN U39397 ( .B(n37353), .A(n31778), .Z(n37351) );
  XNOR U39398 ( .A(\modmult_1/zin[0][515] ), .B(n37354), .Z(n31778) );
  IV U39399 ( .A(n37352), .Z(n37354) );
  XOR U39400 ( .A(n37352), .B(n31779), .Z(n37353) );
  XNOR U39401 ( .A(n37355), .B(n37356), .Z(n31779) );
  ANDN U39402 ( .B(\modmult_1/xin[1023] ), .A(n37357), .Z(n37355) );
  IV U39403 ( .A(n37356), .Z(n37357) );
  XNOR U39404 ( .A(m[516]), .B(n37358), .Z(n37356) );
  NAND U39405 ( .A(n37359), .B(mul_pow), .Z(n37358) );
  XOR U39406 ( .A(m[516]), .B(c[516]), .Z(n37359) );
  XOR U39407 ( .A(n37360), .B(n37361), .Z(n37352) );
  ANDN U39408 ( .B(n37362), .A(n31776), .Z(n37360) );
  XNOR U39409 ( .A(\modmult_1/zin[0][514] ), .B(n37363), .Z(n31776) );
  IV U39410 ( .A(n37361), .Z(n37363) );
  XOR U39411 ( .A(n37361), .B(n31777), .Z(n37362) );
  XNOR U39412 ( .A(n37364), .B(n37365), .Z(n31777) );
  ANDN U39413 ( .B(\modmult_1/xin[1023] ), .A(n37366), .Z(n37364) );
  IV U39414 ( .A(n37365), .Z(n37366) );
  XNOR U39415 ( .A(m[515]), .B(n37367), .Z(n37365) );
  NAND U39416 ( .A(n37368), .B(mul_pow), .Z(n37367) );
  XOR U39417 ( .A(m[515]), .B(c[515]), .Z(n37368) );
  XOR U39418 ( .A(n37369), .B(n37370), .Z(n37361) );
  ANDN U39419 ( .B(n37371), .A(n31774), .Z(n37369) );
  XNOR U39420 ( .A(\modmult_1/zin[0][513] ), .B(n37372), .Z(n31774) );
  IV U39421 ( .A(n37370), .Z(n37372) );
  XOR U39422 ( .A(n37370), .B(n31775), .Z(n37371) );
  XNOR U39423 ( .A(n37373), .B(n37374), .Z(n31775) );
  ANDN U39424 ( .B(\modmult_1/xin[1023] ), .A(n37375), .Z(n37373) );
  IV U39425 ( .A(n37374), .Z(n37375) );
  XNOR U39426 ( .A(m[514]), .B(n37376), .Z(n37374) );
  NAND U39427 ( .A(n37377), .B(mul_pow), .Z(n37376) );
  XOR U39428 ( .A(m[514]), .B(c[514]), .Z(n37377) );
  XOR U39429 ( .A(n37378), .B(n37379), .Z(n37370) );
  ANDN U39430 ( .B(n37380), .A(n31772), .Z(n37378) );
  XNOR U39431 ( .A(\modmult_1/zin[0][512] ), .B(n37381), .Z(n31772) );
  IV U39432 ( .A(n37379), .Z(n37381) );
  XOR U39433 ( .A(n37379), .B(n31773), .Z(n37380) );
  XNOR U39434 ( .A(n37382), .B(n37383), .Z(n31773) );
  ANDN U39435 ( .B(\modmult_1/xin[1023] ), .A(n37384), .Z(n37382) );
  IV U39436 ( .A(n37383), .Z(n37384) );
  XNOR U39437 ( .A(m[513]), .B(n37385), .Z(n37383) );
  NAND U39438 ( .A(n37386), .B(mul_pow), .Z(n37385) );
  XOR U39439 ( .A(m[513]), .B(c[513]), .Z(n37386) );
  XOR U39440 ( .A(n37387), .B(n37388), .Z(n37379) );
  ANDN U39441 ( .B(n37389), .A(n31770), .Z(n37387) );
  XNOR U39442 ( .A(\modmult_1/zin[0][511] ), .B(n37390), .Z(n31770) );
  IV U39443 ( .A(n37388), .Z(n37390) );
  XOR U39444 ( .A(n37388), .B(n31771), .Z(n37389) );
  XNOR U39445 ( .A(n37391), .B(n37392), .Z(n31771) );
  ANDN U39446 ( .B(\modmult_1/xin[1023] ), .A(n37393), .Z(n37391) );
  IV U39447 ( .A(n37392), .Z(n37393) );
  XNOR U39448 ( .A(m[512]), .B(n37394), .Z(n37392) );
  NAND U39449 ( .A(n37395), .B(mul_pow), .Z(n37394) );
  XOR U39450 ( .A(m[512]), .B(c[512]), .Z(n37395) );
  XOR U39451 ( .A(n37396), .B(n37397), .Z(n37388) );
  ANDN U39452 ( .B(n37398), .A(n31768), .Z(n37396) );
  XNOR U39453 ( .A(\modmult_1/zin[0][510] ), .B(n37399), .Z(n31768) );
  IV U39454 ( .A(n37397), .Z(n37399) );
  XOR U39455 ( .A(n37397), .B(n31769), .Z(n37398) );
  XNOR U39456 ( .A(n37400), .B(n37401), .Z(n31769) );
  ANDN U39457 ( .B(\modmult_1/xin[1023] ), .A(n37402), .Z(n37400) );
  IV U39458 ( .A(n37401), .Z(n37402) );
  XNOR U39459 ( .A(m[511]), .B(n37403), .Z(n37401) );
  NAND U39460 ( .A(n37404), .B(mul_pow), .Z(n37403) );
  XOR U39461 ( .A(m[511]), .B(c[511]), .Z(n37404) );
  XOR U39462 ( .A(n37405), .B(n37406), .Z(n37397) );
  ANDN U39463 ( .B(n37407), .A(n31766), .Z(n37405) );
  XNOR U39464 ( .A(\modmult_1/zin[0][509] ), .B(n37408), .Z(n31766) );
  IV U39465 ( .A(n37406), .Z(n37408) );
  XOR U39466 ( .A(n37406), .B(n31767), .Z(n37407) );
  XNOR U39467 ( .A(n37409), .B(n37410), .Z(n31767) );
  ANDN U39468 ( .B(\modmult_1/xin[1023] ), .A(n37411), .Z(n37409) );
  IV U39469 ( .A(n37410), .Z(n37411) );
  XNOR U39470 ( .A(m[510]), .B(n37412), .Z(n37410) );
  NAND U39471 ( .A(n37413), .B(mul_pow), .Z(n37412) );
  XOR U39472 ( .A(m[510]), .B(c[510]), .Z(n37413) );
  XOR U39473 ( .A(n37414), .B(n37415), .Z(n37406) );
  ANDN U39474 ( .B(n37416), .A(n31764), .Z(n37414) );
  XNOR U39475 ( .A(\modmult_1/zin[0][508] ), .B(n37417), .Z(n31764) );
  IV U39476 ( .A(n37415), .Z(n37417) );
  XOR U39477 ( .A(n37415), .B(n31765), .Z(n37416) );
  XNOR U39478 ( .A(n37418), .B(n37419), .Z(n31765) );
  ANDN U39479 ( .B(\modmult_1/xin[1023] ), .A(n37420), .Z(n37418) );
  IV U39480 ( .A(n37419), .Z(n37420) );
  XNOR U39481 ( .A(m[509]), .B(n37421), .Z(n37419) );
  NAND U39482 ( .A(n37422), .B(mul_pow), .Z(n37421) );
  XOR U39483 ( .A(m[509]), .B(c[509]), .Z(n37422) );
  XOR U39484 ( .A(n37423), .B(n37424), .Z(n37415) );
  ANDN U39485 ( .B(n37425), .A(n31762), .Z(n37423) );
  XNOR U39486 ( .A(\modmult_1/zin[0][507] ), .B(n37426), .Z(n31762) );
  IV U39487 ( .A(n37424), .Z(n37426) );
  XOR U39488 ( .A(n37424), .B(n31763), .Z(n37425) );
  XNOR U39489 ( .A(n37427), .B(n37428), .Z(n31763) );
  ANDN U39490 ( .B(\modmult_1/xin[1023] ), .A(n37429), .Z(n37427) );
  IV U39491 ( .A(n37428), .Z(n37429) );
  XNOR U39492 ( .A(m[508]), .B(n37430), .Z(n37428) );
  NAND U39493 ( .A(n37431), .B(mul_pow), .Z(n37430) );
  XOR U39494 ( .A(m[508]), .B(c[508]), .Z(n37431) );
  XOR U39495 ( .A(n37432), .B(n37433), .Z(n37424) );
  ANDN U39496 ( .B(n37434), .A(n31760), .Z(n37432) );
  XNOR U39497 ( .A(\modmult_1/zin[0][506] ), .B(n37435), .Z(n31760) );
  IV U39498 ( .A(n37433), .Z(n37435) );
  XOR U39499 ( .A(n37433), .B(n31761), .Z(n37434) );
  XNOR U39500 ( .A(n37436), .B(n37437), .Z(n31761) );
  ANDN U39501 ( .B(\modmult_1/xin[1023] ), .A(n37438), .Z(n37436) );
  IV U39502 ( .A(n37437), .Z(n37438) );
  XNOR U39503 ( .A(m[507]), .B(n37439), .Z(n37437) );
  NAND U39504 ( .A(n37440), .B(mul_pow), .Z(n37439) );
  XOR U39505 ( .A(m[507]), .B(c[507]), .Z(n37440) );
  XOR U39506 ( .A(n37441), .B(n37442), .Z(n37433) );
  ANDN U39507 ( .B(n37443), .A(n31758), .Z(n37441) );
  XNOR U39508 ( .A(\modmult_1/zin[0][505] ), .B(n37444), .Z(n31758) );
  IV U39509 ( .A(n37442), .Z(n37444) );
  XOR U39510 ( .A(n37442), .B(n31759), .Z(n37443) );
  XNOR U39511 ( .A(n37445), .B(n37446), .Z(n31759) );
  ANDN U39512 ( .B(\modmult_1/xin[1023] ), .A(n37447), .Z(n37445) );
  IV U39513 ( .A(n37446), .Z(n37447) );
  XNOR U39514 ( .A(m[506]), .B(n37448), .Z(n37446) );
  NAND U39515 ( .A(n37449), .B(mul_pow), .Z(n37448) );
  XOR U39516 ( .A(m[506]), .B(c[506]), .Z(n37449) );
  XOR U39517 ( .A(n37450), .B(n37451), .Z(n37442) );
  ANDN U39518 ( .B(n37452), .A(n31756), .Z(n37450) );
  XNOR U39519 ( .A(\modmult_1/zin[0][504] ), .B(n37453), .Z(n31756) );
  IV U39520 ( .A(n37451), .Z(n37453) );
  XOR U39521 ( .A(n37451), .B(n31757), .Z(n37452) );
  XNOR U39522 ( .A(n37454), .B(n37455), .Z(n31757) );
  ANDN U39523 ( .B(\modmult_1/xin[1023] ), .A(n37456), .Z(n37454) );
  IV U39524 ( .A(n37455), .Z(n37456) );
  XNOR U39525 ( .A(m[505]), .B(n37457), .Z(n37455) );
  NAND U39526 ( .A(n37458), .B(mul_pow), .Z(n37457) );
  XOR U39527 ( .A(m[505]), .B(c[505]), .Z(n37458) );
  XOR U39528 ( .A(n37459), .B(n37460), .Z(n37451) );
  ANDN U39529 ( .B(n37461), .A(n31754), .Z(n37459) );
  XNOR U39530 ( .A(\modmult_1/zin[0][503] ), .B(n37462), .Z(n31754) );
  IV U39531 ( .A(n37460), .Z(n37462) );
  XOR U39532 ( .A(n37460), .B(n31755), .Z(n37461) );
  XNOR U39533 ( .A(n37463), .B(n37464), .Z(n31755) );
  ANDN U39534 ( .B(\modmult_1/xin[1023] ), .A(n37465), .Z(n37463) );
  IV U39535 ( .A(n37464), .Z(n37465) );
  XNOR U39536 ( .A(m[504]), .B(n37466), .Z(n37464) );
  NAND U39537 ( .A(n37467), .B(mul_pow), .Z(n37466) );
  XOR U39538 ( .A(m[504]), .B(c[504]), .Z(n37467) );
  XOR U39539 ( .A(n37468), .B(n37469), .Z(n37460) );
  ANDN U39540 ( .B(n37470), .A(n31752), .Z(n37468) );
  XNOR U39541 ( .A(\modmult_1/zin[0][502] ), .B(n37471), .Z(n31752) );
  IV U39542 ( .A(n37469), .Z(n37471) );
  XOR U39543 ( .A(n37469), .B(n31753), .Z(n37470) );
  XNOR U39544 ( .A(n37472), .B(n37473), .Z(n31753) );
  ANDN U39545 ( .B(\modmult_1/xin[1023] ), .A(n37474), .Z(n37472) );
  IV U39546 ( .A(n37473), .Z(n37474) );
  XNOR U39547 ( .A(m[503]), .B(n37475), .Z(n37473) );
  NAND U39548 ( .A(n37476), .B(mul_pow), .Z(n37475) );
  XOR U39549 ( .A(m[503]), .B(c[503]), .Z(n37476) );
  XOR U39550 ( .A(n37477), .B(n37478), .Z(n37469) );
  ANDN U39551 ( .B(n37479), .A(n31750), .Z(n37477) );
  XNOR U39552 ( .A(\modmult_1/zin[0][501] ), .B(n37480), .Z(n31750) );
  IV U39553 ( .A(n37478), .Z(n37480) );
  XOR U39554 ( .A(n37478), .B(n31751), .Z(n37479) );
  XNOR U39555 ( .A(n37481), .B(n37482), .Z(n31751) );
  ANDN U39556 ( .B(\modmult_1/xin[1023] ), .A(n37483), .Z(n37481) );
  IV U39557 ( .A(n37482), .Z(n37483) );
  XNOR U39558 ( .A(m[502]), .B(n37484), .Z(n37482) );
  NAND U39559 ( .A(n37485), .B(mul_pow), .Z(n37484) );
  XOR U39560 ( .A(m[502]), .B(c[502]), .Z(n37485) );
  XOR U39561 ( .A(n37486), .B(n37487), .Z(n37478) );
  ANDN U39562 ( .B(n37488), .A(n31748), .Z(n37486) );
  XNOR U39563 ( .A(\modmult_1/zin[0][500] ), .B(n37489), .Z(n31748) );
  IV U39564 ( .A(n37487), .Z(n37489) );
  XOR U39565 ( .A(n37487), .B(n31749), .Z(n37488) );
  XNOR U39566 ( .A(n37490), .B(n37491), .Z(n31749) );
  ANDN U39567 ( .B(\modmult_1/xin[1023] ), .A(n37492), .Z(n37490) );
  IV U39568 ( .A(n37491), .Z(n37492) );
  XNOR U39569 ( .A(m[501]), .B(n37493), .Z(n37491) );
  NAND U39570 ( .A(n37494), .B(mul_pow), .Z(n37493) );
  XOR U39571 ( .A(m[501]), .B(c[501]), .Z(n37494) );
  XOR U39572 ( .A(n37495), .B(n37496), .Z(n37487) );
  ANDN U39573 ( .B(n37497), .A(n31746), .Z(n37495) );
  XNOR U39574 ( .A(\modmult_1/zin[0][499] ), .B(n37498), .Z(n31746) );
  IV U39575 ( .A(n37496), .Z(n37498) );
  XOR U39576 ( .A(n37496), .B(n31747), .Z(n37497) );
  XNOR U39577 ( .A(n37499), .B(n37500), .Z(n31747) );
  ANDN U39578 ( .B(\modmult_1/xin[1023] ), .A(n37501), .Z(n37499) );
  IV U39579 ( .A(n37500), .Z(n37501) );
  XNOR U39580 ( .A(m[500]), .B(n37502), .Z(n37500) );
  NAND U39581 ( .A(n37503), .B(mul_pow), .Z(n37502) );
  XOR U39582 ( .A(m[500]), .B(c[500]), .Z(n37503) );
  XOR U39583 ( .A(n37504), .B(n37505), .Z(n37496) );
  ANDN U39584 ( .B(n37506), .A(n31744), .Z(n37504) );
  XNOR U39585 ( .A(\modmult_1/zin[0][498] ), .B(n37507), .Z(n31744) );
  IV U39586 ( .A(n37505), .Z(n37507) );
  XOR U39587 ( .A(n37505), .B(n31745), .Z(n37506) );
  XNOR U39588 ( .A(n37508), .B(n37509), .Z(n31745) );
  ANDN U39589 ( .B(\modmult_1/xin[1023] ), .A(n37510), .Z(n37508) );
  IV U39590 ( .A(n37509), .Z(n37510) );
  XNOR U39591 ( .A(m[499]), .B(n37511), .Z(n37509) );
  NAND U39592 ( .A(n37512), .B(mul_pow), .Z(n37511) );
  XOR U39593 ( .A(m[499]), .B(c[499]), .Z(n37512) );
  XOR U39594 ( .A(n37513), .B(n37514), .Z(n37505) );
  ANDN U39595 ( .B(n37515), .A(n31742), .Z(n37513) );
  XNOR U39596 ( .A(\modmult_1/zin[0][497] ), .B(n37516), .Z(n31742) );
  IV U39597 ( .A(n37514), .Z(n37516) );
  XOR U39598 ( .A(n37514), .B(n31743), .Z(n37515) );
  XNOR U39599 ( .A(n37517), .B(n37518), .Z(n31743) );
  ANDN U39600 ( .B(\modmult_1/xin[1023] ), .A(n37519), .Z(n37517) );
  IV U39601 ( .A(n37518), .Z(n37519) );
  XNOR U39602 ( .A(m[498]), .B(n37520), .Z(n37518) );
  NAND U39603 ( .A(n37521), .B(mul_pow), .Z(n37520) );
  XOR U39604 ( .A(m[498]), .B(c[498]), .Z(n37521) );
  XOR U39605 ( .A(n37522), .B(n37523), .Z(n37514) );
  ANDN U39606 ( .B(n37524), .A(n31740), .Z(n37522) );
  XNOR U39607 ( .A(\modmult_1/zin[0][496] ), .B(n37525), .Z(n31740) );
  IV U39608 ( .A(n37523), .Z(n37525) );
  XOR U39609 ( .A(n37523), .B(n31741), .Z(n37524) );
  XNOR U39610 ( .A(n37526), .B(n37527), .Z(n31741) );
  ANDN U39611 ( .B(\modmult_1/xin[1023] ), .A(n37528), .Z(n37526) );
  IV U39612 ( .A(n37527), .Z(n37528) );
  XNOR U39613 ( .A(m[497]), .B(n37529), .Z(n37527) );
  NAND U39614 ( .A(n37530), .B(mul_pow), .Z(n37529) );
  XOR U39615 ( .A(m[497]), .B(c[497]), .Z(n37530) );
  XOR U39616 ( .A(n37531), .B(n37532), .Z(n37523) );
  ANDN U39617 ( .B(n37533), .A(n31738), .Z(n37531) );
  XNOR U39618 ( .A(\modmult_1/zin[0][495] ), .B(n37534), .Z(n31738) );
  IV U39619 ( .A(n37532), .Z(n37534) );
  XOR U39620 ( .A(n37532), .B(n31739), .Z(n37533) );
  XNOR U39621 ( .A(n37535), .B(n37536), .Z(n31739) );
  ANDN U39622 ( .B(\modmult_1/xin[1023] ), .A(n37537), .Z(n37535) );
  IV U39623 ( .A(n37536), .Z(n37537) );
  XNOR U39624 ( .A(m[496]), .B(n37538), .Z(n37536) );
  NAND U39625 ( .A(n37539), .B(mul_pow), .Z(n37538) );
  XOR U39626 ( .A(m[496]), .B(c[496]), .Z(n37539) );
  XOR U39627 ( .A(n37540), .B(n37541), .Z(n37532) );
  ANDN U39628 ( .B(n37542), .A(n31736), .Z(n37540) );
  XNOR U39629 ( .A(\modmult_1/zin[0][494] ), .B(n37543), .Z(n31736) );
  IV U39630 ( .A(n37541), .Z(n37543) );
  XOR U39631 ( .A(n37541), .B(n31737), .Z(n37542) );
  XNOR U39632 ( .A(n37544), .B(n37545), .Z(n31737) );
  ANDN U39633 ( .B(\modmult_1/xin[1023] ), .A(n37546), .Z(n37544) );
  IV U39634 ( .A(n37545), .Z(n37546) );
  XNOR U39635 ( .A(m[495]), .B(n37547), .Z(n37545) );
  NAND U39636 ( .A(n37548), .B(mul_pow), .Z(n37547) );
  XOR U39637 ( .A(m[495]), .B(c[495]), .Z(n37548) );
  XOR U39638 ( .A(n37549), .B(n37550), .Z(n37541) );
  ANDN U39639 ( .B(n37551), .A(n31734), .Z(n37549) );
  XNOR U39640 ( .A(\modmult_1/zin[0][493] ), .B(n37552), .Z(n31734) );
  IV U39641 ( .A(n37550), .Z(n37552) );
  XOR U39642 ( .A(n37550), .B(n31735), .Z(n37551) );
  XNOR U39643 ( .A(n37553), .B(n37554), .Z(n31735) );
  ANDN U39644 ( .B(\modmult_1/xin[1023] ), .A(n37555), .Z(n37553) );
  IV U39645 ( .A(n37554), .Z(n37555) );
  XNOR U39646 ( .A(m[494]), .B(n37556), .Z(n37554) );
  NAND U39647 ( .A(n37557), .B(mul_pow), .Z(n37556) );
  XOR U39648 ( .A(m[494]), .B(c[494]), .Z(n37557) );
  XOR U39649 ( .A(n37558), .B(n37559), .Z(n37550) );
  ANDN U39650 ( .B(n37560), .A(n31732), .Z(n37558) );
  XNOR U39651 ( .A(\modmult_1/zin[0][492] ), .B(n37561), .Z(n31732) );
  IV U39652 ( .A(n37559), .Z(n37561) );
  XOR U39653 ( .A(n37559), .B(n31733), .Z(n37560) );
  XNOR U39654 ( .A(n37562), .B(n37563), .Z(n31733) );
  ANDN U39655 ( .B(\modmult_1/xin[1023] ), .A(n37564), .Z(n37562) );
  IV U39656 ( .A(n37563), .Z(n37564) );
  XNOR U39657 ( .A(m[493]), .B(n37565), .Z(n37563) );
  NAND U39658 ( .A(n37566), .B(mul_pow), .Z(n37565) );
  XOR U39659 ( .A(m[493]), .B(c[493]), .Z(n37566) );
  XOR U39660 ( .A(n37567), .B(n37568), .Z(n37559) );
  ANDN U39661 ( .B(n37569), .A(n31730), .Z(n37567) );
  XNOR U39662 ( .A(\modmult_1/zin[0][491] ), .B(n37570), .Z(n31730) );
  IV U39663 ( .A(n37568), .Z(n37570) );
  XOR U39664 ( .A(n37568), .B(n31731), .Z(n37569) );
  XNOR U39665 ( .A(n37571), .B(n37572), .Z(n31731) );
  ANDN U39666 ( .B(\modmult_1/xin[1023] ), .A(n37573), .Z(n37571) );
  IV U39667 ( .A(n37572), .Z(n37573) );
  XNOR U39668 ( .A(m[492]), .B(n37574), .Z(n37572) );
  NAND U39669 ( .A(n37575), .B(mul_pow), .Z(n37574) );
  XOR U39670 ( .A(m[492]), .B(c[492]), .Z(n37575) );
  XOR U39671 ( .A(n37576), .B(n37577), .Z(n37568) );
  ANDN U39672 ( .B(n37578), .A(n31728), .Z(n37576) );
  XNOR U39673 ( .A(\modmult_1/zin[0][490] ), .B(n37579), .Z(n31728) );
  IV U39674 ( .A(n37577), .Z(n37579) );
  XOR U39675 ( .A(n37577), .B(n31729), .Z(n37578) );
  XNOR U39676 ( .A(n37580), .B(n37581), .Z(n31729) );
  ANDN U39677 ( .B(\modmult_1/xin[1023] ), .A(n37582), .Z(n37580) );
  IV U39678 ( .A(n37581), .Z(n37582) );
  XNOR U39679 ( .A(m[491]), .B(n37583), .Z(n37581) );
  NAND U39680 ( .A(n37584), .B(mul_pow), .Z(n37583) );
  XOR U39681 ( .A(m[491]), .B(c[491]), .Z(n37584) );
  XOR U39682 ( .A(n37585), .B(n37586), .Z(n37577) );
  ANDN U39683 ( .B(n37587), .A(n31726), .Z(n37585) );
  XNOR U39684 ( .A(\modmult_1/zin[0][489] ), .B(n37588), .Z(n31726) );
  IV U39685 ( .A(n37586), .Z(n37588) );
  XOR U39686 ( .A(n37586), .B(n31727), .Z(n37587) );
  XNOR U39687 ( .A(n37589), .B(n37590), .Z(n31727) );
  ANDN U39688 ( .B(\modmult_1/xin[1023] ), .A(n37591), .Z(n37589) );
  IV U39689 ( .A(n37590), .Z(n37591) );
  XNOR U39690 ( .A(m[490]), .B(n37592), .Z(n37590) );
  NAND U39691 ( .A(n37593), .B(mul_pow), .Z(n37592) );
  XOR U39692 ( .A(m[490]), .B(c[490]), .Z(n37593) );
  XOR U39693 ( .A(n37594), .B(n37595), .Z(n37586) );
  ANDN U39694 ( .B(n37596), .A(n31724), .Z(n37594) );
  XNOR U39695 ( .A(\modmult_1/zin[0][488] ), .B(n37597), .Z(n31724) );
  IV U39696 ( .A(n37595), .Z(n37597) );
  XOR U39697 ( .A(n37595), .B(n31725), .Z(n37596) );
  XNOR U39698 ( .A(n37598), .B(n37599), .Z(n31725) );
  ANDN U39699 ( .B(\modmult_1/xin[1023] ), .A(n37600), .Z(n37598) );
  IV U39700 ( .A(n37599), .Z(n37600) );
  XNOR U39701 ( .A(m[489]), .B(n37601), .Z(n37599) );
  NAND U39702 ( .A(n37602), .B(mul_pow), .Z(n37601) );
  XOR U39703 ( .A(m[489]), .B(c[489]), .Z(n37602) );
  XOR U39704 ( .A(n37603), .B(n37604), .Z(n37595) );
  ANDN U39705 ( .B(n37605), .A(n31722), .Z(n37603) );
  XNOR U39706 ( .A(\modmult_1/zin[0][487] ), .B(n37606), .Z(n31722) );
  IV U39707 ( .A(n37604), .Z(n37606) );
  XOR U39708 ( .A(n37604), .B(n31723), .Z(n37605) );
  XNOR U39709 ( .A(n37607), .B(n37608), .Z(n31723) );
  ANDN U39710 ( .B(\modmult_1/xin[1023] ), .A(n37609), .Z(n37607) );
  IV U39711 ( .A(n37608), .Z(n37609) );
  XNOR U39712 ( .A(m[488]), .B(n37610), .Z(n37608) );
  NAND U39713 ( .A(n37611), .B(mul_pow), .Z(n37610) );
  XOR U39714 ( .A(m[488]), .B(c[488]), .Z(n37611) );
  XOR U39715 ( .A(n37612), .B(n37613), .Z(n37604) );
  ANDN U39716 ( .B(n37614), .A(n31720), .Z(n37612) );
  XNOR U39717 ( .A(\modmult_1/zin[0][486] ), .B(n37615), .Z(n31720) );
  IV U39718 ( .A(n37613), .Z(n37615) );
  XOR U39719 ( .A(n37613), .B(n31721), .Z(n37614) );
  XNOR U39720 ( .A(n37616), .B(n37617), .Z(n31721) );
  ANDN U39721 ( .B(\modmult_1/xin[1023] ), .A(n37618), .Z(n37616) );
  IV U39722 ( .A(n37617), .Z(n37618) );
  XNOR U39723 ( .A(m[487]), .B(n37619), .Z(n37617) );
  NAND U39724 ( .A(n37620), .B(mul_pow), .Z(n37619) );
  XOR U39725 ( .A(m[487]), .B(c[487]), .Z(n37620) );
  XOR U39726 ( .A(n37621), .B(n37622), .Z(n37613) );
  ANDN U39727 ( .B(n37623), .A(n31718), .Z(n37621) );
  XNOR U39728 ( .A(\modmult_1/zin[0][485] ), .B(n37624), .Z(n31718) );
  IV U39729 ( .A(n37622), .Z(n37624) );
  XOR U39730 ( .A(n37622), .B(n31719), .Z(n37623) );
  XNOR U39731 ( .A(n37625), .B(n37626), .Z(n31719) );
  ANDN U39732 ( .B(\modmult_1/xin[1023] ), .A(n37627), .Z(n37625) );
  IV U39733 ( .A(n37626), .Z(n37627) );
  XNOR U39734 ( .A(m[486]), .B(n37628), .Z(n37626) );
  NAND U39735 ( .A(n37629), .B(mul_pow), .Z(n37628) );
  XOR U39736 ( .A(m[486]), .B(c[486]), .Z(n37629) );
  XOR U39737 ( .A(n37630), .B(n37631), .Z(n37622) );
  ANDN U39738 ( .B(n37632), .A(n31716), .Z(n37630) );
  XNOR U39739 ( .A(\modmult_1/zin[0][484] ), .B(n37633), .Z(n31716) );
  IV U39740 ( .A(n37631), .Z(n37633) );
  XOR U39741 ( .A(n37631), .B(n31717), .Z(n37632) );
  XNOR U39742 ( .A(n37634), .B(n37635), .Z(n31717) );
  ANDN U39743 ( .B(\modmult_1/xin[1023] ), .A(n37636), .Z(n37634) );
  IV U39744 ( .A(n37635), .Z(n37636) );
  XNOR U39745 ( .A(m[485]), .B(n37637), .Z(n37635) );
  NAND U39746 ( .A(n37638), .B(mul_pow), .Z(n37637) );
  XOR U39747 ( .A(m[485]), .B(c[485]), .Z(n37638) );
  XOR U39748 ( .A(n37639), .B(n37640), .Z(n37631) );
  ANDN U39749 ( .B(n37641), .A(n31714), .Z(n37639) );
  XNOR U39750 ( .A(\modmult_1/zin[0][483] ), .B(n37642), .Z(n31714) );
  IV U39751 ( .A(n37640), .Z(n37642) );
  XOR U39752 ( .A(n37640), .B(n31715), .Z(n37641) );
  XNOR U39753 ( .A(n37643), .B(n37644), .Z(n31715) );
  ANDN U39754 ( .B(\modmult_1/xin[1023] ), .A(n37645), .Z(n37643) );
  IV U39755 ( .A(n37644), .Z(n37645) );
  XNOR U39756 ( .A(m[484]), .B(n37646), .Z(n37644) );
  NAND U39757 ( .A(n37647), .B(mul_pow), .Z(n37646) );
  XOR U39758 ( .A(m[484]), .B(c[484]), .Z(n37647) );
  XOR U39759 ( .A(n37648), .B(n37649), .Z(n37640) );
  ANDN U39760 ( .B(n37650), .A(n31712), .Z(n37648) );
  XNOR U39761 ( .A(\modmult_1/zin[0][482] ), .B(n37651), .Z(n31712) );
  IV U39762 ( .A(n37649), .Z(n37651) );
  XOR U39763 ( .A(n37649), .B(n31713), .Z(n37650) );
  XNOR U39764 ( .A(n37652), .B(n37653), .Z(n31713) );
  ANDN U39765 ( .B(\modmult_1/xin[1023] ), .A(n37654), .Z(n37652) );
  IV U39766 ( .A(n37653), .Z(n37654) );
  XNOR U39767 ( .A(m[483]), .B(n37655), .Z(n37653) );
  NAND U39768 ( .A(n37656), .B(mul_pow), .Z(n37655) );
  XOR U39769 ( .A(m[483]), .B(c[483]), .Z(n37656) );
  XOR U39770 ( .A(n37657), .B(n37658), .Z(n37649) );
  ANDN U39771 ( .B(n37659), .A(n31710), .Z(n37657) );
  XNOR U39772 ( .A(\modmult_1/zin[0][481] ), .B(n37660), .Z(n31710) );
  IV U39773 ( .A(n37658), .Z(n37660) );
  XOR U39774 ( .A(n37658), .B(n31711), .Z(n37659) );
  XNOR U39775 ( .A(n37661), .B(n37662), .Z(n31711) );
  ANDN U39776 ( .B(\modmult_1/xin[1023] ), .A(n37663), .Z(n37661) );
  IV U39777 ( .A(n37662), .Z(n37663) );
  XNOR U39778 ( .A(m[482]), .B(n37664), .Z(n37662) );
  NAND U39779 ( .A(n37665), .B(mul_pow), .Z(n37664) );
  XOR U39780 ( .A(m[482]), .B(c[482]), .Z(n37665) );
  XOR U39781 ( .A(n37666), .B(n37667), .Z(n37658) );
  ANDN U39782 ( .B(n37668), .A(n31708), .Z(n37666) );
  XNOR U39783 ( .A(\modmult_1/zin[0][480] ), .B(n37669), .Z(n31708) );
  IV U39784 ( .A(n37667), .Z(n37669) );
  XOR U39785 ( .A(n37667), .B(n31709), .Z(n37668) );
  XNOR U39786 ( .A(n37670), .B(n37671), .Z(n31709) );
  ANDN U39787 ( .B(\modmult_1/xin[1023] ), .A(n37672), .Z(n37670) );
  IV U39788 ( .A(n37671), .Z(n37672) );
  XNOR U39789 ( .A(m[481]), .B(n37673), .Z(n37671) );
  NAND U39790 ( .A(n37674), .B(mul_pow), .Z(n37673) );
  XOR U39791 ( .A(m[481]), .B(c[481]), .Z(n37674) );
  XOR U39792 ( .A(n37675), .B(n37676), .Z(n37667) );
  ANDN U39793 ( .B(n37677), .A(n31706), .Z(n37675) );
  XNOR U39794 ( .A(\modmult_1/zin[0][479] ), .B(n37678), .Z(n31706) );
  IV U39795 ( .A(n37676), .Z(n37678) );
  XOR U39796 ( .A(n37676), .B(n31707), .Z(n37677) );
  XNOR U39797 ( .A(n37679), .B(n37680), .Z(n31707) );
  ANDN U39798 ( .B(\modmult_1/xin[1023] ), .A(n37681), .Z(n37679) );
  IV U39799 ( .A(n37680), .Z(n37681) );
  XNOR U39800 ( .A(m[480]), .B(n37682), .Z(n37680) );
  NAND U39801 ( .A(n37683), .B(mul_pow), .Z(n37682) );
  XOR U39802 ( .A(m[480]), .B(c[480]), .Z(n37683) );
  XOR U39803 ( .A(n37684), .B(n37685), .Z(n37676) );
  ANDN U39804 ( .B(n37686), .A(n31704), .Z(n37684) );
  XNOR U39805 ( .A(\modmult_1/zin[0][478] ), .B(n37687), .Z(n31704) );
  IV U39806 ( .A(n37685), .Z(n37687) );
  XOR U39807 ( .A(n37685), .B(n31705), .Z(n37686) );
  XNOR U39808 ( .A(n37688), .B(n37689), .Z(n31705) );
  ANDN U39809 ( .B(\modmult_1/xin[1023] ), .A(n37690), .Z(n37688) );
  IV U39810 ( .A(n37689), .Z(n37690) );
  XNOR U39811 ( .A(m[479]), .B(n37691), .Z(n37689) );
  NAND U39812 ( .A(n37692), .B(mul_pow), .Z(n37691) );
  XOR U39813 ( .A(m[479]), .B(c[479]), .Z(n37692) );
  XOR U39814 ( .A(n37693), .B(n37694), .Z(n37685) );
  ANDN U39815 ( .B(n37695), .A(n31702), .Z(n37693) );
  XNOR U39816 ( .A(\modmult_1/zin[0][477] ), .B(n37696), .Z(n31702) );
  IV U39817 ( .A(n37694), .Z(n37696) );
  XOR U39818 ( .A(n37694), .B(n31703), .Z(n37695) );
  XNOR U39819 ( .A(n37697), .B(n37698), .Z(n31703) );
  ANDN U39820 ( .B(\modmult_1/xin[1023] ), .A(n37699), .Z(n37697) );
  IV U39821 ( .A(n37698), .Z(n37699) );
  XNOR U39822 ( .A(m[478]), .B(n37700), .Z(n37698) );
  NAND U39823 ( .A(n37701), .B(mul_pow), .Z(n37700) );
  XOR U39824 ( .A(m[478]), .B(c[478]), .Z(n37701) );
  XOR U39825 ( .A(n37702), .B(n37703), .Z(n37694) );
  ANDN U39826 ( .B(n37704), .A(n31700), .Z(n37702) );
  XNOR U39827 ( .A(\modmult_1/zin[0][476] ), .B(n37705), .Z(n31700) );
  IV U39828 ( .A(n37703), .Z(n37705) );
  XOR U39829 ( .A(n37703), .B(n31701), .Z(n37704) );
  XNOR U39830 ( .A(n37706), .B(n37707), .Z(n31701) );
  ANDN U39831 ( .B(\modmult_1/xin[1023] ), .A(n37708), .Z(n37706) );
  IV U39832 ( .A(n37707), .Z(n37708) );
  XNOR U39833 ( .A(m[477]), .B(n37709), .Z(n37707) );
  NAND U39834 ( .A(n37710), .B(mul_pow), .Z(n37709) );
  XOR U39835 ( .A(m[477]), .B(c[477]), .Z(n37710) );
  XOR U39836 ( .A(n37711), .B(n37712), .Z(n37703) );
  ANDN U39837 ( .B(n37713), .A(n31698), .Z(n37711) );
  XNOR U39838 ( .A(\modmult_1/zin[0][475] ), .B(n37714), .Z(n31698) );
  IV U39839 ( .A(n37712), .Z(n37714) );
  XOR U39840 ( .A(n37712), .B(n31699), .Z(n37713) );
  XNOR U39841 ( .A(n37715), .B(n37716), .Z(n31699) );
  ANDN U39842 ( .B(\modmult_1/xin[1023] ), .A(n37717), .Z(n37715) );
  IV U39843 ( .A(n37716), .Z(n37717) );
  XNOR U39844 ( .A(m[476]), .B(n37718), .Z(n37716) );
  NAND U39845 ( .A(n37719), .B(mul_pow), .Z(n37718) );
  XOR U39846 ( .A(m[476]), .B(c[476]), .Z(n37719) );
  XOR U39847 ( .A(n37720), .B(n37721), .Z(n37712) );
  ANDN U39848 ( .B(n37722), .A(n31696), .Z(n37720) );
  XNOR U39849 ( .A(\modmult_1/zin[0][474] ), .B(n37723), .Z(n31696) );
  IV U39850 ( .A(n37721), .Z(n37723) );
  XOR U39851 ( .A(n37721), .B(n31697), .Z(n37722) );
  XNOR U39852 ( .A(n37724), .B(n37725), .Z(n31697) );
  ANDN U39853 ( .B(\modmult_1/xin[1023] ), .A(n37726), .Z(n37724) );
  IV U39854 ( .A(n37725), .Z(n37726) );
  XNOR U39855 ( .A(m[475]), .B(n37727), .Z(n37725) );
  NAND U39856 ( .A(n37728), .B(mul_pow), .Z(n37727) );
  XOR U39857 ( .A(m[475]), .B(c[475]), .Z(n37728) );
  XOR U39858 ( .A(n37729), .B(n37730), .Z(n37721) );
  ANDN U39859 ( .B(n37731), .A(n31694), .Z(n37729) );
  XNOR U39860 ( .A(\modmult_1/zin[0][473] ), .B(n37732), .Z(n31694) );
  IV U39861 ( .A(n37730), .Z(n37732) );
  XOR U39862 ( .A(n37730), .B(n31695), .Z(n37731) );
  XNOR U39863 ( .A(n37733), .B(n37734), .Z(n31695) );
  ANDN U39864 ( .B(\modmult_1/xin[1023] ), .A(n37735), .Z(n37733) );
  IV U39865 ( .A(n37734), .Z(n37735) );
  XNOR U39866 ( .A(m[474]), .B(n37736), .Z(n37734) );
  NAND U39867 ( .A(n37737), .B(mul_pow), .Z(n37736) );
  XOR U39868 ( .A(m[474]), .B(c[474]), .Z(n37737) );
  XOR U39869 ( .A(n37738), .B(n37739), .Z(n37730) );
  ANDN U39870 ( .B(n37740), .A(n31692), .Z(n37738) );
  XNOR U39871 ( .A(\modmult_1/zin[0][472] ), .B(n37741), .Z(n31692) );
  IV U39872 ( .A(n37739), .Z(n37741) );
  XOR U39873 ( .A(n37739), .B(n31693), .Z(n37740) );
  XNOR U39874 ( .A(n37742), .B(n37743), .Z(n31693) );
  ANDN U39875 ( .B(\modmult_1/xin[1023] ), .A(n37744), .Z(n37742) );
  IV U39876 ( .A(n37743), .Z(n37744) );
  XNOR U39877 ( .A(m[473]), .B(n37745), .Z(n37743) );
  NAND U39878 ( .A(n37746), .B(mul_pow), .Z(n37745) );
  XOR U39879 ( .A(m[473]), .B(c[473]), .Z(n37746) );
  XOR U39880 ( .A(n37747), .B(n37748), .Z(n37739) );
  ANDN U39881 ( .B(n37749), .A(n31690), .Z(n37747) );
  XNOR U39882 ( .A(\modmult_1/zin[0][471] ), .B(n37750), .Z(n31690) );
  IV U39883 ( .A(n37748), .Z(n37750) );
  XOR U39884 ( .A(n37748), .B(n31691), .Z(n37749) );
  XNOR U39885 ( .A(n37751), .B(n37752), .Z(n31691) );
  ANDN U39886 ( .B(\modmult_1/xin[1023] ), .A(n37753), .Z(n37751) );
  IV U39887 ( .A(n37752), .Z(n37753) );
  XNOR U39888 ( .A(m[472]), .B(n37754), .Z(n37752) );
  NAND U39889 ( .A(n37755), .B(mul_pow), .Z(n37754) );
  XOR U39890 ( .A(m[472]), .B(c[472]), .Z(n37755) );
  XOR U39891 ( .A(n37756), .B(n37757), .Z(n37748) );
  ANDN U39892 ( .B(n37758), .A(n31688), .Z(n37756) );
  XNOR U39893 ( .A(\modmult_1/zin[0][470] ), .B(n37759), .Z(n31688) );
  IV U39894 ( .A(n37757), .Z(n37759) );
  XOR U39895 ( .A(n37757), .B(n31689), .Z(n37758) );
  XNOR U39896 ( .A(n37760), .B(n37761), .Z(n31689) );
  ANDN U39897 ( .B(\modmult_1/xin[1023] ), .A(n37762), .Z(n37760) );
  IV U39898 ( .A(n37761), .Z(n37762) );
  XNOR U39899 ( .A(m[471]), .B(n37763), .Z(n37761) );
  NAND U39900 ( .A(n37764), .B(mul_pow), .Z(n37763) );
  XOR U39901 ( .A(m[471]), .B(c[471]), .Z(n37764) );
  XOR U39902 ( .A(n37765), .B(n37766), .Z(n37757) );
  ANDN U39903 ( .B(n37767), .A(n31686), .Z(n37765) );
  XNOR U39904 ( .A(\modmult_1/zin[0][469] ), .B(n37768), .Z(n31686) );
  IV U39905 ( .A(n37766), .Z(n37768) );
  XOR U39906 ( .A(n37766), .B(n31687), .Z(n37767) );
  XNOR U39907 ( .A(n37769), .B(n37770), .Z(n31687) );
  ANDN U39908 ( .B(\modmult_1/xin[1023] ), .A(n37771), .Z(n37769) );
  IV U39909 ( .A(n37770), .Z(n37771) );
  XNOR U39910 ( .A(m[470]), .B(n37772), .Z(n37770) );
  NAND U39911 ( .A(n37773), .B(mul_pow), .Z(n37772) );
  XOR U39912 ( .A(m[470]), .B(c[470]), .Z(n37773) );
  XOR U39913 ( .A(n37774), .B(n37775), .Z(n37766) );
  ANDN U39914 ( .B(n37776), .A(n31684), .Z(n37774) );
  XNOR U39915 ( .A(\modmult_1/zin[0][468] ), .B(n37777), .Z(n31684) );
  IV U39916 ( .A(n37775), .Z(n37777) );
  XOR U39917 ( .A(n37775), .B(n31685), .Z(n37776) );
  XNOR U39918 ( .A(n37778), .B(n37779), .Z(n31685) );
  ANDN U39919 ( .B(\modmult_1/xin[1023] ), .A(n37780), .Z(n37778) );
  IV U39920 ( .A(n37779), .Z(n37780) );
  XNOR U39921 ( .A(m[469]), .B(n37781), .Z(n37779) );
  NAND U39922 ( .A(n37782), .B(mul_pow), .Z(n37781) );
  XOR U39923 ( .A(m[469]), .B(c[469]), .Z(n37782) );
  XOR U39924 ( .A(n37783), .B(n37784), .Z(n37775) );
  ANDN U39925 ( .B(n37785), .A(n31682), .Z(n37783) );
  XNOR U39926 ( .A(\modmult_1/zin[0][467] ), .B(n37786), .Z(n31682) );
  IV U39927 ( .A(n37784), .Z(n37786) );
  XOR U39928 ( .A(n37784), .B(n31683), .Z(n37785) );
  XNOR U39929 ( .A(n37787), .B(n37788), .Z(n31683) );
  ANDN U39930 ( .B(\modmult_1/xin[1023] ), .A(n37789), .Z(n37787) );
  IV U39931 ( .A(n37788), .Z(n37789) );
  XNOR U39932 ( .A(m[468]), .B(n37790), .Z(n37788) );
  NAND U39933 ( .A(n37791), .B(mul_pow), .Z(n37790) );
  XOR U39934 ( .A(m[468]), .B(c[468]), .Z(n37791) );
  XOR U39935 ( .A(n37792), .B(n37793), .Z(n37784) );
  ANDN U39936 ( .B(n37794), .A(n31680), .Z(n37792) );
  XNOR U39937 ( .A(\modmult_1/zin[0][466] ), .B(n37795), .Z(n31680) );
  IV U39938 ( .A(n37793), .Z(n37795) );
  XOR U39939 ( .A(n37793), .B(n31681), .Z(n37794) );
  XNOR U39940 ( .A(n37796), .B(n37797), .Z(n31681) );
  ANDN U39941 ( .B(\modmult_1/xin[1023] ), .A(n37798), .Z(n37796) );
  IV U39942 ( .A(n37797), .Z(n37798) );
  XNOR U39943 ( .A(m[467]), .B(n37799), .Z(n37797) );
  NAND U39944 ( .A(n37800), .B(mul_pow), .Z(n37799) );
  XOR U39945 ( .A(m[467]), .B(c[467]), .Z(n37800) );
  XOR U39946 ( .A(n37801), .B(n37802), .Z(n37793) );
  ANDN U39947 ( .B(n37803), .A(n31678), .Z(n37801) );
  XNOR U39948 ( .A(\modmult_1/zin[0][465] ), .B(n37804), .Z(n31678) );
  IV U39949 ( .A(n37802), .Z(n37804) );
  XOR U39950 ( .A(n37802), .B(n31679), .Z(n37803) );
  XNOR U39951 ( .A(n37805), .B(n37806), .Z(n31679) );
  ANDN U39952 ( .B(\modmult_1/xin[1023] ), .A(n37807), .Z(n37805) );
  IV U39953 ( .A(n37806), .Z(n37807) );
  XNOR U39954 ( .A(m[466]), .B(n37808), .Z(n37806) );
  NAND U39955 ( .A(n37809), .B(mul_pow), .Z(n37808) );
  XOR U39956 ( .A(m[466]), .B(c[466]), .Z(n37809) );
  XOR U39957 ( .A(n37810), .B(n37811), .Z(n37802) );
  ANDN U39958 ( .B(n37812), .A(n31676), .Z(n37810) );
  XNOR U39959 ( .A(\modmult_1/zin[0][464] ), .B(n37813), .Z(n31676) );
  IV U39960 ( .A(n37811), .Z(n37813) );
  XOR U39961 ( .A(n37811), .B(n31677), .Z(n37812) );
  XNOR U39962 ( .A(n37814), .B(n37815), .Z(n31677) );
  ANDN U39963 ( .B(\modmult_1/xin[1023] ), .A(n37816), .Z(n37814) );
  IV U39964 ( .A(n37815), .Z(n37816) );
  XNOR U39965 ( .A(m[465]), .B(n37817), .Z(n37815) );
  NAND U39966 ( .A(n37818), .B(mul_pow), .Z(n37817) );
  XOR U39967 ( .A(m[465]), .B(c[465]), .Z(n37818) );
  XOR U39968 ( .A(n37819), .B(n37820), .Z(n37811) );
  ANDN U39969 ( .B(n37821), .A(n31674), .Z(n37819) );
  XNOR U39970 ( .A(\modmult_1/zin[0][463] ), .B(n37822), .Z(n31674) );
  IV U39971 ( .A(n37820), .Z(n37822) );
  XOR U39972 ( .A(n37820), .B(n31675), .Z(n37821) );
  XNOR U39973 ( .A(n37823), .B(n37824), .Z(n31675) );
  ANDN U39974 ( .B(\modmult_1/xin[1023] ), .A(n37825), .Z(n37823) );
  IV U39975 ( .A(n37824), .Z(n37825) );
  XNOR U39976 ( .A(m[464]), .B(n37826), .Z(n37824) );
  NAND U39977 ( .A(n37827), .B(mul_pow), .Z(n37826) );
  XOR U39978 ( .A(m[464]), .B(c[464]), .Z(n37827) );
  XOR U39979 ( .A(n37828), .B(n37829), .Z(n37820) );
  ANDN U39980 ( .B(n37830), .A(n31672), .Z(n37828) );
  XNOR U39981 ( .A(\modmult_1/zin[0][462] ), .B(n37831), .Z(n31672) );
  IV U39982 ( .A(n37829), .Z(n37831) );
  XOR U39983 ( .A(n37829), .B(n31673), .Z(n37830) );
  XNOR U39984 ( .A(n37832), .B(n37833), .Z(n31673) );
  ANDN U39985 ( .B(\modmult_1/xin[1023] ), .A(n37834), .Z(n37832) );
  IV U39986 ( .A(n37833), .Z(n37834) );
  XNOR U39987 ( .A(m[463]), .B(n37835), .Z(n37833) );
  NAND U39988 ( .A(n37836), .B(mul_pow), .Z(n37835) );
  XOR U39989 ( .A(m[463]), .B(c[463]), .Z(n37836) );
  XOR U39990 ( .A(n37837), .B(n37838), .Z(n37829) );
  ANDN U39991 ( .B(n37839), .A(n31670), .Z(n37837) );
  XNOR U39992 ( .A(\modmult_1/zin[0][461] ), .B(n37840), .Z(n31670) );
  IV U39993 ( .A(n37838), .Z(n37840) );
  XOR U39994 ( .A(n37838), .B(n31671), .Z(n37839) );
  XNOR U39995 ( .A(n37841), .B(n37842), .Z(n31671) );
  ANDN U39996 ( .B(\modmult_1/xin[1023] ), .A(n37843), .Z(n37841) );
  IV U39997 ( .A(n37842), .Z(n37843) );
  XNOR U39998 ( .A(m[462]), .B(n37844), .Z(n37842) );
  NAND U39999 ( .A(n37845), .B(mul_pow), .Z(n37844) );
  XOR U40000 ( .A(m[462]), .B(c[462]), .Z(n37845) );
  XOR U40001 ( .A(n37846), .B(n37847), .Z(n37838) );
  ANDN U40002 ( .B(n37848), .A(n31668), .Z(n37846) );
  XNOR U40003 ( .A(\modmult_1/zin[0][460] ), .B(n37849), .Z(n31668) );
  IV U40004 ( .A(n37847), .Z(n37849) );
  XOR U40005 ( .A(n37847), .B(n31669), .Z(n37848) );
  XNOR U40006 ( .A(n37850), .B(n37851), .Z(n31669) );
  ANDN U40007 ( .B(\modmult_1/xin[1023] ), .A(n37852), .Z(n37850) );
  IV U40008 ( .A(n37851), .Z(n37852) );
  XNOR U40009 ( .A(m[461]), .B(n37853), .Z(n37851) );
  NAND U40010 ( .A(n37854), .B(mul_pow), .Z(n37853) );
  XOR U40011 ( .A(m[461]), .B(c[461]), .Z(n37854) );
  XOR U40012 ( .A(n37855), .B(n37856), .Z(n37847) );
  ANDN U40013 ( .B(n37857), .A(n31666), .Z(n37855) );
  XNOR U40014 ( .A(\modmult_1/zin[0][459] ), .B(n37858), .Z(n31666) );
  IV U40015 ( .A(n37856), .Z(n37858) );
  XOR U40016 ( .A(n37856), .B(n31667), .Z(n37857) );
  XNOR U40017 ( .A(n37859), .B(n37860), .Z(n31667) );
  ANDN U40018 ( .B(\modmult_1/xin[1023] ), .A(n37861), .Z(n37859) );
  IV U40019 ( .A(n37860), .Z(n37861) );
  XNOR U40020 ( .A(m[460]), .B(n37862), .Z(n37860) );
  NAND U40021 ( .A(n37863), .B(mul_pow), .Z(n37862) );
  XOR U40022 ( .A(m[460]), .B(c[460]), .Z(n37863) );
  XOR U40023 ( .A(n37864), .B(n37865), .Z(n37856) );
  ANDN U40024 ( .B(n37866), .A(n31664), .Z(n37864) );
  XNOR U40025 ( .A(\modmult_1/zin[0][458] ), .B(n37867), .Z(n31664) );
  IV U40026 ( .A(n37865), .Z(n37867) );
  XOR U40027 ( .A(n37865), .B(n31665), .Z(n37866) );
  XNOR U40028 ( .A(n37868), .B(n37869), .Z(n31665) );
  ANDN U40029 ( .B(\modmult_1/xin[1023] ), .A(n37870), .Z(n37868) );
  IV U40030 ( .A(n37869), .Z(n37870) );
  XNOR U40031 ( .A(m[459]), .B(n37871), .Z(n37869) );
  NAND U40032 ( .A(n37872), .B(mul_pow), .Z(n37871) );
  XOR U40033 ( .A(m[459]), .B(c[459]), .Z(n37872) );
  XOR U40034 ( .A(n37873), .B(n37874), .Z(n37865) );
  ANDN U40035 ( .B(n37875), .A(n31662), .Z(n37873) );
  XNOR U40036 ( .A(\modmult_1/zin[0][457] ), .B(n37876), .Z(n31662) );
  IV U40037 ( .A(n37874), .Z(n37876) );
  XOR U40038 ( .A(n37874), .B(n31663), .Z(n37875) );
  XNOR U40039 ( .A(n37877), .B(n37878), .Z(n31663) );
  ANDN U40040 ( .B(\modmult_1/xin[1023] ), .A(n37879), .Z(n37877) );
  IV U40041 ( .A(n37878), .Z(n37879) );
  XNOR U40042 ( .A(m[458]), .B(n37880), .Z(n37878) );
  NAND U40043 ( .A(n37881), .B(mul_pow), .Z(n37880) );
  XOR U40044 ( .A(m[458]), .B(c[458]), .Z(n37881) );
  XOR U40045 ( .A(n37882), .B(n37883), .Z(n37874) );
  ANDN U40046 ( .B(n37884), .A(n31660), .Z(n37882) );
  XNOR U40047 ( .A(\modmult_1/zin[0][456] ), .B(n37885), .Z(n31660) );
  IV U40048 ( .A(n37883), .Z(n37885) );
  XOR U40049 ( .A(n37883), .B(n31661), .Z(n37884) );
  XNOR U40050 ( .A(n37886), .B(n37887), .Z(n31661) );
  ANDN U40051 ( .B(\modmult_1/xin[1023] ), .A(n37888), .Z(n37886) );
  IV U40052 ( .A(n37887), .Z(n37888) );
  XNOR U40053 ( .A(m[457]), .B(n37889), .Z(n37887) );
  NAND U40054 ( .A(n37890), .B(mul_pow), .Z(n37889) );
  XOR U40055 ( .A(m[457]), .B(c[457]), .Z(n37890) );
  XOR U40056 ( .A(n37891), .B(n37892), .Z(n37883) );
  ANDN U40057 ( .B(n37893), .A(n31658), .Z(n37891) );
  XNOR U40058 ( .A(\modmult_1/zin[0][455] ), .B(n37894), .Z(n31658) );
  IV U40059 ( .A(n37892), .Z(n37894) );
  XOR U40060 ( .A(n37892), .B(n31659), .Z(n37893) );
  XNOR U40061 ( .A(n37895), .B(n37896), .Z(n31659) );
  ANDN U40062 ( .B(\modmult_1/xin[1023] ), .A(n37897), .Z(n37895) );
  IV U40063 ( .A(n37896), .Z(n37897) );
  XNOR U40064 ( .A(m[456]), .B(n37898), .Z(n37896) );
  NAND U40065 ( .A(n37899), .B(mul_pow), .Z(n37898) );
  XOR U40066 ( .A(m[456]), .B(c[456]), .Z(n37899) );
  XOR U40067 ( .A(n37900), .B(n37901), .Z(n37892) );
  ANDN U40068 ( .B(n37902), .A(n31656), .Z(n37900) );
  XNOR U40069 ( .A(\modmult_1/zin[0][454] ), .B(n37903), .Z(n31656) );
  IV U40070 ( .A(n37901), .Z(n37903) );
  XOR U40071 ( .A(n37901), .B(n31657), .Z(n37902) );
  XNOR U40072 ( .A(n37904), .B(n37905), .Z(n31657) );
  ANDN U40073 ( .B(\modmult_1/xin[1023] ), .A(n37906), .Z(n37904) );
  IV U40074 ( .A(n37905), .Z(n37906) );
  XNOR U40075 ( .A(m[455]), .B(n37907), .Z(n37905) );
  NAND U40076 ( .A(n37908), .B(mul_pow), .Z(n37907) );
  XOR U40077 ( .A(m[455]), .B(c[455]), .Z(n37908) );
  XOR U40078 ( .A(n37909), .B(n37910), .Z(n37901) );
  ANDN U40079 ( .B(n37911), .A(n31654), .Z(n37909) );
  XNOR U40080 ( .A(\modmult_1/zin[0][453] ), .B(n37912), .Z(n31654) );
  IV U40081 ( .A(n37910), .Z(n37912) );
  XOR U40082 ( .A(n37910), .B(n31655), .Z(n37911) );
  XNOR U40083 ( .A(n37913), .B(n37914), .Z(n31655) );
  ANDN U40084 ( .B(\modmult_1/xin[1023] ), .A(n37915), .Z(n37913) );
  IV U40085 ( .A(n37914), .Z(n37915) );
  XNOR U40086 ( .A(m[454]), .B(n37916), .Z(n37914) );
  NAND U40087 ( .A(n37917), .B(mul_pow), .Z(n37916) );
  XOR U40088 ( .A(m[454]), .B(c[454]), .Z(n37917) );
  XOR U40089 ( .A(n37918), .B(n37919), .Z(n37910) );
  ANDN U40090 ( .B(n37920), .A(n31652), .Z(n37918) );
  XNOR U40091 ( .A(\modmult_1/zin[0][452] ), .B(n37921), .Z(n31652) );
  IV U40092 ( .A(n37919), .Z(n37921) );
  XOR U40093 ( .A(n37919), .B(n31653), .Z(n37920) );
  XNOR U40094 ( .A(n37922), .B(n37923), .Z(n31653) );
  ANDN U40095 ( .B(\modmult_1/xin[1023] ), .A(n37924), .Z(n37922) );
  IV U40096 ( .A(n37923), .Z(n37924) );
  XNOR U40097 ( .A(m[453]), .B(n37925), .Z(n37923) );
  NAND U40098 ( .A(n37926), .B(mul_pow), .Z(n37925) );
  XOR U40099 ( .A(m[453]), .B(c[453]), .Z(n37926) );
  XOR U40100 ( .A(n37927), .B(n37928), .Z(n37919) );
  ANDN U40101 ( .B(n37929), .A(n31650), .Z(n37927) );
  XNOR U40102 ( .A(\modmult_1/zin[0][451] ), .B(n37930), .Z(n31650) );
  IV U40103 ( .A(n37928), .Z(n37930) );
  XOR U40104 ( .A(n37928), .B(n31651), .Z(n37929) );
  XNOR U40105 ( .A(n37931), .B(n37932), .Z(n31651) );
  ANDN U40106 ( .B(\modmult_1/xin[1023] ), .A(n37933), .Z(n37931) );
  IV U40107 ( .A(n37932), .Z(n37933) );
  XNOR U40108 ( .A(m[452]), .B(n37934), .Z(n37932) );
  NAND U40109 ( .A(n37935), .B(mul_pow), .Z(n37934) );
  XOR U40110 ( .A(m[452]), .B(c[452]), .Z(n37935) );
  XOR U40111 ( .A(n37936), .B(n37937), .Z(n37928) );
  ANDN U40112 ( .B(n37938), .A(n31648), .Z(n37936) );
  XNOR U40113 ( .A(\modmult_1/zin[0][450] ), .B(n37939), .Z(n31648) );
  IV U40114 ( .A(n37937), .Z(n37939) );
  XOR U40115 ( .A(n37937), .B(n31649), .Z(n37938) );
  XNOR U40116 ( .A(n37940), .B(n37941), .Z(n31649) );
  ANDN U40117 ( .B(\modmult_1/xin[1023] ), .A(n37942), .Z(n37940) );
  IV U40118 ( .A(n37941), .Z(n37942) );
  XNOR U40119 ( .A(m[451]), .B(n37943), .Z(n37941) );
  NAND U40120 ( .A(n37944), .B(mul_pow), .Z(n37943) );
  XOR U40121 ( .A(m[451]), .B(c[451]), .Z(n37944) );
  XOR U40122 ( .A(n37945), .B(n37946), .Z(n37937) );
  ANDN U40123 ( .B(n37947), .A(n31646), .Z(n37945) );
  XNOR U40124 ( .A(\modmult_1/zin[0][449] ), .B(n37948), .Z(n31646) );
  IV U40125 ( .A(n37946), .Z(n37948) );
  XOR U40126 ( .A(n37946), .B(n31647), .Z(n37947) );
  XNOR U40127 ( .A(n37949), .B(n37950), .Z(n31647) );
  ANDN U40128 ( .B(\modmult_1/xin[1023] ), .A(n37951), .Z(n37949) );
  IV U40129 ( .A(n37950), .Z(n37951) );
  XNOR U40130 ( .A(m[450]), .B(n37952), .Z(n37950) );
  NAND U40131 ( .A(n37953), .B(mul_pow), .Z(n37952) );
  XOR U40132 ( .A(m[450]), .B(c[450]), .Z(n37953) );
  XOR U40133 ( .A(n37954), .B(n37955), .Z(n37946) );
  ANDN U40134 ( .B(n37956), .A(n31644), .Z(n37954) );
  XNOR U40135 ( .A(\modmult_1/zin[0][448] ), .B(n37957), .Z(n31644) );
  IV U40136 ( .A(n37955), .Z(n37957) );
  XOR U40137 ( .A(n37955), .B(n31645), .Z(n37956) );
  XNOR U40138 ( .A(n37958), .B(n37959), .Z(n31645) );
  ANDN U40139 ( .B(\modmult_1/xin[1023] ), .A(n37960), .Z(n37958) );
  IV U40140 ( .A(n37959), .Z(n37960) );
  XNOR U40141 ( .A(m[449]), .B(n37961), .Z(n37959) );
  NAND U40142 ( .A(n37962), .B(mul_pow), .Z(n37961) );
  XOR U40143 ( .A(m[449]), .B(c[449]), .Z(n37962) );
  XOR U40144 ( .A(n37963), .B(n37964), .Z(n37955) );
  ANDN U40145 ( .B(n37965), .A(n31642), .Z(n37963) );
  XNOR U40146 ( .A(\modmult_1/zin[0][447] ), .B(n37966), .Z(n31642) );
  IV U40147 ( .A(n37964), .Z(n37966) );
  XOR U40148 ( .A(n37964), .B(n31643), .Z(n37965) );
  XNOR U40149 ( .A(n37967), .B(n37968), .Z(n31643) );
  ANDN U40150 ( .B(\modmult_1/xin[1023] ), .A(n37969), .Z(n37967) );
  IV U40151 ( .A(n37968), .Z(n37969) );
  XNOR U40152 ( .A(m[448]), .B(n37970), .Z(n37968) );
  NAND U40153 ( .A(n37971), .B(mul_pow), .Z(n37970) );
  XOR U40154 ( .A(m[448]), .B(c[448]), .Z(n37971) );
  XOR U40155 ( .A(n37972), .B(n37973), .Z(n37964) );
  ANDN U40156 ( .B(n37974), .A(n31640), .Z(n37972) );
  XNOR U40157 ( .A(\modmult_1/zin[0][446] ), .B(n37975), .Z(n31640) );
  IV U40158 ( .A(n37973), .Z(n37975) );
  XOR U40159 ( .A(n37973), .B(n31641), .Z(n37974) );
  XNOR U40160 ( .A(n37976), .B(n37977), .Z(n31641) );
  ANDN U40161 ( .B(\modmult_1/xin[1023] ), .A(n37978), .Z(n37976) );
  IV U40162 ( .A(n37977), .Z(n37978) );
  XNOR U40163 ( .A(m[447]), .B(n37979), .Z(n37977) );
  NAND U40164 ( .A(n37980), .B(mul_pow), .Z(n37979) );
  XOR U40165 ( .A(m[447]), .B(c[447]), .Z(n37980) );
  XOR U40166 ( .A(n37981), .B(n37982), .Z(n37973) );
  ANDN U40167 ( .B(n37983), .A(n31638), .Z(n37981) );
  XNOR U40168 ( .A(\modmult_1/zin[0][445] ), .B(n37984), .Z(n31638) );
  IV U40169 ( .A(n37982), .Z(n37984) );
  XOR U40170 ( .A(n37982), .B(n31639), .Z(n37983) );
  XNOR U40171 ( .A(n37985), .B(n37986), .Z(n31639) );
  ANDN U40172 ( .B(\modmult_1/xin[1023] ), .A(n37987), .Z(n37985) );
  IV U40173 ( .A(n37986), .Z(n37987) );
  XNOR U40174 ( .A(m[446]), .B(n37988), .Z(n37986) );
  NAND U40175 ( .A(n37989), .B(mul_pow), .Z(n37988) );
  XOR U40176 ( .A(m[446]), .B(c[446]), .Z(n37989) );
  XOR U40177 ( .A(n37990), .B(n37991), .Z(n37982) );
  ANDN U40178 ( .B(n37992), .A(n31636), .Z(n37990) );
  XNOR U40179 ( .A(\modmult_1/zin[0][444] ), .B(n37993), .Z(n31636) );
  IV U40180 ( .A(n37991), .Z(n37993) );
  XOR U40181 ( .A(n37991), .B(n31637), .Z(n37992) );
  XNOR U40182 ( .A(n37994), .B(n37995), .Z(n31637) );
  ANDN U40183 ( .B(\modmult_1/xin[1023] ), .A(n37996), .Z(n37994) );
  IV U40184 ( .A(n37995), .Z(n37996) );
  XNOR U40185 ( .A(m[445]), .B(n37997), .Z(n37995) );
  NAND U40186 ( .A(n37998), .B(mul_pow), .Z(n37997) );
  XOR U40187 ( .A(m[445]), .B(c[445]), .Z(n37998) );
  XOR U40188 ( .A(n37999), .B(n38000), .Z(n37991) );
  ANDN U40189 ( .B(n38001), .A(n31634), .Z(n37999) );
  XNOR U40190 ( .A(\modmult_1/zin[0][443] ), .B(n38002), .Z(n31634) );
  IV U40191 ( .A(n38000), .Z(n38002) );
  XOR U40192 ( .A(n38000), .B(n31635), .Z(n38001) );
  XNOR U40193 ( .A(n38003), .B(n38004), .Z(n31635) );
  ANDN U40194 ( .B(\modmult_1/xin[1023] ), .A(n38005), .Z(n38003) );
  IV U40195 ( .A(n38004), .Z(n38005) );
  XNOR U40196 ( .A(m[444]), .B(n38006), .Z(n38004) );
  NAND U40197 ( .A(n38007), .B(mul_pow), .Z(n38006) );
  XOR U40198 ( .A(m[444]), .B(c[444]), .Z(n38007) );
  XOR U40199 ( .A(n38008), .B(n38009), .Z(n38000) );
  ANDN U40200 ( .B(n38010), .A(n31632), .Z(n38008) );
  XNOR U40201 ( .A(\modmult_1/zin[0][442] ), .B(n38011), .Z(n31632) );
  IV U40202 ( .A(n38009), .Z(n38011) );
  XOR U40203 ( .A(n38009), .B(n31633), .Z(n38010) );
  XNOR U40204 ( .A(n38012), .B(n38013), .Z(n31633) );
  ANDN U40205 ( .B(\modmult_1/xin[1023] ), .A(n38014), .Z(n38012) );
  IV U40206 ( .A(n38013), .Z(n38014) );
  XNOR U40207 ( .A(m[443]), .B(n38015), .Z(n38013) );
  NAND U40208 ( .A(n38016), .B(mul_pow), .Z(n38015) );
  XOR U40209 ( .A(m[443]), .B(c[443]), .Z(n38016) );
  XOR U40210 ( .A(n38017), .B(n38018), .Z(n38009) );
  ANDN U40211 ( .B(n38019), .A(n31630), .Z(n38017) );
  XNOR U40212 ( .A(\modmult_1/zin[0][441] ), .B(n38020), .Z(n31630) );
  IV U40213 ( .A(n38018), .Z(n38020) );
  XOR U40214 ( .A(n38018), .B(n31631), .Z(n38019) );
  XNOR U40215 ( .A(n38021), .B(n38022), .Z(n31631) );
  ANDN U40216 ( .B(\modmult_1/xin[1023] ), .A(n38023), .Z(n38021) );
  IV U40217 ( .A(n38022), .Z(n38023) );
  XNOR U40218 ( .A(m[442]), .B(n38024), .Z(n38022) );
  NAND U40219 ( .A(n38025), .B(mul_pow), .Z(n38024) );
  XOR U40220 ( .A(m[442]), .B(c[442]), .Z(n38025) );
  XOR U40221 ( .A(n38026), .B(n38027), .Z(n38018) );
  ANDN U40222 ( .B(n38028), .A(n31628), .Z(n38026) );
  XNOR U40223 ( .A(\modmult_1/zin[0][440] ), .B(n38029), .Z(n31628) );
  IV U40224 ( .A(n38027), .Z(n38029) );
  XOR U40225 ( .A(n38027), .B(n31629), .Z(n38028) );
  XNOR U40226 ( .A(n38030), .B(n38031), .Z(n31629) );
  ANDN U40227 ( .B(\modmult_1/xin[1023] ), .A(n38032), .Z(n38030) );
  IV U40228 ( .A(n38031), .Z(n38032) );
  XNOR U40229 ( .A(m[441]), .B(n38033), .Z(n38031) );
  NAND U40230 ( .A(n38034), .B(mul_pow), .Z(n38033) );
  XOR U40231 ( .A(m[441]), .B(c[441]), .Z(n38034) );
  XOR U40232 ( .A(n38035), .B(n38036), .Z(n38027) );
  ANDN U40233 ( .B(n38037), .A(n31626), .Z(n38035) );
  XNOR U40234 ( .A(\modmult_1/zin[0][439] ), .B(n38038), .Z(n31626) );
  IV U40235 ( .A(n38036), .Z(n38038) );
  XOR U40236 ( .A(n38036), .B(n31627), .Z(n38037) );
  XNOR U40237 ( .A(n38039), .B(n38040), .Z(n31627) );
  ANDN U40238 ( .B(\modmult_1/xin[1023] ), .A(n38041), .Z(n38039) );
  IV U40239 ( .A(n38040), .Z(n38041) );
  XNOR U40240 ( .A(m[440]), .B(n38042), .Z(n38040) );
  NAND U40241 ( .A(n38043), .B(mul_pow), .Z(n38042) );
  XOR U40242 ( .A(m[440]), .B(c[440]), .Z(n38043) );
  XOR U40243 ( .A(n38044), .B(n38045), .Z(n38036) );
  ANDN U40244 ( .B(n38046), .A(n31624), .Z(n38044) );
  XNOR U40245 ( .A(\modmult_1/zin[0][438] ), .B(n38047), .Z(n31624) );
  IV U40246 ( .A(n38045), .Z(n38047) );
  XOR U40247 ( .A(n38045), .B(n31625), .Z(n38046) );
  XNOR U40248 ( .A(n38048), .B(n38049), .Z(n31625) );
  ANDN U40249 ( .B(\modmult_1/xin[1023] ), .A(n38050), .Z(n38048) );
  IV U40250 ( .A(n38049), .Z(n38050) );
  XNOR U40251 ( .A(m[439]), .B(n38051), .Z(n38049) );
  NAND U40252 ( .A(n38052), .B(mul_pow), .Z(n38051) );
  XOR U40253 ( .A(m[439]), .B(c[439]), .Z(n38052) );
  XOR U40254 ( .A(n38053), .B(n38054), .Z(n38045) );
  ANDN U40255 ( .B(n38055), .A(n31622), .Z(n38053) );
  XNOR U40256 ( .A(\modmult_1/zin[0][437] ), .B(n38056), .Z(n31622) );
  IV U40257 ( .A(n38054), .Z(n38056) );
  XOR U40258 ( .A(n38054), .B(n31623), .Z(n38055) );
  XNOR U40259 ( .A(n38057), .B(n38058), .Z(n31623) );
  ANDN U40260 ( .B(\modmult_1/xin[1023] ), .A(n38059), .Z(n38057) );
  IV U40261 ( .A(n38058), .Z(n38059) );
  XNOR U40262 ( .A(m[438]), .B(n38060), .Z(n38058) );
  NAND U40263 ( .A(n38061), .B(mul_pow), .Z(n38060) );
  XOR U40264 ( .A(m[438]), .B(c[438]), .Z(n38061) );
  XOR U40265 ( .A(n38062), .B(n38063), .Z(n38054) );
  ANDN U40266 ( .B(n38064), .A(n31620), .Z(n38062) );
  XNOR U40267 ( .A(\modmult_1/zin[0][436] ), .B(n38065), .Z(n31620) );
  IV U40268 ( .A(n38063), .Z(n38065) );
  XOR U40269 ( .A(n38063), .B(n31621), .Z(n38064) );
  XNOR U40270 ( .A(n38066), .B(n38067), .Z(n31621) );
  ANDN U40271 ( .B(\modmult_1/xin[1023] ), .A(n38068), .Z(n38066) );
  IV U40272 ( .A(n38067), .Z(n38068) );
  XNOR U40273 ( .A(m[437]), .B(n38069), .Z(n38067) );
  NAND U40274 ( .A(n38070), .B(mul_pow), .Z(n38069) );
  XOR U40275 ( .A(m[437]), .B(c[437]), .Z(n38070) );
  XOR U40276 ( .A(n38071), .B(n38072), .Z(n38063) );
  ANDN U40277 ( .B(n38073), .A(n31618), .Z(n38071) );
  XNOR U40278 ( .A(\modmult_1/zin[0][435] ), .B(n38074), .Z(n31618) );
  IV U40279 ( .A(n38072), .Z(n38074) );
  XOR U40280 ( .A(n38072), .B(n31619), .Z(n38073) );
  XNOR U40281 ( .A(n38075), .B(n38076), .Z(n31619) );
  ANDN U40282 ( .B(\modmult_1/xin[1023] ), .A(n38077), .Z(n38075) );
  IV U40283 ( .A(n38076), .Z(n38077) );
  XNOR U40284 ( .A(m[436]), .B(n38078), .Z(n38076) );
  NAND U40285 ( .A(n38079), .B(mul_pow), .Z(n38078) );
  XOR U40286 ( .A(m[436]), .B(c[436]), .Z(n38079) );
  XOR U40287 ( .A(n38080), .B(n38081), .Z(n38072) );
  ANDN U40288 ( .B(n38082), .A(n31616), .Z(n38080) );
  XNOR U40289 ( .A(\modmult_1/zin[0][434] ), .B(n38083), .Z(n31616) );
  IV U40290 ( .A(n38081), .Z(n38083) );
  XOR U40291 ( .A(n38081), .B(n31617), .Z(n38082) );
  XNOR U40292 ( .A(n38084), .B(n38085), .Z(n31617) );
  ANDN U40293 ( .B(\modmult_1/xin[1023] ), .A(n38086), .Z(n38084) );
  IV U40294 ( .A(n38085), .Z(n38086) );
  XNOR U40295 ( .A(m[435]), .B(n38087), .Z(n38085) );
  NAND U40296 ( .A(n38088), .B(mul_pow), .Z(n38087) );
  XOR U40297 ( .A(m[435]), .B(c[435]), .Z(n38088) );
  XOR U40298 ( .A(n38089), .B(n38090), .Z(n38081) );
  ANDN U40299 ( .B(n38091), .A(n31614), .Z(n38089) );
  XNOR U40300 ( .A(\modmult_1/zin[0][433] ), .B(n38092), .Z(n31614) );
  IV U40301 ( .A(n38090), .Z(n38092) );
  XOR U40302 ( .A(n38090), .B(n31615), .Z(n38091) );
  XNOR U40303 ( .A(n38093), .B(n38094), .Z(n31615) );
  ANDN U40304 ( .B(\modmult_1/xin[1023] ), .A(n38095), .Z(n38093) );
  IV U40305 ( .A(n38094), .Z(n38095) );
  XNOR U40306 ( .A(m[434]), .B(n38096), .Z(n38094) );
  NAND U40307 ( .A(n38097), .B(mul_pow), .Z(n38096) );
  XOR U40308 ( .A(m[434]), .B(c[434]), .Z(n38097) );
  XOR U40309 ( .A(n38098), .B(n38099), .Z(n38090) );
  ANDN U40310 ( .B(n38100), .A(n31612), .Z(n38098) );
  XNOR U40311 ( .A(\modmult_1/zin[0][432] ), .B(n38101), .Z(n31612) );
  IV U40312 ( .A(n38099), .Z(n38101) );
  XOR U40313 ( .A(n38099), .B(n31613), .Z(n38100) );
  XNOR U40314 ( .A(n38102), .B(n38103), .Z(n31613) );
  ANDN U40315 ( .B(\modmult_1/xin[1023] ), .A(n38104), .Z(n38102) );
  IV U40316 ( .A(n38103), .Z(n38104) );
  XNOR U40317 ( .A(m[433]), .B(n38105), .Z(n38103) );
  NAND U40318 ( .A(n38106), .B(mul_pow), .Z(n38105) );
  XOR U40319 ( .A(m[433]), .B(c[433]), .Z(n38106) );
  XOR U40320 ( .A(n38107), .B(n38108), .Z(n38099) );
  ANDN U40321 ( .B(n38109), .A(n31610), .Z(n38107) );
  XNOR U40322 ( .A(\modmult_1/zin[0][431] ), .B(n38110), .Z(n31610) );
  IV U40323 ( .A(n38108), .Z(n38110) );
  XOR U40324 ( .A(n38108), .B(n31611), .Z(n38109) );
  XNOR U40325 ( .A(n38111), .B(n38112), .Z(n31611) );
  ANDN U40326 ( .B(\modmult_1/xin[1023] ), .A(n38113), .Z(n38111) );
  IV U40327 ( .A(n38112), .Z(n38113) );
  XNOR U40328 ( .A(m[432]), .B(n38114), .Z(n38112) );
  NAND U40329 ( .A(n38115), .B(mul_pow), .Z(n38114) );
  XOR U40330 ( .A(m[432]), .B(c[432]), .Z(n38115) );
  XOR U40331 ( .A(n38116), .B(n38117), .Z(n38108) );
  ANDN U40332 ( .B(n38118), .A(n31608), .Z(n38116) );
  XNOR U40333 ( .A(\modmult_1/zin[0][430] ), .B(n38119), .Z(n31608) );
  IV U40334 ( .A(n38117), .Z(n38119) );
  XOR U40335 ( .A(n38117), .B(n31609), .Z(n38118) );
  XNOR U40336 ( .A(n38120), .B(n38121), .Z(n31609) );
  ANDN U40337 ( .B(\modmult_1/xin[1023] ), .A(n38122), .Z(n38120) );
  IV U40338 ( .A(n38121), .Z(n38122) );
  XNOR U40339 ( .A(m[431]), .B(n38123), .Z(n38121) );
  NAND U40340 ( .A(n38124), .B(mul_pow), .Z(n38123) );
  XOR U40341 ( .A(m[431]), .B(c[431]), .Z(n38124) );
  XOR U40342 ( .A(n38125), .B(n38126), .Z(n38117) );
  ANDN U40343 ( .B(n38127), .A(n31606), .Z(n38125) );
  XNOR U40344 ( .A(\modmult_1/zin[0][429] ), .B(n38128), .Z(n31606) );
  IV U40345 ( .A(n38126), .Z(n38128) );
  XOR U40346 ( .A(n38126), .B(n31607), .Z(n38127) );
  XNOR U40347 ( .A(n38129), .B(n38130), .Z(n31607) );
  ANDN U40348 ( .B(\modmult_1/xin[1023] ), .A(n38131), .Z(n38129) );
  IV U40349 ( .A(n38130), .Z(n38131) );
  XNOR U40350 ( .A(m[430]), .B(n38132), .Z(n38130) );
  NAND U40351 ( .A(n38133), .B(mul_pow), .Z(n38132) );
  XOR U40352 ( .A(m[430]), .B(c[430]), .Z(n38133) );
  XOR U40353 ( .A(n38134), .B(n38135), .Z(n38126) );
  ANDN U40354 ( .B(n38136), .A(n31604), .Z(n38134) );
  XNOR U40355 ( .A(\modmult_1/zin[0][428] ), .B(n38137), .Z(n31604) );
  IV U40356 ( .A(n38135), .Z(n38137) );
  XOR U40357 ( .A(n38135), .B(n31605), .Z(n38136) );
  XNOR U40358 ( .A(n38138), .B(n38139), .Z(n31605) );
  ANDN U40359 ( .B(\modmult_1/xin[1023] ), .A(n38140), .Z(n38138) );
  IV U40360 ( .A(n38139), .Z(n38140) );
  XNOR U40361 ( .A(m[429]), .B(n38141), .Z(n38139) );
  NAND U40362 ( .A(n38142), .B(mul_pow), .Z(n38141) );
  XOR U40363 ( .A(m[429]), .B(c[429]), .Z(n38142) );
  XOR U40364 ( .A(n38143), .B(n38144), .Z(n38135) );
  ANDN U40365 ( .B(n38145), .A(n31602), .Z(n38143) );
  XNOR U40366 ( .A(\modmult_1/zin[0][427] ), .B(n38146), .Z(n31602) );
  IV U40367 ( .A(n38144), .Z(n38146) );
  XOR U40368 ( .A(n38144), .B(n31603), .Z(n38145) );
  XNOR U40369 ( .A(n38147), .B(n38148), .Z(n31603) );
  ANDN U40370 ( .B(\modmult_1/xin[1023] ), .A(n38149), .Z(n38147) );
  IV U40371 ( .A(n38148), .Z(n38149) );
  XNOR U40372 ( .A(m[428]), .B(n38150), .Z(n38148) );
  NAND U40373 ( .A(n38151), .B(mul_pow), .Z(n38150) );
  XOR U40374 ( .A(m[428]), .B(c[428]), .Z(n38151) );
  XOR U40375 ( .A(n38152), .B(n38153), .Z(n38144) );
  ANDN U40376 ( .B(n38154), .A(n31600), .Z(n38152) );
  XNOR U40377 ( .A(\modmult_1/zin[0][426] ), .B(n38155), .Z(n31600) );
  IV U40378 ( .A(n38153), .Z(n38155) );
  XOR U40379 ( .A(n38153), .B(n31601), .Z(n38154) );
  XNOR U40380 ( .A(n38156), .B(n38157), .Z(n31601) );
  ANDN U40381 ( .B(\modmult_1/xin[1023] ), .A(n38158), .Z(n38156) );
  IV U40382 ( .A(n38157), .Z(n38158) );
  XNOR U40383 ( .A(m[427]), .B(n38159), .Z(n38157) );
  NAND U40384 ( .A(n38160), .B(mul_pow), .Z(n38159) );
  XOR U40385 ( .A(m[427]), .B(c[427]), .Z(n38160) );
  XOR U40386 ( .A(n38161), .B(n38162), .Z(n38153) );
  ANDN U40387 ( .B(n38163), .A(n31598), .Z(n38161) );
  XNOR U40388 ( .A(\modmult_1/zin[0][425] ), .B(n38164), .Z(n31598) );
  IV U40389 ( .A(n38162), .Z(n38164) );
  XOR U40390 ( .A(n38162), .B(n31599), .Z(n38163) );
  XNOR U40391 ( .A(n38165), .B(n38166), .Z(n31599) );
  ANDN U40392 ( .B(\modmult_1/xin[1023] ), .A(n38167), .Z(n38165) );
  IV U40393 ( .A(n38166), .Z(n38167) );
  XNOR U40394 ( .A(m[426]), .B(n38168), .Z(n38166) );
  NAND U40395 ( .A(n38169), .B(mul_pow), .Z(n38168) );
  XOR U40396 ( .A(m[426]), .B(c[426]), .Z(n38169) );
  XOR U40397 ( .A(n38170), .B(n38171), .Z(n38162) );
  ANDN U40398 ( .B(n38172), .A(n31596), .Z(n38170) );
  XNOR U40399 ( .A(\modmult_1/zin[0][424] ), .B(n38173), .Z(n31596) );
  IV U40400 ( .A(n38171), .Z(n38173) );
  XOR U40401 ( .A(n38171), .B(n31597), .Z(n38172) );
  XNOR U40402 ( .A(n38174), .B(n38175), .Z(n31597) );
  ANDN U40403 ( .B(\modmult_1/xin[1023] ), .A(n38176), .Z(n38174) );
  IV U40404 ( .A(n38175), .Z(n38176) );
  XNOR U40405 ( .A(m[425]), .B(n38177), .Z(n38175) );
  NAND U40406 ( .A(n38178), .B(mul_pow), .Z(n38177) );
  XOR U40407 ( .A(m[425]), .B(c[425]), .Z(n38178) );
  XOR U40408 ( .A(n38179), .B(n38180), .Z(n38171) );
  ANDN U40409 ( .B(n38181), .A(n31594), .Z(n38179) );
  XNOR U40410 ( .A(\modmult_1/zin[0][423] ), .B(n38182), .Z(n31594) );
  IV U40411 ( .A(n38180), .Z(n38182) );
  XOR U40412 ( .A(n38180), .B(n31595), .Z(n38181) );
  XNOR U40413 ( .A(n38183), .B(n38184), .Z(n31595) );
  ANDN U40414 ( .B(\modmult_1/xin[1023] ), .A(n38185), .Z(n38183) );
  IV U40415 ( .A(n38184), .Z(n38185) );
  XNOR U40416 ( .A(m[424]), .B(n38186), .Z(n38184) );
  NAND U40417 ( .A(n38187), .B(mul_pow), .Z(n38186) );
  XOR U40418 ( .A(m[424]), .B(c[424]), .Z(n38187) );
  XOR U40419 ( .A(n38188), .B(n38189), .Z(n38180) );
  ANDN U40420 ( .B(n38190), .A(n31592), .Z(n38188) );
  XNOR U40421 ( .A(\modmult_1/zin[0][422] ), .B(n38191), .Z(n31592) );
  IV U40422 ( .A(n38189), .Z(n38191) );
  XOR U40423 ( .A(n38189), .B(n31593), .Z(n38190) );
  XNOR U40424 ( .A(n38192), .B(n38193), .Z(n31593) );
  ANDN U40425 ( .B(\modmult_1/xin[1023] ), .A(n38194), .Z(n38192) );
  IV U40426 ( .A(n38193), .Z(n38194) );
  XNOR U40427 ( .A(m[423]), .B(n38195), .Z(n38193) );
  NAND U40428 ( .A(n38196), .B(mul_pow), .Z(n38195) );
  XOR U40429 ( .A(m[423]), .B(c[423]), .Z(n38196) );
  XOR U40430 ( .A(n38197), .B(n38198), .Z(n38189) );
  ANDN U40431 ( .B(n38199), .A(n31590), .Z(n38197) );
  XNOR U40432 ( .A(\modmult_1/zin[0][421] ), .B(n38200), .Z(n31590) );
  IV U40433 ( .A(n38198), .Z(n38200) );
  XOR U40434 ( .A(n38198), .B(n31591), .Z(n38199) );
  XNOR U40435 ( .A(n38201), .B(n38202), .Z(n31591) );
  ANDN U40436 ( .B(\modmult_1/xin[1023] ), .A(n38203), .Z(n38201) );
  IV U40437 ( .A(n38202), .Z(n38203) );
  XNOR U40438 ( .A(m[422]), .B(n38204), .Z(n38202) );
  NAND U40439 ( .A(n38205), .B(mul_pow), .Z(n38204) );
  XOR U40440 ( .A(m[422]), .B(c[422]), .Z(n38205) );
  XOR U40441 ( .A(n38206), .B(n38207), .Z(n38198) );
  ANDN U40442 ( .B(n38208), .A(n31588), .Z(n38206) );
  XNOR U40443 ( .A(\modmult_1/zin[0][420] ), .B(n38209), .Z(n31588) );
  IV U40444 ( .A(n38207), .Z(n38209) );
  XOR U40445 ( .A(n38207), .B(n31589), .Z(n38208) );
  XNOR U40446 ( .A(n38210), .B(n38211), .Z(n31589) );
  ANDN U40447 ( .B(\modmult_1/xin[1023] ), .A(n38212), .Z(n38210) );
  IV U40448 ( .A(n38211), .Z(n38212) );
  XNOR U40449 ( .A(m[421]), .B(n38213), .Z(n38211) );
  NAND U40450 ( .A(n38214), .B(mul_pow), .Z(n38213) );
  XOR U40451 ( .A(m[421]), .B(c[421]), .Z(n38214) );
  XOR U40452 ( .A(n38215), .B(n38216), .Z(n38207) );
  ANDN U40453 ( .B(n38217), .A(n31586), .Z(n38215) );
  XNOR U40454 ( .A(\modmult_1/zin[0][419] ), .B(n38218), .Z(n31586) );
  IV U40455 ( .A(n38216), .Z(n38218) );
  XOR U40456 ( .A(n38216), .B(n31587), .Z(n38217) );
  XNOR U40457 ( .A(n38219), .B(n38220), .Z(n31587) );
  ANDN U40458 ( .B(\modmult_1/xin[1023] ), .A(n38221), .Z(n38219) );
  IV U40459 ( .A(n38220), .Z(n38221) );
  XNOR U40460 ( .A(m[420]), .B(n38222), .Z(n38220) );
  NAND U40461 ( .A(n38223), .B(mul_pow), .Z(n38222) );
  XOR U40462 ( .A(m[420]), .B(c[420]), .Z(n38223) );
  XOR U40463 ( .A(n38224), .B(n38225), .Z(n38216) );
  ANDN U40464 ( .B(n38226), .A(n31584), .Z(n38224) );
  XNOR U40465 ( .A(\modmult_1/zin[0][418] ), .B(n38227), .Z(n31584) );
  IV U40466 ( .A(n38225), .Z(n38227) );
  XOR U40467 ( .A(n38225), .B(n31585), .Z(n38226) );
  XNOR U40468 ( .A(n38228), .B(n38229), .Z(n31585) );
  ANDN U40469 ( .B(\modmult_1/xin[1023] ), .A(n38230), .Z(n38228) );
  IV U40470 ( .A(n38229), .Z(n38230) );
  XNOR U40471 ( .A(m[419]), .B(n38231), .Z(n38229) );
  NAND U40472 ( .A(n38232), .B(mul_pow), .Z(n38231) );
  XOR U40473 ( .A(m[419]), .B(c[419]), .Z(n38232) );
  XOR U40474 ( .A(n38233), .B(n38234), .Z(n38225) );
  ANDN U40475 ( .B(n38235), .A(n31582), .Z(n38233) );
  XNOR U40476 ( .A(\modmult_1/zin[0][417] ), .B(n38236), .Z(n31582) );
  IV U40477 ( .A(n38234), .Z(n38236) );
  XOR U40478 ( .A(n38234), .B(n31583), .Z(n38235) );
  XNOR U40479 ( .A(n38237), .B(n38238), .Z(n31583) );
  ANDN U40480 ( .B(\modmult_1/xin[1023] ), .A(n38239), .Z(n38237) );
  IV U40481 ( .A(n38238), .Z(n38239) );
  XNOR U40482 ( .A(m[418]), .B(n38240), .Z(n38238) );
  NAND U40483 ( .A(n38241), .B(mul_pow), .Z(n38240) );
  XOR U40484 ( .A(m[418]), .B(c[418]), .Z(n38241) );
  XOR U40485 ( .A(n38242), .B(n38243), .Z(n38234) );
  ANDN U40486 ( .B(n38244), .A(n31580), .Z(n38242) );
  XNOR U40487 ( .A(\modmult_1/zin[0][416] ), .B(n38245), .Z(n31580) );
  IV U40488 ( .A(n38243), .Z(n38245) );
  XOR U40489 ( .A(n38243), .B(n31581), .Z(n38244) );
  XNOR U40490 ( .A(n38246), .B(n38247), .Z(n31581) );
  ANDN U40491 ( .B(\modmult_1/xin[1023] ), .A(n38248), .Z(n38246) );
  IV U40492 ( .A(n38247), .Z(n38248) );
  XNOR U40493 ( .A(m[417]), .B(n38249), .Z(n38247) );
  NAND U40494 ( .A(n38250), .B(mul_pow), .Z(n38249) );
  XOR U40495 ( .A(m[417]), .B(c[417]), .Z(n38250) );
  XOR U40496 ( .A(n38251), .B(n38252), .Z(n38243) );
  ANDN U40497 ( .B(n38253), .A(n31578), .Z(n38251) );
  XNOR U40498 ( .A(\modmult_1/zin[0][415] ), .B(n38254), .Z(n31578) );
  IV U40499 ( .A(n38252), .Z(n38254) );
  XOR U40500 ( .A(n38252), .B(n31579), .Z(n38253) );
  XNOR U40501 ( .A(n38255), .B(n38256), .Z(n31579) );
  ANDN U40502 ( .B(\modmult_1/xin[1023] ), .A(n38257), .Z(n38255) );
  IV U40503 ( .A(n38256), .Z(n38257) );
  XNOR U40504 ( .A(m[416]), .B(n38258), .Z(n38256) );
  NAND U40505 ( .A(n38259), .B(mul_pow), .Z(n38258) );
  XOR U40506 ( .A(m[416]), .B(c[416]), .Z(n38259) );
  XOR U40507 ( .A(n38260), .B(n38261), .Z(n38252) );
  ANDN U40508 ( .B(n38262), .A(n31576), .Z(n38260) );
  XNOR U40509 ( .A(\modmult_1/zin[0][414] ), .B(n38263), .Z(n31576) );
  IV U40510 ( .A(n38261), .Z(n38263) );
  XOR U40511 ( .A(n38261), .B(n31577), .Z(n38262) );
  XNOR U40512 ( .A(n38264), .B(n38265), .Z(n31577) );
  ANDN U40513 ( .B(\modmult_1/xin[1023] ), .A(n38266), .Z(n38264) );
  IV U40514 ( .A(n38265), .Z(n38266) );
  XNOR U40515 ( .A(m[415]), .B(n38267), .Z(n38265) );
  NAND U40516 ( .A(n38268), .B(mul_pow), .Z(n38267) );
  XOR U40517 ( .A(m[415]), .B(c[415]), .Z(n38268) );
  XOR U40518 ( .A(n38269), .B(n38270), .Z(n38261) );
  ANDN U40519 ( .B(n38271), .A(n31574), .Z(n38269) );
  XNOR U40520 ( .A(\modmult_1/zin[0][413] ), .B(n38272), .Z(n31574) );
  IV U40521 ( .A(n38270), .Z(n38272) );
  XOR U40522 ( .A(n38270), .B(n31575), .Z(n38271) );
  XNOR U40523 ( .A(n38273), .B(n38274), .Z(n31575) );
  ANDN U40524 ( .B(\modmult_1/xin[1023] ), .A(n38275), .Z(n38273) );
  IV U40525 ( .A(n38274), .Z(n38275) );
  XNOR U40526 ( .A(m[414]), .B(n38276), .Z(n38274) );
  NAND U40527 ( .A(n38277), .B(mul_pow), .Z(n38276) );
  XOR U40528 ( .A(m[414]), .B(c[414]), .Z(n38277) );
  XOR U40529 ( .A(n38278), .B(n38279), .Z(n38270) );
  ANDN U40530 ( .B(n38280), .A(n31572), .Z(n38278) );
  XNOR U40531 ( .A(\modmult_1/zin[0][412] ), .B(n38281), .Z(n31572) );
  IV U40532 ( .A(n38279), .Z(n38281) );
  XOR U40533 ( .A(n38279), .B(n31573), .Z(n38280) );
  XNOR U40534 ( .A(n38282), .B(n38283), .Z(n31573) );
  ANDN U40535 ( .B(\modmult_1/xin[1023] ), .A(n38284), .Z(n38282) );
  IV U40536 ( .A(n38283), .Z(n38284) );
  XNOR U40537 ( .A(m[413]), .B(n38285), .Z(n38283) );
  NAND U40538 ( .A(n38286), .B(mul_pow), .Z(n38285) );
  XOR U40539 ( .A(m[413]), .B(c[413]), .Z(n38286) );
  XOR U40540 ( .A(n38287), .B(n38288), .Z(n38279) );
  ANDN U40541 ( .B(n38289), .A(n31570), .Z(n38287) );
  XNOR U40542 ( .A(\modmult_1/zin[0][411] ), .B(n38290), .Z(n31570) );
  IV U40543 ( .A(n38288), .Z(n38290) );
  XOR U40544 ( .A(n38288), .B(n31571), .Z(n38289) );
  XNOR U40545 ( .A(n38291), .B(n38292), .Z(n31571) );
  ANDN U40546 ( .B(\modmult_1/xin[1023] ), .A(n38293), .Z(n38291) );
  IV U40547 ( .A(n38292), .Z(n38293) );
  XNOR U40548 ( .A(m[412]), .B(n38294), .Z(n38292) );
  NAND U40549 ( .A(n38295), .B(mul_pow), .Z(n38294) );
  XOR U40550 ( .A(m[412]), .B(c[412]), .Z(n38295) );
  XOR U40551 ( .A(n38296), .B(n38297), .Z(n38288) );
  ANDN U40552 ( .B(n38298), .A(n31568), .Z(n38296) );
  XNOR U40553 ( .A(\modmult_1/zin[0][410] ), .B(n38299), .Z(n31568) );
  IV U40554 ( .A(n38297), .Z(n38299) );
  XOR U40555 ( .A(n38297), .B(n31569), .Z(n38298) );
  XNOR U40556 ( .A(n38300), .B(n38301), .Z(n31569) );
  ANDN U40557 ( .B(\modmult_1/xin[1023] ), .A(n38302), .Z(n38300) );
  IV U40558 ( .A(n38301), .Z(n38302) );
  XNOR U40559 ( .A(m[411]), .B(n38303), .Z(n38301) );
  NAND U40560 ( .A(n38304), .B(mul_pow), .Z(n38303) );
  XOR U40561 ( .A(m[411]), .B(c[411]), .Z(n38304) );
  XOR U40562 ( .A(n38305), .B(n38306), .Z(n38297) );
  ANDN U40563 ( .B(n38307), .A(n31566), .Z(n38305) );
  XNOR U40564 ( .A(\modmult_1/zin[0][409] ), .B(n38308), .Z(n31566) );
  IV U40565 ( .A(n38306), .Z(n38308) );
  XOR U40566 ( .A(n38306), .B(n31567), .Z(n38307) );
  XNOR U40567 ( .A(n38309), .B(n38310), .Z(n31567) );
  ANDN U40568 ( .B(\modmult_1/xin[1023] ), .A(n38311), .Z(n38309) );
  IV U40569 ( .A(n38310), .Z(n38311) );
  XNOR U40570 ( .A(m[410]), .B(n38312), .Z(n38310) );
  NAND U40571 ( .A(n38313), .B(mul_pow), .Z(n38312) );
  XOR U40572 ( .A(m[410]), .B(c[410]), .Z(n38313) );
  XOR U40573 ( .A(n38314), .B(n38315), .Z(n38306) );
  ANDN U40574 ( .B(n38316), .A(n31564), .Z(n38314) );
  XNOR U40575 ( .A(\modmult_1/zin[0][408] ), .B(n38317), .Z(n31564) );
  IV U40576 ( .A(n38315), .Z(n38317) );
  XOR U40577 ( .A(n38315), .B(n31565), .Z(n38316) );
  XNOR U40578 ( .A(n38318), .B(n38319), .Z(n31565) );
  ANDN U40579 ( .B(\modmult_1/xin[1023] ), .A(n38320), .Z(n38318) );
  IV U40580 ( .A(n38319), .Z(n38320) );
  XNOR U40581 ( .A(m[409]), .B(n38321), .Z(n38319) );
  NAND U40582 ( .A(n38322), .B(mul_pow), .Z(n38321) );
  XOR U40583 ( .A(m[409]), .B(c[409]), .Z(n38322) );
  XOR U40584 ( .A(n38323), .B(n38324), .Z(n38315) );
  ANDN U40585 ( .B(n38325), .A(n31562), .Z(n38323) );
  XNOR U40586 ( .A(\modmult_1/zin[0][407] ), .B(n38326), .Z(n31562) );
  IV U40587 ( .A(n38324), .Z(n38326) );
  XOR U40588 ( .A(n38324), .B(n31563), .Z(n38325) );
  XNOR U40589 ( .A(n38327), .B(n38328), .Z(n31563) );
  ANDN U40590 ( .B(\modmult_1/xin[1023] ), .A(n38329), .Z(n38327) );
  IV U40591 ( .A(n38328), .Z(n38329) );
  XNOR U40592 ( .A(m[408]), .B(n38330), .Z(n38328) );
  NAND U40593 ( .A(n38331), .B(mul_pow), .Z(n38330) );
  XOR U40594 ( .A(m[408]), .B(c[408]), .Z(n38331) );
  XOR U40595 ( .A(n38332), .B(n38333), .Z(n38324) );
  ANDN U40596 ( .B(n38334), .A(n31560), .Z(n38332) );
  XNOR U40597 ( .A(\modmult_1/zin[0][406] ), .B(n38335), .Z(n31560) );
  IV U40598 ( .A(n38333), .Z(n38335) );
  XOR U40599 ( .A(n38333), .B(n31561), .Z(n38334) );
  XNOR U40600 ( .A(n38336), .B(n38337), .Z(n31561) );
  ANDN U40601 ( .B(\modmult_1/xin[1023] ), .A(n38338), .Z(n38336) );
  IV U40602 ( .A(n38337), .Z(n38338) );
  XNOR U40603 ( .A(m[407]), .B(n38339), .Z(n38337) );
  NAND U40604 ( .A(n38340), .B(mul_pow), .Z(n38339) );
  XOR U40605 ( .A(m[407]), .B(c[407]), .Z(n38340) );
  XOR U40606 ( .A(n38341), .B(n38342), .Z(n38333) );
  ANDN U40607 ( .B(n38343), .A(n31558), .Z(n38341) );
  XNOR U40608 ( .A(\modmult_1/zin[0][405] ), .B(n38344), .Z(n31558) );
  IV U40609 ( .A(n38342), .Z(n38344) );
  XOR U40610 ( .A(n38342), .B(n31559), .Z(n38343) );
  XNOR U40611 ( .A(n38345), .B(n38346), .Z(n31559) );
  ANDN U40612 ( .B(\modmult_1/xin[1023] ), .A(n38347), .Z(n38345) );
  IV U40613 ( .A(n38346), .Z(n38347) );
  XNOR U40614 ( .A(m[406]), .B(n38348), .Z(n38346) );
  NAND U40615 ( .A(n38349), .B(mul_pow), .Z(n38348) );
  XOR U40616 ( .A(m[406]), .B(c[406]), .Z(n38349) );
  XOR U40617 ( .A(n38350), .B(n38351), .Z(n38342) );
  ANDN U40618 ( .B(n38352), .A(n31556), .Z(n38350) );
  XNOR U40619 ( .A(\modmult_1/zin[0][404] ), .B(n38353), .Z(n31556) );
  IV U40620 ( .A(n38351), .Z(n38353) );
  XOR U40621 ( .A(n38351), .B(n31557), .Z(n38352) );
  XNOR U40622 ( .A(n38354), .B(n38355), .Z(n31557) );
  ANDN U40623 ( .B(\modmult_1/xin[1023] ), .A(n38356), .Z(n38354) );
  IV U40624 ( .A(n38355), .Z(n38356) );
  XNOR U40625 ( .A(m[405]), .B(n38357), .Z(n38355) );
  NAND U40626 ( .A(n38358), .B(mul_pow), .Z(n38357) );
  XOR U40627 ( .A(m[405]), .B(c[405]), .Z(n38358) );
  XOR U40628 ( .A(n38359), .B(n38360), .Z(n38351) );
  ANDN U40629 ( .B(n38361), .A(n31554), .Z(n38359) );
  XNOR U40630 ( .A(\modmult_1/zin[0][403] ), .B(n38362), .Z(n31554) );
  IV U40631 ( .A(n38360), .Z(n38362) );
  XOR U40632 ( .A(n38360), .B(n31555), .Z(n38361) );
  XNOR U40633 ( .A(n38363), .B(n38364), .Z(n31555) );
  ANDN U40634 ( .B(\modmult_1/xin[1023] ), .A(n38365), .Z(n38363) );
  IV U40635 ( .A(n38364), .Z(n38365) );
  XNOR U40636 ( .A(m[404]), .B(n38366), .Z(n38364) );
  NAND U40637 ( .A(n38367), .B(mul_pow), .Z(n38366) );
  XOR U40638 ( .A(m[404]), .B(c[404]), .Z(n38367) );
  XOR U40639 ( .A(n38368), .B(n38369), .Z(n38360) );
  ANDN U40640 ( .B(n38370), .A(n31552), .Z(n38368) );
  XNOR U40641 ( .A(\modmult_1/zin[0][402] ), .B(n38371), .Z(n31552) );
  IV U40642 ( .A(n38369), .Z(n38371) );
  XOR U40643 ( .A(n38369), .B(n31553), .Z(n38370) );
  XNOR U40644 ( .A(n38372), .B(n38373), .Z(n31553) );
  ANDN U40645 ( .B(\modmult_1/xin[1023] ), .A(n38374), .Z(n38372) );
  IV U40646 ( .A(n38373), .Z(n38374) );
  XNOR U40647 ( .A(m[403]), .B(n38375), .Z(n38373) );
  NAND U40648 ( .A(n38376), .B(mul_pow), .Z(n38375) );
  XOR U40649 ( .A(m[403]), .B(c[403]), .Z(n38376) );
  XOR U40650 ( .A(n38377), .B(n38378), .Z(n38369) );
  ANDN U40651 ( .B(n38379), .A(n31550), .Z(n38377) );
  XNOR U40652 ( .A(\modmult_1/zin[0][401] ), .B(n38380), .Z(n31550) );
  IV U40653 ( .A(n38378), .Z(n38380) );
  XOR U40654 ( .A(n38378), .B(n31551), .Z(n38379) );
  XNOR U40655 ( .A(n38381), .B(n38382), .Z(n31551) );
  ANDN U40656 ( .B(\modmult_1/xin[1023] ), .A(n38383), .Z(n38381) );
  IV U40657 ( .A(n38382), .Z(n38383) );
  XNOR U40658 ( .A(m[402]), .B(n38384), .Z(n38382) );
  NAND U40659 ( .A(n38385), .B(mul_pow), .Z(n38384) );
  XOR U40660 ( .A(m[402]), .B(c[402]), .Z(n38385) );
  XOR U40661 ( .A(n38386), .B(n38387), .Z(n38378) );
  ANDN U40662 ( .B(n38388), .A(n31548), .Z(n38386) );
  XNOR U40663 ( .A(\modmult_1/zin[0][400] ), .B(n38389), .Z(n31548) );
  IV U40664 ( .A(n38387), .Z(n38389) );
  XOR U40665 ( .A(n38387), .B(n31549), .Z(n38388) );
  XNOR U40666 ( .A(n38390), .B(n38391), .Z(n31549) );
  ANDN U40667 ( .B(\modmult_1/xin[1023] ), .A(n38392), .Z(n38390) );
  IV U40668 ( .A(n38391), .Z(n38392) );
  XNOR U40669 ( .A(m[401]), .B(n38393), .Z(n38391) );
  NAND U40670 ( .A(n38394), .B(mul_pow), .Z(n38393) );
  XOR U40671 ( .A(m[401]), .B(c[401]), .Z(n38394) );
  XOR U40672 ( .A(n38395), .B(n38396), .Z(n38387) );
  ANDN U40673 ( .B(n38397), .A(n31546), .Z(n38395) );
  XNOR U40674 ( .A(\modmult_1/zin[0][399] ), .B(n38398), .Z(n31546) );
  IV U40675 ( .A(n38396), .Z(n38398) );
  XOR U40676 ( .A(n38396), .B(n31547), .Z(n38397) );
  XNOR U40677 ( .A(n38399), .B(n38400), .Z(n31547) );
  ANDN U40678 ( .B(\modmult_1/xin[1023] ), .A(n38401), .Z(n38399) );
  IV U40679 ( .A(n38400), .Z(n38401) );
  XNOR U40680 ( .A(m[400]), .B(n38402), .Z(n38400) );
  NAND U40681 ( .A(n38403), .B(mul_pow), .Z(n38402) );
  XOR U40682 ( .A(m[400]), .B(c[400]), .Z(n38403) );
  XOR U40683 ( .A(n38404), .B(n38405), .Z(n38396) );
  ANDN U40684 ( .B(n38406), .A(n31544), .Z(n38404) );
  XNOR U40685 ( .A(\modmult_1/zin[0][398] ), .B(n38407), .Z(n31544) );
  IV U40686 ( .A(n38405), .Z(n38407) );
  XOR U40687 ( .A(n38405), .B(n31545), .Z(n38406) );
  XNOR U40688 ( .A(n38408), .B(n38409), .Z(n31545) );
  ANDN U40689 ( .B(\modmult_1/xin[1023] ), .A(n38410), .Z(n38408) );
  IV U40690 ( .A(n38409), .Z(n38410) );
  XNOR U40691 ( .A(m[399]), .B(n38411), .Z(n38409) );
  NAND U40692 ( .A(n38412), .B(mul_pow), .Z(n38411) );
  XOR U40693 ( .A(m[399]), .B(c[399]), .Z(n38412) );
  XOR U40694 ( .A(n38413), .B(n38414), .Z(n38405) );
  ANDN U40695 ( .B(n38415), .A(n31542), .Z(n38413) );
  XNOR U40696 ( .A(\modmult_1/zin[0][397] ), .B(n38416), .Z(n31542) );
  IV U40697 ( .A(n38414), .Z(n38416) );
  XOR U40698 ( .A(n38414), .B(n31543), .Z(n38415) );
  XNOR U40699 ( .A(n38417), .B(n38418), .Z(n31543) );
  ANDN U40700 ( .B(\modmult_1/xin[1023] ), .A(n38419), .Z(n38417) );
  IV U40701 ( .A(n38418), .Z(n38419) );
  XNOR U40702 ( .A(m[398]), .B(n38420), .Z(n38418) );
  NAND U40703 ( .A(n38421), .B(mul_pow), .Z(n38420) );
  XOR U40704 ( .A(m[398]), .B(c[398]), .Z(n38421) );
  XOR U40705 ( .A(n38422), .B(n38423), .Z(n38414) );
  ANDN U40706 ( .B(n38424), .A(n31540), .Z(n38422) );
  XNOR U40707 ( .A(\modmult_1/zin[0][396] ), .B(n38425), .Z(n31540) );
  IV U40708 ( .A(n38423), .Z(n38425) );
  XOR U40709 ( .A(n38423), .B(n31541), .Z(n38424) );
  XNOR U40710 ( .A(n38426), .B(n38427), .Z(n31541) );
  ANDN U40711 ( .B(\modmult_1/xin[1023] ), .A(n38428), .Z(n38426) );
  IV U40712 ( .A(n38427), .Z(n38428) );
  XNOR U40713 ( .A(m[397]), .B(n38429), .Z(n38427) );
  NAND U40714 ( .A(n38430), .B(mul_pow), .Z(n38429) );
  XOR U40715 ( .A(m[397]), .B(c[397]), .Z(n38430) );
  XOR U40716 ( .A(n38431), .B(n38432), .Z(n38423) );
  ANDN U40717 ( .B(n38433), .A(n31538), .Z(n38431) );
  XNOR U40718 ( .A(\modmult_1/zin[0][395] ), .B(n38434), .Z(n31538) );
  IV U40719 ( .A(n38432), .Z(n38434) );
  XOR U40720 ( .A(n38432), .B(n31539), .Z(n38433) );
  XNOR U40721 ( .A(n38435), .B(n38436), .Z(n31539) );
  ANDN U40722 ( .B(\modmult_1/xin[1023] ), .A(n38437), .Z(n38435) );
  IV U40723 ( .A(n38436), .Z(n38437) );
  XNOR U40724 ( .A(m[396]), .B(n38438), .Z(n38436) );
  NAND U40725 ( .A(n38439), .B(mul_pow), .Z(n38438) );
  XOR U40726 ( .A(m[396]), .B(c[396]), .Z(n38439) );
  XOR U40727 ( .A(n38440), .B(n38441), .Z(n38432) );
  ANDN U40728 ( .B(n38442), .A(n31536), .Z(n38440) );
  XNOR U40729 ( .A(\modmult_1/zin[0][394] ), .B(n38443), .Z(n31536) );
  IV U40730 ( .A(n38441), .Z(n38443) );
  XOR U40731 ( .A(n38441), .B(n31537), .Z(n38442) );
  XNOR U40732 ( .A(n38444), .B(n38445), .Z(n31537) );
  ANDN U40733 ( .B(\modmult_1/xin[1023] ), .A(n38446), .Z(n38444) );
  IV U40734 ( .A(n38445), .Z(n38446) );
  XNOR U40735 ( .A(m[395]), .B(n38447), .Z(n38445) );
  NAND U40736 ( .A(n38448), .B(mul_pow), .Z(n38447) );
  XOR U40737 ( .A(m[395]), .B(c[395]), .Z(n38448) );
  XOR U40738 ( .A(n38449), .B(n38450), .Z(n38441) );
  ANDN U40739 ( .B(n38451), .A(n31534), .Z(n38449) );
  XNOR U40740 ( .A(\modmult_1/zin[0][393] ), .B(n38452), .Z(n31534) );
  IV U40741 ( .A(n38450), .Z(n38452) );
  XOR U40742 ( .A(n38450), .B(n31535), .Z(n38451) );
  XNOR U40743 ( .A(n38453), .B(n38454), .Z(n31535) );
  ANDN U40744 ( .B(\modmult_1/xin[1023] ), .A(n38455), .Z(n38453) );
  IV U40745 ( .A(n38454), .Z(n38455) );
  XNOR U40746 ( .A(m[394]), .B(n38456), .Z(n38454) );
  NAND U40747 ( .A(n38457), .B(mul_pow), .Z(n38456) );
  XOR U40748 ( .A(m[394]), .B(c[394]), .Z(n38457) );
  XOR U40749 ( .A(n38458), .B(n38459), .Z(n38450) );
  ANDN U40750 ( .B(n38460), .A(n31532), .Z(n38458) );
  XNOR U40751 ( .A(\modmult_1/zin[0][392] ), .B(n38461), .Z(n31532) );
  IV U40752 ( .A(n38459), .Z(n38461) );
  XOR U40753 ( .A(n38459), .B(n31533), .Z(n38460) );
  XNOR U40754 ( .A(n38462), .B(n38463), .Z(n31533) );
  ANDN U40755 ( .B(\modmult_1/xin[1023] ), .A(n38464), .Z(n38462) );
  IV U40756 ( .A(n38463), .Z(n38464) );
  XNOR U40757 ( .A(m[393]), .B(n38465), .Z(n38463) );
  NAND U40758 ( .A(n38466), .B(mul_pow), .Z(n38465) );
  XOR U40759 ( .A(m[393]), .B(c[393]), .Z(n38466) );
  XOR U40760 ( .A(n38467), .B(n38468), .Z(n38459) );
  ANDN U40761 ( .B(n38469), .A(n31530), .Z(n38467) );
  XNOR U40762 ( .A(\modmult_1/zin[0][391] ), .B(n38470), .Z(n31530) );
  IV U40763 ( .A(n38468), .Z(n38470) );
  XOR U40764 ( .A(n38468), .B(n31531), .Z(n38469) );
  XNOR U40765 ( .A(n38471), .B(n38472), .Z(n31531) );
  ANDN U40766 ( .B(\modmult_1/xin[1023] ), .A(n38473), .Z(n38471) );
  IV U40767 ( .A(n38472), .Z(n38473) );
  XNOR U40768 ( .A(m[392]), .B(n38474), .Z(n38472) );
  NAND U40769 ( .A(n38475), .B(mul_pow), .Z(n38474) );
  XOR U40770 ( .A(m[392]), .B(c[392]), .Z(n38475) );
  XOR U40771 ( .A(n38476), .B(n38477), .Z(n38468) );
  ANDN U40772 ( .B(n38478), .A(n31528), .Z(n38476) );
  XNOR U40773 ( .A(\modmult_1/zin[0][390] ), .B(n38479), .Z(n31528) );
  IV U40774 ( .A(n38477), .Z(n38479) );
  XOR U40775 ( .A(n38477), .B(n31529), .Z(n38478) );
  XNOR U40776 ( .A(n38480), .B(n38481), .Z(n31529) );
  ANDN U40777 ( .B(\modmult_1/xin[1023] ), .A(n38482), .Z(n38480) );
  IV U40778 ( .A(n38481), .Z(n38482) );
  XNOR U40779 ( .A(m[391]), .B(n38483), .Z(n38481) );
  NAND U40780 ( .A(n38484), .B(mul_pow), .Z(n38483) );
  XOR U40781 ( .A(m[391]), .B(c[391]), .Z(n38484) );
  XOR U40782 ( .A(n38485), .B(n38486), .Z(n38477) );
  ANDN U40783 ( .B(n38487), .A(n31526), .Z(n38485) );
  XNOR U40784 ( .A(\modmult_1/zin[0][389] ), .B(n38488), .Z(n31526) );
  IV U40785 ( .A(n38486), .Z(n38488) );
  XOR U40786 ( .A(n38486), .B(n31527), .Z(n38487) );
  XNOR U40787 ( .A(n38489), .B(n38490), .Z(n31527) );
  ANDN U40788 ( .B(\modmult_1/xin[1023] ), .A(n38491), .Z(n38489) );
  IV U40789 ( .A(n38490), .Z(n38491) );
  XNOR U40790 ( .A(m[390]), .B(n38492), .Z(n38490) );
  NAND U40791 ( .A(n38493), .B(mul_pow), .Z(n38492) );
  XOR U40792 ( .A(m[390]), .B(c[390]), .Z(n38493) );
  XOR U40793 ( .A(n38494), .B(n38495), .Z(n38486) );
  ANDN U40794 ( .B(n38496), .A(n31524), .Z(n38494) );
  XNOR U40795 ( .A(\modmult_1/zin[0][388] ), .B(n38497), .Z(n31524) );
  IV U40796 ( .A(n38495), .Z(n38497) );
  XOR U40797 ( .A(n38495), .B(n31525), .Z(n38496) );
  XNOR U40798 ( .A(n38498), .B(n38499), .Z(n31525) );
  ANDN U40799 ( .B(\modmult_1/xin[1023] ), .A(n38500), .Z(n38498) );
  IV U40800 ( .A(n38499), .Z(n38500) );
  XNOR U40801 ( .A(m[389]), .B(n38501), .Z(n38499) );
  NAND U40802 ( .A(n38502), .B(mul_pow), .Z(n38501) );
  XOR U40803 ( .A(m[389]), .B(c[389]), .Z(n38502) );
  XOR U40804 ( .A(n38503), .B(n38504), .Z(n38495) );
  ANDN U40805 ( .B(n38505), .A(n31522), .Z(n38503) );
  XNOR U40806 ( .A(\modmult_1/zin[0][387] ), .B(n38506), .Z(n31522) );
  IV U40807 ( .A(n38504), .Z(n38506) );
  XOR U40808 ( .A(n38504), .B(n31523), .Z(n38505) );
  XNOR U40809 ( .A(n38507), .B(n38508), .Z(n31523) );
  ANDN U40810 ( .B(\modmult_1/xin[1023] ), .A(n38509), .Z(n38507) );
  IV U40811 ( .A(n38508), .Z(n38509) );
  XNOR U40812 ( .A(m[388]), .B(n38510), .Z(n38508) );
  NAND U40813 ( .A(n38511), .B(mul_pow), .Z(n38510) );
  XOR U40814 ( .A(m[388]), .B(c[388]), .Z(n38511) );
  XOR U40815 ( .A(n38512), .B(n38513), .Z(n38504) );
  ANDN U40816 ( .B(n38514), .A(n31520), .Z(n38512) );
  XNOR U40817 ( .A(\modmult_1/zin[0][386] ), .B(n38515), .Z(n31520) );
  IV U40818 ( .A(n38513), .Z(n38515) );
  XOR U40819 ( .A(n38513), .B(n31521), .Z(n38514) );
  XNOR U40820 ( .A(n38516), .B(n38517), .Z(n31521) );
  ANDN U40821 ( .B(\modmult_1/xin[1023] ), .A(n38518), .Z(n38516) );
  IV U40822 ( .A(n38517), .Z(n38518) );
  XNOR U40823 ( .A(m[387]), .B(n38519), .Z(n38517) );
  NAND U40824 ( .A(n38520), .B(mul_pow), .Z(n38519) );
  XOR U40825 ( .A(m[387]), .B(c[387]), .Z(n38520) );
  XOR U40826 ( .A(n38521), .B(n38522), .Z(n38513) );
  ANDN U40827 ( .B(n38523), .A(n31518), .Z(n38521) );
  XNOR U40828 ( .A(\modmult_1/zin[0][385] ), .B(n38524), .Z(n31518) );
  IV U40829 ( .A(n38522), .Z(n38524) );
  XOR U40830 ( .A(n38522), .B(n31519), .Z(n38523) );
  XNOR U40831 ( .A(n38525), .B(n38526), .Z(n31519) );
  ANDN U40832 ( .B(\modmult_1/xin[1023] ), .A(n38527), .Z(n38525) );
  IV U40833 ( .A(n38526), .Z(n38527) );
  XNOR U40834 ( .A(m[386]), .B(n38528), .Z(n38526) );
  NAND U40835 ( .A(n38529), .B(mul_pow), .Z(n38528) );
  XOR U40836 ( .A(m[386]), .B(c[386]), .Z(n38529) );
  XOR U40837 ( .A(n38530), .B(n38531), .Z(n38522) );
  ANDN U40838 ( .B(n38532), .A(n31516), .Z(n38530) );
  XNOR U40839 ( .A(\modmult_1/zin[0][384] ), .B(n38533), .Z(n31516) );
  IV U40840 ( .A(n38531), .Z(n38533) );
  XOR U40841 ( .A(n38531), .B(n31517), .Z(n38532) );
  XNOR U40842 ( .A(n38534), .B(n38535), .Z(n31517) );
  ANDN U40843 ( .B(\modmult_1/xin[1023] ), .A(n38536), .Z(n38534) );
  IV U40844 ( .A(n38535), .Z(n38536) );
  XNOR U40845 ( .A(m[385]), .B(n38537), .Z(n38535) );
  NAND U40846 ( .A(n38538), .B(mul_pow), .Z(n38537) );
  XOR U40847 ( .A(m[385]), .B(c[385]), .Z(n38538) );
  XOR U40848 ( .A(n38539), .B(n38540), .Z(n38531) );
  ANDN U40849 ( .B(n38541), .A(n31514), .Z(n38539) );
  XNOR U40850 ( .A(\modmult_1/zin[0][383] ), .B(n38542), .Z(n31514) );
  IV U40851 ( .A(n38540), .Z(n38542) );
  XOR U40852 ( .A(n38540), .B(n31515), .Z(n38541) );
  XNOR U40853 ( .A(n38543), .B(n38544), .Z(n31515) );
  ANDN U40854 ( .B(\modmult_1/xin[1023] ), .A(n38545), .Z(n38543) );
  IV U40855 ( .A(n38544), .Z(n38545) );
  XNOR U40856 ( .A(m[384]), .B(n38546), .Z(n38544) );
  NAND U40857 ( .A(n38547), .B(mul_pow), .Z(n38546) );
  XOR U40858 ( .A(m[384]), .B(c[384]), .Z(n38547) );
  XOR U40859 ( .A(n38548), .B(n38549), .Z(n38540) );
  ANDN U40860 ( .B(n38550), .A(n31512), .Z(n38548) );
  XNOR U40861 ( .A(\modmult_1/zin[0][382] ), .B(n38551), .Z(n31512) );
  IV U40862 ( .A(n38549), .Z(n38551) );
  XOR U40863 ( .A(n38549), .B(n31513), .Z(n38550) );
  XNOR U40864 ( .A(n38552), .B(n38553), .Z(n31513) );
  ANDN U40865 ( .B(\modmult_1/xin[1023] ), .A(n38554), .Z(n38552) );
  IV U40866 ( .A(n38553), .Z(n38554) );
  XNOR U40867 ( .A(m[383]), .B(n38555), .Z(n38553) );
  NAND U40868 ( .A(n38556), .B(mul_pow), .Z(n38555) );
  XOR U40869 ( .A(m[383]), .B(c[383]), .Z(n38556) );
  XOR U40870 ( .A(n38557), .B(n38558), .Z(n38549) );
  ANDN U40871 ( .B(n38559), .A(n31510), .Z(n38557) );
  XNOR U40872 ( .A(\modmult_1/zin[0][381] ), .B(n38560), .Z(n31510) );
  IV U40873 ( .A(n38558), .Z(n38560) );
  XOR U40874 ( .A(n38558), .B(n31511), .Z(n38559) );
  XNOR U40875 ( .A(n38561), .B(n38562), .Z(n31511) );
  ANDN U40876 ( .B(\modmult_1/xin[1023] ), .A(n38563), .Z(n38561) );
  IV U40877 ( .A(n38562), .Z(n38563) );
  XNOR U40878 ( .A(m[382]), .B(n38564), .Z(n38562) );
  NAND U40879 ( .A(n38565), .B(mul_pow), .Z(n38564) );
  XOR U40880 ( .A(m[382]), .B(c[382]), .Z(n38565) );
  XOR U40881 ( .A(n38566), .B(n38567), .Z(n38558) );
  ANDN U40882 ( .B(n38568), .A(n31508), .Z(n38566) );
  XNOR U40883 ( .A(\modmult_1/zin[0][380] ), .B(n38569), .Z(n31508) );
  IV U40884 ( .A(n38567), .Z(n38569) );
  XOR U40885 ( .A(n38567), .B(n31509), .Z(n38568) );
  XNOR U40886 ( .A(n38570), .B(n38571), .Z(n31509) );
  ANDN U40887 ( .B(\modmult_1/xin[1023] ), .A(n38572), .Z(n38570) );
  IV U40888 ( .A(n38571), .Z(n38572) );
  XNOR U40889 ( .A(m[381]), .B(n38573), .Z(n38571) );
  NAND U40890 ( .A(n38574), .B(mul_pow), .Z(n38573) );
  XOR U40891 ( .A(m[381]), .B(c[381]), .Z(n38574) );
  XOR U40892 ( .A(n38575), .B(n38576), .Z(n38567) );
  ANDN U40893 ( .B(n38577), .A(n31506), .Z(n38575) );
  XNOR U40894 ( .A(\modmult_1/zin[0][379] ), .B(n38578), .Z(n31506) );
  IV U40895 ( .A(n38576), .Z(n38578) );
  XOR U40896 ( .A(n38576), .B(n31507), .Z(n38577) );
  XNOR U40897 ( .A(n38579), .B(n38580), .Z(n31507) );
  ANDN U40898 ( .B(\modmult_1/xin[1023] ), .A(n38581), .Z(n38579) );
  IV U40899 ( .A(n38580), .Z(n38581) );
  XNOR U40900 ( .A(m[380]), .B(n38582), .Z(n38580) );
  NAND U40901 ( .A(n38583), .B(mul_pow), .Z(n38582) );
  XOR U40902 ( .A(m[380]), .B(c[380]), .Z(n38583) );
  XOR U40903 ( .A(n38584), .B(n38585), .Z(n38576) );
  ANDN U40904 ( .B(n38586), .A(n31504), .Z(n38584) );
  XNOR U40905 ( .A(\modmult_1/zin[0][378] ), .B(n38587), .Z(n31504) );
  IV U40906 ( .A(n38585), .Z(n38587) );
  XOR U40907 ( .A(n38585), .B(n31505), .Z(n38586) );
  XNOR U40908 ( .A(n38588), .B(n38589), .Z(n31505) );
  ANDN U40909 ( .B(\modmult_1/xin[1023] ), .A(n38590), .Z(n38588) );
  IV U40910 ( .A(n38589), .Z(n38590) );
  XNOR U40911 ( .A(m[379]), .B(n38591), .Z(n38589) );
  NAND U40912 ( .A(n38592), .B(mul_pow), .Z(n38591) );
  XOR U40913 ( .A(m[379]), .B(c[379]), .Z(n38592) );
  XOR U40914 ( .A(n38593), .B(n38594), .Z(n38585) );
  ANDN U40915 ( .B(n38595), .A(n31502), .Z(n38593) );
  XNOR U40916 ( .A(\modmult_1/zin[0][377] ), .B(n38596), .Z(n31502) );
  IV U40917 ( .A(n38594), .Z(n38596) );
  XOR U40918 ( .A(n38594), .B(n31503), .Z(n38595) );
  XNOR U40919 ( .A(n38597), .B(n38598), .Z(n31503) );
  ANDN U40920 ( .B(\modmult_1/xin[1023] ), .A(n38599), .Z(n38597) );
  IV U40921 ( .A(n38598), .Z(n38599) );
  XNOR U40922 ( .A(m[378]), .B(n38600), .Z(n38598) );
  NAND U40923 ( .A(n38601), .B(mul_pow), .Z(n38600) );
  XOR U40924 ( .A(m[378]), .B(c[378]), .Z(n38601) );
  XOR U40925 ( .A(n38602), .B(n38603), .Z(n38594) );
  ANDN U40926 ( .B(n38604), .A(n31500), .Z(n38602) );
  XNOR U40927 ( .A(\modmult_1/zin[0][376] ), .B(n38605), .Z(n31500) );
  IV U40928 ( .A(n38603), .Z(n38605) );
  XOR U40929 ( .A(n38603), .B(n31501), .Z(n38604) );
  XNOR U40930 ( .A(n38606), .B(n38607), .Z(n31501) );
  ANDN U40931 ( .B(\modmult_1/xin[1023] ), .A(n38608), .Z(n38606) );
  IV U40932 ( .A(n38607), .Z(n38608) );
  XNOR U40933 ( .A(m[377]), .B(n38609), .Z(n38607) );
  NAND U40934 ( .A(n38610), .B(mul_pow), .Z(n38609) );
  XOR U40935 ( .A(m[377]), .B(c[377]), .Z(n38610) );
  XOR U40936 ( .A(n38611), .B(n38612), .Z(n38603) );
  ANDN U40937 ( .B(n38613), .A(n31498), .Z(n38611) );
  XNOR U40938 ( .A(\modmult_1/zin[0][375] ), .B(n38614), .Z(n31498) );
  IV U40939 ( .A(n38612), .Z(n38614) );
  XOR U40940 ( .A(n38612), .B(n31499), .Z(n38613) );
  XNOR U40941 ( .A(n38615), .B(n38616), .Z(n31499) );
  ANDN U40942 ( .B(\modmult_1/xin[1023] ), .A(n38617), .Z(n38615) );
  IV U40943 ( .A(n38616), .Z(n38617) );
  XNOR U40944 ( .A(m[376]), .B(n38618), .Z(n38616) );
  NAND U40945 ( .A(n38619), .B(mul_pow), .Z(n38618) );
  XOR U40946 ( .A(m[376]), .B(c[376]), .Z(n38619) );
  XOR U40947 ( .A(n38620), .B(n38621), .Z(n38612) );
  ANDN U40948 ( .B(n38622), .A(n31496), .Z(n38620) );
  XNOR U40949 ( .A(\modmult_1/zin[0][374] ), .B(n38623), .Z(n31496) );
  IV U40950 ( .A(n38621), .Z(n38623) );
  XOR U40951 ( .A(n38621), .B(n31497), .Z(n38622) );
  XNOR U40952 ( .A(n38624), .B(n38625), .Z(n31497) );
  ANDN U40953 ( .B(\modmult_1/xin[1023] ), .A(n38626), .Z(n38624) );
  IV U40954 ( .A(n38625), .Z(n38626) );
  XNOR U40955 ( .A(m[375]), .B(n38627), .Z(n38625) );
  NAND U40956 ( .A(n38628), .B(mul_pow), .Z(n38627) );
  XOR U40957 ( .A(m[375]), .B(c[375]), .Z(n38628) );
  XOR U40958 ( .A(n38629), .B(n38630), .Z(n38621) );
  ANDN U40959 ( .B(n38631), .A(n31494), .Z(n38629) );
  XNOR U40960 ( .A(\modmult_1/zin[0][373] ), .B(n38632), .Z(n31494) );
  IV U40961 ( .A(n38630), .Z(n38632) );
  XOR U40962 ( .A(n38630), .B(n31495), .Z(n38631) );
  XNOR U40963 ( .A(n38633), .B(n38634), .Z(n31495) );
  ANDN U40964 ( .B(\modmult_1/xin[1023] ), .A(n38635), .Z(n38633) );
  IV U40965 ( .A(n38634), .Z(n38635) );
  XNOR U40966 ( .A(m[374]), .B(n38636), .Z(n38634) );
  NAND U40967 ( .A(n38637), .B(mul_pow), .Z(n38636) );
  XOR U40968 ( .A(m[374]), .B(c[374]), .Z(n38637) );
  XOR U40969 ( .A(n38638), .B(n38639), .Z(n38630) );
  ANDN U40970 ( .B(n38640), .A(n31492), .Z(n38638) );
  XNOR U40971 ( .A(\modmult_1/zin[0][372] ), .B(n38641), .Z(n31492) );
  IV U40972 ( .A(n38639), .Z(n38641) );
  XOR U40973 ( .A(n38639), .B(n31493), .Z(n38640) );
  XNOR U40974 ( .A(n38642), .B(n38643), .Z(n31493) );
  ANDN U40975 ( .B(\modmult_1/xin[1023] ), .A(n38644), .Z(n38642) );
  IV U40976 ( .A(n38643), .Z(n38644) );
  XNOR U40977 ( .A(m[373]), .B(n38645), .Z(n38643) );
  NAND U40978 ( .A(n38646), .B(mul_pow), .Z(n38645) );
  XOR U40979 ( .A(m[373]), .B(c[373]), .Z(n38646) );
  XOR U40980 ( .A(n38647), .B(n38648), .Z(n38639) );
  ANDN U40981 ( .B(n38649), .A(n31490), .Z(n38647) );
  XNOR U40982 ( .A(\modmult_1/zin[0][371] ), .B(n38650), .Z(n31490) );
  IV U40983 ( .A(n38648), .Z(n38650) );
  XOR U40984 ( .A(n38648), .B(n31491), .Z(n38649) );
  XNOR U40985 ( .A(n38651), .B(n38652), .Z(n31491) );
  ANDN U40986 ( .B(\modmult_1/xin[1023] ), .A(n38653), .Z(n38651) );
  IV U40987 ( .A(n38652), .Z(n38653) );
  XNOR U40988 ( .A(m[372]), .B(n38654), .Z(n38652) );
  NAND U40989 ( .A(n38655), .B(mul_pow), .Z(n38654) );
  XOR U40990 ( .A(m[372]), .B(c[372]), .Z(n38655) );
  XOR U40991 ( .A(n38656), .B(n38657), .Z(n38648) );
  ANDN U40992 ( .B(n38658), .A(n31488), .Z(n38656) );
  XNOR U40993 ( .A(\modmult_1/zin[0][370] ), .B(n38659), .Z(n31488) );
  IV U40994 ( .A(n38657), .Z(n38659) );
  XOR U40995 ( .A(n38657), .B(n31489), .Z(n38658) );
  XNOR U40996 ( .A(n38660), .B(n38661), .Z(n31489) );
  ANDN U40997 ( .B(\modmult_1/xin[1023] ), .A(n38662), .Z(n38660) );
  IV U40998 ( .A(n38661), .Z(n38662) );
  XNOR U40999 ( .A(m[371]), .B(n38663), .Z(n38661) );
  NAND U41000 ( .A(n38664), .B(mul_pow), .Z(n38663) );
  XOR U41001 ( .A(m[371]), .B(c[371]), .Z(n38664) );
  XOR U41002 ( .A(n38665), .B(n38666), .Z(n38657) );
  ANDN U41003 ( .B(n38667), .A(n31486), .Z(n38665) );
  XNOR U41004 ( .A(\modmult_1/zin[0][369] ), .B(n38668), .Z(n31486) );
  IV U41005 ( .A(n38666), .Z(n38668) );
  XOR U41006 ( .A(n38666), .B(n31487), .Z(n38667) );
  XNOR U41007 ( .A(n38669), .B(n38670), .Z(n31487) );
  ANDN U41008 ( .B(\modmult_1/xin[1023] ), .A(n38671), .Z(n38669) );
  IV U41009 ( .A(n38670), .Z(n38671) );
  XNOR U41010 ( .A(m[370]), .B(n38672), .Z(n38670) );
  NAND U41011 ( .A(n38673), .B(mul_pow), .Z(n38672) );
  XOR U41012 ( .A(m[370]), .B(c[370]), .Z(n38673) );
  XOR U41013 ( .A(n38674), .B(n38675), .Z(n38666) );
  ANDN U41014 ( .B(n38676), .A(n31484), .Z(n38674) );
  XNOR U41015 ( .A(\modmult_1/zin[0][368] ), .B(n38677), .Z(n31484) );
  IV U41016 ( .A(n38675), .Z(n38677) );
  XOR U41017 ( .A(n38675), .B(n31485), .Z(n38676) );
  XNOR U41018 ( .A(n38678), .B(n38679), .Z(n31485) );
  ANDN U41019 ( .B(\modmult_1/xin[1023] ), .A(n38680), .Z(n38678) );
  IV U41020 ( .A(n38679), .Z(n38680) );
  XNOR U41021 ( .A(m[369]), .B(n38681), .Z(n38679) );
  NAND U41022 ( .A(n38682), .B(mul_pow), .Z(n38681) );
  XOR U41023 ( .A(m[369]), .B(c[369]), .Z(n38682) );
  XOR U41024 ( .A(n38683), .B(n38684), .Z(n38675) );
  ANDN U41025 ( .B(n38685), .A(n31482), .Z(n38683) );
  XNOR U41026 ( .A(\modmult_1/zin[0][367] ), .B(n38686), .Z(n31482) );
  IV U41027 ( .A(n38684), .Z(n38686) );
  XOR U41028 ( .A(n38684), .B(n31483), .Z(n38685) );
  XNOR U41029 ( .A(n38687), .B(n38688), .Z(n31483) );
  ANDN U41030 ( .B(\modmult_1/xin[1023] ), .A(n38689), .Z(n38687) );
  IV U41031 ( .A(n38688), .Z(n38689) );
  XNOR U41032 ( .A(m[368]), .B(n38690), .Z(n38688) );
  NAND U41033 ( .A(n38691), .B(mul_pow), .Z(n38690) );
  XOR U41034 ( .A(m[368]), .B(c[368]), .Z(n38691) );
  XOR U41035 ( .A(n38692), .B(n38693), .Z(n38684) );
  ANDN U41036 ( .B(n38694), .A(n31480), .Z(n38692) );
  XNOR U41037 ( .A(\modmult_1/zin[0][366] ), .B(n38695), .Z(n31480) );
  IV U41038 ( .A(n38693), .Z(n38695) );
  XOR U41039 ( .A(n38693), .B(n31481), .Z(n38694) );
  XNOR U41040 ( .A(n38696), .B(n38697), .Z(n31481) );
  ANDN U41041 ( .B(\modmult_1/xin[1023] ), .A(n38698), .Z(n38696) );
  IV U41042 ( .A(n38697), .Z(n38698) );
  XNOR U41043 ( .A(m[367]), .B(n38699), .Z(n38697) );
  NAND U41044 ( .A(n38700), .B(mul_pow), .Z(n38699) );
  XOR U41045 ( .A(m[367]), .B(c[367]), .Z(n38700) );
  XOR U41046 ( .A(n38701), .B(n38702), .Z(n38693) );
  ANDN U41047 ( .B(n38703), .A(n31478), .Z(n38701) );
  XNOR U41048 ( .A(\modmult_1/zin[0][365] ), .B(n38704), .Z(n31478) );
  IV U41049 ( .A(n38702), .Z(n38704) );
  XOR U41050 ( .A(n38702), .B(n31479), .Z(n38703) );
  XNOR U41051 ( .A(n38705), .B(n38706), .Z(n31479) );
  ANDN U41052 ( .B(\modmult_1/xin[1023] ), .A(n38707), .Z(n38705) );
  IV U41053 ( .A(n38706), .Z(n38707) );
  XNOR U41054 ( .A(m[366]), .B(n38708), .Z(n38706) );
  NAND U41055 ( .A(n38709), .B(mul_pow), .Z(n38708) );
  XOR U41056 ( .A(m[366]), .B(c[366]), .Z(n38709) );
  XOR U41057 ( .A(n38710), .B(n38711), .Z(n38702) );
  ANDN U41058 ( .B(n38712), .A(n31476), .Z(n38710) );
  XNOR U41059 ( .A(\modmult_1/zin[0][364] ), .B(n38713), .Z(n31476) );
  IV U41060 ( .A(n38711), .Z(n38713) );
  XOR U41061 ( .A(n38711), .B(n31477), .Z(n38712) );
  XNOR U41062 ( .A(n38714), .B(n38715), .Z(n31477) );
  ANDN U41063 ( .B(\modmult_1/xin[1023] ), .A(n38716), .Z(n38714) );
  IV U41064 ( .A(n38715), .Z(n38716) );
  XNOR U41065 ( .A(m[365]), .B(n38717), .Z(n38715) );
  NAND U41066 ( .A(n38718), .B(mul_pow), .Z(n38717) );
  XOR U41067 ( .A(m[365]), .B(c[365]), .Z(n38718) );
  XOR U41068 ( .A(n38719), .B(n38720), .Z(n38711) );
  ANDN U41069 ( .B(n38721), .A(n31474), .Z(n38719) );
  XNOR U41070 ( .A(\modmult_1/zin[0][363] ), .B(n38722), .Z(n31474) );
  IV U41071 ( .A(n38720), .Z(n38722) );
  XOR U41072 ( .A(n38720), .B(n31475), .Z(n38721) );
  XNOR U41073 ( .A(n38723), .B(n38724), .Z(n31475) );
  ANDN U41074 ( .B(\modmult_1/xin[1023] ), .A(n38725), .Z(n38723) );
  IV U41075 ( .A(n38724), .Z(n38725) );
  XNOR U41076 ( .A(m[364]), .B(n38726), .Z(n38724) );
  NAND U41077 ( .A(n38727), .B(mul_pow), .Z(n38726) );
  XOR U41078 ( .A(m[364]), .B(c[364]), .Z(n38727) );
  XOR U41079 ( .A(n38728), .B(n38729), .Z(n38720) );
  ANDN U41080 ( .B(n38730), .A(n31472), .Z(n38728) );
  XNOR U41081 ( .A(\modmult_1/zin[0][362] ), .B(n38731), .Z(n31472) );
  IV U41082 ( .A(n38729), .Z(n38731) );
  XOR U41083 ( .A(n38729), .B(n31473), .Z(n38730) );
  XNOR U41084 ( .A(n38732), .B(n38733), .Z(n31473) );
  ANDN U41085 ( .B(\modmult_1/xin[1023] ), .A(n38734), .Z(n38732) );
  IV U41086 ( .A(n38733), .Z(n38734) );
  XNOR U41087 ( .A(m[363]), .B(n38735), .Z(n38733) );
  NAND U41088 ( .A(n38736), .B(mul_pow), .Z(n38735) );
  XOR U41089 ( .A(m[363]), .B(c[363]), .Z(n38736) );
  XOR U41090 ( .A(n38737), .B(n38738), .Z(n38729) );
  ANDN U41091 ( .B(n38739), .A(n31470), .Z(n38737) );
  XNOR U41092 ( .A(\modmult_1/zin[0][361] ), .B(n38740), .Z(n31470) );
  IV U41093 ( .A(n38738), .Z(n38740) );
  XOR U41094 ( .A(n38738), .B(n31471), .Z(n38739) );
  XNOR U41095 ( .A(n38741), .B(n38742), .Z(n31471) );
  ANDN U41096 ( .B(\modmult_1/xin[1023] ), .A(n38743), .Z(n38741) );
  IV U41097 ( .A(n38742), .Z(n38743) );
  XNOR U41098 ( .A(m[362]), .B(n38744), .Z(n38742) );
  NAND U41099 ( .A(n38745), .B(mul_pow), .Z(n38744) );
  XOR U41100 ( .A(m[362]), .B(c[362]), .Z(n38745) );
  XOR U41101 ( .A(n38746), .B(n38747), .Z(n38738) );
  ANDN U41102 ( .B(n38748), .A(n31468), .Z(n38746) );
  XNOR U41103 ( .A(\modmult_1/zin[0][360] ), .B(n38749), .Z(n31468) );
  IV U41104 ( .A(n38747), .Z(n38749) );
  XOR U41105 ( .A(n38747), .B(n31469), .Z(n38748) );
  XNOR U41106 ( .A(n38750), .B(n38751), .Z(n31469) );
  ANDN U41107 ( .B(\modmult_1/xin[1023] ), .A(n38752), .Z(n38750) );
  IV U41108 ( .A(n38751), .Z(n38752) );
  XNOR U41109 ( .A(m[361]), .B(n38753), .Z(n38751) );
  NAND U41110 ( .A(n38754), .B(mul_pow), .Z(n38753) );
  XOR U41111 ( .A(m[361]), .B(c[361]), .Z(n38754) );
  XOR U41112 ( .A(n38755), .B(n38756), .Z(n38747) );
  ANDN U41113 ( .B(n38757), .A(n31466), .Z(n38755) );
  XNOR U41114 ( .A(\modmult_1/zin[0][359] ), .B(n38758), .Z(n31466) );
  IV U41115 ( .A(n38756), .Z(n38758) );
  XOR U41116 ( .A(n38756), .B(n31467), .Z(n38757) );
  XNOR U41117 ( .A(n38759), .B(n38760), .Z(n31467) );
  ANDN U41118 ( .B(\modmult_1/xin[1023] ), .A(n38761), .Z(n38759) );
  IV U41119 ( .A(n38760), .Z(n38761) );
  XNOR U41120 ( .A(m[360]), .B(n38762), .Z(n38760) );
  NAND U41121 ( .A(n38763), .B(mul_pow), .Z(n38762) );
  XOR U41122 ( .A(m[360]), .B(c[360]), .Z(n38763) );
  XOR U41123 ( .A(n38764), .B(n38765), .Z(n38756) );
  ANDN U41124 ( .B(n38766), .A(n31464), .Z(n38764) );
  XNOR U41125 ( .A(\modmult_1/zin[0][358] ), .B(n38767), .Z(n31464) );
  IV U41126 ( .A(n38765), .Z(n38767) );
  XOR U41127 ( .A(n38765), .B(n31465), .Z(n38766) );
  XNOR U41128 ( .A(n38768), .B(n38769), .Z(n31465) );
  ANDN U41129 ( .B(\modmult_1/xin[1023] ), .A(n38770), .Z(n38768) );
  IV U41130 ( .A(n38769), .Z(n38770) );
  XNOR U41131 ( .A(m[359]), .B(n38771), .Z(n38769) );
  NAND U41132 ( .A(n38772), .B(mul_pow), .Z(n38771) );
  XOR U41133 ( .A(m[359]), .B(c[359]), .Z(n38772) );
  XOR U41134 ( .A(n38773), .B(n38774), .Z(n38765) );
  ANDN U41135 ( .B(n38775), .A(n31462), .Z(n38773) );
  XNOR U41136 ( .A(\modmult_1/zin[0][357] ), .B(n38776), .Z(n31462) );
  IV U41137 ( .A(n38774), .Z(n38776) );
  XOR U41138 ( .A(n38774), .B(n31463), .Z(n38775) );
  XNOR U41139 ( .A(n38777), .B(n38778), .Z(n31463) );
  ANDN U41140 ( .B(\modmult_1/xin[1023] ), .A(n38779), .Z(n38777) );
  IV U41141 ( .A(n38778), .Z(n38779) );
  XNOR U41142 ( .A(m[358]), .B(n38780), .Z(n38778) );
  NAND U41143 ( .A(n38781), .B(mul_pow), .Z(n38780) );
  XOR U41144 ( .A(m[358]), .B(c[358]), .Z(n38781) );
  XOR U41145 ( .A(n38782), .B(n38783), .Z(n38774) );
  ANDN U41146 ( .B(n38784), .A(n31460), .Z(n38782) );
  XNOR U41147 ( .A(\modmult_1/zin[0][356] ), .B(n38785), .Z(n31460) );
  IV U41148 ( .A(n38783), .Z(n38785) );
  XOR U41149 ( .A(n38783), .B(n31461), .Z(n38784) );
  XNOR U41150 ( .A(n38786), .B(n38787), .Z(n31461) );
  ANDN U41151 ( .B(\modmult_1/xin[1023] ), .A(n38788), .Z(n38786) );
  IV U41152 ( .A(n38787), .Z(n38788) );
  XNOR U41153 ( .A(m[357]), .B(n38789), .Z(n38787) );
  NAND U41154 ( .A(n38790), .B(mul_pow), .Z(n38789) );
  XOR U41155 ( .A(m[357]), .B(c[357]), .Z(n38790) );
  XOR U41156 ( .A(n38791), .B(n38792), .Z(n38783) );
  ANDN U41157 ( .B(n38793), .A(n31458), .Z(n38791) );
  XNOR U41158 ( .A(\modmult_1/zin[0][355] ), .B(n38794), .Z(n31458) );
  IV U41159 ( .A(n38792), .Z(n38794) );
  XOR U41160 ( .A(n38792), .B(n31459), .Z(n38793) );
  XNOR U41161 ( .A(n38795), .B(n38796), .Z(n31459) );
  ANDN U41162 ( .B(\modmult_1/xin[1023] ), .A(n38797), .Z(n38795) );
  IV U41163 ( .A(n38796), .Z(n38797) );
  XNOR U41164 ( .A(m[356]), .B(n38798), .Z(n38796) );
  NAND U41165 ( .A(n38799), .B(mul_pow), .Z(n38798) );
  XOR U41166 ( .A(m[356]), .B(c[356]), .Z(n38799) );
  XOR U41167 ( .A(n38800), .B(n38801), .Z(n38792) );
  ANDN U41168 ( .B(n38802), .A(n31456), .Z(n38800) );
  XNOR U41169 ( .A(\modmult_1/zin[0][354] ), .B(n38803), .Z(n31456) );
  IV U41170 ( .A(n38801), .Z(n38803) );
  XOR U41171 ( .A(n38801), .B(n31457), .Z(n38802) );
  XNOR U41172 ( .A(n38804), .B(n38805), .Z(n31457) );
  ANDN U41173 ( .B(\modmult_1/xin[1023] ), .A(n38806), .Z(n38804) );
  IV U41174 ( .A(n38805), .Z(n38806) );
  XNOR U41175 ( .A(m[355]), .B(n38807), .Z(n38805) );
  NAND U41176 ( .A(n38808), .B(mul_pow), .Z(n38807) );
  XOR U41177 ( .A(m[355]), .B(c[355]), .Z(n38808) );
  XOR U41178 ( .A(n38809), .B(n38810), .Z(n38801) );
  ANDN U41179 ( .B(n38811), .A(n31454), .Z(n38809) );
  XNOR U41180 ( .A(\modmult_1/zin[0][353] ), .B(n38812), .Z(n31454) );
  IV U41181 ( .A(n38810), .Z(n38812) );
  XOR U41182 ( .A(n38810), .B(n31455), .Z(n38811) );
  XNOR U41183 ( .A(n38813), .B(n38814), .Z(n31455) );
  ANDN U41184 ( .B(\modmult_1/xin[1023] ), .A(n38815), .Z(n38813) );
  IV U41185 ( .A(n38814), .Z(n38815) );
  XNOR U41186 ( .A(m[354]), .B(n38816), .Z(n38814) );
  NAND U41187 ( .A(n38817), .B(mul_pow), .Z(n38816) );
  XOR U41188 ( .A(m[354]), .B(c[354]), .Z(n38817) );
  XOR U41189 ( .A(n38818), .B(n38819), .Z(n38810) );
  ANDN U41190 ( .B(n38820), .A(n31452), .Z(n38818) );
  XNOR U41191 ( .A(\modmult_1/zin[0][352] ), .B(n38821), .Z(n31452) );
  IV U41192 ( .A(n38819), .Z(n38821) );
  XOR U41193 ( .A(n38819), .B(n31453), .Z(n38820) );
  XNOR U41194 ( .A(n38822), .B(n38823), .Z(n31453) );
  ANDN U41195 ( .B(\modmult_1/xin[1023] ), .A(n38824), .Z(n38822) );
  IV U41196 ( .A(n38823), .Z(n38824) );
  XNOR U41197 ( .A(m[353]), .B(n38825), .Z(n38823) );
  NAND U41198 ( .A(n38826), .B(mul_pow), .Z(n38825) );
  XOR U41199 ( .A(m[353]), .B(c[353]), .Z(n38826) );
  XOR U41200 ( .A(n38827), .B(n38828), .Z(n38819) );
  ANDN U41201 ( .B(n38829), .A(n31450), .Z(n38827) );
  XNOR U41202 ( .A(\modmult_1/zin[0][351] ), .B(n38830), .Z(n31450) );
  IV U41203 ( .A(n38828), .Z(n38830) );
  XOR U41204 ( .A(n38828), .B(n31451), .Z(n38829) );
  XNOR U41205 ( .A(n38831), .B(n38832), .Z(n31451) );
  ANDN U41206 ( .B(\modmult_1/xin[1023] ), .A(n38833), .Z(n38831) );
  IV U41207 ( .A(n38832), .Z(n38833) );
  XNOR U41208 ( .A(m[352]), .B(n38834), .Z(n38832) );
  NAND U41209 ( .A(n38835), .B(mul_pow), .Z(n38834) );
  XOR U41210 ( .A(m[352]), .B(c[352]), .Z(n38835) );
  XOR U41211 ( .A(n38836), .B(n38837), .Z(n38828) );
  ANDN U41212 ( .B(n38838), .A(n31448), .Z(n38836) );
  XNOR U41213 ( .A(\modmult_1/zin[0][350] ), .B(n38839), .Z(n31448) );
  IV U41214 ( .A(n38837), .Z(n38839) );
  XOR U41215 ( .A(n38837), .B(n31449), .Z(n38838) );
  XNOR U41216 ( .A(n38840), .B(n38841), .Z(n31449) );
  ANDN U41217 ( .B(\modmult_1/xin[1023] ), .A(n38842), .Z(n38840) );
  IV U41218 ( .A(n38841), .Z(n38842) );
  XNOR U41219 ( .A(m[351]), .B(n38843), .Z(n38841) );
  NAND U41220 ( .A(n38844), .B(mul_pow), .Z(n38843) );
  XOR U41221 ( .A(m[351]), .B(c[351]), .Z(n38844) );
  XOR U41222 ( .A(n38845), .B(n38846), .Z(n38837) );
  ANDN U41223 ( .B(n38847), .A(n31446), .Z(n38845) );
  XNOR U41224 ( .A(\modmult_1/zin[0][349] ), .B(n38848), .Z(n31446) );
  IV U41225 ( .A(n38846), .Z(n38848) );
  XOR U41226 ( .A(n38846), .B(n31447), .Z(n38847) );
  XNOR U41227 ( .A(n38849), .B(n38850), .Z(n31447) );
  ANDN U41228 ( .B(\modmult_1/xin[1023] ), .A(n38851), .Z(n38849) );
  IV U41229 ( .A(n38850), .Z(n38851) );
  XNOR U41230 ( .A(m[350]), .B(n38852), .Z(n38850) );
  NAND U41231 ( .A(n38853), .B(mul_pow), .Z(n38852) );
  XOR U41232 ( .A(m[350]), .B(c[350]), .Z(n38853) );
  XOR U41233 ( .A(n38854), .B(n38855), .Z(n38846) );
  ANDN U41234 ( .B(n38856), .A(n31444), .Z(n38854) );
  XNOR U41235 ( .A(\modmult_1/zin[0][348] ), .B(n38857), .Z(n31444) );
  IV U41236 ( .A(n38855), .Z(n38857) );
  XOR U41237 ( .A(n38855), .B(n31445), .Z(n38856) );
  XNOR U41238 ( .A(n38858), .B(n38859), .Z(n31445) );
  ANDN U41239 ( .B(\modmult_1/xin[1023] ), .A(n38860), .Z(n38858) );
  IV U41240 ( .A(n38859), .Z(n38860) );
  XNOR U41241 ( .A(m[349]), .B(n38861), .Z(n38859) );
  NAND U41242 ( .A(n38862), .B(mul_pow), .Z(n38861) );
  XOR U41243 ( .A(m[349]), .B(c[349]), .Z(n38862) );
  XOR U41244 ( .A(n38863), .B(n38864), .Z(n38855) );
  ANDN U41245 ( .B(n38865), .A(n31442), .Z(n38863) );
  XNOR U41246 ( .A(\modmult_1/zin[0][347] ), .B(n38866), .Z(n31442) );
  IV U41247 ( .A(n38864), .Z(n38866) );
  XOR U41248 ( .A(n38864), .B(n31443), .Z(n38865) );
  XNOR U41249 ( .A(n38867), .B(n38868), .Z(n31443) );
  ANDN U41250 ( .B(\modmult_1/xin[1023] ), .A(n38869), .Z(n38867) );
  IV U41251 ( .A(n38868), .Z(n38869) );
  XNOR U41252 ( .A(m[348]), .B(n38870), .Z(n38868) );
  NAND U41253 ( .A(n38871), .B(mul_pow), .Z(n38870) );
  XOR U41254 ( .A(m[348]), .B(c[348]), .Z(n38871) );
  XOR U41255 ( .A(n38872), .B(n38873), .Z(n38864) );
  ANDN U41256 ( .B(n38874), .A(n31440), .Z(n38872) );
  XNOR U41257 ( .A(\modmult_1/zin[0][346] ), .B(n38875), .Z(n31440) );
  IV U41258 ( .A(n38873), .Z(n38875) );
  XOR U41259 ( .A(n38873), .B(n31441), .Z(n38874) );
  XNOR U41260 ( .A(n38876), .B(n38877), .Z(n31441) );
  ANDN U41261 ( .B(\modmult_1/xin[1023] ), .A(n38878), .Z(n38876) );
  IV U41262 ( .A(n38877), .Z(n38878) );
  XNOR U41263 ( .A(m[347]), .B(n38879), .Z(n38877) );
  NAND U41264 ( .A(n38880), .B(mul_pow), .Z(n38879) );
  XOR U41265 ( .A(m[347]), .B(c[347]), .Z(n38880) );
  XOR U41266 ( .A(n38881), .B(n38882), .Z(n38873) );
  ANDN U41267 ( .B(n38883), .A(n31438), .Z(n38881) );
  XNOR U41268 ( .A(\modmult_1/zin[0][345] ), .B(n38884), .Z(n31438) );
  IV U41269 ( .A(n38882), .Z(n38884) );
  XOR U41270 ( .A(n38882), .B(n31439), .Z(n38883) );
  XNOR U41271 ( .A(n38885), .B(n38886), .Z(n31439) );
  ANDN U41272 ( .B(\modmult_1/xin[1023] ), .A(n38887), .Z(n38885) );
  IV U41273 ( .A(n38886), .Z(n38887) );
  XNOR U41274 ( .A(m[346]), .B(n38888), .Z(n38886) );
  NAND U41275 ( .A(n38889), .B(mul_pow), .Z(n38888) );
  XOR U41276 ( .A(m[346]), .B(c[346]), .Z(n38889) );
  XOR U41277 ( .A(n38890), .B(n38891), .Z(n38882) );
  ANDN U41278 ( .B(n38892), .A(n31436), .Z(n38890) );
  XNOR U41279 ( .A(\modmult_1/zin[0][344] ), .B(n38893), .Z(n31436) );
  IV U41280 ( .A(n38891), .Z(n38893) );
  XOR U41281 ( .A(n38891), .B(n31437), .Z(n38892) );
  XNOR U41282 ( .A(n38894), .B(n38895), .Z(n31437) );
  ANDN U41283 ( .B(\modmult_1/xin[1023] ), .A(n38896), .Z(n38894) );
  IV U41284 ( .A(n38895), .Z(n38896) );
  XNOR U41285 ( .A(m[345]), .B(n38897), .Z(n38895) );
  NAND U41286 ( .A(n38898), .B(mul_pow), .Z(n38897) );
  XOR U41287 ( .A(m[345]), .B(c[345]), .Z(n38898) );
  XOR U41288 ( .A(n38899), .B(n38900), .Z(n38891) );
  ANDN U41289 ( .B(n38901), .A(n31434), .Z(n38899) );
  XNOR U41290 ( .A(\modmult_1/zin[0][343] ), .B(n38902), .Z(n31434) );
  IV U41291 ( .A(n38900), .Z(n38902) );
  XOR U41292 ( .A(n38900), .B(n31435), .Z(n38901) );
  XNOR U41293 ( .A(n38903), .B(n38904), .Z(n31435) );
  ANDN U41294 ( .B(\modmult_1/xin[1023] ), .A(n38905), .Z(n38903) );
  IV U41295 ( .A(n38904), .Z(n38905) );
  XNOR U41296 ( .A(m[344]), .B(n38906), .Z(n38904) );
  NAND U41297 ( .A(n38907), .B(mul_pow), .Z(n38906) );
  XOR U41298 ( .A(m[344]), .B(c[344]), .Z(n38907) );
  XOR U41299 ( .A(n38908), .B(n38909), .Z(n38900) );
  ANDN U41300 ( .B(n38910), .A(n31432), .Z(n38908) );
  XNOR U41301 ( .A(\modmult_1/zin[0][342] ), .B(n38911), .Z(n31432) );
  IV U41302 ( .A(n38909), .Z(n38911) );
  XOR U41303 ( .A(n38909), .B(n31433), .Z(n38910) );
  XNOR U41304 ( .A(n38912), .B(n38913), .Z(n31433) );
  ANDN U41305 ( .B(\modmult_1/xin[1023] ), .A(n38914), .Z(n38912) );
  IV U41306 ( .A(n38913), .Z(n38914) );
  XNOR U41307 ( .A(m[343]), .B(n38915), .Z(n38913) );
  NAND U41308 ( .A(n38916), .B(mul_pow), .Z(n38915) );
  XOR U41309 ( .A(m[343]), .B(c[343]), .Z(n38916) );
  XOR U41310 ( .A(n38917), .B(n38918), .Z(n38909) );
  ANDN U41311 ( .B(n38919), .A(n31430), .Z(n38917) );
  XNOR U41312 ( .A(\modmult_1/zin[0][341] ), .B(n38920), .Z(n31430) );
  IV U41313 ( .A(n38918), .Z(n38920) );
  XOR U41314 ( .A(n38918), .B(n31431), .Z(n38919) );
  XNOR U41315 ( .A(n38921), .B(n38922), .Z(n31431) );
  ANDN U41316 ( .B(\modmult_1/xin[1023] ), .A(n38923), .Z(n38921) );
  IV U41317 ( .A(n38922), .Z(n38923) );
  XNOR U41318 ( .A(m[342]), .B(n38924), .Z(n38922) );
  NAND U41319 ( .A(n38925), .B(mul_pow), .Z(n38924) );
  XOR U41320 ( .A(m[342]), .B(c[342]), .Z(n38925) );
  XOR U41321 ( .A(n38926), .B(n38927), .Z(n38918) );
  ANDN U41322 ( .B(n38928), .A(n31428), .Z(n38926) );
  XNOR U41323 ( .A(\modmult_1/zin[0][340] ), .B(n38929), .Z(n31428) );
  IV U41324 ( .A(n38927), .Z(n38929) );
  XOR U41325 ( .A(n38927), .B(n31429), .Z(n38928) );
  XNOR U41326 ( .A(n38930), .B(n38931), .Z(n31429) );
  ANDN U41327 ( .B(\modmult_1/xin[1023] ), .A(n38932), .Z(n38930) );
  IV U41328 ( .A(n38931), .Z(n38932) );
  XNOR U41329 ( .A(m[341]), .B(n38933), .Z(n38931) );
  NAND U41330 ( .A(n38934), .B(mul_pow), .Z(n38933) );
  XOR U41331 ( .A(m[341]), .B(c[341]), .Z(n38934) );
  XOR U41332 ( .A(n38935), .B(n38936), .Z(n38927) );
  ANDN U41333 ( .B(n38937), .A(n31426), .Z(n38935) );
  XNOR U41334 ( .A(\modmult_1/zin[0][339] ), .B(n38938), .Z(n31426) );
  IV U41335 ( .A(n38936), .Z(n38938) );
  XOR U41336 ( .A(n38936), .B(n31427), .Z(n38937) );
  XNOR U41337 ( .A(n38939), .B(n38940), .Z(n31427) );
  ANDN U41338 ( .B(\modmult_1/xin[1023] ), .A(n38941), .Z(n38939) );
  IV U41339 ( .A(n38940), .Z(n38941) );
  XNOR U41340 ( .A(m[340]), .B(n38942), .Z(n38940) );
  NAND U41341 ( .A(n38943), .B(mul_pow), .Z(n38942) );
  XOR U41342 ( .A(m[340]), .B(c[340]), .Z(n38943) );
  XOR U41343 ( .A(n38944), .B(n38945), .Z(n38936) );
  ANDN U41344 ( .B(n38946), .A(n31424), .Z(n38944) );
  XNOR U41345 ( .A(\modmult_1/zin[0][338] ), .B(n38947), .Z(n31424) );
  IV U41346 ( .A(n38945), .Z(n38947) );
  XOR U41347 ( .A(n38945), .B(n31425), .Z(n38946) );
  XNOR U41348 ( .A(n38948), .B(n38949), .Z(n31425) );
  ANDN U41349 ( .B(\modmult_1/xin[1023] ), .A(n38950), .Z(n38948) );
  IV U41350 ( .A(n38949), .Z(n38950) );
  XNOR U41351 ( .A(m[339]), .B(n38951), .Z(n38949) );
  NAND U41352 ( .A(n38952), .B(mul_pow), .Z(n38951) );
  XOR U41353 ( .A(m[339]), .B(c[339]), .Z(n38952) );
  XOR U41354 ( .A(n38953), .B(n38954), .Z(n38945) );
  ANDN U41355 ( .B(n38955), .A(n31422), .Z(n38953) );
  XNOR U41356 ( .A(\modmult_1/zin[0][337] ), .B(n38956), .Z(n31422) );
  IV U41357 ( .A(n38954), .Z(n38956) );
  XOR U41358 ( .A(n38954), .B(n31423), .Z(n38955) );
  XNOR U41359 ( .A(n38957), .B(n38958), .Z(n31423) );
  ANDN U41360 ( .B(\modmult_1/xin[1023] ), .A(n38959), .Z(n38957) );
  IV U41361 ( .A(n38958), .Z(n38959) );
  XNOR U41362 ( .A(m[338]), .B(n38960), .Z(n38958) );
  NAND U41363 ( .A(n38961), .B(mul_pow), .Z(n38960) );
  XOR U41364 ( .A(m[338]), .B(c[338]), .Z(n38961) );
  XOR U41365 ( .A(n38962), .B(n38963), .Z(n38954) );
  ANDN U41366 ( .B(n38964), .A(n31420), .Z(n38962) );
  XNOR U41367 ( .A(\modmult_1/zin[0][336] ), .B(n38965), .Z(n31420) );
  IV U41368 ( .A(n38963), .Z(n38965) );
  XOR U41369 ( .A(n38963), .B(n31421), .Z(n38964) );
  XNOR U41370 ( .A(n38966), .B(n38967), .Z(n31421) );
  ANDN U41371 ( .B(\modmult_1/xin[1023] ), .A(n38968), .Z(n38966) );
  IV U41372 ( .A(n38967), .Z(n38968) );
  XNOR U41373 ( .A(m[337]), .B(n38969), .Z(n38967) );
  NAND U41374 ( .A(n38970), .B(mul_pow), .Z(n38969) );
  XOR U41375 ( .A(m[337]), .B(c[337]), .Z(n38970) );
  XOR U41376 ( .A(n38971), .B(n38972), .Z(n38963) );
  ANDN U41377 ( .B(n38973), .A(n31418), .Z(n38971) );
  XNOR U41378 ( .A(\modmult_1/zin[0][335] ), .B(n38974), .Z(n31418) );
  IV U41379 ( .A(n38972), .Z(n38974) );
  XOR U41380 ( .A(n38972), .B(n31419), .Z(n38973) );
  XNOR U41381 ( .A(n38975), .B(n38976), .Z(n31419) );
  ANDN U41382 ( .B(\modmult_1/xin[1023] ), .A(n38977), .Z(n38975) );
  IV U41383 ( .A(n38976), .Z(n38977) );
  XNOR U41384 ( .A(m[336]), .B(n38978), .Z(n38976) );
  NAND U41385 ( .A(n38979), .B(mul_pow), .Z(n38978) );
  XOR U41386 ( .A(m[336]), .B(c[336]), .Z(n38979) );
  XOR U41387 ( .A(n38980), .B(n38981), .Z(n38972) );
  ANDN U41388 ( .B(n38982), .A(n31416), .Z(n38980) );
  XNOR U41389 ( .A(\modmult_1/zin[0][334] ), .B(n38983), .Z(n31416) );
  IV U41390 ( .A(n38981), .Z(n38983) );
  XOR U41391 ( .A(n38981), .B(n31417), .Z(n38982) );
  XNOR U41392 ( .A(n38984), .B(n38985), .Z(n31417) );
  ANDN U41393 ( .B(\modmult_1/xin[1023] ), .A(n38986), .Z(n38984) );
  IV U41394 ( .A(n38985), .Z(n38986) );
  XNOR U41395 ( .A(m[335]), .B(n38987), .Z(n38985) );
  NAND U41396 ( .A(n38988), .B(mul_pow), .Z(n38987) );
  XOR U41397 ( .A(m[335]), .B(c[335]), .Z(n38988) );
  XOR U41398 ( .A(n38989), .B(n38990), .Z(n38981) );
  ANDN U41399 ( .B(n38991), .A(n31414), .Z(n38989) );
  XNOR U41400 ( .A(\modmult_1/zin[0][333] ), .B(n38992), .Z(n31414) );
  IV U41401 ( .A(n38990), .Z(n38992) );
  XOR U41402 ( .A(n38990), .B(n31415), .Z(n38991) );
  XNOR U41403 ( .A(n38993), .B(n38994), .Z(n31415) );
  ANDN U41404 ( .B(\modmult_1/xin[1023] ), .A(n38995), .Z(n38993) );
  IV U41405 ( .A(n38994), .Z(n38995) );
  XNOR U41406 ( .A(m[334]), .B(n38996), .Z(n38994) );
  NAND U41407 ( .A(n38997), .B(mul_pow), .Z(n38996) );
  XOR U41408 ( .A(m[334]), .B(c[334]), .Z(n38997) );
  XOR U41409 ( .A(n38998), .B(n38999), .Z(n38990) );
  ANDN U41410 ( .B(n39000), .A(n31412), .Z(n38998) );
  XNOR U41411 ( .A(\modmult_1/zin[0][332] ), .B(n39001), .Z(n31412) );
  IV U41412 ( .A(n38999), .Z(n39001) );
  XOR U41413 ( .A(n38999), .B(n31413), .Z(n39000) );
  XNOR U41414 ( .A(n39002), .B(n39003), .Z(n31413) );
  ANDN U41415 ( .B(\modmult_1/xin[1023] ), .A(n39004), .Z(n39002) );
  IV U41416 ( .A(n39003), .Z(n39004) );
  XNOR U41417 ( .A(m[333]), .B(n39005), .Z(n39003) );
  NAND U41418 ( .A(n39006), .B(mul_pow), .Z(n39005) );
  XOR U41419 ( .A(m[333]), .B(c[333]), .Z(n39006) );
  XOR U41420 ( .A(n39007), .B(n39008), .Z(n38999) );
  ANDN U41421 ( .B(n39009), .A(n31410), .Z(n39007) );
  XNOR U41422 ( .A(\modmult_1/zin[0][331] ), .B(n39010), .Z(n31410) );
  IV U41423 ( .A(n39008), .Z(n39010) );
  XOR U41424 ( .A(n39008), .B(n31411), .Z(n39009) );
  XNOR U41425 ( .A(n39011), .B(n39012), .Z(n31411) );
  ANDN U41426 ( .B(\modmult_1/xin[1023] ), .A(n39013), .Z(n39011) );
  IV U41427 ( .A(n39012), .Z(n39013) );
  XNOR U41428 ( .A(m[332]), .B(n39014), .Z(n39012) );
  NAND U41429 ( .A(n39015), .B(mul_pow), .Z(n39014) );
  XOR U41430 ( .A(m[332]), .B(c[332]), .Z(n39015) );
  XOR U41431 ( .A(n39016), .B(n39017), .Z(n39008) );
  ANDN U41432 ( .B(n39018), .A(n31408), .Z(n39016) );
  XNOR U41433 ( .A(\modmult_1/zin[0][330] ), .B(n39019), .Z(n31408) );
  IV U41434 ( .A(n39017), .Z(n39019) );
  XOR U41435 ( .A(n39017), .B(n31409), .Z(n39018) );
  XNOR U41436 ( .A(n39020), .B(n39021), .Z(n31409) );
  ANDN U41437 ( .B(\modmult_1/xin[1023] ), .A(n39022), .Z(n39020) );
  IV U41438 ( .A(n39021), .Z(n39022) );
  XNOR U41439 ( .A(m[331]), .B(n39023), .Z(n39021) );
  NAND U41440 ( .A(n39024), .B(mul_pow), .Z(n39023) );
  XOR U41441 ( .A(m[331]), .B(c[331]), .Z(n39024) );
  XOR U41442 ( .A(n39025), .B(n39026), .Z(n39017) );
  ANDN U41443 ( .B(n39027), .A(n31406), .Z(n39025) );
  XNOR U41444 ( .A(\modmult_1/zin[0][329] ), .B(n39028), .Z(n31406) );
  IV U41445 ( .A(n39026), .Z(n39028) );
  XOR U41446 ( .A(n39026), .B(n31407), .Z(n39027) );
  XNOR U41447 ( .A(n39029), .B(n39030), .Z(n31407) );
  ANDN U41448 ( .B(\modmult_1/xin[1023] ), .A(n39031), .Z(n39029) );
  IV U41449 ( .A(n39030), .Z(n39031) );
  XNOR U41450 ( .A(m[330]), .B(n39032), .Z(n39030) );
  NAND U41451 ( .A(n39033), .B(mul_pow), .Z(n39032) );
  XOR U41452 ( .A(m[330]), .B(c[330]), .Z(n39033) );
  XOR U41453 ( .A(n39034), .B(n39035), .Z(n39026) );
  ANDN U41454 ( .B(n39036), .A(n31404), .Z(n39034) );
  XNOR U41455 ( .A(\modmult_1/zin[0][328] ), .B(n39037), .Z(n31404) );
  IV U41456 ( .A(n39035), .Z(n39037) );
  XOR U41457 ( .A(n39035), .B(n31405), .Z(n39036) );
  XNOR U41458 ( .A(n39038), .B(n39039), .Z(n31405) );
  ANDN U41459 ( .B(\modmult_1/xin[1023] ), .A(n39040), .Z(n39038) );
  IV U41460 ( .A(n39039), .Z(n39040) );
  XNOR U41461 ( .A(m[329]), .B(n39041), .Z(n39039) );
  NAND U41462 ( .A(n39042), .B(mul_pow), .Z(n39041) );
  XOR U41463 ( .A(m[329]), .B(c[329]), .Z(n39042) );
  XOR U41464 ( .A(n39043), .B(n39044), .Z(n39035) );
  ANDN U41465 ( .B(n39045), .A(n31402), .Z(n39043) );
  XNOR U41466 ( .A(\modmult_1/zin[0][327] ), .B(n39046), .Z(n31402) );
  IV U41467 ( .A(n39044), .Z(n39046) );
  XOR U41468 ( .A(n39044), .B(n31403), .Z(n39045) );
  XNOR U41469 ( .A(n39047), .B(n39048), .Z(n31403) );
  ANDN U41470 ( .B(\modmult_1/xin[1023] ), .A(n39049), .Z(n39047) );
  IV U41471 ( .A(n39048), .Z(n39049) );
  XNOR U41472 ( .A(m[328]), .B(n39050), .Z(n39048) );
  NAND U41473 ( .A(n39051), .B(mul_pow), .Z(n39050) );
  XOR U41474 ( .A(m[328]), .B(c[328]), .Z(n39051) );
  XOR U41475 ( .A(n39052), .B(n39053), .Z(n39044) );
  ANDN U41476 ( .B(n39054), .A(n31400), .Z(n39052) );
  XNOR U41477 ( .A(\modmult_1/zin[0][326] ), .B(n39055), .Z(n31400) );
  IV U41478 ( .A(n39053), .Z(n39055) );
  XOR U41479 ( .A(n39053), .B(n31401), .Z(n39054) );
  XNOR U41480 ( .A(n39056), .B(n39057), .Z(n31401) );
  ANDN U41481 ( .B(\modmult_1/xin[1023] ), .A(n39058), .Z(n39056) );
  IV U41482 ( .A(n39057), .Z(n39058) );
  XNOR U41483 ( .A(m[327]), .B(n39059), .Z(n39057) );
  NAND U41484 ( .A(n39060), .B(mul_pow), .Z(n39059) );
  XOR U41485 ( .A(m[327]), .B(c[327]), .Z(n39060) );
  XOR U41486 ( .A(n39061), .B(n39062), .Z(n39053) );
  ANDN U41487 ( .B(n39063), .A(n31398), .Z(n39061) );
  XNOR U41488 ( .A(\modmult_1/zin[0][325] ), .B(n39064), .Z(n31398) );
  IV U41489 ( .A(n39062), .Z(n39064) );
  XOR U41490 ( .A(n39062), .B(n31399), .Z(n39063) );
  XNOR U41491 ( .A(n39065), .B(n39066), .Z(n31399) );
  ANDN U41492 ( .B(\modmult_1/xin[1023] ), .A(n39067), .Z(n39065) );
  IV U41493 ( .A(n39066), .Z(n39067) );
  XNOR U41494 ( .A(m[326]), .B(n39068), .Z(n39066) );
  NAND U41495 ( .A(n39069), .B(mul_pow), .Z(n39068) );
  XOR U41496 ( .A(m[326]), .B(c[326]), .Z(n39069) );
  XOR U41497 ( .A(n39070), .B(n39071), .Z(n39062) );
  ANDN U41498 ( .B(n39072), .A(n31396), .Z(n39070) );
  XNOR U41499 ( .A(\modmult_1/zin[0][324] ), .B(n39073), .Z(n31396) );
  IV U41500 ( .A(n39071), .Z(n39073) );
  XOR U41501 ( .A(n39071), .B(n31397), .Z(n39072) );
  XNOR U41502 ( .A(n39074), .B(n39075), .Z(n31397) );
  ANDN U41503 ( .B(\modmult_1/xin[1023] ), .A(n39076), .Z(n39074) );
  IV U41504 ( .A(n39075), .Z(n39076) );
  XNOR U41505 ( .A(m[325]), .B(n39077), .Z(n39075) );
  NAND U41506 ( .A(n39078), .B(mul_pow), .Z(n39077) );
  XOR U41507 ( .A(m[325]), .B(c[325]), .Z(n39078) );
  XOR U41508 ( .A(n39079), .B(n39080), .Z(n39071) );
  ANDN U41509 ( .B(n39081), .A(n31394), .Z(n39079) );
  XNOR U41510 ( .A(\modmult_1/zin[0][323] ), .B(n39082), .Z(n31394) );
  IV U41511 ( .A(n39080), .Z(n39082) );
  XOR U41512 ( .A(n39080), .B(n31395), .Z(n39081) );
  XNOR U41513 ( .A(n39083), .B(n39084), .Z(n31395) );
  ANDN U41514 ( .B(\modmult_1/xin[1023] ), .A(n39085), .Z(n39083) );
  IV U41515 ( .A(n39084), .Z(n39085) );
  XNOR U41516 ( .A(m[324]), .B(n39086), .Z(n39084) );
  NAND U41517 ( .A(n39087), .B(mul_pow), .Z(n39086) );
  XOR U41518 ( .A(m[324]), .B(c[324]), .Z(n39087) );
  XOR U41519 ( .A(n39088), .B(n39089), .Z(n39080) );
  ANDN U41520 ( .B(n39090), .A(n31392), .Z(n39088) );
  XNOR U41521 ( .A(\modmult_1/zin[0][322] ), .B(n39091), .Z(n31392) );
  IV U41522 ( .A(n39089), .Z(n39091) );
  XOR U41523 ( .A(n39089), .B(n31393), .Z(n39090) );
  XNOR U41524 ( .A(n39092), .B(n39093), .Z(n31393) );
  ANDN U41525 ( .B(\modmult_1/xin[1023] ), .A(n39094), .Z(n39092) );
  IV U41526 ( .A(n39093), .Z(n39094) );
  XNOR U41527 ( .A(m[323]), .B(n39095), .Z(n39093) );
  NAND U41528 ( .A(n39096), .B(mul_pow), .Z(n39095) );
  XOR U41529 ( .A(m[323]), .B(c[323]), .Z(n39096) );
  XOR U41530 ( .A(n39097), .B(n39098), .Z(n39089) );
  ANDN U41531 ( .B(n39099), .A(n31390), .Z(n39097) );
  XNOR U41532 ( .A(\modmult_1/zin[0][321] ), .B(n39100), .Z(n31390) );
  IV U41533 ( .A(n39098), .Z(n39100) );
  XOR U41534 ( .A(n39098), .B(n31391), .Z(n39099) );
  XNOR U41535 ( .A(n39101), .B(n39102), .Z(n31391) );
  ANDN U41536 ( .B(\modmult_1/xin[1023] ), .A(n39103), .Z(n39101) );
  IV U41537 ( .A(n39102), .Z(n39103) );
  XNOR U41538 ( .A(m[322]), .B(n39104), .Z(n39102) );
  NAND U41539 ( .A(n39105), .B(mul_pow), .Z(n39104) );
  XOR U41540 ( .A(m[322]), .B(c[322]), .Z(n39105) );
  XOR U41541 ( .A(n39106), .B(n39107), .Z(n39098) );
  ANDN U41542 ( .B(n39108), .A(n31388), .Z(n39106) );
  XNOR U41543 ( .A(\modmult_1/zin[0][320] ), .B(n39109), .Z(n31388) );
  IV U41544 ( .A(n39107), .Z(n39109) );
  XOR U41545 ( .A(n39107), .B(n31389), .Z(n39108) );
  XNOR U41546 ( .A(n39110), .B(n39111), .Z(n31389) );
  ANDN U41547 ( .B(\modmult_1/xin[1023] ), .A(n39112), .Z(n39110) );
  IV U41548 ( .A(n39111), .Z(n39112) );
  XNOR U41549 ( .A(m[321]), .B(n39113), .Z(n39111) );
  NAND U41550 ( .A(n39114), .B(mul_pow), .Z(n39113) );
  XOR U41551 ( .A(m[321]), .B(c[321]), .Z(n39114) );
  XOR U41552 ( .A(n39115), .B(n39116), .Z(n39107) );
  ANDN U41553 ( .B(n39117), .A(n31386), .Z(n39115) );
  XNOR U41554 ( .A(\modmult_1/zin[0][319] ), .B(n39118), .Z(n31386) );
  IV U41555 ( .A(n39116), .Z(n39118) );
  XOR U41556 ( .A(n39116), .B(n31387), .Z(n39117) );
  XNOR U41557 ( .A(n39119), .B(n39120), .Z(n31387) );
  ANDN U41558 ( .B(\modmult_1/xin[1023] ), .A(n39121), .Z(n39119) );
  IV U41559 ( .A(n39120), .Z(n39121) );
  XNOR U41560 ( .A(m[320]), .B(n39122), .Z(n39120) );
  NAND U41561 ( .A(n39123), .B(mul_pow), .Z(n39122) );
  XOR U41562 ( .A(m[320]), .B(c[320]), .Z(n39123) );
  XOR U41563 ( .A(n39124), .B(n39125), .Z(n39116) );
  ANDN U41564 ( .B(n39126), .A(n31384), .Z(n39124) );
  XNOR U41565 ( .A(\modmult_1/zin[0][318] ), .B(n39127), .Z(n31384) );
  IV U41566 ( .A(n39125), .Z(n39127) );
  XOR U41567 ( .A(n39125), .B(n31385), .Z(n39126) );
  XNOR U41568 ( .A(n39128), .B(n39129), .Z(n31385) );
  ANDN U41569 ( .B(\modmult_1/xin[1023] ), .A(n39130), .Z(n39128) );
  IV U41570 ( .A(n39129), .Z(n39130) );
  XNOR U41571 ( .A(m[319]), .B(n39131), .Z(n39129) );
  NAND U41572 ( .A(n39132), .B(mul_pow), .Z(n39131) );
  XOR U41573 ( .A(m[319]), .B(c[319]), .Z(n39132) );
  XOR U41574 ( .A(n39133), .B(n39134), .Z(n39125) );
  ANDN U41575 ( .B(n39135), .A(n31382), .Z(n39133) );
  XNOR U41576 ( .A(\modmult_1/zin[0][317] ), .B(n39136), .Z(n31382) );
  IV U41577 ( .A(n39134), .Z(n39136) );
  XOR U41578 ( .A(n39134), .B(n31383), .Z(n39135) );
  XNOR U41579 ( .A(n39137), .B(n39138), .Z(n31383) );
  ANDN U41580 ( .B(\modmult_1/xin[1023] ), .A(n39139), .Z(n39137) );
  IV U41581 ( .A(n39138), .Z(n39139) );
  XNOR U41582 ( .A(m[318]), .B(n39140), .Z(n39138) );
  NAND U41583 ( .A(n39141), .B(mul_pow), .Z(n39140) );
  XOR U41584 ( .A(m[318]), .B(c[318]), .Z(n39141) );
  XOR U41585 ( .A(n39142), .B(n39143), .Z(n39134) );
  ANDN U41586 ( .B(n39144), .A(n31380), .Z(n39142) );
  XNOR U41587 ( .A(\modmult_1/zin[0][316] ), .B(n39145), .Z(n31380) );
  IV U41588 ( .A(n39143), .Z(n39145) );
  XOR U41589 ( .A(n39143), .B(n31381), .Z(n39144) );
  XNOR U41590 ( .A(n39146), .B(n39147), .Z(n31381) );
  ANDN U41591 ( .B(\modmult_1/xin[1023] ), .A(n39148), .Z(n39146) );
  IV U41592 ( .A(n39147), .Z(n39148) );
  XNOR U41593 ( .A(m[317]), .B(n39149), .Z(n39147) );
  NAND U41594 ( .A(n39150), .B(mul_pow), .Z(n39149) );
  XOR U41595 ( .A(m[317]), .B(c[317]), .Z(n39150) );
  XOR U41596 ( .A(n39151), .B(n39152), .Z(n39143) );
  ANDN U41597 ( .B(n39153), .A(n31378), .Z(n39151) );
  XNOR U41598 ( .A(\modmult_1/zin[0][315] ), .B(n39154), .Z(n31378) );
  IV U41599 ( .A(n39152), .Z(n39154) );
  XOR U41600 ( .A(n39152), .B(n31379), .Z(n39153) );
  XNOR U41601 ( .A(n39155), .B(n39156), .Z(n31379) );
  ANDN U41602 ( .B(\modmult_1/xin[1023] ), .A(n39157), .Z(n39155) );
  IV U41603 ( .A(n39156), .Z(n39157) );
  XNOR U41604 ( .A(m[316]), .B(n39158), .Z(n39156) );
  NAND U41605 ( .A(n39159), .B(mul_pow), .Z(n39158) );
  XOR U41606 ( .A(m[316]), .B(c[316]), .Z(n39159) );
  XOR U41607 ( .A(n39160), .B(n39161), .Z(n39152) );
  ANDN U41608 ( .B(n39162), .A(n31376), .Z(n39160) );
  XNOR U41609 ( .A(\modmult_1/zin[0][314] ), .B(n39163), .Z(n31376) );
  IV U41610 ( .A(n39161), .Z(n39163) );
  XOR U41611 ( .A(n39161), .B(n31377), .Z(n39162) );
  XNOR U41612 ( .A(n39164), .B(n39165), .Z(n31377) );
  ANDN U41613 ( .B(\modmult_1/xin[1023] ), .A(n39166), .Z(n39164) );
  IV U41614 ( .A(n39165), .Z(n39166) );
  XNOR U41615 ( .A(m[315]), .B(n39167), .Z(n39165) );
  NAND U41616 ( .A(n39168), .B(mul_pow), .Z(n39167) );
  XOR U41617 ( .A(m[315]), .B(c[315]), .Z(n39168) );
  XOR U41618 ( .A(n39169), .B(n39170), .Z(n39161) );
  ANDN U41619 ( .B(n39171), .A(n31374), .Z(n39169) );
  XNOR U41620 ( .A(\modmult_1/zin[0][313] ), .B(n39172), .Z(n31374) );
  IV U41621 ( .A(n39170), .Z(n39172) );
  XOR U41622 ( .A(n39170), .B(n31375), .Z(n39171) );
  XNOR U41623 ( .A(n39173), .B(n39174), .Z(n31375) );
  ANDN U41624 ( .B(\modmult_1/xin[1023] ), .A(n39175), .Z(n39173) );
  IV U41625 ( .A(n39174), .Z(n39175) );
  XNOR U41626 ( .A(m[314]), .B(n39176), .Z(n39174) );
  NAND U41627 ( .A(n39177), .B(mul_pow), .Z(n39176) );
  XOR U41628 ( .A(m[314]), .B(c[314]), .Z(n39177) );
  XOR U41629 ( .A(n39178), .B(n39179), .Z(n39170) );
  ANDN U41630 ( .B(n39180), .A(n31372), .Z(n39178) );
  XNOR U41631 ( .A(\modmult_1/zin[0][312] ), .B(n39181), .Z(n31372) );
  IV U41632 ( .A(n39179), .Z(n39181) );
  XOR U41633 ( .A(n39179), .B(n31373), .Z(n39180) );
  XNOR U41634 ( .A(n39182), .B(n39183), .Z(n31373) );
  ANDN U41635 ( .B(\modmult_1/xin[1023] ), .A(n39184), .Z(n39182) );
  IV U41636 ( .A(n39183), .Z(n39184) );
  XNOR U41637 ( .A(m[313]), .B(n39185), .Z(n39183) );
  NAND U41638 ( .A(n39186), .B(mul_pow), .Z(n39185) );
  XOR U41639 ( .A(m[313]), .B(c[313]), .Z(n39186) );
  XOR U41640 ( .A(n39187), .B(n39188), .Z(n39179) );
  ANDN U41641 ( .B(n39189), .A(n31370), .Z(n39187) );
  XNOR U41642 ( .A(\modmult_1/zin[0][311] ), .B(n39190), .Z(n31370) );
  IV U41643 ( .A(n39188), .Z(n39190) );
  XOR U41644 ( .A(n39188), .B(n31371), .Z(n39189) );
  XNOR U41645 ( .A(n39191), .B(n39192), .Z(n31371) );
  ANDN U41646 ( .B(\modmult_1/xin[1023] ), .A(n39193), .Z(n39191) );
  IV U41647 ( .A(n39192), .Z(n39193) );
  XNOR U41648 ( .A(m[312]), .B(n39194), .Z(n39192) );
  NAND U41649 ( .A(n39195), .B(mul_pow), .Z(n39194) );
  XOR U41650 ( .A(m[312]), .B(c[312]), .Z(n39195) );
  XOR U41651 ( .A(n39196), .B(n39197), .Z(n39188) );
  ANDN U41652 ( .B(n39198), .A(n31368), .Z(n39196) );
  XNOR U41653 ( .A(\modmult_1/zin[0][310] ), .B(n39199), .Z(n31368) );
  IV U41654 ( .A(n39197), .Z(n39199) );
  XOR U41655 ( .A(n39197), .B(n31369), .Z(n39198) );
  XNOR U41656 ( .A(n39200), .B(n39201), .Z(n31369) );
  ANDN U41657 ( .B(\modmult_1/xin[1023] ), .A(n39202), .Z(n39200) );
  IV U41658 ( .A(n39201), .Z(n39202) );
  XNOR U41659 ( .A(m[311]), .B(n39203), .Z(n39201) );
  NAND U41660 ( .A(n39204), .B(mul_pow), .Z(n39203) );
  XOR U41661 ( .A(m[311]), .B(c[311]), .Z(n39204) );
  XOR U41662 ( .A(n39205), .B(n39206), .Z(n39197) );
  ANDN U41663 ( .B(n39207), .A(n31366), .Z(n39205) );
  XNOR U41664 ( .A(\modmult_1/zin[0][309] ), .B(n39208), .Z(n31366) );
  IV U41665 ( .A(n39206), .Z(n39208) );
  XOR U41666 ( .A(n39206), .B(n31367), .Z(n39207) );
  XNOR U41667 ( .A(n39209), .B(n39210), .Z(n31367) );
  ANDN U41668 ( .B(\modmult_1/xin[1023] ), .A(n39211), .Z(n39209) );
  IV U41669 ( .A(n39210), .Z(n39211) );
  XNOR U41670 ( .A(m[310]), .B(n39212), .Z(n39210) );
  NAND U41671 ( .A(n39213), .B(mul_pow), .Z(n39212) );
  XOR U41672 ( .A(m[310]), .B(c[310]), .Z(n39213) );
  XOR U41673 ( .A(n39214), .B(n39215), .Z(n39206) );
  ANDN U41674 ( .B(n39216), .A(n31364), .Z(n39214) );
  XNOR U41675 ( .A(\modmult_1/zin[0][308] ), .B(n39217), .Z(n31364) );
  IV U41676 ( .A(n39215), .Z(n39217) );
  XOR U41677 ( .A(n39215), .B(n31365), .Z(n39216) );
  XNOR U41678 ( .A(n39218), .B(n39219), .Z(n31365) );
  ANDN U41679 ( .B(\modmult_1/xin[1023] ), .A(n39220), .Z(n39218) );
  IV U41680 ( .A(n39219), .Z(n39220) );
  XNOR U41681 ( .A(m[309]), .B(n39221), .Z(n39219) );
  NAND U41682 ( .A(n39222), .B(mul_pow), .Z(n39221) );
  XOR U41683 ( .A(m[309]), .B(c[309]), .Z(n39222) );
  XOR U41684 ( .A(n39223), .B(n39224), .Z(n39215) );
  ANDN U41685 ( .B(n39225), .A(n31362), .Z(n39223) );
  XNOR U41686 ( .A(\modmult_1/zin[0][307] ), .B(n39226), .Z(n31362) );
  IV U41687 ( .A(n39224), .Z(n39226) );
  XOR U41688 ( .A(n39224), .B(n31363), .Z(n39225) );
  XNOR U41689 ( .A(n39227), .B(n39228), .Z(n31363) );
  ANDN U41690 ( .B(\modmult_1/xin[1023] ), .A(n39229), .Z(n39227) );
  IV U41691 ( .A(n39228), .Z(n39229) );
  XNOR U41692 ( .A(m[308]), .B(n39230), .Z(n39228) );
  NAND U41693 ( .A(n39231), .B(mul_pow), .Z(n39230) );
  XOR U41694 ( .A(m[308]), .B(c[308]), .Z(n39231) );
  XOR U41695 ( .A(n39232), .B(n39233), .Z(n39224) );
  ANDN U41696 ( .B(n39234), .A(n31360), .Z(n39232) );
  XNOR U41697 ( .A(\modmult_1/zin[0][306] ), .B(n39235), .Z(n31360) );
  IV U41698 ( .A(n39233), .Z(n39235) );
  XOR U41699 ( .A(n39233), .B(n31361), .Z(n39234) );
  XNOR U41700 ( .A(n39236), .B(n39237), .Z(n31361) );
  ANDN U41701 ( .B(\modmult_1/xin[1023] ), .A(n39238), .Z(n39236) );
  IV U41702 ( .A(n39237), .Z(n39238) );
  XNOR U41703 ( .A(m[307]), .B(n39239), .Z(n39237) );
  NAND U41704 ( .A(n39240), .B(mul_pow), .Z(n39239) );
  XOR U41705 ( .A(m[307]), .B(c[307]), .Z(n39240) );
  XOR U41706 ( .A(n39241), .B(n39242), .Z(n39233) );
  ANDN U41707 ( .B(n39243), .A(n31358), .Z(n39241) );
  XNOR U41708 ( .A(\modmult_1/zin[0][305] ), .B(n39244), .Z(n31358) );
  IV U41709 ( .A(n39242), .Z(n39244) );
  XOR U41710 ( .A(n39242), .B(n31359), .Z(n39243) );
  XNOR U41711 ( .A(n39245), .B(n39246), .Z(n31359) );
  ANDN U41712 ( .B(\modmult_1/xin[1023] ), .A(n39247), .Z(n39245) );
  IV U41713 ( .A(n39246), .Z(n39247) );
  XNOR U41714 ( .A(m[306]), .B(n39248), .Z(n39246) );
  NAND U41715 ( .A(n39249), .B(mul_pow), .Z(n39248) );
  XOR U41716 ( .A(m[306]), .B(c[306]), .Z(n39249) );
  XOR U41717 ( .A(n39250), .B(n39251), .Z(n39242) );
  ANDN U41718 ( .B(n39252), .A(n31356), .Z(n39250) );
  XNOR U41719 ( .A(\modmult_1/zin[0][304] ), .B(n39253), .Z(n31356) );
  IV U41720 ( .A(n39251), .Z(n39253) );
  XOR U41721 ( .A(n39251), .B(n31357), .Z(n39252) );
  XNOR U41722 ( .A(n39254), .B(n39255), .Z(n31357) );
  ANDN U41723 ( .B(\modmult_1/xin[1023] ), .A(n39256), .Z(n39254) );
  IV U41724 ( .A(n39255), .Z(n39256) );
  XNOR U41725 ( .A(m[305]), .B(n39257), .Z(n39255) );
  NAND U41726 ( .A(n39258), .B(mul_pow), .Z(n39257) );
  XOR U41727 ( .A(m[305]), .B(c[305]), .Z(n39258) );
  XOR U41728 ( .A(n39259), .B(n39260), .Z(n39251) );
  ANDN U41729 ( .B(n39261), .A(n31354), .Z(n39259) );
  XNOR U41730 ( .A(\modmult_1/zin[0][303] ), .B(n39262), .Z(n31354) );
  IV U41731 ( .A(n39260), .Z(n39262) );
  XOR U41732 ( .A(n39260), .B(n31355), .Z(n39261) );
  XNOR U41733 ( .A(n39263), .B(n39264), .Z(n31355) );
  ANDN U41734 ( .B(\modmult_1/xin[1023] ), .A(n39265), .Z(n39263) );
  IV U41735 ( .A(n39264), .Z(n39265) );
  XNOR U41736 ( .A(m[304]), .B(n39266), .Z(n39264) );
  NAND U41737 ( .A(n39267), .B(mul_pow), .Z(n39266) );
  XOR U41738 ( .A(m[304]), .B(c[304]), .Z(n39267) );
  XOR U41739 ( .A(n39268), .B(n39269), .Z(n39260) );
  ANDN U41740 ( .B(n39270), .A(n31352), .Z(n39268) );
  XNOR U41741 ( .A(\modmult_1/zin[0][302] ), .B(n39271), .Z(n31352) );
  IV U41742 ( .A(n39269), .Z(n39271) );
  XOR U41743 ( .A(n39269), .B(n31353), .Z(n39270) );
  XNOR U41744 ( .A(n39272), .B(n39273), .Z(n31353) );
  ANDN U41745 ( .B(\modmult_1/xin[1023] ), .A(n39274), .Z(n39272) );
  IV U41746 ( .A(n39273), .Z(n39274) );
  XNOR U41747 ( .A(m[303]), .B(n39275), .Z(n39273) );
  NAND U41748 ( .A(n39276), .B(mul_pow), .Z(n39275) );
  XOR U41749 ( .A(m[303]), .B(c[303]), .Z(n39276) );
  XOR U41750 ( .A(n39277), .B(n39278), .Z(n39269) );
  ANDN U41751 ( .B(n39279), .A(n31350), .Z(n39277) );
  XNOR U41752 ( .A(\modmult_1/zin[0][301] ), .B(n39280), .Z(n31350) );
  IV U41753 ( .A(n39278), .Z(n39280) );
  XOR U41754 ( .A(n39278), .B(n31351), .Z(n39279) );
  XNOR U41755 ( .A(n39281), .B(n39282), .Z(n31351) );
  ANDN U41756 ( .B(\modmult_1/xin[1023] ), .A(n39283), .Z(n39281) );
  IV U41757 ( .A(n39282), .Z(n39283) );
  XNOR U41758 ( .A(m[302]), .B(n39284), .Z(n39282) );
  NAND U41759 ( .A(n39285), .B(mul_pow), .Z(n39284) );
  XOR U41760 ( .A(m[302]), .B(c[302]), .Z(n39285) );
  XOR U41761 ( .A(n39286), .B(n39287), .Z(n39278) );
  ANDN U41762 ( .B(n39288), .A(n31348), .Z(n39286) );
  XNOR U41763 ( .A(\modmult_1/zin[0][300] ), .B(n39289), .Z(n31348) );
  IV U41764 ( .A(n39287), .Z(n39289) );
  XOR U41765 ( .A(n39287), .B(n31349), .Z(n39288) );
  XNOR U41766 ( .A(n39290), .B(n39291), .Z(n31349) );
  ANDN U41767 ( .B(\modmult_1/xin[1023] ), .A(n39292), .Z(n39290) );
  IV U41768 ( .A(n39291), .Z(n39292) );
  XNOR U41769 ( .A(m[301]), .B(n39293), .Z(n39291) );
  NAND U41770 ( .A(n39294), .B(mul_pow), .Z(n39293) );
  XOR U41771 ( .A(m[301]), .B(c[301]), .Z(n39294) );
  XOR U41772 ( .A(n39295), .B(n39296), .Z(n39287) );
  ANDN U41773 ( .B(n39297), .A(n31346), .Z(n39295) );
  XNOR U41774 ( .A(\modmult_1/zin[0][299] ), .B(n39298), .Z(n31346) );
  IV U41775 ( .A(n39296), .Z(n39298) );
  XOR U41776 ( .A(n39296), .B(n31347), .Z(n39297) );
  XNOR U41777 ( .A(n39299), .B(n39300), .Z(n31347) );
  ANDN U41778 ( .B(\modmult_1/xin[1023] ), .A(n39301), .Z(n39299) );
  IV U41779 ( .A(n39300), .Z(n39301) );
  XNOR U41780 ( .A(m[300]), .B(n39302), .Z(n39300) );
  NAND U41781 ( .A(n39303), .B(mul_pow), .Z(n39302) );
  XOR U41782 ( .A(m[300]), .B(c[300]), .Z(n39303) );
  XOR U41783 ( .A(n39304), .B(n39305), .Z(n39296) );
  ANDN U41784 ( .B(n39306), .A(n31344), .Z(n39304) );
  XNOR U41785 ( .A(\modmult_1/zin[0][298] ), .B(n39307), .Z(n31344) );
  IV U41786 ( .A(n39305), .Z(n39307) );
  XOR U41787 ( .A(n39305), .B(n31345), .Z(n39306) );
  XNOR U41788 ( .A(n39308), .B(n39309), .Z(n31345) );
  ANDN U41789 ( .B(\modmult_1/xin[1023] ), .A(n39310), .Z(n39308) );
  IV U41790 ( .A(n39309), .Z(n39310) );
  XNOR U41791 ( .A(m[299]), .B(n39311), .Z(n39309) );
  NAND U41792 ( .A(n39312), .B(mul_pow), .Z(n39311) );
  XOR U41793 ( .A(m[299]), .B(c[299]), .Z(n39312) );
  XOR U41794 ( .A(n39313), .B(n39314), .Z(n39305) );
  ANDN U41795 ( .B(n39315), .A(n31342), .Z(n39313) );
  XNOR U41796 ( .A(\modmult_1/zin[0][297] ), .B(n39316), .Z(n31342) );
  IV U41797 ( .A(n39314), .Z(n39316) );
  XOR U41798 ( .A(n39314), .B(n31343), .Z(n39315) );
  XNOR U41799 ( .A(n39317), .B(n39318), .Z(n31343) );
  ANDN U41800 ( .B(\modmult_1/xin[1023] ), .A(n39319), .Z(n39317) );
  IV U41801 ( .A(n39318), .Z(n39319) );
  XNOR U41802 ( .A(m[298]), .B(n39320), .Z(n39318) );
  NAND U41803 ( .A(n39321), .B(mul_pow), .Z(n39320) );
  XOR U41804 ( .A(m[298]), .B(c[298]), .Z(n39321) );
  XOR U41805 ( .A(n39322), .B(n39323), .Z(n39314) );
  ANDN U41806 ( .B(n39324), .A(n31340), .Z(n39322) );
  XNOR U41807 ( .A(\modmult_1/zin[0][296] ), .B(n39325), .Z(n31340) );
  IV U41808 ( .A(n39323), .Z(n39325) );
  XOR U41809 ( .A(n39323), .B(n31341), .Z(n39324) );
  XNOR U41810 ( .A(n39326), .B(n39327), .Z(n31341) );
  ANDN U41811 ( .B(\modmult_1/xin[1023] ), .A(n39328), .Z(n39326) );
  IV U41812 ( .A(n39327), .Z(n39328) );
  XNOR U41813 ( .A(m[297]), .B(n39329), .Z(n39327) );
  NAND U41814 ( .A(n39330), .B(mul_pow), .Z(n39329) );
  XOR U41815 ( .A(m[297]), .B(c[297]), .Z(n39330) );
  XOR U41816 ( .A(n39331), .B(n39332), .Z(n39323) );
  ANDN U41817 ( .B(n39333), .A(n31338), .Z(n39331) );
  XNOR U41818 ( .A(\modmult_1/zin[0][295] ), .B(n39334), .Z(n31338) );
  IV U41819 ( .A(n39332), .Z(n39334) );
  XOR U41820 ( .A(n39332), .B(n31339), .Z(n39333) );
  XNOR U41821 ( .A(n39335), .B(n39336), .Z(n31339) );
  ANDN U41822 ( .B(\modmult_1/xin[1023] ), .A(n39337), .Z(n39335) );
  IV U41823 ( .A(n39336), .Z(n39337) );
  XNOR U41824 ( .A(m[296]), .B(n39338), .Z(n39336) );
  NAND U41825 ( .A(n39339), .B(mul_pow), .Z(n39338) );
  XOR U41826 ( .A(m[296]), .B(c[296]), .Z(n39339) );
  XOR U41827 ( .A(n39340), .B(n39341), .Z(n39332) );
  ANDN U41828 ( .B(n39342), .A(n31336), .Z(n39340) );
  XNOR U41829 ( .A(\modmult_1/zin[0][294] ), .B(n39343), .Z(n31336) );
  IV U41830 ( .A(n39341), .Z(n39343) );
  XOR U41831 ( .A(n39341), .B(n31337), .Z(n39342) );
  XNOR U41832 ( .A(n39344), .B(n39345), .Z(n31337) );
  ANDN U41833 ( .B(\modmult_1/xin[1023] ), .A(n39346), .Z(n39344) );
  IV U41834 ( .A(n39345), .Z(n39346) );
  XNOR U41835 ( .A(m[295]), .B(n39347), .Z(n39345) );
  NAND U41836 ( .A(n39348), .B(mul_pow), .Z(n39347) );
  XOR U41837 ( .A(m[295]), .B(c[295]), .Z(n39348) );
  XOR U41838 ( .A(n39349), .B(n39350), .Z(n39341) );
  ANDN U41839 ( .B(n39351), .A(n31334), .Z(n39349) );
  XNOR U41840 ( .A(\modmult_1/zin[0][293] ), .B(n39352), .Z(n31334) );
  IV U41841 ( .A(n39350), .Z(n39352) );
  XOR U41842 ( .A(n39350), .B(n31335), .Z(n39351) );
  XNOR U41843 ( .A(n39353), .B(n39354), .Z(n31335) );
  ANDN U41844 ( .B(\modmult_1/xin[1023] ), .A(n39355), .Z(n39353) );
  IV U41845 ( .A(n39354), .Z(n39355) );
  XNOR U41846 ( .A(m[294]), .B(n39356), .Z(n39354) );
  NAND U41847 ( .A(n39357), .B(mul_pow), .Z(n39356) );
  XOR U41848 ( .A(m[294]), .B(c[294]), .Z(n39357) );
  XOR U41849 ( .A(n39358), .B(n39359), .Z(n39350) );
  ANDN U41850 ( .B(n39360), .A(n31332), .Z(n39358) );
  XNOR U41851 ( .A(\modmult_1/zin[0][292] ), .B(n39361), .Z(n31332) );
  IV U41852 ( .A(n39359), .Z(n39361) );
  XOR U41853 ( .A(n39359), .B(n31333), .Z(n39360) );
  XNOR U41854 ( .A(n39362), .B(n39363), .Z(n31333) );
  ANDN U41855 ( .B(\modmult_1/xin[1023] ), .A(n39364), .Z(n39362) );
  IV U41856 ( .A(n39363), .Z(n39364) );
  XNOR U41857 ( .A(m[293]), .B(n39365), .Z(n39363) );
  NAND U41858 ( .A(n39366), .B(mul_pow), .Z(n39365) );
  XOR U41859 ( .A(m[293]), .B(c[293]), .Z(n39366) );
  XOR U41860 ( .A(n39367), .B(n39368), .Z(n39359) );
  ANDN U41861 ( .B(n39369), .A(n31330), .Z(n39367) );
  XNOR U41862 ( .A(\modmult_1/zin[0][291] ), .B(n39370), .Z(n31330) );
  IV U41863 ( .A(n39368), .Z(n39370) );
  XOR U41864 ( .A(n39368), .B(n31331), .Z(n39369) );
  XNOR U41865 ( .A(n39371), .B(n39372), .Z(n31331) );
  ANDN U41866 ( .B(\modmult_1/xin[1023] ), .A(n39373), .Z(n39371) );
  IV U41867 ( .A(n39372), .Z(n39373) );
  XNOR U41868 ( .A(m[292]), .B(n39374), .Z(n39372) );
  NAND U41869 ( .A(n39375), .B(mul_pow), .Z(n39374) );
  XOR U41870 ( .A(m[292]), .B(c[292]), .Z(n39375) );
  XOR U41871 ( .A(n39376), .B(n39377), .Z(n39368) );
  ANDN U41872 ( .B(n39378), .A(n31328), .Z(n39376) );
  XNOR U41873 ( .A(\modmult_1/zin[0][290] ), .B(n39379), .Z(n31328) );
  IV U41874 ( .A(n39377), .Z(n39379) );
  XOR U41875 ( .A(n39377), .B(n31329), .Z(n39378) );
  XNOR U41876 ( .A(n39380), .B(n39381), .Z(n31329) );
  ANDN U41877 ( .B(\modmult_1/xin[1023] ), .A(n39382), .Z(n39380) );
  IV U41878 ( .A(n39381), .Z(n39382) );
  XNOR U41879 ( .A(m[291]), .B(n39383), .Z(n39381) );
  NAND U41880 ( .A(n39384), .B(mul_pow), .Z(n39383) );
  XOR U41881 ( .A(m[291]), .B(c[291]), .Z(n39384) );
  XOR U41882 ( .A(n39385), .B(n39386), .Z(n39377) );
  ANDN U41883 ( .B(n39387), .A(n31326), .Z(n39385) );
  XNOR U41884 ( .A(\modmult_1/zin[0][289] ), .B(n39388), .Z(n31326) );
  IV U41885 ( .A(n39386), .Z(n39388) );
  XOR U41886 ( .A(n39386), .B(n31327), .Z(n39387) );
  XNOR U41887 ( .A(n39389), .B(n39390), .Z(n31327) );
  ANDN U41888 ( .B(\modmult_1/xin[1023] ), .A(n39391), .Z(n39389) );
  IV U41889 ( .A(n39390), .Z(n39391) );
  XNOR U41890 ( .A(m[290]), .B(n39392), .Z(n39390) );
  NAND U41891 ( .A(n39393), .B(mul_pow), .Z(n39392) );
  XOR U41892 ( .A(m[290]), .B(c[290]), .Z(n39393) );
  XOR U41893 ( .A(n39394), .B(n39395), .Z(n39386) );
  ANDN U41894 ( .B(n39396), .A(n31324), .Z(n39394) );
  XNOR U41895 ( .A(\modmult_1/zin[0][288] ), .B(n39397), .Z(n31324) );
  IV U41896 ( .A(n39395), .Z(n39397) );
  XOR U41897 ( .A(n39395), .B(n31325), .Z(n39396) );
  XNOR U41898 ( .A(n39398), .B(n39399), .Z(n31325) );
  ANDN U41899 ( .B(\modmult_1/xin[1023] ), .A(n39400), .Z(n39398) );
  IV U41900 ( .A(n39399), .Z(n39400) );
  XNOR U41901 ( .A(m[289]), .B(n39401), .Z(n39399) );
  NAND U41902 ( .A(n39402), .B(mul_pow), .Z(n39401) );
  XOR U41903 ( .A(m[289]), .B(c[289]), .Z(n39402) );
  XOR U41904 ( .A(n39403), .B(n39404), .Z(n39395) );
  ANDN U41905 ( .B(n39405), .A(n31322), .Z(n39403) );
  XNOR U41906 ( .A(\modmult_1/zin[0][287] ), .B(n39406), .Z(n31322) );
  IV U41907 ( .A(n39404), .Z(n39406) );
  XOR U41908 ( .A(n39404), .B(n31323), .Z(n39405) );
  XNOR U41909 ( .A(n39407), .B(n39408), .Z(n31323) );
  ANDN U41910 ( .B(\modmult_1/xin[1023] ), .A(n39409), .Z(n39407) );
  IV U41911 ( .A(n39408), .Z(n39409) );
  XNOR U41912 ( .A(m[288]), .B(n39410), .Z(n39408) );
  NAND U41913 ( .A(n39411), .B(mul_pow), .Z(n39410) );
  XOR U41914 ( .A(m[288]), .B(c[288]), .Z(n39411) );
  XOR U41915 ( .A(n39412), .B(n39413), .Z(n39404) );
  ANDN U41916 ( .B(n39414), .A(n31320), .Z(n39412) );
  XNOR U41917 ( .A(\modmult_1/zin[0][286] ), .B(n39415), .Z(n31320) );
  IV U41918 ( .A(n39413), .Z(n39415) );
  XOR U41919 ( .A(n39413), .B(n31321), .Z(n39414) );
  XNOR U41920 ( .A(n39416), .B(n39417), .Z(n31321) );
  ANDN U41921 ( .B(\modmult_1/xin[1023] ), .A(n39418), .Z(n39416) );
  IV U41922 ( .A(n39417), .Z(n39418) );
  XNOR U41923 ( .A(m[287]), .B(n39419), .Z(n39417) );
  NAND U41924 ( .A(n39420), .B(mul_pow), .Z(n39419) );
  XOR U41925 ( .A(m[287]), .B(c[287]), .Z(n39420) );
  XOR U41926 ( .A(n39421), .B(n39422), .Z(n39413) );
  ANDN U41927 ( .B(n39423), .A(n31318), .Z(n39421) );
  XNOR U41928 ( .A(\modmult_1/zin[0][285] ), .B(n39424), .Z(n31318) );
  IV U41929 ( .A(n39422), .Z(n39424) );
  XOR U41930 ( .A(n39422), .B(n31319), .Z(n39423) );
  XNOR U41931 ( .A(n39425), .B(n39426), .Z(n31319) );
  ANDN U41932 ( .B(\modmult_1/xin[1023] ), .A(n39427), .Z(n39425) );
  IV U41933 ( .A(n39426), .Z(n39427) );
  XNOR U41934 ( .A(m[286]), .B(n39428), .Z(n39426) );
  NAND U41935 ( .A(n39429), .B(mul_pow), .Z(n39428) );
  XOR U41936 ( .A(m[286]), .B(c[286]), .Z(n39429) );
  XOR U41937 ( .A(n39430), .B(n39431), .Z(n39422) );
  ANDN U41938 ( .B(n39432), .A(n31316), .Z(n39430) );
  XNOR U41939 ( .A(\modmult_1/zin[0][284] ), .B(n39433), .Z(n31316) );
  IV U41940 ( .A(n39431), .Z(n39433) );
  XOR U41941 ( .A(n39431), .B(n31317), .Z(n39432) );
  XNOR U41942 ( .A(n39434), .B(n39435), .Z(n31317) );
  ANDN U41943 ( .B(\modmult_1/xin[1023] ), .A(n39436), .Z(n39434) );
  IV U41944 ( .A(n39435), .Z(n39436) );
  XNOR U41945 ( .A(m[285]), .B(n39437), .Z(n39435) );
  NAND U41946 ( .A(n39438), .B(mul_pow), .Z(n39437) );
  XOR U41947 ( .A(m[285]), .B(c[285]), .Z(n39438) );
  XOR U41948 ( .A(n39439), .B(n39440), .Z(n39431) );
  ANDN U41949 ( .B(n39441), .A(n31314), .Z(n39439) );
  XNOR U41950 ( .A(\modmult_1/zin[0][283] ), .B(n39442), .Z(n31314) );
  IV U41951 ( .A(n39440), .Z(n39442) );
  XOR U41952 ( .A(n39440), .B(n31315), .Z(n39441) );
  XNOR U41953 ( .A(n39443), .B(n39444), .Z(n31315) );
  ANDN U41954 ( .B(\modmult_1/xin[1023] ), .A(n39445), .Z(n39443) );
  IV U41955 ( .A(n39444), .Z(n39445) );
  XNOR U41956 ( .A(m[284]), .B(n39446), .Z(n39444) );
  NAND U41957 ( .A(n39447), .B(mul_pow), .Z(n39446) );
  XOR U41958 ( .A(m[284]), .B(c[284]), .Z(n39447) );
  XOR U41959 ( .A(n39448), .B(n39449), .Z(n39440) );
  ANDN U41960 ( .B(n39450), .A(n31312), .Z(n39448) );
  XNOR U41961 ( .A(\modmult_1/zin[0][282] ), .B(n39451), .Z(n31312) );
  IV U41962 ( .A(n39449), .Z(n39451) );
  XOR U41963 ( .A(n39449), .B(n31313), .Z(n39450) );
  XNOR U41964 ( .A(n39452), .B(n39453), .Z(n31313) );
  ANDN U41965 ( .B(\modmult_1/xin[1023] ), .A(n39454), .Z(n39452) );
  IV U41966 ( .A(n39453), .Z(n39454) );
  XNOR U41967 ( .A(m[283]), .B(n39455), .Z(n39453) );
  NAND U41968 ( .A(n39456), .B(mul_pow), .Z(n39455) );
  XOR U41969 ( .A(m[283]), .B(c[283]), .Z(n39456) );
  XOR U41970 ( .A(n39457), .B(n39458), .Z(n39449) );
  ANDN U41971 ( .B(n39459), .A(n31310), .Z(n39457) );
  XNOR U41972 ( .A(\modmult_1/zin[0][281] ), .B(n39460), .Z(n31310) );
  IV U41973 ( .A(n39458), .Z(n39460) );
  XOR U41974 ( .A(n39458), .B(n31311), .Z(n39459) );
  XNOR U41975 ( .A(n39461), .B(n39462), .Z(n31311) );
  ANDN U41976 ( .B(\modmult_1/xin[1023] ), .A(n39463), .Z(n39461) );
  IV U41977 ( .A(n39462), .Z(n39463) );
  XNOR U41978 ( .A(m[282]), .B(n39464), .Z(n39462) );
  NAND U41979 ( .A(n39465), .B(mul_pow), .Z(n39464) );
  XOR U41980 ( .A(m[282]), .B(c[282]), .Z(n39465) );
  XOR U41981 ( .A(n39466), .B(n39467), .Z(n39458) );
  ANDN U41982 ( .B(n39468), .A(n31308), .Z(n39466) );
  XNOR U41983 ( .A(\modmult_1/zin[0][280] ), .B(n39469), .Z(n31308) );
  IV U41984 ( .A(n39467), .Z(n39469) );
  XOR U41985 ( .A(n39467), .B(n31309), .Z(n39468) );
  XNOR U41986 ( .A(n39470), .B(n39471), .Z(n31309) );
  ANDN U41987 ( .B(\modmult_1/xin[1023] ), .A(n39472), .Z(n39470) );
  IV U41988 ( .A(n39471), .Z(n39472) );
  XNOR U41989 ( .A(m[281]), .B(n39473), .Z(n39471) );
  NAND U41990 ( .A(n39474), .B(mul_pow), .Z(n39473) );
  XOR U41991 ( .A(m[281]), .B(c[281]), .Z(n39474) );
  XOR U41992 ( .A(n39475), .B(n39476), .Z(n39467) );
  ANDN U41993 ( .B(n39477), .A(n31306), .Z(n39475) );
  XNOR U41994 ( .A(\modmult_1/zin[0][279] ), .B(n39478), .Z(n31306) );
  IV U41995 ( .A(n39476), .Z(n39478) );
  XOR U41996 ( .A(n39476), .B(n31307), .Z(n39477) );
  XNOR U41997 ( .A(n39479), .B(n39480), .Z(n31307) );
  ANDN U41998 ( .B(\modmult_1/xin[1023] ), .A(n39481), .Z(n39479) );
  IV U41999 ( .A(n39480), .Z(n39481) );
  XNOR U42000 ( .A(m[280]), .B(n39482), .Z(n39480) );
  NAND U42001 ( .A(n39483), .B(mul_pow), .Z(n39482) );
  XOR U42002 ( .A(m[280]), .B(c[280]), .Z(n39483) );
  XOR U42003 ( .A(n39484), .B(n39485), .Z(n39476) );
  ANDN U42004 ( .B(n39486), .A(n31304), .Z(n39484) );
  XNOR U42005 ( .A(\modmult_1/zin[0][278] ), .B(n39487), .Z(n31304) );
  IV U42006 ( .A(n39485), .Z(n39487) );
  XOR U42007 ( .A(n39485), .B(n31305), .Z(n39486) );
  XNOR U42008 ( .A(n39488), .B(n39489), .Z(n31305) );
  ANDN U42009 ( .B(\modmult_1/xin[1023] ), .A(n39490), .Z(n39488) );
  IV U42010 ( .A(n39489), .Z(n39490) );
  XNOR U42011 ( .A(m[279]), .B(n39491), .Z(n39489) );
  NAND U42012 ( .A(n39492), .B(mul_pow), .Z(n39491) );
  XOR U42013 ( .A(m[279]), .B(c[279]), .Z(n39492) );
  XOR U42014 ( .A(n39493), .B(n39494), .Z(n39485) );
  ANDN U42015 ( .B(n39495), .A(n31302), .Z(n39493) );
  XNOR U42016 ( .A(\modmult_1/zin[0][277] ), .B(n39496), .Z(n31302) );
  IV U42017 ( .A(n39494), .Z(n39496) );
  XOR U42018 ( .A(n39494), .B(n31303), .Z(n39495) );
  XNOR U42019 ( .A(n39497), .B(n39498), .Z(n31303) );
  ANDN U42020 ( .B(\modmult_1/xin[1023] ), .A(n39499), .Z(n39497) );
  IV U42021 ( .A(n39498), .Z(n39499) );
  XNOR U42022 ( .A(m[278]), .B(n39500), .Z(n39498) );
  NAND U42023 ( .A(n39501), .B(mul_pow), .Z(n39500) );
  XOR U42024 ( .A(m[278]), .B(c[278]), .Z(n39501) );
  XOR U42025 ( .A(n39502), .B(n39503), .Z(n39494) );
  ANDN U42026 ( .B(n39504), .A(n31300), .Z(n39502) );
  XNOR U42027 ( .A(\modmult_1/zin[0][276] ), .B(n39505), .Z(n31300) );
  IV U42028 ( .A(n39503), .Z(n39505) );
  XOR U42029 ( .A(n39503), .B(n31301), .Z(n39504) );
  XNOR U42030 ( .A(n39506), .B(n39507), .Z(n31301) );
  ANDN U42031 ( .B(\modmult_1/xin[1023] ), .A(n39508), .Z(n39506) );
  IV U42032 ( .A(n39507), .Z(n39508) );
  XNOR U42033 ( .A(m[277]), .B(n39509), .Z(n39507) );
  NAND U42034 ( .A(n39510), .B(mul_pow), .Z(n39509) );
  XOR U42035 ( .A(m[277]), .B(c[277]), .Z(n39510) );
  XOR U42036 ( .A(n39511), .B(n39512), .Z(n39503) );
  ANDN U42037 ( .B(n39513), .A(n31298), .Z(n39511) );
  XNOR U42038 ( .A(\modmult_1/zin[0][275] ), .B(n39514), .Z(n31298) );
  IV U42039 ( .A(n39512), .Z(n39514) );
  XOR U42040 ( .A(n39512), .B(n31299), .Z(n39513) );
  XNOR U42041 ( .A(n39515), .B(n39516), .Z(n31299) );
  ANDN U42042 ( .B(\modmult_1/xin[1023] ), .A(n39517), .Z(n39515) );
  IV U42043 ( .A(n39516), .Z(n39517) );
  XNOR U42044 ( .A(m[276]), .B(n39518), .Z(n39516) );
  NAND U42045 ( .A(n39519), .B(mul_pow), .Z(n39518) );
  XOR U42046 ( .A(m[276]), .B(c[276]), .Z(n39519) );
  XOR U42047 ( .A(n39520), .B(n39521), .Z(n39512) );
  ANDN U42048 ( .B(n39522), .A(n31296), .Z(n39520) );
  XNOR U42049 ( .A(\modmult_1/zin[0][274] ), .B(n39523), .Z(n31296) );
  IV U42050 ( .A(n39521), .Z(n39523) );
  XOR U42051 ( .A(n39521), .B(n31297), .Z(n39522) );
  XNOR U42052 ( .A(n39524), .B(n39525), .Z(n31297) );
  ANDN U42053 ( .B(\modmult_1/xin[1023] ), .A(n39526), .Z(n39524) );
  IV U42054 ( .A(n39525), .Z(n39526) );
  XNOR U42055 ( .A(m[275]), .B(n39527), .Z(n39525) );
  NAND U42056 ( .A(n39528), .B(mul_pow), .Z(n39527) );
  XOR U42057 ( .A(m[275]), .B(c[275]), .Z(n39528) );
  XOR U42058 ( .A(n39529), .B(n39530), .Z(n39521) );
  ANDN U42059 ( .B(n39531), .A(n31294), .Z(n39529) );
  XNOR U42060 ( .A(\modmult_1/zin[0][273] ), .B(n39532), .Z(n31294) );
  IV U42061 ( .A(n39530), .Z(n39532) );
  XOR U42062 ( .A(n39530), .B(n31295), .Z(n39531) );
  XNOR U42063 ( .A(n39533), .B(n39534), .Z(n31295) );
  ANDN U42064 ( .B(\modmult_1/xin[1023] ), .A(n39535), .Z(n39533) );
  IV U42065 ( .A(n39534), .Z(n39535) );
  XNOR U42066 ( .A(m[274]), .B(n39536), .Z(n39534) );
  NAND U42067 ( .A(n39537), .B(mul_pow), .Z(n39536) );
  XOR U42068 ( .A(m[274]), .B(c[274]), .Z(n39537) );
  XOR U42069 ( .A(n39538), .B(n39539), .Z(n39530) );
  ANDN U42070 ( .B(n39540), .A(n31292), .Z(n39538) );
  XNOR U42071 ( .A(\modmult_1/zin[0][272] ), .B(n39541), .Z(n31292) );
  IV U42072 ( .A(n39539), .Z(n39541) );
  XOR U42073 ( .A(n39539), .B(n31293), .Z(n39540) );
  XNOR U42074 ( .A(n39542), .B(n39543), .Z(n31293) );
  ANDN U42075 ( .B(\modmult_1/xin[1023] ), .A(n39544), .Z(n39542) );
  IV U42076 ( .A(n39543), .Z(n39544) );
  XNOR U42077 ( .A(m[273]), .B(n39545), .Z(n39543) );
  NAND U42078 ( .A(n39546), .B(mul_pow), .Z(n39545) );
  XOR U42079 ( .A(m[273]), .B(c[273]), .Z(n39546) );
  XOR U42080 ( .A(n39547), .B(n39548), .Z(n39539) );
  ANDN U42081 ( .B(n39549), .A(n31290), .Z(n39547) );
  XNOR U42082 ( .A(\modmult_1/zin[0][271] ), .B(n39550), .Z(n31290) );
  IV U42083 ( .A(n39548), .Z(n39550) );
  XOR U42084 ( .A(n39548), .B(n31291), .Z(n39549) );
  XNOR U42085 ( .A(n39551), .B(n39552), .Z(n31291) );
  ANDN U42086 ( .B(\modmult_1/xin[1023] ), .A(n39553), .Z(n39551) );
  IV U42087 ( .A(n39552), .Z(n39553) );
  XNOR U42088 ( .A(m[272]), .B(n39554), .Z(n39552) );
  NAND U42089 ( .A(n39555), .B(mul_pow), .Z(n39554) );
  XOR U42090 ( .A(m[272]), .B(c[272]), .Z(n39555) );
  XOR U42091 ( .A(n39556), .B(n39557), .Z(n39548) );
  ANDN U42092 ( .B(n39558), .A(n31288), .Z(n39556) );
  XNOR U42093 ( .A(\modmult_1/zin[0][270] ), .B(n39559), .Z(n31288) );
  IV U42094 ( .A(n39557), .Z(n39559) );
  XOR U42095 ( .A(n39557), .B(n31289), .Z(n39558) );
  XNOR U42096 ( .A(n39560), .B(n39561), .Z(n31289) );
  ANDN U42097 ( .B(\modmult_1/xin[1023] ), .A(n39562), .Z(n39560) );
  IV U42098 ( .A(n39561), .Z(n39562) );
  XNOR U42099 ( .A(m[271]), .B(n39563), .Z(n39561) );
  NAND U42100 ( .A(n39564), .B(mul_pow), .Z(n39563) );
  XOR U42101 ( .A(m[271]), .B(c[271]), .Z(n39564) );
  XOR U42102 ( .A(n39565), .B(n39566), .Z(n39557) );
  ANDN U42103 ( .B(n39567), .A(n31286), .Z(n39565) );
  XNOR U42104 ( .A(\modmult_1/zin[0][269] ), .B(n39568), .Z(n31286) );
  IV U42105 ( .A(n39566), .Z(n39568) );
  XOR U42106 ( .A(n39566), .B(n31287), .Z(n39567) );
  XNOR U42107 ( .A(n39569), .B(n39570), .Z(n31287) );
  ANDN U42108 ( .B(\modmult_1/xin[1023] ), .A(n39571), .Z(n39569) );
  IV U42109 ( .A(n39570), .Z(n39571) );
  XNOR U42110 ( .A(m[270]), .B(n39572), .Z(n39570) );
  NAND U42111 ( .A(n39573), .B(mul_pow), .Z(n39572) );
  XOR U42112 ( .A(m[270]), .B(c[270]), .Z(n39573) );
  XOR U42113 ( .A(n39574), .B(n39575), .Z(n39566) );
  ANDN U42114 ( .B(n39576), .A(n31284), .Z(n39574) );
  XNOR U42115 ( .A(\modmult_1/zin[0][268] ), .B(n39577), .Z(n31284) );
  IV U42116 ( .A(n39575), .Z(n39577) );
  XOR U42117 ( .A(n39575), .B(n31285), .Z(n39576) );
  XNOR U42118 ( .A(n39578), .B(n39579), .Z(n31285) );
  ANDN U42119 ( .B(\modmult_1/xin[1023] ), .A(n39580), .Z(n39578) );
  IV U42120 ( .A(n39579), .Z(n39580) );
  XNOR U42121 ( .A(m[269]), .B(n39581), .Z(n39579) );
  NAND U42122 ( .A(n39582), .B(mul_pow), .Z(n39581) );
  XOR U42123 ( .A(m[269]), .B(c[269]), .Z(n39582) );
  XOR U42124 ( .A(n39583), .B(n39584), .Z(n39575) );
  ANDN U42125 ( .B(n39585), .A(n31282), .Z(n39583) );
  XNOR U42126 ( .A(\modmult_1/zin[0][267] ), .B(n39586), .Z(n31282) );
  IV U42127 ( .A(n39584), .Z(n39586) );
  XOR U42128 ( .A(n39584), .B(n31283), .Z(n39585) );
  XNOR U42129 ( .A(n39587), .B(n39588), .Z(n31283) );
  ANDN U42130 ( .B(\modmult_1/xin[1023] ), .A(n39589), .Z(n39587) );
  IV U42131 ( .A(n39588), .Z(n39589) );
  XNOR U42132 ( .A(m[268]), .B(n39590), .Z(n39588) );
  NAND U42133 ( .A(n39591), .B(mul_pow), .Z(n39590) );
  XOR U42134 ( .A(m[268]), .B(c[268]), .Z(n39591) );
  XOR U42135 ( .A(n39592), .B(n39593), .Z(n39584) );
  ANDN U42136 ( .B(n39594), .A(n31280), .Z(n39592) );
  XNOR U42137 ( .A(\modmult_1/zin[0][266] ), .B(n39595), .Z(n31280) );
  IV U42138 ( .A(n39593), .Z(n39595) );
  XOR U42139 ( .A(n39593), .B(n31281), .Z(n39594) );
  XNOR U42140 ( .A(n39596), .B(n39597), .Z(n31281) );
  ANDN U42141 ( .B(\modmult_1/xin[1023] ), .A(n39598), .Z(n39596) );
  IV U42142 ( .A(n39597), .Z(n39598) );
  XNOR U42143 ( .A(m[267]), .B(n39599), .Z(n39597) );
  NAND U42144 ( .A(n39600), .B(mul_pow), .Z(n39599) );
  XOR U42145 ( .A(m[267]), .B(c[267]), .Z(n39600) );
  XOR U42146 ( .A(n39601), .B(n39602), .Z(n39593) );
  ANDN U42147 ( .B(n39603), .A(n31278), .Z(n39601) );
  XNOR U42148 ( .A(\modmult_1/zin[0][265] ), .B(n39604), .Z(n31278) );
  IV U42149 ( .A(n39602), .Z(n39604) );
  XOR U42150 ( .A(n39602), .B(n31279), .Z(n39603) );
  XNOR U42151 ( .A(n39605), .B(n39606), .Z(n31279) );
  ANDN U42152 ( .B(\modmult_1/xin[1023] ), .A(n39607), .Z(n39605) );
  IV U42153 ( .A(n39606), .Z(n39607) );
  XNOR U42154 ( .A(m[266]), .B(n39608), .Z(n39606) );
  NAND U42155 ( .A(n39609), .B(mul_pow), .Z(n39608) );
  XOR U42156 ( .A(m[266]), .B(c[266]), .Z(n39609) );
  XOR U42157 ( .A(n39610), .B(n39611), .Z(n39602) );
  ANDN U42158 ( .B(n39612), .A(n31276), .Z(n39610) );
  XNOR U42159 ( .A(\modmult_1/zin[0][264] ), .B(n39613), .Z(n31276) );
  IV U42160 ( .A(n39611), .Z(n39613) );
  XOR U42161 ( .A(n39611), .B(n31277), .Z(n39612) );
  XNOR U42162 ( .A(n39614), .B(n39615), .Z(n31277) );
  ANDN U42163 ( .B(\modmult_1/xin[1023] ), .A(n39616), .Z(n39614) );
  IV U42164 ( .A(n39615), .Z(n39616) );
  XNOR U42165 ( .A(m[265]), .B(n39617), .Z(n39615) );
  NAND U42166 ( .A(n39618), .B(mul_pow), .Z(n39617) );
  XOR U42167 ( .A(m[265]), .B(c[265]), .Z(n39618) );
  XOR U42168 ( .A(n39619), .B(n39620), .Z(n39611) );
  ANDN U42169 ( .B(n39621), .A(n31274), .Z(n39619) );
  XNOR U42170 ( .A(\modmult_1/zin[0][263] ), .B(n39622), .Z(n31274) );
  IV U42171 ( .A(n39620), .Z(n39622) );
  XOR U42172 ( .A(n39620), .B(n31275), .Z(n39621) );
  XNOR U42173 ( .A(n39623), .B(n39624), .Z(n31275) );
  ANDN U42174 ( .B(\modmult_1/xin[1023] ), .A(n39625), .Z(n39623) );
  IV U42175 ( .A(n39624), .Z(n39625) );
  XNOR U42176 ( .A(m[264]), .B(n39626), .Z(n39624) );
  NAND U42177 ( .A(n39627), .B(mul_pow), .Z(n39626) );
  XOR U42178 ( .A(m[264]), .B(c[264]), .Z(n39627) );
  XOR U42179 ( .A(n39628), .B(n39629), .Z(n39620) );
  ANDN U42180 ( .B(n39630), .A(n31272), .Z(n39628) );
  XNOR U42181 ( .A(\modmult_1/zin[0][262] ), .B(n39631), .Z(n31272) );
  IV U42182 ( .A(n39629), .Z(n39631) );
  XOR U42183 ( .A(n39629), .B(n31273), .Z(n39630) );
  XNOR U42184 ( .A(n39632), .B(n39633), .Z(n31273) );
  ANDN U42185 ( .B(\modmult_1/xin[1023] ), .A(n39634), .Z(n39632) );
  IV U42186 ( .A(n39633), .Z(n39634) );
  XNOR U42187 ( .A(m[263]), .B(n39635), .Z(n39633) );
  NAND U42188 ( .A(n39636), .B(mul_pow), .Z(n39635) );
  XOR U42189 ( .A(m[263]), .B(c[263]), .Z(n39636) );
  XOR U42190 ( .A(n39637), .B(n39638), .Z(n39629) );
  ANDN U42191 ( .B(n39639), .A(n31270), .Z(n39637) );
  XNOR U42192 ( .A(\modmult_1/zin[0][261] ), .B(n39640), .Z(n31270) );
  IV U42193 ( .A(n39638), .Z(n39640) );
  XOR U42194 ( .A(n39638), .B(n31271), .Z(n39639) );
  XNOR U42195 ( .A(n39641), .B(n39642), .Z(n31271) );
  ANDN U42196 ( .B(\modmult_1/xin[1023] ), .A(n39643), .Z(n39641) );
  IV U42197 ( .A(n39642), .Z(n39643) );
  XNOR U42198 ( .A(m[262]), .B(n39644), .Z(n39642) );
  NAND U42199 ( .A(n39645), .B(mul_pow), .Z(n39644) );
  XOR U42200 ( .A(m[262]), .B(c[262]), .Z(n39645) );
  XOR U42201 ( .A(n39646), .B(n39647), .Z(n39638) );
  ANDN U42202 ( .B(n39648), .A(n31268), .Z(n39646) );
  XNOR U42203 ( .A(\modmult_1/zin[0][260] ), .B(n39649), .Z(n31268) );
  IV U42204 ( .A(n39647), .Z(n39649) );
  XOR U42205 ( .A(n39647), .B(n31269), .Z(n39648) );
  XNOR U42206 ( .A(n39650), .B(n39651), .Z(n31269) );
  ANDN U42207 ( .B(\modmult_1/xin[1023] ), .A(n39652), .Z(n39650) );
  IV U42208 ( .A(n39651), .Z(n39652) );
  XNOR U42209 ( .A(m[261]), .B(n39653), .Z(n39651) );
  NAND U42210 ( .A(n39654), .B(mul_pow), .Z(n39653) );
  XOR U42211 ( .A(m[261]), .B(c[261]), .Z(n39654) );
  XOR U42212 ( .A(n39655), .B(n39656), .Z(n39647) );
  ANDN U42213 ( .B(n39657), .A(n31266), .Z(n39655) );
  XNOR U42214 ( .A(\modmult_1/zin[0][259] ), .B(n39658), .Z(n31266) );
  IV U42215 ( .A(n39656), .Z(n39658) );
  XOR U42216 ( .A(n39656), .B(n31267), .Z(n39657) );
  XNOR U42217 ( .A(n39659), .B(n39660), .Z(n31267) );
  ANDN U42218 ( .B(\modmult_1/xin[1023] ), .A(n39661), .Z(n39659) );
  IV U42219 ( .A(n39660), .Z(n39661) );
  XNOR U42220 ( .A(m[260]), .B(n39662), .Z(n39660) );
  NAND U42221 ( .A(n39663), .B(mul_pow), .Z(n39662) );
  XOR U42222 ( .A(m[260]), .B(c[260]), .Z(n39663) );
  XOR U42223 ( .A(n39664), .B(n39665), .Z(n39656) );
  ANDN U42224 ( .B(n39666), .A(n31264), .Z(n39664) );
  XNOR U42225 ( .A(\modmult_1/zin[0][258] ), .B(n39667), .Z(n31264) );
  IV U42226 ( .A(n39665), .Z(n39667) );
  XOR U42227 ( .A(n39665), .B(n31265), .Z(n39666) );
  XNOR U42228 ( .A(n39668), .B(n39669), .Z(n31265) );
  ANDN U42229 ( .B(\modmult_1/xin[1023] ), .A(n39670), .Z(n39668) );
  IV U42230 ( .A(n39669), .Z(n39670) );
  XNOR U42231 ( .A(m[259]), .B(n39671), .Z(n39669) );
  NAND U42232 ( .A(n39672), .B(mul_pow), .Z(n39671) );
  XOR U42233 ( .A(m[259]), .B(c[259]), .Z(n39672) );
  XOR U42234 ( .A(n39673), .B(n39674), .Z(n39665) );
  ANDN U42235 ( .B(n39675), .A(n31262), .Z(n39673) );
  XNOR U42236 ( .A(\modmult_1/zin[0][257] ), .B(n39676), .Z(n31262) );
  IV U42237 ( .A(n39674), .Z(n39676) );
  XOR U42238 ( .A(n39674), .B(n31263), .Z(n39675) );
  XNOR U42239 ( .A(n39677), .B(n39678), .Z(n31263) );
  ANDN U42240 ( .B(\modmult_1/xin[1023] ), .A(n39679), .Z(n39677) );
  IV U42241 ( .A(n39678), .Z(n39679) );
  XNOR U42242 ( .A(m[258]), .B(n39680), .Z(n39678) );
  NAND U42243 ( .A(n39681), .B(mul_pow), .Z(n39680) );
  XOR U42244 ( .A(m[258]), .B(c[258]), .Z(n39681) );
  XOR U42245 ( .A(n39682), .B(n39683), .Z(n39674) );
  ANDN U42246 ( .B(n39684), .A(n31260), .Z(n39682) );
  XNOR U42247 ( .A(\modmult_1/zin[0][256] ), .B(n39685), .Z(n31260) );
  IV U42248 ( .A(n39683), .Z(n39685) );
  XOR U42249 ( .A(n39683), .B(n31261), .Z(n39684) );
  XNOR U42250 ( .A(n39686), .B(n39687), .Z(n31261) );
  ANDN U42251 ( .B(\modmult_1/xin[1023] ), .A(n39688), .Z(n39686) );
  IV U42252 ( .A(n39687), .Z(n39688) );
  XNOR U42253 ( .A(m[257]), .B(n39689), .Z(n39687) );
  NAND U42254 ( .A(n39690), .B(mul_pow), .Z(n39689) );
  XOR U42255 ( .A(m[257]), .B(c[257]), .Z(n39690) );
  XOR U42256 ( .A(n39691), .B(n39692), .Z(n39683) );
  ANDN U42257 ( .B(n39693), .A(n31258), .Z(n39691) );
  XNOR U42258 ( .A(\modmult_1/zin[0][255] ), .B(n39694), .Z(n31258) );
  IV U42259 ( .A(n39692), .Z(n39694) );
  XOR U42260 ( .A(n39692), .B(n31259), .Z(n39693) );
  XNOR U42261 ( .A(n39695), .B(n39696), .Z(n31259) );
  ANDN U42262 ( .B(\modmult_1/xin[1023] ), .A(n39697), .Z(n39695) );
  IV U42263 ( .A(n39696), .Z(n39697) );
  XNOR U42264 ( .A(m[256]), .B(n39698), .Z(n39696) );
  NAND U42265 ( .A(n39699), .B(mul_pow), .Z(n39698) );
  XOR U42266 ( .A(m[256]), .B(c[256]), .Z(n39699) );
  XOR U42267 ( .A(n39700), .B(n39701), .Z(n39692) );
  ANDN U42268 ( .B(n39702), .A(n31256), .Z(n39700) );
  XNOR U42269 ( .A(\modmult_1/zin[0][254] ), .B(n39703), .Z(n31256) );
  IV U42270 ( .A(n39701), .Z(n39703) );
  XOR U42271 ( .A(n39701), .B(n31257), .Z(n39702) );
  XNOR U42272 ( .A(n39704), .B(n39705), .Z(n31257) );
  ANDN U42273 ( .B(\modmult_1/xin[1023] ), .A(n39706), .Z(n39704) );
  IV U42274 ( .A(n39705), .Z(n39706) );
  XNOR U42275 ( .A(m[255]), .B(n39707), .Z(n39705) );
  NAND U42276 ( .A(n39708), .B(mul_pow), .Z(n39707) );
  XOR U42277 ( .A(m[255]), .B(c[255]), .Z(n39708) );
  XOR U42278 ( .A(n39709), .B(n39710), .Z(n39701) );
  ANDN U42279 ( .B(n39711), .A(n31254), .Z(n39709) );
  XNOR U42280 ( .A(\modmult_1/zin[0][253] ), .B(n39712), .Z(n31254) );
  IV U42281 ( .A(n39710), .Z(n39712) );
  XOR U42282 ( .A(n39710), .B(n31255), .Z(n39711) );
  XNOR U42283 ( .A(n39713), .B(n39714), .Z(n31255) );
  ANDN U42284 ( .B(\modmult_1/xin[1023] ), .A(n39715), .Z(n39713) );
  IV U42285 ( .A(n39714), .Z(n39715) );
  XNOR U42286 ( .A(m[254]), .B(n39716), .Z(n39714) );
  NAND U42287 ( .A(n39717), .B(mul_pow), .Z(n39716) );
  XOR U42288 ( .A(m[254]), .B(c[254]), .Z(n39717) );
  XOR U42289 ( .A(n39718), .B(n39719), .Z(n39710) );
  ANDN U42290 ( .B(n39720), .A(n31252), .Z(n39718) );
  XNOR U42291 ( .A(\modmult_1/zin[0][252] ), .B(n39721), .Z(n31252) );
  IV U42292 ( .A(n39719), .Z(n39721) );
  XOR U42293 ( .A(n39719), .B(n31253), .Z(n39720) );
  XNOR U42294 ( .A(n39722), .B(n39723), .Z(n31253) );
  ANDN U42295 ( .B(\modmult_1/xin[1023] ), .A(n39724), .Z(n39722) );
  IV U42296 ( .A(n39723), .Z(n39724) );
  XNOR U42297 ( .A(m[253]), .B(n39725), .Z(n39723) );
  NAND U42298 ( .A(n39726), .B(mul_pow), .Z(n39725) );
  XOR U42299 ( .A(m[253]), .B(c[253]), .Z(n39726) );
  XOR U42300 ( .A(n39727), .B(n39728), .Z(n39719) );
  ANDN U42301 ( .B(n39729), .A(n31250), .Z(n39727) );
  XNOR U42302 ( .A(\modmult_1/zin[0][251] ), .B(n39730), .Z(n31250) );
  IV U42303 ( .A(n39728), .Z(n39730) );
  XOR U42304 ( .A(n39728), .B(n31251), .Z(n39729) );
  XNOR U42305 ( .A(n39731), .B(n39732), .Z(n31251) );
  ANDN U42306 ( .B(\modmult_1/xin[1023] ), .A(n39733), .Z(n39731) );
  IV U42307 ( .A(n39732), .Z(n39733) );
  XNOR U42308 ( .A(m[252]), .B(n39734), .Z(n39732) );
  NAND U42309 ( .A(n39735), .B(mul_pow), .Z(n39734) );
  XOR U42310 ( .A(m[252]), .B(c[252]), .Z(n39735) );
  XOR U42311 ( .A(n39736), .B(n39737), .Z(n39728) );
  ANDN U42312 ( .B(n39738), .A(n31248), .Z(n39736) );
  XNOR U42313 ( .A(\modmult_1/zin[0][250] ), .B(n39739), .Z(n31248) );
  IV U42314 ( .A(n39737), .Z(n39739) );
  XOR U42315 ( .A(n39737), .B(n31249), .Z(n39738) );
  XNOR U42316 ( .A(n39740), .B(n39741), .Z(n31249) );
  ANDN U42317 ( .B(\modmult_1/xin[1023] ), .A(n39742), .Z(n39740) );
  IV U42318 ( .A(n39741), .Z(n39742) );
  XNOR U42319 ( .A(m[251]), .B(n39743), .Z(n39741) );
  NAND U42320 ( .A(n39744), .B(mul_pow), .Z(n39743) );
  XOR U42321 ( .A(m[251]), .B(c[251]), .Z(n39744) );
  XOR U42322 ( .A(n39745), .B(n39746), .Z(n39737) );
  ANDN U42323 ( .B(n39747), .A(n31246), .Z(n39745) );
  XNOR U42324 ( .A(\modmult_1/zin[0][249] ), .B(n39748), .Z(n31246) );
  IV U42325 ( .A(n39746), .Z(n39748) );
  XOR U42326 ( .A(n39746), .B(n31247), .Z(n39747) );
  XNOR U42327 ( .A(n39749), .B(n39750), .Z(n31247) );
  ANDN U42328 ( .B(\modmult_1/xin[1023] ), .A(n39751), .Z(n39749) );
  IV U42329 ( .A(n39750), .Z(n39751) );
  XNOR U42330 ( .A(m[250]), .B(n39752), .Z(n39750) );
  NAND U42331 ( .A(n39753), .B(mul_pow), .Z(n39752) );
  XOR U42332 ( .A(m[250]), .B(c[250]), .Z(n39753) );
  XOR U42333 ( .A(n39754), .B(n39755), .Z(n39746) );
  ANDN U42334 ( .B(n39756), .A(n31244), .Z(n39754) );
  XNOR U42335 ( .A(\modmult_1/zin[0][248] ), .B(n39757), .Z(n31244) );
  IV U42336 ( .A(n39755), .Z(n39757) );
  XOR U42337 ( .A(n39755), .B(n31245), .Z(n39756) );
  XNOR U42338 ( .A(n39758), .B(n39759), .Z(n31245) );
  ANDN U42339 ( .B(\modmult_1/xin[1023] ), .A(n39760), .Z(n39758) );
  IV U42340 ( .A(n39759), .Z(n39760) );
  XNOR U42341 ( .A(m[249]), .B(n39761), .Z(n39759) );
  NAND U42342 ( .A(n39762), .B(mul_pow), .Z(n39761) );
  XOR U42343 ( .A(m[249]), .B(c[249]), .Z(n39762) );
  XOR U42344 ( .A(n39763), .B(n39764), .Z(n39755) );
  ANDN U42345 ( .B(n39765), .A(n31242), .Z(n39763) );
  XNOR U42346 ( .A(\modmult_1/zin[0][247] ), .B(n39766), .Z(n31242) );
  IV U42347 ( .A(n39764), .Z(n39766) );
  XOR U42348 ( .A(n39764), .B(n31243), .Z(n39765) );
  XNOR U42349 ( .A(n39767), .B(n39768), .Z(n31243) );
  ANDN U42350 ( .B(\modmult_1/xin[1023] ), .A(n39769), .Z(n39767) );
  IV U42351 ( .A(n39768), .Z(n39769) );
  XNOR U42352 ( .A(m[248]), .B(n39770), .Z(n39768) );
  NAND U42353 ( .A(n39771), .B(mul_pow), .Z(n39770) );
  XOR U42354 ( .A(m[248]), .B(c[248]), .Z(n39771) );
  XOR U42355 ( .A(n39772), .B(n39773), .Z(n39764) );
  ANDN U42356 ( .B(n39774), .A(n31240), .Z(n39772) );
  XNOR U42357 ( .A(\modmult_1/zin[0][246] ), .B(n39775), .Z(n31240) );
  IV U42358 ( .A(n39773), .Z(n39775) );
  XOR U42359 ( .A(n39773), .B(n31241), .Z(n39774) );
  XNOR U42360 ( .A(n39776), .B(n39777), .Z(n31241) );
  ANDN U42361 ( .B(\modmult_1/xin[1023] ), .A(n39778), .Z(n39776) );
  IV U42362 ( .A(n39777), .Z(n39778) );
  XNOR U42363 ( .A(m[247]), .B(n39779), .Z(n39777) );
  NAND U42364 ( .A(n39780), .B(mul_pow), .Z(n39779) );
  XOR U42365 ( .A(m[247]), .B(c[247]), .Z(n39780) );
  XOR U42366 ( .A(n39781), .B(n39782), .Z(n39773) );
  ANDN U42367 ( .B(n39783), .A(n31238), .Z(n39781) );
  XNOR U42368 ( .A(\modmult_1/zin[0][245] ), .B(n39784), .Z(n31238) );
  IV U42369 ( .A(n39782), .Z(n39784) );
  XOR U42370 ( .A(n39782), .B(n31239), .Z(n39783) );
  XNOR U42371 ( .A(n39785), .B(n39786), .Z(n31239) );
  ANDN U42372 ( .B(\modmult_1/xin[1023] ), .A(n39787), .Z(n39785) );
  IV U42373 ( .A(n39786), .Z(n39787) );
  XNOR U42374 ( .A(m[246]), .B(n39788), .Z(n39786) );
  NAND U42375 ( .A(n39789), .B(mul_pow), .Z(n39788) );
  XOR U42376 ( .A(m[246]), .B(c[246]), .Z(n39789) );
  XOR U42377 ( .A(n39790), .B(n39791), .Z(n39782) );
  ANDN U42378 ( .B(n39792), .A(n31236), .Z(n39790) );
  XNOR U42379 ( .A(\modmult_1/zin[0][244] ), .B(n39793), .Z(n31236) );
  IV U42380 ( .A(n39791), .Z(n39793) );
  XOR U42381 ( .A(n39791), .B(n31237), .Z(n39792) );
  XNOR U42382 ( .A(n39794), .B(n39795), .Z(n31237) );
  ANDN U42383 ( .B(\modmult_1/xin[1023] ), .A(n39796), .Z(n39794) );
  IV U42384 ( .A(n39795), .Z(n39796) );
  XNOR U42385 ( .A(m[245]), .B(n39797), .Z(n39795) );
  NAND U42386 ( .A(n39798), .B(mul_pow), .Z(n39797) );
  XOR U42387 ( .A(m[245]), .B(c[245]), .Z(n39798) );
  XOR U42388 ( .A(n39799), .B(n39800), .Z(n39791) );
  ANDN U42389 ( .B(n39801), .A(n31234), .Z(n39799) );
  XNOR U42390 ( .A(\modmult_1/zin[0][243] ), .B(n39802), .Z(n31234) );
  IV U42391 ( .A(n39800), .Z(n39802) );
  XOR U42392 ( .A(n39800), .B(n31235), .Z(n39801) );
  XNOR U42393 ( .A(n39803), .B(n39804), .Z(n31235) );
  ANDN U42394 ( .B(\modmult_1/xin[1023] ), .A(n39805), .Z(n39803) );
  IV U42395 ( .A(n39804), .Z(n39805) );
  XNOR U42396 ( .A(m[244]), .B(n39806), .Z(n39804) );
  NAND U42397 ( .A(n39807), .B(mul_pow), .Z(n39806) );
  XOR U42398 ( .A(m[244]), .B(c[244]), .Z(n39807) );
  XOR U42399 ( .A(n39808), .B(n39809), .Z(n39800) );
  ANDN U42400 ( .B(n39810), .A(n31232), .Z(n39808) );
  XNOR U42401 ( .A(\modmult_1/zin[0][242] ), .B(n39811), .Z(n31232) );
  IV U42402 ( .A(n39809), .Z(n39811) );
  XOR U42403 ( .A(n39809), .B(n31233), .Z(n39810) );
  XNOR U42404 ( .A(n39812), .B(n39813), .Z(n31233) );
  ANDN U42405 ( .B(\modmult_1/xin[1023] ), .A(n39814), .Z(n39812) );
  IV U42406 ( .A(n39813), .Z(n39814) );
  XNOR U42407 ( .A(m[243]), .B(n39815), .Z(n39813) );
  NAND U42408 ( .A(n39816), .B(mul_pow), .Z(n39815) );
  XOR U42409 ( .A(m[243]), .B(c[243]), .Z(n39816) );
  XOR U42410 ( .A(n39817), .B(n39818), .Z(n39809) );
  ANDN U42411 ( .B(n39819), .A(n31230), .Z(n39817) );
  XNOR U42412 ( .A(\modmult_1/zin[0][241] ), .B(n39820), .Z(n31230) );
  IV U42413 ( .A(n39818), .Z(n39820) );
  XOR U42414 ( .A(n39818), .B(n31231), .Z(n39819) );
  XNOR U42415 ( .A(n39821), .B(n39822), .Z(n31231) );
  ANDN U42416 ( .B(\modmult_1/xin[1023] ), .A(n39823), .Z(n39821) );
  IV U42417 ( .A(n39822), .Z(n39823) );
  XNOR U42418 ( .A(m[242]), .B(n39824), .Z(n39822) );
  NAND U42419 ( .A(n39825), .B(mul_pow), .Z(n39824) );
  XOR U42420 ( .A(m[242]), .B(c[242]), .Z(n39825) );
  XOR U42421 ( .A(n39826), .B(n39827), .Z(n39818) );
  ANDN U42422 ( .B(n39828), .A(n31228), .Z(n39826) );
  XNOR U42423 ( .A(\modmult_1/zin[0][240] ), .B(n39829), .Z(n31228) );
  IV U42424 ( .A(n39827), .Z(n39829) );
  XOR U42425 ( .A(n39827), .B(n31229), .Z(n39828) );
  XNOR U42426 ( .A(n39830), .B(n39831), .Z(n31229) );
  ANDN U42427 ( .B(\modmult_1/xin[1023] ), .A(n39832), .Z(n39830) );
  IV U42428 ( .A(n39831), .Z(n39832) );
  XNOR U42429 ( .A(m[241]), .B(n39833), .Z(n39831) );
  NAND U42430 ( .A(n39834), .B(mul_pow), .Z(n39833) );
  XOR U42431 ( .A(m[241]), .B(c[241]), .Z(n39834) );
  XOR U42432 ( .A(n39835), .B(n39836), .Z(n39827) );
  ANDN U42433 ( .B(n39837), .A(n31226), .Z(n39835) );
  XNOR U42434 ( .A(\modmult_1/zin[0][239] ), .B(n39838), .Z(n31226) );
  IV U42435 ( .A(n39836), .Z(n39838) );
  XOR U42436 ( .A(n39836), .B(n31227), .Z(n39837) );
  XNOR U42437 ( .A(n39839), .B(n39840), .Z(n31227) );
  ANDN U42438 ( .B(\modmult_1/xin[1023] ), .A(n39841), .Z(n39839) );
  IV U42439 ( .A(n39840), .Z(n39841) );
  XNOR U42440 ( .A(m[240]), .B(n39842), .Z(n39840) );
  NAND U42441 ( .A(n39843), .B(mul_pow), .Z(n39842) );
  XOR U42442 ( .A(m[240]), .B(c[240]), .Z(n39843) );
  XOR U42443 ( .A(n39844), .B(n39845), .Z(n39836) );
  ANDN U42444 ( .B(n39846), .A(n31224), .Z(n39844) );
  XNOR U42445 ( .A(\modmult_1/zin[0][238] ), .B(n39847), .Z(n31224) );
  IV U42446 ( .A(n39845), .Z(n39847) );
  XOR U42447 ( .A(n39845), .B(n31225), .Z(n39846) );
  XNOR U42448 ( .A(n39848), .B(n39849), .Z(n31225) );
  ANDN U42449 ( .B(\modmult_1/xin[1023] ), .A(n39850), .Z(n39848) );
  IV U42450 ( .A(n39849), .Z(n39850) );
  XNOR U42451 ( .A(m[239]), .B(n39851), .Z(n39849) );
  NAND U42452 ( .A(n39852), .B(mul_pow), .Z(n39851) );
  XOR U42453 ( .A(m[239]), .B(c[239]), .Z(n39852) );
  XOR U42454 ( .A(n39853), .B(n39854), .Z(n39845) );
  ANDN U42455 ( .B(n39855), .A(n31222), .Z(n39853) );
  XNOR U42456 ( .A(\modmult_1/zin[0][237] ), .B(n39856), .Z(n31222) );
  IV U42457 ( .A(n39854), .Z(n39856) );
  XOR U42458 ( .A(n39854), .B(n31223), .Z(n39855) );
  XNOR U42459 ( .A(n39857), .B(n39858), .Z(n31223) );
  ANDN U42460 ( .B(\modmult_1/xin[1023] ), .A(n39859), .Z(n39857) );
  IV U42461 ( .A(n39858), .Z(n39859) );
  XNOR U42462 ( .A(m[238]), .B(n39860), .Z(n39858) );
  NAND U42463 ( .A(n39861), .B(mul_pow), .Z(n39860) );
  XOR U42464 ( .A(m[238]), .B(c[238]), .Z(n39861) );
  XOR U42465 ( .A(n39862), .B(n39863), .Z(n39854) );
  ANDN U42466 ( .B(n39864), .A(n31220), .Z(n39862) );
  XNOR U42467 ( .A(\modmult_1/zin[0][236] ), .B(n39865), .Z(n31220) );
  IV U42468 ( .A(n39863), .Z(n39865) );
  XOR U42469 ( .A(n39863), .B(n31221), .Z(n39864) );
  XNOR U42470 ( .A(n39866), .B(n39867), .Z(n31221) );
  ANDN U42471 ( .B(\modmult_1/xin[1023] ), .A(n39868), .Z(n39866) );
  IV U42472 ( .A(n39867), .Z(n39868) );
  XNOR U42473 ( .A(m[237]), .B(n39869), .Z(n39867) );
  NAND U42474 ( .A(n39870), .B(mul_pow), .Z(n39869) );
  XOR U42475 ( .A(m[237]), .B(c[237]), .Z(n39870) );
  XOR U42476 ( .A(n39871), .B(n39872), .Z(n39863) );
  ANDN U42477 ( .B(n39873), .A(n31218), .Z(n39871) );
  XNOR U42478 ( .A(\modmult_1/zin[0][235] ), .B(n39874), .Z(n31218) );
  IV U42479 ( .A(n39872), .Z(n39874) );
  XOR U42480 ( .A(n39872), .B(n31219), .Z(n39873) );
  XNOR U42481 ( .A(n39875), .B(n39876), .Z(n31219) );
  ANDN U42482 ( .B(\modmult_1/xin[1023] ), .A(n39877), .Z(n39875) );
  IV U42483 ( .A(n39876), .Z(n39877) );
  XNOR U42484 ( .A(m[236]), .B(n39878), .Z(n39876) );
  NAND U42485 ( .A(n39879), .B(mul_pow), .Z(n39878) );
  XOR U42486 ( .A(m[236]), .B(c[236]), .Z(n39879) );
  XOR U42487 ( .A(n39880), .B(n39881), .Z(n39872) );
  ANDN U42488 ( .B(n39882), .A(n31216), .Z(n39880) );
  XNOR U42489 ( .A(\modmult_1/zin[0][234] ), .B(n39883), .Z(n31216) );
  IV U42490 ( .A(n39881), .Z(n39883) );
  XOR U42491 ( .A(n39881), .B(n31217), .Z(n39882) );
  XNOR U42492 ( .A(n39884), .B(n39885), .Z(n31217) );
  ANDN U42493 ( .B(\modmult_1/xin[1023] ), .A(n39886), .Z(n39884) );
  IV U42494 ( .A(n39885), .Z(n39886) );
  XNOR U42495 ( .A(m[235]), .B(n39887), .Z(n39885) );
  NAND U42496 ( .A(n39888), .B(mul_pow), .Z(n39887) );
  XOR U42497 ( .A(m[235]), .B(c[235]), .Z(n39888) );
  XOR U42498 ( .A(n39889), .B(n39890), .Z(n39881) );
  ANDN U42499 ( .B(n39891), .A(n31214), .Z(n39889) );
  XNOR U42500 ( .A(\modmult_1/zin[0][233] ), .B(n39892), .Z(n31214) );
  IV U42501 ( .A(n39890), .Z(n39892) );
  XOR U42502 ( .A(n39890), .B(n31215), .Z(n39891) );
  XNOR U42503 ( .A(n39893), .B(n39894), .Z(n31215) );
  ANDN U42504 ( .B(\modmult_1/xin[1023] ), .A(n39895), .Z(n39893) );
  IV U42505 ( .A(n39894), .Z(n39895) );
  XNOR U42506 ( .A(m[234]), .B(n39896), .Z(n39894) );
  NAND U42507 ( .A(n39897), .B(mul_pow), .Z(n39896) );
  XOR U42508 ( .A(m[234]), .B(c[234]), .Z(n39897) );
  XOR U42509 ( .A(n39898), .B(n39899), .Z(n39890) );
  ANDN U42510 ( .B(n39900), .A(n31212), .Z(n39898) );
  XNOR U42511 ( .A(\modmult_1/zin[0][232] ), .B(n39901), .Z(n31212) );
  IV U42512 ( .A(n39899), .Z(n39901) );
  XOR U42513 ( .A(n39899), .B(n31213), .Z(n39900) );
  XNOR U42514 ( .A(n39902), .B(n39903), .Z(n31213) );
  ANDN U42515 ( .B(\modmult_1/xin[1023] ), .A(n39904), .Z(n39902) );
  IV U42516 ( .A(n39903), .Z(n39904) );
  XNOR U42517 ( .A(m[233]), .B(n39905), .Z(n39903) );
  NAND U42518 ( .A(n39906), .B(mul_pow), .Z(n39905) );
  XOR U42519 ( .A(m[233]), .B(c[233]), .Z(n39906) );
  XOR U42520 ( .A(n39907), .B(n39908), .Z(n39899) );
  ANDN U42521 ( .B(n39909), .A(n31210), .Z(n39907) );
  XNOR U42522 ( .A(\modmult_1/zin[0][231] ), .B(n39910), .Z(n31210) );
  IV U42523 ( .A(n39908), .Z(n39910) );
  XOR U42524 ( .A(n39908), .B(n31211), .Z(n39909) );
  XNOR U42525 ( .A(n39911), .B(n39912), .Z(n31211) );
  ANDN U42526 ( .B(\modmult_1/xin[1023] ), .A(n39913), .Z(n39911) );
  IV U42527 ( .A(n39912), .Z(n39913) );
  XNOR U42528 ( .A(m[232]), .B(n39914), .Z(n39912) );
  NAND U42529 ( .A(n39915), .B(mul_pow), .Z(n39914) );
  XOR U42530 ( .A(m[232]), .B(c[232]), .Z(n39915) );
  XOR U42531 ( .A(n39916), .B(n39917), .Z(n39908) );
  ANDN U42532 ( .B(n39918), .A(n31208), .Z(n39916) );
  XNOR U42533 ( .A(\modmult_1/zin[0][230] ), .B(n39919), .Z(n31208) );
  IV U42534 ( .A(n39917), .Z(n39919) );
  XOR U42535 ( .A(n39917), .B(n31209), .Z(n39918) );
  XNOR U42536 ( .A(n39920), .B(n39921), .Z(n31209) );
  ANDN U42537 ( .B(\modmult_1/xin[1023] ), .A(n39922), .Z(n39920) );
  IV U42538 ( .A(n39921), .Z(n39922) );
  XNOR U42539 ( .A(m[231]), .B(n39923), .Z(n39921) );
  NAND U42540 ( .A(n39924), .B(mul_pow), .Z(n39923) );
  XOR U42541 ( .A(m[231]), .B(c[231]), .Z(n39924) );
  XOR U42542 ( .A(n39925), .B(n39926), .Z(n39917) );
  ANDN U42543 ( .B(n39927), .A(n31206), .Z(n39925) );
  XNOR U42544 ( .A(\modmult_1/zin[0][229] ), .B(n39928), .Z(n31206) );
  IV U42545 ( .A(n39926), .Z(n39928) );
  XOR U42546 ( .A(n39926), .B(n31207), .Z(n39927) );
  XNOR U42547 ( .A(n39929), .B(n39930), .Z(n31207) );
  ANDN U42548 ( .B(\modmult_1/xin[1023] ), .A(n39931), .Z(n39929) );
  IV U42549 ( .A(n39930), .Z(n39931) );
  XNOR U42550 ( .A(m[230]), .B(n39932), .Z(n39930) );
  NAND U42551 ( .A(n39933), .B(mul_pow), .Z(n39932) );
  XOR U42552 ( .A(m[230]), .B(c[230]), .Z(n39933) );
  XOR U42553 ( .A(n39934), .B(n39935), .Z(n39926) );
  ANDN U42554 ( .B(n39936), .A(n31204), .Z(n39934) );
  XNOR U42555 ( .A(\modmult_1/zin[0][228] ), .B(n39937), .Z(n31204) );
  IV U42556 ( .A(n39935), .Z(n39937) );
  XOR U42557 ( .A(n39935), .B(n31205), .Z(n39936) );
  XNOR U42558 ( .A(n39938), .B(n39939), .Z(n31205) );
  ANDN U42559 ( .B(\modmult_1/xin[1023] ), .A(n39940), .Z(n39938) );
  IV U42560 ( .A(n39939), .Z(n39940) );
  XNOR U42561 ( .A(m[229]), .B(n39941), .Z(n39939) );
  NAND U42562 ( .A(n39942), .B(mul_pow), .Z(n39941) );
  XOR U42563 ( .A(m[229]), .B(c[229]), .Z(n39942) );
  XOR U42564 ( .A(n39943), .B(n39944), .Z(n39935) );
  ANDN U42565 ( .B(n39945), .A(n31202), .Z(n39943) );
  XNOR U42566 ( .A(\modmult_1/zin[0][227] ), .B(n39946), .Z(n31202) );
  IV U42567 ( .A(n39944), .Z(n39946) );
  XOR U42568 ( .A(n39944), .B(n31203), .Z(n39945) );
  XNOR U42569 ( .A(n39947), .B(n39948), .Z(n31203) );
  ANDN U42570 ( .B(\modmult_1/xin[1023] ), .A(n39949), .Z(n39947) );
  IV U42571 ( .A(n39948), .Z(n39949) );
  XNOR U42572 ( .A(m[228]), .B(n39950), .Z(n39948) );
  NAND U42573 ( .A(n39951), .B(mul_pow), .Z(n39950) );
  XOR U42574 ( .A(m[228]), .B(c[228]), .Z(n39951) );
  XOR U42575 ( .A(n39952), .B(n39953), .Z(n39944) );
  ANDN U42576 ( .B(n39954), .A(n31200), .Z(n39952) );
  XNOR U42577 ( .A(\modmult_1/zin[0][226] ), .B(n39955), .Z(n31200) );
  IV U42578 ( .A(n39953), .Z(n39955) );
  XOR U42579 ( .A(n39953), .B(n31201), .Z(n39954) );
  XNOR U42580 ( .A(n39956), .B(n39957), .Z(n31201) );
  ANDN U42581 ( .B(\modmult_1/xin[1023] ), .A(n39958), .Z(n39956) );
  IV U42582 ( .A(n39957), .Z(n39958) );
  XNOR U42583 ( .A(m[227]), .B(n39959), .Z(n39957) );
  NAND U42584 ( .A(n39960), .B(mul_pow), .Z(n39959) );
  XOR U42585 ( .A(m[227]), .B(c[227]), .Z(n39960) );
  XOR U42586 ( .A(n39961), .B(n39962), .Z(n39953) );
  ANDN U42587 ( .B(n39963), .A(n31198), .Z(n39961) );
  XNOR U42588 ( .A(\modmult_1/zin[0][225] ), .B(n39964), .Z(n31198) );
  IV U42589 ( .A(n39962), .Z(n39964) );
  XOR U42590 ( .A(n39962), .B(n31199), .Z(n39963) );
  XNOR U42591 ( .A(n39965), .B(n39966), .Z(n31199) );
  ANDN U42592 ( .B(\modmult_1/xin[1023] ), .A(n39967), .Z(n39965) );
  IV U42593 ( .A(n39966), .Z(n39967) );
  XNOR U42594 ( .A(m[226]), .B(n39968), .Z(n39966) );
  NAND U42595 ( .A(n39969), .B(mul_pow), .Z(n39968) );
  XOR U42596 ( .A(m[226]), .B(c[226]), .Z(n39969) );
  XOR U42597 ( .A(n39970), .B(n39971), .Z(n39962) );
  ANDN U42598 ( .B(n39972), .A(n31196), .Z(n39970) );
  XNOR U42599 ( .A(\modmult_1/zin[0][224] ), .B(n39973), .Z(n31196) );
  IV U42600 ( .A(n39971), .Z(n39973) );
  XOR U42601 ( .A(n39971), .B(n31197), .Z(n39972) );
  XNOR U42602 ( .A(n39974), .B(n39975), .Z(n31197) );
  ANDN U42603 ( .B(\modmult_1/xin[1023] ), .A(n39976), .Z(n39974) );
  IV U42604 ( .A(n39975), .Z(n39976) );
  XNOR U42605 ( .A(m[225]), .B(n39977), .Z(n39975) );
  NAND U42606 ( .A(n39978), .B(mul_pow), .Z(n39977) );
  XOR U42607 ( .A(m[225]), .B(c[225]), .Z(n39978) );
  XOR U42608 ( .A(n39979), .B(n39980), .Z(n39971) );
  ANDN U42609 ( .B(n39981), .A(n31194), .Z(n39979) );
  XNOR U42610 ( .A(\modmult_1/zin[0][223] ), .B(n39982), .Z(n31194) );
  IV U42611 ( .A(n39980), .Z(n39982) );
  XOR U42612 ( .A(n39980), .B(n31195), .Z(n39981) );
  XNOR U42613 ( .A(n39983), .B(n39984), .Z(n31195) );
  ANDN U42614 ( .B(\modmult_1/xin[1023] ), .A(n39985), .Z(n39983) );
  IV U42615 ( .A(n39984), .Z(n39985) );
  XNOR U42616 ( .A(m[224]), .B(n39986), .Z(n39984) );
  NAND U42617 ( .A(n39987), .B(mul_pow), .Z(n39986) );
  XOR U42618 ( .A(m[224]), .B(c[224]), .Z(n39987) );
  XOR U42619 ( .A(n39988), .B(n39989), .Z(n39980) );
  ANDN U42620 ( .B(n39990), .A(n31192), .Z(n39988) );
  XNOR U42621 ( .A(\modmult_1/zin[0][222] ), .B(n39991), .Z(n31192) );
  IV U42622 ( .A(n39989), .Z(n39991) );
  XOR U42623 ( .A(n39989), .B(n31193), .Z(n39990) );
  XNOR U42624 ( .A(n39992), .B(n39993), .Z(n31193) );
  ANDN U42625 ( .B(\modmult_1/xin[1023] ), .A(n39994), .Z(n39992) );
  IV U42626 ( .A(n39993), .Z(n39994) );
  XNOR U42627 ( .A(m[223]), .B(n39995), .Z(n39993) );
  NAND U42628 ( .A(n39996), .B(mul_pow), .Z(n39995) );
  XOR U42629 ( .A(m[223]), .B(c[223]), .Z(n39996) );
  XOR U42630 ( .A(n39997), .B(n39998), .Z(n39989) );
  ANDN U42631 ( .B(n39999), .A(n31190), .Z(n39997) );
  XNOR U42632 ( .A(\modmult_1/zin[0][221] ), .B(n40000), .Z(n31190) );
  IV U42633 ( .A(n39998), .Z(n40000) );
  XOR U42634 ( .A(n39998), .B(n31191), .Z(n39999) );
  XNOR U42635 ( .A(n40001), .B(n40002), .Z(n31191) );
  ANDN U42636 ( .B(\modmult_1/xin[1023] ), .A(n40003), .Z(n40001) );
  IV U42637 ( .A(n40002), .Z(n40003) );
  XNOR U42638 ( .A(m[222]), .B(n40004), .Z(n40002) );
  NAND U42639 ( .A(n40005), .B(mul_pow), .Z(n40004) );
  XOR U42640 ( .A(m[222]), .B(c[222]), .Z(n40005) );
  XOR U42641 ( .A(n40006), .B(n40007), .Z(n39998) );
  ANDN U42642 ( .B(n40008), .A(n31188), .Z(n40006) );
  XNOR U42643 ( .A(\modmult_1/zin[0][220] ), .B(n40009), .Z(n31188) );
  IV U42644 ( .A(n40007), .Z(n40009) );
  XOR U42645 ( .A(n40007), .B(n31189), .Z(n40008) );
  XNOR U42646 ( .A(n40010), .B(n40011), .Z(n31189) );
  ANDN U42647 ( .B(\modmult_1/xin[1023] ), .A(n40012), .Z(n40010) );
  IV U42648 ( .A(n40011), .Z(n40012) );
  XNOR U42649 ( .A(m[221]), .B(n40013), .Z(n40011) );
  NAND U42650 ( .A(n40014), .B(mul_pow), .Z(n40013) );
  XOR U42651 ( .A(m[221]), .B(c[221]), .Z(n40014) );
  XOR U42652 ( .A(n40015), .B(n40016), .Z(n40007) );
  ANDN U42653 ( .B(n40017), .A(n31186), .Z(n40015) );
  XNOR U42654 ( .A(\modmult_1/zin[0][219] ), .B(n40018), .Z(n31186) );
  IV U42655 ( .A(n40016), .Z(n40018) );
  XOR U42656 ( .A(n40016), .B(n31187), .Z(n40017) );
  XNOR U42657 ( .A(n40019), .B(n40020), .Z(n31187) );
  ANDN U42658 ( .B(\modmult_1/xin[1023] ), .A(n40021), .Z(n40019) );
  IV U42659 ( .A(n40020), .Z(n40021) );
  XNOR U42660 ( .A(m[220]), .B(n40022), .Z(n40020) );
  NAND U42661 ( .A(n40023), .B(mul_pow), .Z(n40022) );
  XOR U42662 ( .A(m[220]), .B(c[220]), .Z(n40023) );
  XOR U42663 ( .A(n40024), .B(n40025), .Z(n40016) );
  ANDN U42664 ( .B(n40026), .A(n31184), .Z(n40024) );
  XNOR U42665 ( .A(\modmult_1/zin[0][218] ), .B(n40027), .Z(n31184) );
  IV U42666 ( .A(n40025), .Z(n40027) );
  XOR U42667 ( .A(n40025), .B(n31185), .Z(n40026) );
  XNOR U42668 ( .A(n40028), .B(n40029), .Z(n31185) );
  ANDN U42669 ( .B(\modmult_1/xin[1023] ), .A(n40030), .Z(n40028) );
  IV U42670 ( .A(n40029), .Z(n40030) );
  XNOR U42671 ( .A(m[219]), .B(n40031), .Z(n40029) );
  NAND U42672 ( .A(n40032), .B(mul_pow), .Z(n40031) );
  XOR U42673 ( .A(m[219]), .B(c[219]), .Z(n40032) );
  XOR U42674 ( .A(n40033), .B(n40034), .Z(n40025) );
  ANDN U42675 ( .B(n40035), .A(n31182), .Z(n40033) );
  XNOR U42676 ( .A(\modmult_1/zin[0][217] ), .B(n40036), .Z(n31182) );
  IV U42677 ( .A(n40034), .Z(n40036) );
  XOR U42678 ( .A(n40034), .B(n31183), .Z(n40035) );
  XNOR U42679 ( .A(n40037), .B(n40038), .Z(n31183) );
  ANDN U42680 ( .B(\modmult_1/xin[1023] ), .A(n40039), .Z(n40037) );
  IV U42681 ( .A(n40038), .Z(n40039) );
  XNOR U42682 ( .A(m[218]), .B(n40040), .Z(n40038) );
  NAND U42683 ( .A(n40041), .B(mul_pow), .Z(n40040) );
  XOR U42684 ( .A(m[218]), .B(c[218]), .Z(n40041) );
  XOR U42685 ( .A(n40042), .B(n40043), .Z(n40034) );
  ANDN U42686 ( .B(n40044), .A(n31180), .Z(n40042) );
  XNOR U42687 ( .A(\modmult_1/zin[0][216] ), .B(n40045), .Z(n31180) );
  IV U42688 ( .A(n40043), .Z(n40045) );
  XOR U42689 ( .A(n40043), .B(n31181), .Z(n40044) );
  XNOR U42690 ( .A(n40046), .B(n40047), .Z(n31181) );
  ANDN U42691 ( .B(\modmult_1/xin[1023] ), .A(n40048), .Z(n40046) );
  IV U42692 ( .A(n40047), .Z(n40048) );
  XNOR U42693 ( .A(m[217]), .B(n40049), .Z(n40047) );
  NAND U42694 ( .A(n40050), .B(mul_pow), .Z(n40049) );
  XOR U42695 ( .A(m[217]), .B(c[217]), .Z(n40050) );
  XOR U42696 ( .A(n40051), .B(n40052), .Z(n40043) );
  ANDN U42697 ( .B(n40053), .A(n31178), .Z(n40051) );
  XNOR U42698 ( .A(\modmult_1/zin[0][215] ), .B(n40054), .Z(n31178) );
  IV U42699 ( .A(n40052), .Z(n40054) );
  XOR U42700 ( .A(n40052), .B(n31179), .Z(n40053) );
  XNOR U42701 ( .A(n40055), .B(n40056), .Z(n31179) );
  ANDN U42702 ( .B(\modmult_1/xin[1023] ), .A(n40057), .Z(n40055) );
  IV U42703 ( .A(n40056), .Z(n40057) );
  XNOR U42704 ( .A(m[216]), .B(n40058), .Z(n40056) );
  NAND U42705 ( .A(n40059), .B(mul_pow), .Z(n40058) );
  XOR U42706 ( .A(m[216]), .B(c[216]), .Z(n40059) );
  XOR U42707 ( .A(n40060), .B(n40061), .Z(n40052) );
  ANDN U42708 ( .B(n40062), .A(n31176), .Z(n40060) );
  XNOR U42709 ( .A(\modmult_1/zin[0][214] ), .B(n40063), .Z(n31176) );
  IV U42710 ( .A(n40061), .Z(n40063) );
  XOR U42711 ( .A(n40061), .B(n31177), .Z(n40062) );
  XNOR U42712 ( .A(n40064), .B(n40065), .Z(n31177) );
  ANDN U42713 ( .B(\modmult_1/xin[1023] ), .A(n40066), .Z(n40064) );
  IV U42714 ( .A(n40065), .Z(n40066) );
  XNOR U42715 ( .A(m[215]), .B(n40067), .Z(n40065) );
  NAND U42716 ( .A(n40068), .B(mul_pow), .Z(n40067) );
  XOR U42717 ( .A(m[215]), .B(c[215]), .Z(n40068) );
  XOR U42718 ( .A(n40069), .B(n40070), .Z(n40061) );
  ANDN U42719 ( .B(n40071), .A(n31174), .Z(n40069) );
  XNOR U42720 ( .A(\modmult_1/zin[0][213] ), .B(n40072), .Z(n31174) );
  IV U42721 ( .A(n40070), .Z(n40072) );
  XOR U42722 ( .A(n40070), .B(n31175), .Z(n40071) );
  XNOR U42723 ( .A(n40073), .B(n40074), .Z(n31175) );
  ANDN U42724 ( .B(\modmult_1/xin[1023] ), .A(n40075), .Z(n40073) );
  IV U42725 ( .A(n40074), .Z(n40075) );
  XNOR U42726 ( .A(m[214]), .B(n40076), .Z(n40074) );
  NAND U42727 ( .A(n40077), .B(mul_pow), .Z(n40076) );
  XOR U42728 ( .A(m[214]), .B(c[214]), .Z(n40077) );
  XOR U42729 ( .A(n40078), .B(n40079), .Z(n40070) );
  ANDN U42730 ( .B(n40080), .A(n31172), .Z(n40078) );
  XNOR U42731 ( .A(\modmult_1/zin[0][212] ), .B(n40081), .Z(n31172) );
  IV U42732 ( .A(n40079), .Z(n40081) );
  XOR U42733 ( .A(n40079), .B(n31173), .Z(n40080) );
  XNOR U42734 ( .A(n40082), .B(n40083), .Z(n31173) );
  ANDN U42735 ( .B(\modmult_1/xin[1023] ), .A(n40084), .Z(n40082) );
  IV U42736 ( .A(n40083), .Z(n40084) );
  XNOR U42737 ( .A(m[213]), .B(n40085), .Z(n40083) );
  NAND U42738 ( .A(n40086), .B(mul_pow), .Z(n40085) );
  XOR U42739 ( .A(m[213]), .B(c[213]), .Z(n40086) );
  XOR U42740 ( .A(n40087), .B(n40088), .Z(n40079) );
  ANDN U42741 ( .B(n40089), .A(n31170), .Z(n40087) );
  XNOR U42742 ( .A(\modmult_1/zin[0][211] ), .B(n40090), .Z(n31170) );
  IV U42743 ( .A(n40088), .Z(n40090) );
  XOR U42744 ( .A(n40088), .B(n31171), .Z(n40089) );
  XNOR U42745 ( .A(n40091), .B(n40092), .Z(n31171) );
  ANDN U42746 ( .B(\modmult_1/xin[1023] ), .A(n40093), .Z(n40091) );
  IV U42747 ( .A(n40092), .Z(n40093) );
  XNOR U42748 ( .A(m[212]), .B(n40094), .Z(n40092) );
  NAND U42749 ( .A(n40095), .B(mul_pow), .Z(n40094) );
  XOR U42750 ( .A(m[212]), .B(c[212]), .Z(n40095) );
  XOR U42751 ( .A(n40096), .B(n40097), .Z(n40088) );
  ANDN U42752 ( .B(n40098), .A(n31168), .Z(n40096) );
  XNOR U42753 ( .A(\modmult_1/zin[0][210] ), .B(n40099), .Z(n31168) );
  IV U42754 ( .A(n40097), .Z(n40099) );
  XOR U42755 ( .A(n40097), .B(n31169), .Z(n40098) );
  XNOR U42756 ( .A(n40100), .B(n40101), .Z(n31169) );
  ANDN U42757 ( .B(\modmult_1/xin[1023] ), .A(n40102), .Z(n40100) );
  IV U42758 ( .A(n40101), .Z(n40102) );
  XNOR U42759 ( .A(m[211]), .B(n40103), .Z(n40101) );
  NAND U42760 ( .A(n40104), .B(mul_pow), .Z(n40103) );
  XOR U42761 ( .A(m[211]), .B(c[211]), .Z(n40104) );
  XOR U42762 ( .A(n40105), .B(n40106), .Z(n40097) );
  ANDN U42763 ( .B(n40107), .A(n31166), .Z(n40105) );
  XNOR U42764 ( .A(\modmult_1/zin[0][209] ), .B(n40108), .Z(n31166) );
  IV U42765 ( .A(n40106), .Z(n40108) );
  XOR U42766 ( .A(n40106), .B(n31167), .Z(n40107) );
  XNOR U42767 ( .A(n40109), .B(n40110), .Z(n31167) );
  ANDN U42768 ( .B(\modmult_1/xin[1023] ), .A(n40111), .Z(n40109) );
  IV U42769 ( .A(n40110), .Z(n40111) );
  XNOR U42770 ( .A(m[210]), .B(n40112), .Z(n40110) );
  NAND U42771 ( .A(n40113), .B(mul_pow), .Z(n40112) );
  XOR U42772 ( .A(m[210]), .B(c[210]), .Z(n40113) );
  XOR U42773 ( .A(n40114), .B(n40115), .Z(n40106) );
  ANDN U42774 ( .B(n40116), .A(n31164), .Z(n40114) );
  XNOR U42775 ( .A(\modmult_1/zin[0][208] ), .B(n40117), .Z(n31164) );
  IV U42776 ( .A(n40115), .Z(n40117) );
  XOR U42777 ( .A(n40115), .B(n31165), .Z(n40116) );
  XNOR U42778 ( .A(n40118), .B(n40119), .Z(n31165) );
  ANDN U42779 ( .B(\modmult_1/xin[1023] ), .A(n40120), .Z(n40118) );
  IV U42780 ( .A(n40119), .Z(n40120) );
  XNOR U42781 ( .A(m[209]), .B(n40121), .Z(n40119) );
  NAND U42782 ( .A(n40122), .B(mul_pow), .Z(n40121) );
  XOR U42783 ( .A(m[209]), .B(c[209]), .Z(n40122) );
  XOR U42784 ( .A(n40123), .B(n40124), .Z(n40115) );
  ANDN U42785 ( .B(n40125), .A(n31162), .Z(n40123) );
  XNOR U42786 ( .A(\modmult_1/zin[0][207] ), .B(n40126), .Z(n31162) );
  IV U42787 ( .A(n40124), .Z(n40126) );
  XOR U42788 ( .A(n40124), .B(n31163), .Z(n40125) );
  XNOR U42789 ( .A(n40127), .B(n40128), .Z(n31163) );
  ANDN U42790 ( .B(\modmult_1/xin[1023] ), .A(n40129), .Z(n40127) );
  IV U42791 ( .A(n40128), .Z(n40129) );
  XNOR U42792 ( .A(m[208]), .B(n40130), .Z(n40128) );
  NAND U42793 ( .A(n40131), .B(mul_pow), .Z(n40130) );
  XOR U42794 ( .A(m[208]), .B(c[208]), .Z(n40131) );
  XOR U42795 ( .A(n40132), .B(n40133), .Z(n40124) );
  ANDN U42796 ( .B(n40134), .A(n31160), .Z(n40132) );
  XNOR U42797 ( .A(\modmult_1/zin[0][206] ), .B(n40135), .Z(n31160) );
  IV U42798 ( .A(n40133), .Z(n40135) );
  XOR U42799 ( .A(n40133), .B(n31161), .Z(n40134) );
  XNOR U42800 ( .A(n40136), .B(n40137), .Z(n31161) );
  ANDN U42801 ( .B(\modmult_1/xin[1023] ), .A(n40138), .Z(n40136) );
  IV U42802 ( .A(n40137), .Z(n40138) );
  XNOR U42803 ( .A(m[207]), .B(n40139), .Z(n40137) );
  NAND U42804 ( .A(n40140), .B(mul_pow), .Z(n40139) );
  XOR U42805 ( .A(m[207]), .B(c[207]), .Z(n40140) );
  XOR U42806 ( .A(n40141), .B(n40142), .Z(n40133) );
  ANDN U42807 ( .B(n40143), .A(n31158), .Z(n40141) );
  XNOR U42808 ( .A(\modmult_1/zin[0][205] ), .B(n40144), .Z(n31158) );
  IV U42809 ( .A(n40142), .Z(n40144) );
  XOR U42810 ( .A(n40142), .B(n31159), .Z(n40143) );
  XNOR U42811 ( .A(n40145), .B(n40146), .Z(n31159) );
  ANDN U42812 ( .B(\modmult_1/xin[1023] ), .A(n40147), .Z(n40145) );
  IV U42813 ( .A(n40146), .Z(n40147) );
  XNOR U42814 ( .A(m[206]), .B(n40148), .Z(n40146) );
  NAND U42815 ( .A(n40149), .B(mul_pow), .Z(n40148) );
  XOR U42816 ( .A(m[206]), .B(c[206]), .Z(n40149) );
  XOR U42817 ( .A(n40150), .B(n40151), .Z(n40142) );
  ANDN U42818 ( .B(n40152), .A(n31156), .Z(n40150) );
  XNOR U42819 ( .A(\modmult_1/zin[0][204] ), .B(n40153), .Z(n31156) );
  IV U42820 ( .A(n40151), .Z(n40153) );
  XOR U42821 ( .A(n40151), .B(n31157), .Z(n40152) );
  XNOR U42822 ( .A(n40154), .B(n40155), .Z(n31157) );
  ANDN U42823 ( .B(\modmult_1/xin[1023] ), .A(n40156), .Z(n40154) );
  IV U42824 ( .A(n40155), .Z(n40156) );
  XNOR U42825 ( .A(m[205]), .B(n40157), .Z(n40155) );
  NAND U42826 ( .A(n40158), .B(mul_pow), .Z(n40157) );
  XOR U42827 ( .A(m[205]), .B(c[205]), .Z(n40158) );
  XOR U42828 ( .A(n40159), .B(n40160), .Z(n40151) );
  ANDN U42829 ( .B(n40161), .A(n31154), .Z(n40159) );
  XNOR U42830 ( .A(\modmult_1/zin[0][203] ), .B(n40162), .Z(n31154) );
  IV U42831 ( .A(n40160), .Z(n40162) );
  XOR U42832 ( .A(n40160), .B(n31155), .Z(n40161) );
  XNOR U42833 ( .A(n40163), .B(n40164), .Z(n31155) );
  ANDN U42834 ( .B(\modmult_1/xin[1023] ), .A(n40165), .Z(n40163) );
  IV U42835 ( .A(n40164), .Z(n40165) );
  XNOR U42836 ( .A(m[204]), .B(n40166), .Z(n40164) );
  NAND U42837 ( .A(n40167), .B(mul_pow), .Z(n40166) );
  XOR U42838 ( .A(m[204]), .B(c[204]), .Z(n40167) );
  XOR U42839 ( .A(n40168), .B(n40169), .Z(n40160) );
  ANDN U42840 ( .B(n40170), .A(n31152), .Z(n40168) );
  XNOR U42841 ( .A(\modmult_1/zin[0][202] ), .B(n40171), .Z(n31152) );
  IV U42842 ( .A(n40169), .Z(n40171) );
  XOR U42843 ( .A(n40169), .B(n31153), .Z(n40170) );
  XNOR U42844 ( .A(n40172), .B(n40173), .Z(n31153) );
  ANDN U42845 ( .B(\modmult_1/xin[1023] ), .A(n40174), .Z(n40172) );
  IV U42846 ( .A(n40173), .Z(n40174) );
  XNOR U42847 ( .A(m[203]), .B(n40175), .Z(n40173) );
  NAND U42848 ( .A(n40176), .B(mul_pow), .Z(n40175) );
  XOR U42849 ( .A(m[203]), .B(c[203]), .Z(n40176) );
  XOR U42850 ( .A(n40177), .B(n40178), .Z(n40169) );
  ANDN U42851 ( .B(n40179), .A(n31150), .Z(n40177) );
  XNOR U42852 ( .A(\modmult_1/zin[0][201] ), .B(n40180), .Z(n31150) );
  IV U42853 ( .A(n40178), .Z(n40180) );
  XOR U42854 ( .A(n40178), .B(n31151), .Z(n40179) );
  XNOR U42855 ( .A(n40181), .B(n40182), .Z(n31151) );
  ANDN U42856 ( .B(\modmult_1/xin[1023] ), .A(n40183), .Z(n40181) );
  IV U42857 ( .A(n40182), .Z(n40183) );
  XNOR U42858 ( .A(m[202]), .B(n40184), .Z(n40182) );
  NAND U42859 ( .A(n40185), .B(mul_pow), .Z(n40184) );
  XOR U42860 ( .A(m[202]), .B(c[202]), .Z(n40185) );
  XOR U42861 ( .A(n40186), .B(n40187), .Z(n40178) );
  ANDN U42862 ( .B(n40188), .A(n31148), .Z(n40186) );
  XNOR U42863 ( .A(\modmult_1/zin[0][200] ), .B(n40189), .Z(n31148) );
  IV U42864 ( .A(n40187), .Z(n40189) );
  XOR U42865 ( .A(n40187), .B(n31149), .Z(n40188) );
  XNOR U42866 ( .A(n40190), .B(n40191), .Z(n31149) );
  ANDN U42867 ( .B(\modmult_1/xin[1023] ), .A(n40192), .Z(n40190) );
  IV U42868 ( .A(n40191), .Z(n40192) );
  XNOR U42869 ( .A(m[201]), .B(n40193), .Z(n40191) );
  NAND U42870 ( .A(n40194), .B(mul_pow), .Z(n40193) );
  XOR U42871 ( .A(m[201]), .B(c[201]), .Z(n40194) );
  XOR U42872 ( .A(n40195), .B(n40196), .Z(n40187) );
  ANDN U42873 ( .B(n40197), .A(n31146), .Z(n40195) );
  XNOR U42874 ( .A(\modmult_1/zin[0][199] ), .B(n40198), .Z(n31146) );
  IV U42875 ( .A(n40196), .Z(n40198) );
  XOR U42876 ( .A(n40196), .B(n31147), .Z(n40197) );
  XNOR U42877 ( .A(n40199), .B(n40200), .Z(n31147) );
  ANDN U42878 ( .B(\modmult_1/xin[1023] ), .A(n40201), .Z(n40199) );
  IV U42879 ( .A(n40200), .Z(n40201) );
  XNOR U42880 ( .A(m[200]), .B(n40202), .Z(n40200) );
  NAND U42881 ( .A(n40203), .B(mul_pow), .Z(n40202) );
  XOR U42882 ( .A(m[200]), .B(c[200]), .Z(n40203) );
  XOR U42883 ( .A(n40204), .B(n40205), .Z(n40196) );
  ANDN U42884 ( .B(n40206), .A(n31144), .Z(n40204) );
  XNOR U42885 ( .A(\modmult_1/zin[0][198] ), .B(n40207), .Z(n31144) );
  IV U42886 ( .A(n40205), .Z(n40207) );
  XOR U42887 ( .A(n40205), .B(n31145), .Z(n40206) );
  XNOR U42888 ( .A(n40208), .B(n40209), .Z(n31145) );
  ANDN U42889 ( .B(\modmult_1/xin[1023] ), .A(n40210), .Z(n40208) );
  IV U42890 ( .A(n40209), .Z(n40210) );
  XNOR U42891 ( .A(m[199]), .B(n40211), .Z(n40209) );
  NAND U42892 ( .A(n40212), .B(mul_pow), .Z(n40211) );
  XOR U42893 ( .A(m[199]), .B(c[199]), .Z(n40212) );
  XOR U42894 ( .A(n40213), .B(n40214), .Z(n40205) );
  ANDN U42895 ( .B(n40215), .A(n31142), .Z(n40213) );
  XNOR U42896 ( .A(\modmult_1/zin[0][197] ), .B(n40216), .Z(n31142) );
  IV U42897 ( .A(n40214), .Z(n40216) );
  XOR U42898 ( .A(n40214), .B(n31143), .Z(n40215) );
  XNOR U42899 ( .A(n40217), .B(n40218), .Z(n31143) );
  ANDN U42900 ( .B(\modmult_1/xin[1023] ), .A(n40219), .Z(n40217) );
  IV U42901 ( .A(n40218), .Z(n40219) );
  XNOR U42902 ( .A(m[198]), .B(n40220), .Z(n40218) );
  NAND U42903 ( .A(n40221), .B(mul_pow), .Z(n40220) );
  XOR U42904 ( .A(m[198]), .B(c[198]), .Z(n40221) );
  XOR U42905 ( .A(n40222), .B(n40223), .Z(n40214) );
  ANDN U42906 ( .B(n40224), .A(n31140), .Z(n40222) );
  XNOR U42907 ( .A(\modmult_1/zin[0][196] ), .B(n40225), .Z(n31140) );
  IV U42908 ( .A(n40223), .Z(n40225) );
  XOR U42909 ( .A(n40223), .B(n31141), .Z(n40224) );
  XNOR U42910 ( .A(n40226), .B(n40227), .Z(n31141) );
  ANDN U42911 ( .B(\modmult_1/xin[1023] ), .A(n40228), .Z(n40226) );
  IV U42912 ( .A(n40227), .Z(n40228) );
  XNOR U42913 ( .A(m[197]), .B(n40229), .Z(n40227) );
  NAND U42914 ( .A(n40230), .B(mul_pow), .Z(n40229) );
  XOR U42915 ( .A(m[197]), .B(c[197]), .Z(n40230) );
  XOR U42916 ( .A(n40231), .B(n40232), .Z(n40223) );
  ANDN U42917 ( .B(n40233), .A(n31138), .Z(n40231) );
  XNOR U42918 ( .A(\modmult_1/zin[0][195] ), .B(n40234), .Z(n31138) );
  IV U42919 ( .A(n40232), .Z(n40234) );
  XOR U42920 ( .A(n40232), .B(n31139), .Z(n40233) );
  XNOR U42921 ( .A(n40235), .B(n40236), .Z(n31139) );
  ANDN U42922 ( .B(\modmult_1/xin[1023] ), .A(n40237), .Z(n40235) );
  IV U42923 ( .A(n40236), .Z(n40237) );
  XNOR U42924 ( .A(m[196]), .B(n40238), .Z(n40236) );
  NAND U42925 ( .A(n40239), .B(mul_pow), .Z(n40238) );
  XOR U42926 ( .A(m[196]), .B(c[196]), .Z(n40239) );
  XOR U42927 ( .A(n40240), .B(n40241), .Z(n40232) );
  ANDN U42928 ( .B(n40242), .A(n31136), .Z(n40240) );
  XNOR U42929 ( .A(\modmult_1/zin[0][194] ), .B(n40243), .Z(n31136) );
  IV U42930 ( .A(n40241), .Z(n40243) );
  XOR U42931 ( .A(n40241), .B(n31137), .Z(n40242) );
  XNOR U42932 ( .A(n40244), .B(n40245), .Z(n31137) );
  ANDN U42933 ( .B(\modmult_1/xin[1023] ), .A(n40246), .Z(n40244) );
  IV U42934 ( .A(n40245), .Z(n40246) );
  XNOR U42935 ( .A(m[195]), .B(n40247), .Z(n40245) );
  NAND U42936 ( .A(n40248), .B(mul_pow), .Z(n40247) );
  XOR U42937 ( .A(m[195]), .B(c[195]), .Z(n40248) );
  XOR U42938 ( .A(n40249), .B(n40250), .Z(n40241) );
  ANDN U42939 ( .B(n40251), .A(n31134), .Z(n40249) );
  XNOR U42940 ( .A(\modmult_1/zin[0][193] ), .B(n40252), .Z(n31134) );
  IV U42941 ( .A(n40250), .Z(n40252) );
  XOR U42942 ( .A(n40250), .B(n31135), .Z(n40251) );
  XNOR U42943 ( .A(n40253), .B(n40254), .Z(n31135) );
  ANDN U42944 ( .B(\modmult_1/xin[1023] ), .A(n40255), .Z(n40253) );
  IV U42945 ( .A(n40254), .Z(n40255) );
  XNOR U42946 ( .A(m[194]), .B(n40256), .Z(n40254) );
  NAND U42947 ( .A(n40257), .B(mul_pow), .Z(n40256) );
  XOR U42948 ( .A(m[194]), .B(c[194]), .Z(n40257) );
  XOR U42949 ( .A(n40258), .B(n40259), .Z(n40250) );
  ANDN U42950 ( .B(n40260), .A(n31132), .Z(n40258) );
  XNOR U42951 ( .A(\modmult_1/zin[0][192] ), .B(n40261), .Z(n31132) );
  IV U42952 ( .A(n40259), .Z(n40261) );
  XOR U42953 ( .A(n40259), .B(n31133), .Z(n40260) );
  XNOR U42954 ( .A(n40262), .B(n40263), .Z(n31133) );
  ANDN U42955 ( .B(\modmult_1/xin[1023] ), .A(n40264), .Z(n40262) );
  IV U42956 ( .A(n40263), .Z(n40264) );
  XNOR U42957 ( .A(m[193]), .B(n40265), .Z(n40263) );
  NAND U42958 ( .A(n40266), .B(mul_pow), .Z(n40265) );
  XOR U42959 ( .A(m[193]), .B(c[193]), .Z(n40266) );
  XOR U42960 ( .A(n40267), .B(n40268), .Z(n40259) );
  ANDN U42961 ( .B(n40269), .A(n31130), .Z(n40267) );
  XNOR U42962 ( .A(\modmult_1/zin[0][191] ), .B(n40270), .Z(n31130) );
  IV U42963 ( .A(n40268), .Z(n40270) );
  XOR U42964 ( .A(n40268), .B(n31131), .Z(n40269) );
  XNOR U42965 ( .A(n40271), .B(n40272), .Z(n31131) );
  ANDN U42966 ( .B(\modmult_1/xin[1023] ), .A(n40273), .Z(n40271) );
  IV U42967 ( .A(n40272), .Z(n40273) );
  XNOR U42968 ( .A(m[192]), .B(n40274), .Z(n40272) );
  NAND U42969 ( .A(n40275), .B(mul_pow), .Z(n40274) );
  XOR U42970 ( .A(m[192]), .B(c[192]), .Z(n40275) );
  XOR U42971 ( .A(n40276), .B(n40277), .Z(n40268) );
  ANDN U42972 ( .B(n40278), .A(n31128), .Z(n40276) );
  XNOR U42973 ( .A(\modmult_1/zin[0][190] ), .B(n40279), .Z(n31128) );
  IV U42974 ( .A(n40277), .Z(n40279) );
  XOR U42975 ( .A(n40277), .B(n31129), .Z(n40278) );
  XNOR U42976 ( .A(n40280), .B(n40281), .Z(n31129) );
  ANDN U42977 ( .B(\modmult_1/xin[1023] ), .A(n40282), .Z(n40280) );
  IV U42978 ( .A(n40281), .Z(n40282) );
  XNOR U42979 ( .A(m[191]), .B(n40283), .Z(n40281) );
  NAND U42980 ( .A(n40284), .B(mul_pow), .Z(n40283) );
  XOR U42981 ( .A(m[191]), .B(c[191]), .Z(n40284) );
  XOR U42982 ( .A(n40285), .B(n40286), .Z(n40277) );
  ANDN U42983 ( .B(n40287), .A(n31126), .Z(n40285) );
  XNOR U42984 ( .A(\modmult_1/zin[0][189] ), .B(n40288), .Z(n31126) );
  IV U42985 ( .A(n40286), .Z(n40288) );
  XOR U42986 ( .A(n40286), .B(n31127), .Z(n40287) );
  XNOR U42987 ( .A(n40289), .B(n40290), .Z(n31127) );
  ANDN U42988 ( .B(\modmult_1/xin[1023] ), .A(n40291), .Z(n40289) );
  IV U42989 ( .A(n40290), .Z(n40291) );
  XNOR U42990 ( .A(m[190]), .B(n40292), .Z(n40290) );
  NAND U42991 ( .A(n40293), .B(mul_pow), .Z(n40292) );
  XOR U42992 ( .A(m[190]), .B(c[190]), .Z(n40293) );
  XOR U42993 ( .A(n40294), .B(n40295), .Z(n40286) );
  ANDN U42994 ( .B(n40296), .A(n31124), .Z(n40294) );
  XNOR U42995 ( .A(\modmult_1/zin[0][188] ), .B(n40297), .Z(n31124) );
  IV U42996 ( .A(n40295), .Z(n40297) );
  XOR U42997 ( .A(n40295), .B(n31125), .Z(n40296) );
  XNOR U42998 ( .A(n40298), .B(n40299), .Z(n31125) );
  ANDN U42999 ( .B(\modmult_1/xin[1023] ), .A(n40300), .Z(n40298) );
  IV U43000 ( .A(n40299), .Z(n40300) );
  XNOR U43001 ( .A(m[189]), .B(n40301), .Z(n40299) );
  NAND U43002 ( .A(n40302), .B(mul_pow), .Z(n40301) );
  XOR U43003 ( .A(m[189]), .B(c[189]), .Z(n40302) );
  XOR U43004 ( .A(n40303), .B(n40304), .Z(n40295) );
  ANDN U43005 ( .B(n40305), .A(n31122), .Z(n40303) );
  XNOR U43006 ( .A(\modmult_1/zin[0][187] ), .B(n40306), .Z(n31122) );
  IV U43007 ( .A(n40304), .Z(n40306) );
  XOR U43008 ( .A(n40304), .B(n31123), .Z(n40305) );
  XNOR U43009 ( .A(n40307), .B(n40308), .Z(n31123) );
  ANDN U43010 ( .B(\modmult_1/xin[1023] ), .A(n40309), .Z(n40307) );
  IV U43011 ( .A(n40308), .Z(n40309) );
  XNOR U43012 ( .A(m[188]), .B(n40310), .Z(n40308) );
  NAND U43013 ( .A(n40311), .B(mul_pow), .Z(n40310) );
  XOR U43014 ( .A(m[188]), .B(c[188]), .Z(n40311) );
  XOR U43015 ( .A(n40312), .B(n40313), .Z(n40304) );
  ANDN U43016 ( .B(n40314), .A(n31120), .Z(n40312) );
  XNOR U43017 ( .A(\modmult_1/zin[0][186] ), .B(n40315), .Z(n31120) );
  IV U43018 ( .A(n40313), .Z(n40315) );
  XOR U43019 ( .A(n40313), .B(n31121), .Z(n40314) );
  XNOR U43020 ( .A(n40316), .B(n40317), .Z(n31121) );
  ANDN U43021 ( .B(\modmult_1/xin[1023] ), .A(n40318), .Z(n40316) );
  IV U43022 ( .A(n40317), .Z(n40318) );
  XNOR U43023 ( .A(m[187]), .B(n40319), .Z(n40317) );
  NAND U43024 ( .A(n40320), .B(mul_pow), .Z(n40319) );
  XOR U43025 ( .A(m[187]), .B(c[187]), .Z(n40320) );
  XOR U43026 ( .A(n40321), .B(n40322), .Z(n40313) );
  ANDN U43027 ( .B(n40323), .A(n31118), .Z(n40321) );
  XNOR U43028 ( .A(\modmult_1/zin[0][185] ), .B(n40324), .Z(n31118) );
  IV U43029 ( .A(n40322), .Z(n40324) );
  XOR U43030 ( .A(n40322), .B(n31119), .Z(n40323) );
  XNOR U43031 ( .A(n40325), .B(n40326), .Z(n31119) );
  ANDN U43032 ( .B(\modmult_1/xin[1023] ), .A(n40327), .Z(n40325) );
  IV U43033 ( .A(n40326), .Z(n40327) );
  XNOR U43034 ( .A(m[186]), .B(n40328), .Z(n40326) );
  NAND U43035 ( .A(n40329), .B(mul_pow), .Z(n40328) );
  XOR U43036 ( .A(m[186]), .B(c[186]), .Z(n40329) );
  XOR U43037 ( .A(n40330), .B(n40331), .Z(n40322) );
  ANDN U43038 ( .B(n40332), .A(n31116), .Z(n40330) );
  XNOR U43039 ( .A(\modmult_1/zin[0][184] ), .B(n40333), .Z(n31116) );
  IV U43040 ( .A(n40331), .Z(n40333) );
  XOR U43041 ( .A(n40331), .B(n31117), .Z(n40332) );
  XNOR U43042 ( .A(n40334), .B(n40335), .Z(n31117) );
  ANDN U43043 ( .B(\modmult_1/xin[1023] ), .A(n40336), .Z(n40334) );
  IV U43044 ( .A(n40335), .Z(n40336) );
  XNOR U43045 ( .A(m[185]), .B(n40337), .Z(n40335) );
  NAND U43046 ( .A(n40338), .B(mul_pow), .Z(n40337) );
  XOR U43047 ( .A(m[185]), .B(c[185]), .Z(n40338) );
  XOR U43048 ( .A(n40339), .B(n40340), .Z(n40331) );
  ANDN U43049 ( .B(n40341), .A(n31114), .Z(n40339) );
  XNOR U43050 ( .A(\modmult_1/zin[0][183] ), .B(n40342), .Z(n31114) );
  IV U43051 ( .A(n40340), .Z(n40342) );
  XOR U43052 ( .A(n40340), .B(n31115), .Z(n40341) );
  XNOR U43053 ( .A(n40343), .B(n40344), .Z(n31115) );
  ANDN U43054 ( .B(\modmult_1/xin[1023] ), .A(n40345), .Z(n40343) );
  IV U43055 ( .A(n40344), .Z(n40345) );
  XNOR U43056 ( .A(m[184]), .B(n40346), .Z(n40344) );
  NAND U43057 ( .A(n40347), .B(mul_pow), .Z(n40346) );
  XOR U43058 ( .A(m[184]), .B(c[184]), .Z(n40347) );
  XOR U43059 ( .A(n40348), .B(n40349), .Z(n40340) );
  ANDN U43060 ( .B(n40350), .A(n31112), .Z(n40348) );
  XNOR U43061 ( .A(\modmult_1/zin[0][182] ), .B(n40351), .Z(n31112) );
  IV U43062 ( .A(n40349), .Z(n40351) );
  XOR U43063 ( .A(n40349), .B(n31113), .Z(n40350) );
  XNOR U43064 ( .A(n40352), .B(n40353), .Z(n31113) );
  ANDN U43065 ( .B(\modmult_1/xin[1023] ), .A(n40354), .Z(n40352) );
  IV U43066 ( .A(n40353), .Z(n40354) );
  XNOR U43067 ( .A(m[183]), .B(n40355), .Z(n40353) );
  NAND U43068 ( .A(n40356), .B(mul_pow), .Z(n40355) );
  XOR U43069 ( .A(m[183]), .B(c[183]), .Z(n40356) );
  XOR U43070 ( .A(n40357), .B(n40358), .Z(n40349) );
  ANDN U43071 ( .B(n40359), .A(n31110), .Z(n40357) );
  XNOR U43072 ( .A(\modmult_1/zin[0][181] ), .B(n40360), .Z(n31110) );
  IV U43073 ( .A(n40358), .Z(n40360) );
  XOR U43074 ( .A(n40358), .B(n31111), .Z(n40359) );
  XNOR U43075 ( .A(n40361), .B(n40362), .Z(n31111) );
  ANDN U43076 ( .B(\modmult_1/xin[1023] ), .A(n40363), .Z(n40361) );
  IV U43077 ( .A(n40362), .Z(n40363) );
  XNOR U43078 ( .A(m[182]), .B(n40364), .Z(n40362) );
  NAND U43079 ( .A(n40365), .B(mul_pow), .Z(n40364) );
  XOR U43080 ( .A(m[182]), .B(c[182]), .Z(n40365) );
  XOR U43081 ( .A(n40366), .B(n40367), .Z(n40358) );
  ANDN U43082 ( .B(n40368), .A(n31108), .Z(n40366) );
  XNOR U43083 ( .A(\modmult_1/zin[0][180] ), .B(n40369), .Z(n31108) );
  IV U43084 ( .A(n40367), .Z(n40369) );
  XOR U43085 ( .A(n40367), .B(n31109), .Z(n40368) );
  XNOR U43086 ( .A(n40370), .B(n40371), .Z(n31109) );
  ANDN U43087 ( .B(\modmult_1/xin[1023] ), .A(n40372), .Z(n40370) );
  IV U43088 ( .A(n40371), .Z(n40372) );
  XNOR U43089 ( .A(m[181]), .B(n40373), .Z(n40371) );
  NAND U43090 ( .A(n40374), .B(mul_pow), .Z(n40373) );
  XOR U43091 ( .A(m[181]), .B(c[181]), .Z(n40374) );
  XOR U43092 ( .A(n40375), .B(n40376), .Z(n40367) );
  ANDN U43093 ( .B(n40377), .A(n31106), .Z(n40375) );
  XNOR U43094 ( .A(\modmult_1/zin[0][179] ), .B(n40378), .Z(n31106) );
  IV U43095 ( .A(n40376), .Z(n40378) );
  XOR U43096 ( .A(n40376), .B(n31107), .Z(n40377) );
  XNOR U43097 ( .A(n40379), .B(n40380), .Z(n31107) );
  ANDN U43098 ( .B(\modmult_1/xin[1023] ), .A(n40381), .Z(n40379) );
  IV U43099 ( .A(n40380), .Z(n40381) );
  XNOR U43100 ( .A(m[180]), .B(n40382), .Z(n40380) );
  NAND U43101 ( .A(n40383), .B(mul_pow), .Z(n40382) );
  XOR U43102 ( .A(m[180]), .B(c[180]), .Z(n40383) );
  XOR U43103 ( .A(n40384), .B(n40385), .Z(n40376) );
  ANDN U43104 ( .B(n40386), .A(n31104), .Z(n40384) );
  XNOR U43105 ( .A(\modmult_1/zin[0][178] ), .B(n40387), .Z(n31104) );
  IV U43106 ( .A(n40385), .Z(n40387) );
  XOR U43107 ( .A(n40385), .B(n31105), .Z(n40386) );
  XNOR U43108 ( .A(n40388), .B(n40389), .Z(n31105) );
  ANDN U43109 ( .B(\modmult_1/xin[1023] ), .A(n40390), .Z(n40388) );
  IV U43110 ( .A(n40389), .Z(n40390) );
  XNOR U43111 ( .A(m[179]), .B(n40391), .Z(n40389) );
  NAND U43112 ( .A(n40392), .B(mul_pow), .Z(n40391) );
  XOR U43113 ( .A(m[179]), .B(c[179]), .Z(n40392) );
  XOR U43114 ( .A(n40393), .B(n40394), .Z(n40385) );
  ANDN U43115 ( .B(n40395), .A(n31102), .Z(n40393) );
  XNOR U43116 ( .A(\modmult_1/zin[0][177] ), .B(n40396), .Z(n31102) );
  IV U43117 ( .A(n40394), .Z(n40396) );
  XOR U43118 ( .A(n40394), .B(n31103), .Z(n40395) );
  XNOR U43119 ( .A(n40397), .B(n40398), .Z(n31103) );
  ANDN U43120 ( .B(\modmult_1/xin[1023] ), .A(n40399), .Z(n40397) );
  IV U43121 ( .A(n40398), .Z(n40399) );
  XNOR U43122 ( .A(m[178]), .B(n40400), .Z(n40398) );
  NAND U43123 ( .A(n40401), .B(mul_pow), .Z(n40400) );
  XOR U43124 ( .A(m[178]), .B(c[178]), .Z(n40401) );
  XOR U43125 ( .A(n40402), .B(n40403), .Z(n40394) );
  ANDN U43126 ( .B(n40404), .A(n31100), .Z(n40402) );
  XNOR U43127 ( .A(\modmult_1/zin[0][176] ), .B(n40405), .Z(n31100) );
  IV U43128 ( .A(n40403), .Z(n40405) );
  XOR U43129 ( .A(n40403), .B(n31101), .Z(n40404) );
  XNOR U43130 ( .A(n40406), .B(n40407), .Z(n31101) );
  ANDN U43131 ( .B(\modmult_1/xin[1023] ), .A(n40408), .Z(n40406) );
  IV U43132 ( .A(n40407), .Z(n40408) );
  XNOR U43133 ( .A(m[177]), .B(n40409), .Z(n40407) );
  NAND U43134 ( .A(n40410), .B(mul_pow), .Z(n40409) );
  XOR U43135 ( .A(m[177]), .B(c[177]), .Z(n40410) );
  XOR U43136 ( .A(n40411), .B(n40412), .Z(n40403) );
  ANDN U43137 ( .B(n40413), .A(n31098), .Z(n40411) );
  XNOR U43138 ( .A(\modmult_1/zin[0][175] ), .B(n40414), .Z(n31098) );
  IV U43139 ( .A(n40412), .Z(n40414) );
  XOR U43140 ( .A(n40412), .B(n31099), .Z(n40413) );
  XNOR U43141 ( .A(n40415), .B(n40416), .Z(n31099) );
  ANDN U43142 ( .B(\modmult_1/xin[1023] ), .A(n40417), .Z(n40415) );
  IV U43143 ( .A(n40416), .Z(n40417) );
  XNOR U43144 ( .A(m[176]), .B(n40418), .Z(n40416) );
  NAND U43145 ( .A(n40419), .B(mul_pow), .Z(n40418) );
  XOR U43146 ( .A(m[176]), .B(c[176]), .Z(n40419) );
  XOR U43147 ( .A(n40420), .B(n40421), .Z(n40412) );
  ANDN U43148 ( .B(n40422), .A(n31096), .Z(n40420) );
  XNOR U43149 ( .A(\modmult_1/zin[0][174] ), .B(n40423), .Z(n31096) );
  IV U43150 ( .A(n40421), .Z(n40423) );
  XOR U43151 ( .A(n40421), .B(n31097), .Z(n40422) );
  XNOR U43152 ( .A(n40424), .B(n40425), .Z(n31097) );
  ANDN U43153 ( .B(\modmult_1/xin[1023] ), .A(n40426), .Z(n40424) );
  IV U43154 ( .A(n40425), .Z(n40426) );
  XNOR U43155 ( .A(m[175]), .B(n40427), .Z(n40425) );
  NAND U43156 ( .A(n40428), .B(mul_pow), .Z(n40427) );
  XOR U43157 ( .A(m[175]), .B(c[175]), .Z(n40428) );
  XOR U43158 ( .A(n40429), .B(n40430), .Z(n40421) );
  ANDN U43159 ( .B(n40431), .A(n31094), .Z(n40429) );
  XNOR U43160 ( .A(\modmult_1/zin[0][173] ), .B(n40432), .Z(n31094) );
  IV U43161 ( .A(n40430), .Z(n40432) );
  XOR U43162 ( .A(n40430), .B(n31095), .Z(n40431) );
  XNOR U43163 ( .A(n40433), .B(n40434), .Z(n31095) );
  ANDN U43164 ( .B(\modmult_1/xin[1023] ), .A(n40435), .Z(n40433) );
  IV U43165 ( .A(n40434), .Z(n40435) );
  XNOR U43166 ( .A(m[174]), .B(n40436), .Z(n40434) );
  NAND U43167 ( .A(n40437), .B(mul_pow), .Z(n40436) );
  XOR U43168 ( .A(m[174]), .B(c[174]), .Z(n40437) );
  XOR U43169 ( .A(n40438), .B(n40439), .Z(n40430) );
  ANDN U43170 ( .B(n40440), .A(n31092), .Z(n40438) );
  XNOR U43171 ( .A(\modmult_1/zin[0][172] ), .B(n40441), .Z(n31092) );
  IV U43172 ( .A(n40439), .Z(n40441) );
  XOR U43173 ( .A(n40439), .B(n31093), .Z(n40440) );
  XNOR U43174 ( .A(n40442), .B(n40443), .Z(n31093) );
  ANDN U43175 ( .B(\modmult_1/xin[1023] ), .A(n40444), .Z(n40442) );
  IV U43176 ( .A(n40443), .Z(n40444) );
  XNOR U43177 ( .A(m[173]), .B(n40445), .Z(n40443) );
  NAND U43178 ( .A(n40446), .B(mul_pow), .Z(n40445) );
  XOR U43179 ( .A(m[173]), .B(c[173]), .Z(n40446) );
  XOR U43180 ( .A(n40447), .B(n40448), .Z(n40439) );
  ANDN U43181 ( .B(n40449), .A(n31090), .Z(n40447) );
  XNOR U43182 ( .A(\modmult_1/zin[0][171] ), .B(n40450), .Z(n31090) );
  IV U43183 ( .A(n40448), .Z(n40450) );
  XOR U43184 ( .A(n40448), .B(n31091), .Z(n40449) );
  XNOR U43185 ( .A(n40451), .B(n40452), .Z(n31091) );
  ANDN U43186 ( .B(\modmult_1/xin[1023] ), .A(n40453), .Z(n40451) );
  IV U43187 ( .A(n40452), .Z(n40453) );
  XNOR U43188 ( .A(m[172]), .B(n40454), .Z(n40452) );
  NAND U43189 ( .A(n40455), .B(mul_pow), .Z(n40454) );
  XOR U43190 ( .A(m[172]), .B(c[172]), .Z(n40455) );
  XOR U43191 ( .A(n40456), .B(n40457), .Z(n40448) );
  ANDN U43192 ( .B(n40458), .A(n31088), .Z(n40456) );
  XNOR U43193 ( .A(\modmult_1/zin[0][170] ), .B(n40459), .Z(n31088) );
  IV U43194 ( .A(n40457), .Z(n40459) );
  XOR U43195 ( .A(n40457), .B(n31089), .Z(n40458) );
  XNOR U43196 ( .A(n40460), .B(n40461), .Z(n31089) );
  ANDN U43197 ( .B(\modmult_1/xin[1023] ), .A(n40462), .Z(n40460) );
  IV U43198 ( .A(n40461), .Z(n40462) );
  XNOR U43199 ( .A(m[171]), .B(n40463), .Z(n40461) );
  NAND U43200 ( .A(n40464), .B(mul_pow), .Z(n40463) );
  XOR U43201 ( .A(m[171]), .B(c[171]), .Z(n40464) );
  XOR U43202 ( .A(n40465), .B(n40466), .Z(n40457) );
  ANDN U43203 ( .B(n40467), .A(n31086), .Z(n40465) );
  XNOR U43204 ( .A(\modmult_1/zin[0][169] ), .B(n40468), .Z(n31086) );
  IV U43205 ( .A(n40466), .Z(n40468) );
  XOR U43206 ( .A(n40466), .B(n31087), .Z(n40467) );
  XNOR U43207 ( .A(n40469), .B(n40470), .Z(n31087) );
  ANDN U43208 ( .B(\modmult_1/xin[1023] ), .A(n40471), .Z(n40469) );
  IV U43209 ( .A(n40470), .Z(n40471) );
  XNOR U43210 ( .A(m[170]), .B(n40472), .Z(n40470) );
  NAND U43211 ( .A(n40473), .B(mul_pow), .Z(n40472) );
  XOR U43212 ( .A(m[170]), .B(c[170]), .Z(n40473) );
  XOR U43213 ( .A(n40474), .B(n40475), .Z(n40466) );
  ANDN U43214 ( .B(n40476), .A(n31084), .Z(n40474) );
  XNOR U43215 ( .A(\modmult_1/zin[0][168] ), .B(n40477), .Z(n31084) );
  IV U43216 ( .A(n40475), .Z(n40477) );
  XOR U43217 ( .A(n40475), .B(n31085), .Z(n40476) );
  XNOR U43218 ( .A(n40478), .B(n40479), .Z(n31085) );
  ANDN U43219 ( .B(\modmult_1/xin[1023] ), .A(n40480), .Z(n40478) );
  IV U43220 ( .A(n40479), .Z(n40480) );
  XNOR U43221 ( .A(m[169]), .B(n40481), .Z(n40479) );
  NAND U43222 ( .A(n40482), .B(mul_pow), .Z(n40481) );
  XOR U43223 ( .A(m[169]), .B(c[169]), .Z(n40482) );
  XOR U43224 ( .A(n40483), .B(n40484), .Z(n40475) );
  ANDN U43225 ( .B(n40485), .A(n31082), .Z(n40483) );
  XNOR U43226 ( .A(\modmult_1/zin[0][167] ), .B(n40486), .Z(n31082) );
  IV U43227 ( .A(n40484), .Z(n40486) );
  XOR U43228 ( .A(n40484), .B(n31083), .Z(n40485) );
  XNOR U43229 ( .A(n40487), .B(n40488), .Z(n31083) );
  ANDN U43230 ( .B(\modmult_1/xin[1023] ), .A(n40489), .Z(n40487) );
  IV U43231 ( .A(n40488), .Z(n40489) );
  XNOR U43232 ( .A(m[168]), .B(n40490), .Z(n40488) );
  NAND U43233 ( .A(n40491), .B(mul_pow), .Z(n40490) );
  XOR U43234 ( .A(m[168]), .B(c[168]), .Z(n40491) );
  XOR U43235 ( .A(n40492), .B(n40493), .Z(n40484) );
  ANDN U43236 ( .B(n40494), .A(n31080), .Z(n40492) );
  XNOR U43237 ( .A(\modmult_1/zin[0][166] ), .B(n40495), .Z(n31080) );
  IV U43238 ( .A(n40493), .Z(n40495) );
  XOR U43239 ( .A(n40493), .B(n31081), .Z(n40494) );
  XNOR U43240 ( .A(n40496), .B(n40497), .Z(n31081) );
  ANDN U43241 ( .B(\modmult_1/xin[1023] ), .A(n40498), .Z(n40496) );
  IV U43242 ( .A(n40497), .Z(n40498) );
  XNOR U43243 ( .A(m[167]), .B(n40499), .Z(n40497) );
  NAND U43244 ( .A(n40500), .B(mul_pow), .Z(n40499) );
  XOR U43245 ( .A(m[167]), .B(c[167]), .Z(n40500) );
  XOR U43246 ( .A(n40501), .B(n40502), .Z(n40493) );
  ANDN U43247 ( .B(n40503), .A(n31078), .Z(n40501) );
  XNOR U43248 ( .A(\modmult_1/zin[0][165] ), .B(n40504), .Z(n31078) );
  IV U43249 ( .A(n40502), .Z(n40504) );
  XOR U43250 ( .A(n40502), .B(n31079), .Z(n40503) );
  XNOR U43251 ( .A(n40505), .B(n40506), .Z(n31079) );
  ANDN U43252 ( .B(\modmult_1/xin[1023] ), .A(n40507), .Z(n40505) );
  IV U43253 ( .A(n40506), .Z(n40507) );
  XNOR U43254 ( .A(m[166]), .B(n40508), .Z(n40506) );
  NAND U43255 ( .A(n40509), .B(mul_pow), .Z(n40508) );
  XOR U43256 ( .A(m[166]), .B(c[166]), .Z(n40509) );
  XOR U43257 ( .A(n40510), .B(n40511), .Z(n40502) );
  ANDN U43258 ( .B(n40512), .A(n31076), .Z(n40510) );
  XNOR U43259 ( .A(\modmult_1/zin[0][164] ), .B(n40513), .Z(n31076) );
  IV U43260 ( .A(n40511), .Z(n40513) );
  XOR U43261 ( .A(n40511), .B(n31077), .Z(n40512) );
  XNOR U43262 ( .A(n40514), .B(n40515), .Z(n31077) );
  ANDN U43263 ( .B(\modmult_1/xin[1023] ), .A(n40516), .Z(n40514) );
  IV U43264 ( .A(n40515), .Z(n40516) );
  XNOR U43265 ( .A(m[165]), .B(n40517), .Z(n40515) );
  NAND U43266 ( .A(n40518), .B(mul_pow), .Z(n40517) );
  XOR U43267 ( .A(m[165]), .B(c[165]), .Z(n40518) );
  XOR U43268 ( .A(n40519), .B(n40520), .Z(n40511) );
  ANDN U43269 ( .B(n40521), .A(n31074), .Z(n40519) );
  XNOR U43270 ( .A(\modmult_1/zin[0][163] ), .B(n40522), .Z(n31074) );
  IV U43271 ( .A(n40520), .Z(n40522) );
  XOR U43272 ( .A(n40520), .B(n31075), .Z(n40521) );
  XNOR U43273 ( .A(n40523), .B(n40524), .Z(n31075) );
  ANDN U43274 ( .B(\modmult_1/xin[1023] ), .A(n40525), .Z(n40523) );
  IV U43275 ( .A(n40524), .Z(n40525) );
  XNOR U43276 ( .A(m[164]), .B(n40526), .Z(n40524) );
  NAND U43277 ( .A(n40527), .B(mul_pow), .Z(n40526) );
  XOR U43278 ( .A(m[164]), .B(c[164]), .Z(n40527) );
  XOR U43279 ( .A(n40528), .B(n40529), .Z(n40520) );
  ANDN U43280 ( .B(n40530), .A(n31072), .Z(n40528) );
  XNOR U43281 ( .A(\modmult_1/zin[0][162] ), .B(n40531), .Z(n31072) );
  IV U43282 ( .A(n40529), .Z(n40531) );
  XOR U43283 ( .A(n40529), .B(n31073), .Z(n40530) );
  XNOR U43284 ( .A(n40532), .B(n40533), .Z(n31073) );
  ANDN U43285 ( .B(\modmult_1/xin[1023] ), .A(n40534), .Z(n40532) );
  IV U43286 ( .A(n40533), .Z(n40534) );
  XNOR U43287 ( .A(m[163]), .B(n40535), .Z(n40533) );
  NAND U43288 ( .A(n40536), .B(mul_pow), .Z(n40535) );
  XOR U43289 ( .A(m[163]), .B(c[163]), .Z(n40536) );
  XOR U43290 ( .A(n40537), .B(n40538), .Z(n40529) );
  ANDN U43291 ( .B(n40539), .A(n31070), .Z(n40537) );
  XNOR U43292 ( .A(\modmult_1/zin[0][161] ), .B(n40540), .Z(n31070) );
  IV U43293 ( .A(n40538), .Z(n40540) );
  XOR U43294 ( .A(n40538), .B(n31071), .Z(n40539) );
  XNOR U43295 ( .A(n40541), .B(n40542), .Z(n31071) );
  ANDN U43296 ( .B(\modmult_1/xin[1023] ), .A(n40543), .Z(n40541) );
  IV U43297 ( .A(n40542), .Z(n40543) );
  XNOR U43298 ( .A(m[162]), .B(n40544), .Z(n40542) );
  NAND U43299 ( .A(n40545), .B(mul_pow), .Z(n40544) );
  XOR U43300 ( .A(m[162]), .B(c[162]), .Z(n40545) );
  XOR U43301 ( .A(n40546), .B(n40547), .Z(n40538) );
  ANDN U43302 ( .B(n40548), .A(n31068), .Z(n40546) );
  XNOR U43303 ( .A(\modmult_1/zin[0][160] ), .B(n40549), .Z(n31068) );
  IV U43304 ( .A(n40547), .Z(n40549) );
  XOR U43305 ( .A(n40547), .B(n31069), .Z(n40548) );
  XNOR U43306 ( .A(n40550), .B(n40551), .Z(n31069) );
  ANDN U43307 ( .B(\modmult_1/xin[1023] ), .A(n40552), .Z(n40550) );
  IV U43308 ( .A(n40551), .Z(n40552) );
  XNOR U43309 ( .A(m[161]), .B(n40553), .Z(n40551) );
  NAND U43310 ( .A(n40554), .B(mul_pow), .Z(n40553) );
  XOR U43311 ( .A(m[161]), .B(c[161]), .Z(n40554) );
  XOR U43312 ( .A(n40555), .B(n40556), .Z(n40547) );
  ANDN U43313 ( .B(n40557), .A(n31066), .Z(n40555) );
  XNOR U43314 ( .A(\modmult_1/zin[0][159] ), .B(n40558), .Z(n31066) );
  IV U43315 ( .A(n40556), .Z(n40558) );
  XOR U43316 ( .A(n40556), .B(n31067), .Z(n40557) );
  XNOR U43317 ( .A(n40559), .B(n40560), .Z(n31067) );
  ANDN U43318 ( .B(\modmult_1/xin[1023] ), .A(n40561), .Z(n40559) );
  IV U43319 ( .A(n40560), .Z(n40561) );
  XNOR U43320 ( .A(m[160]), .B(n40562), .Z(n40560) );
  NAND U43321 ( .A(n40563), .B(mul_pow), .Z(n40562) );
  XOR U43322 ( .A(m[160]), .B(c[160]), .Z(n40563) );
  XOR U43323 ( .A(n40564), .B(n40565), .Z(n40556) );
  ANDN U43324 ( .B(n40566), .A(n31064), .Z(n40564) );
  XNOR U43325 ( .A(\modmult_1/zin[0][158] ), .B(n40567), .Z(n31064) );
  IV U43326 ( .A(n40565), .Z(n40567) );
  XOR U43327 ( .A(n40565), .B(n31065), .Z(n40566) );
  XNOR U43328 ( .A(n40568), .B(n40569), .Z(n31065) );
  ANDN U43329 ( .B(\modmult_1/xin[1023] ), .A(n40570), .Z(n40568) );
  IV U43330 ( .A(n40569), .Z(n40570) );
  XNOR U43331 ( .A(m[159]), .B(n40571), .Z(n40569) );
  NAND U43332 ( .A(n40572), .B(mul_pow), .Z(n40571) );
  XOR U43333 ( .A(m[159]), .B(c[159]), .Z(n40572) );
  XOR U43334 ( .A(n40573), .B(n40574), .Z(n40565) );
  ANDN U43335 ( .B(n40575), .A(n31062), .Z(n40573) );
  XNOR U43336 ( .A(\modmult_1/zin[0][157] ), .B(n40576), .Z(n31062) );
  IV U43337 ( .A(n40574), .Z(n40576) );
  XOR U43338 ( .A(n40574), .B(n31063), .Z(n40575) );
  XNOR U43339 ( .A(n40577), .B(n40578), .Z(n31063) );
  ANDN U43340 ( .B(\modmult_1/xin[1023] ), .A(n40579), .Z(n40577) );
  IV U43341 ( .A(n40578), .Z(n40579) );
  XNOR U43342 ( .A(m[158]), .B(n40580), .Z(n40578) );
  NAND U43343 ( .A(n40581), .B(mul_pow), .Z(n40580) );
  XOR U43344 ( .A(m[158]), .B(c[158]), .Z(n40581) );
  XOR U43345 ( .A(n40582), .B(n40583), .Z(n40574) );
  ANDN U43346 ( .B(n40584), .A(n31060), .Z(n40582) );
  XNOR U43347 ( .A(\modmult_1/zin[0][156] ), .B(n40585), .Z(n31060) );
  IV U43348 ( .A(n40583), .Z(n40585) );
  XOR U43349 ( .A(n40583), .B(n31061), .Z(n40584) );
  XNOR U43350 ( .A(n40586), .B(n40587), .Z(n31061) );
  ANDN U43351 ( .B(\modmult_1/xin[1023] ), .A(n40588), .Z(n40586) );
  IV U43352 ( .A(n40587), .Z(n40588) );
  XNOR U43353 ( .A(m[157]), .B(n40589), .Z(n40587) );
  NAND U43354 ( .A(n40590), .B(mul_pow), .Z(n40589) );
  XOR U43355 ( .A(m[157]), .B(c[157]), .Z(n40590) );
  XOR U43356 ( .A(n40591), .B(n40592), .Z(n40583) );
  ANDN U43357 ( .B(n40593), .A(n31058), .Z(n40591) );
  XNOR U43358 ( .A(\modmult_1/zin[0][155] ), .B(n40594), .Z(n31058) );
  IV U43359 ( .A(n40592), .Z(n40594) );
  XOR U43360 ( .A(n40592), .B(n31059), .Z(n40593) );
  XNOR U43361 ( .A(n40595), .B(n40596), .Z(n31059) );
  ANDN U43362 ( .B(\modmult_1/xin[1023] ), .A(n40597), .Z(n40595) );
  IV U43363 ( .A(n40596), .Z(n40597) );
  XNOR U43364 ( .A(m[156]), .B(n40598), .Z(n40596) );
  NAND U43365 ( .A(n40599), .B(mul_pow), .Z(n40598) );
  XOR U43366 ( .A(m[156]), .B(c[156]), .Z(n40599) );
  XOR U43367 ( .A(n40600), .B(n40601), .Z(n40592) );
  ANDN U43368 ( .B(n40602), .A(n31056), .Z(n40600) );
  XNOR U43369 ( .A(\modmult_1/zin[0][154] ), .B(n40603), .Z(n31056) );
  IV U43370 ( .A(n40601), .Z(n40603) );
  XOR U43371 ( .A(n40601), .B(n31057), .Z(n40602) );
  XNOR U43372 ( .A(n40604), .B(n40605), .Z(n31057) );
  ANDN U43373 ( .B(\modmult_1/xin[1023] ), .A(n40606), .Z(n40604) );
  IV U43374 ( .A(n40605), .Z(n40606) );
  XNOR U43375 ( .A(m[155]), .B(n40607), .Z(n40605) );
  NAND U43376 ( .A(n40608), .B(mul_pow), .Z(n40607) );
  XOR U43377 ( .A(m[155]), .B(c[155]), .Z(n40608) );
  XOR U43378 ( .A(n40609), .B(n40610), .Z(n40601) );
  ANDN U43379 ( .B(n40611), .A(n31054), .Z(n40609) );
  XNOR U43380 ( .A(\modmult_1/zin[0][153] ), .B(n40612), .Z(n31054) );
  IV U43381 ( .A(n40610), .Z(n40612) );
  XOR U43382 ( .A(n40610), .B(n31055), .Z(n40611) );
  XNOR U43383 ( .A(n40613), .B(n40614), .Z(n31055) );
  ANDN U43384 ( .B(\modmult_1/xin[1023] ), .A(n40615), .Z(n40613) );
  IV U43385 ( .A(n40614), .Z(n40615) );
  XNOR U43386 ( .A(m[154]), .B(n40616), .Z(n40614) );
  NAND U43387 ( .A(n40617), .B(mul_pow), .Z(n40616) );
  XOR U43388 ( .A(m[154]), .B(c[154]), .Z(n40617) );
  XOR U43389 ( .A(n40618), .B(n40619), .Z(n40610) );
  ANDN U43390 ( .B(n40620), .A(n31052), .Z(n40618) );
  XNOR U43391 ( .A(\modmult_1/zin[0][152] ), .B(n40621), .Z(n31052) );
  IV U43392 ( .A(n40619), .Z(n40621) );
  XOR U43393 ( .A(n40619), .B(n31053), .Z(n40620) );
  XNOR U43394 ( .A(n40622), .B(n40623), .Z(n31053) );
  ANDN U43395 ( .B(\modmult_1/xin[1023] ), .A(n40624), .Z(n40622) );
  IV U43396 ( .A(n40623), .Z(n40624) );
  XNOR U43397 ( .A(m[153]), .B(n40625), .Z(n40623) );
  NAND U43398 ( .A(n40626), .B(mul_pow), .Z(n40625) );
  XOR U43399 ( .A(m[153]), .B(c[153]), .Z(n40626) );
  XOR U43400 ( .A(n40627), .B(n40628), .Z(n40619) );
  ANDN U43401 ( .B(n40629), .A(n31050), .Z(n40627) );
  XNOR U43402 ( .A(\modmult_1/zin[0][151] ), .B(n40630), .Z(n31050) );
  IV U43403 ( .A(n40628), .Z(n40630) );
  XOR U43404 ( .A(n40628), .B(n31051), .Z(n40629) );
  XNOR U43405 ( .A(n40631), .B(n40632), .Z(n31051) );
  ANDN U43406 ( .B(\modmult_1/xin[1023] ), .A(n40633), .Z(n40631) );
  IV U43407 ( .A(n40632), .Z(n40633) );
  XNOR U43408 ( .A(m[152]), .B(n40634), .Z(n40632) );
  NAND U43409 ( .A(n40635), .B(mul_pow), .Z(n40634) );
  XOR U43410 ( .A(m[152]), .B(c[152]), .Z(n40635) );
  XOR U43411 ( .A(n40636), .B(n40637), .Z(n40628) );
  ANDN U43412 ( .B(n40638), .A(n31048), .Z(n40636) );
  XNOR U43413 ( .A(\modmult_1/zin[0][150] ), .B(n40639), .Z(n31048) );
  IV U43414 ( .A(n40637), .Z(n40639) );
  XOR U43415 ( .A(n40637), .B(n31049), .Z(n40638) );
  XNOR U43416 ( .A(n40640), .B(n40641), .Z(n31049) );
  ANDN U43417 ( .B(\modmult_1/xin[1023] ), .A(n40642), .Z(n40640) );
  IV U43418 ( .A(n40641), .Z(n40642) );
  XNOR U43419 ( .A(m[151]), .B(n40643), .Z(n40641) );
  NAND U43420 ( .A(n40644), .B(mul_pow), .Z(n40643) );
  XOR U43421 ( .A(m[151]), .B(c[151]), .Z(n40644) );
  XOR U43422 ( .A(n40645), .B(n40646), .Z(n40637) );
  ANDN U43423 ( .B(n40647), .A(n31046), .Z(n40645) );
  XNOR U43424 ( .A(\modmult_1/zin[0][149] ), .B(n40648), .Z(n31046) );
  IV U43425 ( .A(n40646), .Z(n40648) );
  XOR U43426 ( .A(n40646), .B(n31047), .Z(n40647) );
  XNOR U43427 ( .A(n40649), .B(n40650), .Z(n31047) );
  ANDN U43428 ( .B(\modmult_1/xin[1023] ), .A(n40651), .Z(n40649) );
  IV U43429 ( .A(n40650), .Z(n40651) );
  XNOR U43430 ( .A(m[150]), .B(n40652), .Z(n40650) );
  NAND U43431 ( .A(n40653), .B(mul_pow), .Z(n40652) );
  XOR U43432 ( .A(m[150]), .B(c[150]), .Z(n40653) );
  XOR U43433 ( .A(n40654), .B(n40655), .Z(n40646) );
  ANDN U43434 ( .B(n40656), .A(n31044), .Z(n40654) );
  XNOR U43435 ( .A(\modmult_1/zin[0][148] ), .B(n40657), .Z(n31044) );
  IV U43436 ( .A(n40655), .Z(n40657) );
  XOR U43437 ( .A(n40655), .B(n31045), .Z(n40656) );
  XNOR U43438 ( .A(n40658), .B(n40659), .Z(n31045) );
  ANDN U43439 ( .B(\modmult_1/xin[1023] ), .A(n40660), .Z(n40658) );
  IV U43440 ( .A(n40659), .Z(n40660) );
  XNOR U43441 ( .A(m[149]), .B(n40661), .Z(n40659) );
  NAND U43442 ( .A(n40662), .B(mul_pow), .Z(n40661) );
  XOR U43443 ( .A(m[149]), .B(c[149]), .Z(n40662) );
  XOR U43444 ( .A(n40663), .B(n40664), .Z(n40655) );
  ANDN U43445 ( .B(n40665), .A(n31042), .Z(n40663) );
  XNOR U43446 ( .A(\modmult_1/zin[0][147] ), .B(n40666), .Z(n31042) );
  IV U43447 ( .A(n40664), .Z(n40666) );
  XOR U43448 ( .A(n40664), .B(n31043), .Z(n40665) );
  XNOR U43449 ( .A(n40667), .B(n40668), .Z(n31043) );
  ANDN U43450 ( .B(\modmult_1/xin[1023] ), .A(n40669), .Z(n40667) );
  IV U43451 ( .A(n40668), .Z(n40669) );
  XNOR U43452 ( .A(m[148]), .B(n40670), .Z(n40668) );
  NAND U43453 ( .A(n40671), .B(mul_pow), .Z(n40670) );
  XOR U43454 ( .A(m[148]), .B(c[148]), .Z(n40671) );
  XOR U43455 ( .A(n40672), .B(n40673), .Z(n40664) );
  ANDN U43456 ( .B(n40674), .A(n31040), .Z(n40672) );
  XNOR U43457 ( .A(\modmult_1/zin[0][146] ), .B(n40675), .Z(n31040) );
  IV U43458 ( .A(n40673), .Z(n40675) );
  XOR U43459 ( .A(n40673), .B(n31041), .Z(n40674) );
  XNOR U43460 ( .A(n40676), .B(n40677), .Z(n31041) );
  ANDN U43461 ( .B(\modmult_1/xin[1023] ), .A(n40678), .Z(n40676) );
  IV U43462 ( .A(n40677), .Z(n40678) );
  XNOR U43463 ( .A(m[147]), .B(n40679), .Z(n40677) );
  NAND U43464 ( .A(n40680), .B(mul_pow), .Z(n40679) );
  XOR U43465 ( .A(m[147]), .B(c[147]), .Z(n40680) );
  XOR U43466 ( .A(n40681), .B(n40682), .Z(n40673) );
  ANDN U43467 ( .B(n40683), .A(n31038), .Z(n40681) );
  XNOR U43468 ( .A(\modmult_1/zin[0][145] ), .B(n40684), .Z(n31038) );
  IV U43469 ( .A(n40682), .Z(n40684) );
  XOR U43470 ( .A(n40682), .B(n31039), .Z(n40683) );
  XNOR U43471 ( .A(n40685), .B(n40686), .Z(n31039) );
  ANDN U43472 ( .B(\modmult_1/xin[1023] ), .A(n40687), .Z(n40685) );
  IV U43473 ( .A(n40686), .Z(n40687) );
  XNOR U43474 ( .A(m[146]), .B(n40688), .Z(n40686) );
  NAND U43475 ( .A(n40689), .B(mul_pow), .Z(n40688) );
  XOR U43476 ( .A(m[146]), .B(c[146]), .Z(n40689) );
  XOR U43477 ( .A(n40690), .B(n40691), .Z(n40682) );
  ANDN U43478 ( .B(n40692), .A(n31036), .Z(n40690) );
  XNOR U43479 ( .A(\modmult_1/zin[0][144] ), .B(n40693), .Z(n31036) );
  IV U43480 ( .A(n40691), .Z(n40693) );
  XOR U43481 ( .A(n40691), .B(n31037), .Z(n40692) );
  XNOR U43482 ( .A(n40694), .B(n40695), .Z(n31037) );
  ANDN U43483 ( .B(\modmult_1/xin[1023] ), .A(n40696), .Z(n40694) );
  IV U43484 ( .A(n40695), .Z(n40696) );
  XNOR U43485 ( .A(m[145]), .B(n40697), .Z(n40695) );
  NAND U43486 ( .A(n40698), .B(mul_pow), .Z(n40697) );
  XOR U43487 ( .A(m[145]), .B(c[145]), .Z(n40698) );
  XOR U43488 ( .A(n40699), .B(n40700), .Z(n40691) );
  ANDN U43489 ( .B(n40701), .A(n31034), .Z(n40699) );
  XNOR U43490 ( .A(\modmult_1/zin[0][143] ), .B(n40702), .Z(n31034) );
  IV U43491 ( .A(n40700), .Z(n40702) );
  XOR U43492 ( .A(n40700), .B(n31035), .Z(n40701) );
  XNOR U43493 ( .A(n40703), .B(n40704), .Z(n31035) );
  ANDN U43494 ( .B(\modmult_1/xin[1023] ), .A(n40705), .Z(n40703) );
  IV U43495 ( .A(n40704), .Z(n40705) );
  XNOR U43496 ( .A(m[144]), .B(n40706), .Z(n40704) );
  NAND U43497 ( .A(n40707), .B(mul_pow), .Z(n40706) );
  XOR U43498 ( .A(m[144]), .B(c[144]), .Z(n40707) );
  XOR U43499 ( .A(n40708), .B(n40709), .Z(n40700) );
  ANDN U43500 ( .B(n40710), .A(n31032), .Z(n40708) );
  XNOR U43501 ( .A(\modmult_1/zin[0][142] ), .B(n40711), .Z(n31032) );
  IV U43502 ( .A(n40709), .Z(n40711) );
  XOR U43503 ( .A(n40709), .B(n31033), .Z(n40710) );
  XNOR U43504 ( .A(n40712), .B(n40713), .Z(n31033) );
  ANDN U43505 ( .B(\modmult_1/xin[1023] ), .A(n40714), .Z(n40712) );
  IV U43506 ( .A(n40713), .Z(n40714) );
  XNOR U43507 ( .A(m[143]), .B(n40715), .Z(n40713) );
  NAND U43508 ( .A(n40716), .B(mul_pow), .Z(n40715) );
  XOR U43509 ( .A(m[143]), .B(c[143]), .Z(n40716) );
  XOR U43510 ( .A(n40717), .B(n40718), .Z(n40709) );
  ANDN U43511 ( .B(n40719), .A(n31030), .Z(n40717) );
  XNOR U43512 ( .A(\modmult_1/zin[0][141] ), .B(n40720), .Z(n31030) );
  IV U43513 ( .A(n40718), .Z(n40720) );
  XOR U43514 ( .A(n40718), .B(n31031), .Z(n40719) );
  XNOR U43515 ( .A(n40721), .B(n40722), .Z(n31031) );
  ANDN U43516 ( .B(\modmult_1/xin[1023] ), .A(n40723), .Z(n40721) );
  IV U43517 ( .A(n40722), .Z(n40723) );
  XNOR U43518 ( .A(m[142]), .B(n40724), .Z(n40722) );
  NAND U43519 ( .A(n40725), .B(mul_pow), .Z(n40724) );
  XOR U43520 ( .A(m[142]), .B(c[142]), .Z(n40725) );
  XOR U43521 ( .A(n40726), .B(n40727), .Z(n40718) );
  ANDN U43522 ( .B(n40728), .A(n31028), .Z(n40726) );
  XNOR U43523 ( .A(\modmult_1/zin[0][140] ), .B(n40729), .Z(n31028) );
  IV U43524 ( .A(n40727), .Z(n40729) );
  XOR U43525 ( .A(n40727), .B(n31029), .Z(n40728) );
  XNOR U43526 ( .A(n40730), .B(n40731), .Z(n31029) );
  ANDN U43527 ( .B(\modmult_1/xin[1023] ), .A(n40732), .Z(n40730) );
  IV U43528 ( .A(n40731), .Z(n40732) );
  XNOR U43529 ( .A(m[141]), .B(n40733), .Z(n40731) );
  NAND U43530 ( .A(n40734), .B(mul_pow), .Z(n40733) );
  XOR U43531 ( .A(m[141]), .B(c[141]), .Z(n40734) );
  XOR U43532 ( .A(n40735), .B(n40736), .Z(n40727) );
  ANDN U43533 ( .B(n40737), .A(n31026), .Z(n40735) );
  XNOR U43534 ( .A(\modmult_1/zin[0][139] ), .B(n40738), .Z(n31026) );
  IV U43535 ( .A(n40736), .Z(n40738) );
  XOR U43536 ( .A(n40736), .B(n31027), .Z(n40737) );
  XNOR U43537 ( .A(n40739), .B(n40740), .Z(n31027) );
  ANDN U43538 ( .B(\modmult_1/xin[1023] ), .A(n40741), .Z(n40739) );
  IV U43539 ( .A(n40740), .Z(n40741) );
  XNOR U43540 ( .A(m[140]), .B(n40742), .Z(n40740) );
  NAND U43541 ( .A(n40743), .B(mul_pow), .Z(n40742) );
  XOR U43542 ( .A(m[140]), .B(c[140]), .Z(n40743) );
  XOR U43543 ( .A(n40744), .B(n40745), .Z(n40736) );
  ANDN U43544 ( .B(n40746), .A(n31024), .Z(n40744) );
  XNOR U43545 ( .A(\modmult_1/zin[0][138] ), .B(n40747), .Z(n31024) );
  IV U43546 ( .A(n40745), .Z(n40747) );
  XOR U43547 ( .A(n40745), .B(n31025), .Z(n40746) );
  XNOR U43548 ( .A(n40748), .B(n40749), .Z(n31025) );
  ANDN U43549 ( .B(\modmult_1/xin[1023] ), .A(n40750), .Z(n40748) );
  IV U43550 ( .A(n40749), .Z(n40750) );
  XNOR U43551 ( .A(m[139]), .B(n40751), .Z(n40749) );
  NAND U43552 ( .A(n40752), .B(mul_pow), .Z(n40751) );
  XOR U43553 ( .A(m[139]), .B(c[139]), .Z(n40752) );
  XOR U43554 ( .A(n40753), .B(n40754), .Z(n40745) );
  ANDN U43555 ( .B(n40755), .A(n31022), .Z(n40753) );
  XNOR U43556 ( .A(\modmult_1/zin[0][137] ), .B(n40756), .Z(n31022) );
  IV U43557 ( .A(n40754), .Z(n40756) );
  XOR U43558 ( .A(n40754), .B(n31023), .Z(n40755) );
  XNOR U43559 ( .A(n40757), .B(n40758), .Z(n31023) );
  ANDN U43560 ( .B(\modmult_1/xin[1023] ), .A(n40759), .Z(n40757) );
  IV U43561 ( .A(n40758), .Z(n40759) );
  XNOR U43562 ( .A(m[138]), .B(n40760), .Z(n40758) );
  NAND U43563 ( .A(n40761), .B(mul_pow), .Z(n40760) );
  XOR U43564 ( .A(m[138]), .B(c[138]), .Z(n40761) );
  XOR U43565 ( .A(n40762), .B(n40763), .Z(n40754) );
  ANDN U43566 ( .B(n40764), .A(n31020), .Z(n40762) );
  XNOR U43567 ( .A(\modmult_1/zin[0][136] ), .B(n40765), .Z(n31020) );
  IV U43568 ( .A(n40763), .Z(n40765) );
  XOR U43569 ( .A(n40763), .B(n31021), .Z(n40764) );
  XNOR U43570 ( .A(n40766), .B(n40767), .Z(n31021) );
  ANDN U43571 ( .B(\modmult_1/xin[1023] ), .A(n40768), .Z(n40766) );
  IV U43572 ( .A(n40767), .Z(n40768) );
  XNOR U43573 ( .A(m[137]), .B(n40769), .Z(n40767) );
  NAND U43574 ( .A(n40770), .B(mul_pow), .Z(n40769) );
  XOR U43575 ( .A(m[137]), .B(c[137]), .Z(n40770) );
  XOR U43576 ( .A(n40771), .B(n40772), .Z(n40763) );
  ANDN U43577 ( .B(n40773), .A(n31018), .Z(n40771) );
  XNOR U43578 ( .A(\modmult_1/zin[0][135] ), .B(n40774), .Z(n31018) );
  IV U43579 ( .A(n40772), .Z(n40774) );
  XOR U43580 ( .A(n40772), .B(n31019), .Z(n40773) );
  XNOR U43581 ( .A(n40775), .B(n40776), .Z(n31019) );
  ANDN U43582 ( .B(\modmult_1/xin[1023] ), .A(n40777), .Z(n40775) );
  IV U43583 ( .A(n40776), .Z(n40777) );
  XNOR U43584 ( .A(m[136]), .B(n40778), .Z(n40776) );
  NAND U43585 ( .A(n40779), .B(mul_pow), .Z(n40778) );
  XOR U43586 ( .A(m[136]), .B(c[136]), .Z(n40779) );
  XOR U43587 ( .A(n40780), .B(n40781), .Z(n40772) );
  ANDN U43588 ( .B(n40782), .A(n31016), .Z(n40780) );
  XNOR U43589 ( .A(\modmult_1/zin[0][134] ), .B(n40783), .Z(n31016) );
  IV U43590 ( .A(n40781), .Z(n40783) );
  XOR U43591 ( .A(n40781), .B(n31017), .Z(n40782) );
  XNOR U43592 ( .A(n40784), .B(n40785), .Z(n31017) );
  ANDN U43593 ( .B(\modmult_1/xin[1023] ), .A(n40786), .Z(n40784) );
  IV U43594 ( .A(n40785), .Z(n40786) );
  XNOR U43595 ( .A(m[135]), .B(n40787), .Z(n40785) );
  NAND U43596 ( .A(n40788), .B(mul_pow), .Z(n40787) );
  XOR U43597 ( .A(m[135]), .B(c[135]), .Z(n40788) );
  XOR U43598 ( .A(n40789), .B(n40790), .Z(n40781) );
  ANDN U43599 ( .B(n40791), .A(n31014), .Z(n40789) );
  XNOR U43600 ( .A(\modmult_1/zin[0][133] ), .B(n40792), .Z(n31014) );
  IV U43601 ( .A(n40790), .Z(n40792) );
  XOR U43602 ( .A(n40790), .B(n31015), .Z(n40791) );
  XNOR U43603 ( .A(n40793), .B(n40794), .Z(n31015) );
  ANDN U43604 ( .B(\modmult_1/xin[1023] ), .A(n40795), .Z(n40793) );
  IV U43605 ( .A(n40794), .Z(n40795) );
  XNOR U43606 ( .A(m[134]), .B(n40796), .Z(n40794) );
  NAND U43607 ( .A(n40797), .B(mul_pow), .Z(n40796) );
  XOR U43608 ( .A(m[134]), .B(c[134]), .Z(n40797) );
  XOR U43609 ( .A(n40798), .B(n40799), .Z(n40790) );
  ANDN U43610 ( .B(n40800), .A(n31012), .Z(n40798) );
  XNOR U43611 ( .A(\modmult_1/zin[0][132] ), .B(n40801), .Z(n31012) );
  IV U43612 ( .A(n40799), .Z(n40801) );
  XOR U43613 ( .A(n40799), .B(n31013), .Z(n40800) );
  XNOR U43614 ( .A(n40802), .B(n40803), .Z(n31013) );
  ANDN U43615 ( .B(\modmult_1/xin[1023] ), .A(n40804), .Z(n40802) );
  IV U43616 ( .A(n40803), .Z(n40804) );
  XNOR U43617 ( .A(m[133]), .B(n40805), .Z(n40803) );
  NAND U43618 ( .A(n40806), .B(mul_pow), .Z(n40805) );
  XOR U43619 ( .A(m[133]), .B(c[133]), .Z(n40806) );
  XOR U43620 ( .A(n40807), .B(n40808), .Z(n40799) );
  ANDN U43621 ( .B(n40809), .A(n31010), .Z(n40807) );
  XNOR U43622 ( .A(\modmult_1/zin[0][131] ), .B(n40810), .Z(n31010) );
  IV U43623 ( .A(n40808), .Z(n40810) );
  XOR U43624 ( .A(n40808), .B(n31011), .Z(n40809) );
  XNOR U43625 ( .A(n40811), .B(n40812), .Z(n31011) );
  ANDN U43626 ( .B(\modmult_1/xin[1023] ), .A(n40813), .Z(n40811) );
  IV U43627 ( .A(n40812), .Z(n40813) );
  XNOR U43628 ( .A(m[132]), .B(n40814), .Z(n40812) );
  NAND U43629 ( .A(n40815), .B(mul_pow), .Z(n40814) );
  XOR U43630 ( .A(m[132]), .B(c[132]), .Z(n40815) );
  XOR U43631 ( .A(n40816), .B(n40817), .Z(n40808) );
  ANDN U43632 ( .B(n40818), .A(n31008), .Z(n40816) );
  XNOR U43633 ( .A(\modmult_1/zin[0][130] ), .B(n40819), .Z(n31008) );
  IV U43634 ( .A(n40817), .Z(n40819) );
  XOR U43635 ( .A(n40817), .B(n31009), .Z(n40818) );
  XNOR U43636 ( .A(n40820), .B(n40821), .Z(n31009) );
  ANDN U43637 ( .B(\modmult_1/xin[1023] ), .A(n40822), .Z(n40820) );
  IV U43638 ( .A(n40821), .Z(n40822) );
  XNOR U43639 ( .A(m[131]), .B(n40823), .Z(n40821) );
  NAND U43640 ( .A(n40824), .B(mul_pow), .Z(n40823) );
  XOR U43641 ( .A(m[131]), .B(c[131]), .Z(n40824) );
  XOR U43642 ( .A(n40825), .B(n40826), .Z(n40817) );
  ANDN U43643 ( .B(n40827), .A(n31006), .Z(n40825) );
  XNOR U43644 ( .A(\modmult_1/zin[0][129] ), .B(n40828), .Z(n31006) );
  IV U43645 ( .A(n40826), .Z(n40828) );
  XOR U43646 ( .A(n40826), .B(n31007), .Z(n40827) );
  XNOR U43647 ( .A(n40829), .B(n40830), .Z(n31007) );
  ANDN U43648 ( .B(\modmult_1/xin[1023] ), .A(n40831), .Z(n40829) );
  IV U43649 ( .A(n40830), .Z(n40831) );
  XNOR U43650 ( .A(m[130]), .B(n40832), .Z(n40830) );
  NAND U43651 ( .A(n40833), .B(mul_pow), .Z(n40832) );
  XOR U43652 ( .A(m[130]), .B(c[130]), .Z(n40833) );
  XOR U43653 ( .A(n40834), .B(n40835), .Z(n40826) );
  ANDN U43654 ( .B(n40836), .A(n31004), .Z(n40834) );
  XNOR U43655 ( .A(\modmult_1/zin[0][128] ), .B(n40837), .Z(n31004) );
  IV U43656 ( .A(n40835), .Z(n40837) );
  XOR U43657 ( .A(n40835), .B(n31005), .Z(n40836) );
  XNOR U43658 ( .A(n40838), .B(n40839), .Z(n31005) );
  ANDN U43659 ( .B(\modmult_1/xin[1023] ), .A(n40840), .Z(n40838) );
  IV U43660 ( .A(n40839), .Z(n40840) );
  XNOR U43661 ( .A(m[129]), .B(n40841), .Z(n40839) );
  NAND U43662 ( .A(n40842), .B(mul_pow), .Z(n40841) );
  XOR U43663 ( .A(m[129]), .B(c[129]), .Z(n40842) );
  XOR U43664 ( .A(n40843), .B(n40844), .Z(n40835) );
  ANDN U43665 ( .B(n40845), .A(n31002), .Z(n40843) );
  XNOR U43666 ( .A(\modmult_1/zin[0][127] ), .B(n40846), .Z(n31002) );
  IV U43667 ( .A(n40844), .Z(n40846) );
  XOR U43668 ( .A(n40844), .B(n31003), .Z(n40845) );
  XNOR U43669 ( .A(n40847), .B(n40848), .Z(n31003) );
  ANDN U43670 ( .B(\modmult_1/xin[1023] ), .A(n40849), .Z(n40847) );
  IV U43671 ( .A(n40848), .Z(n40849) );
  XNOR U43672 ( .A(m[128]), .B(n40850), .Z(n40848) );
  NAND U43673 ( .A(n40851), .B(mul_pow), .Z(n40850) );
  XOR U43674 ( .A(m[128]), .B(c[128]), .Z(n40851) );
  XOR U43675 ( .A(n40852), .B(n40853), .Z(n40844) );
  ANDN U43676 ( .B(n40854), .A(n31000), .Z(n40852) );
  XNOR U43677 ( .A(\modmult_1/zin[0][126] ), .B(n40855), .Z(n31000) );
  IV U43678 ( .A(n40853), .Z(n40855) );
  XOR U43679 ( .A(n40853), .B(n31001), .Z(n40854) );
  XNOR U43680 ( .A(n40856), .B(n40857), .Z(n31001) );
  ANDN U43681 ( .B(\modmult_1/xin[1023] ), .A(n40858), .Z(n40856) );
  IV U43682 ( .A(n40857), .Z(n40858) );
  XNOR U43683 ( .A(m[127]), .B(n40859), .Z(n40857) );
  NAND U43684 ( .A(n40860), .B(mul_pow), .Z(n40859) );
  XOR U43685 ( .A(m[127]), .B(c[127]), .Z(n40860) );
  XOR U43686 ( .A(n40861), .B(n40862), .Z(n40853) );
  ANDN U43687 ( .B(n40863), .A(n30998), .Z(n40861) );
  XNOR U43688 ( .A(\modmult_1/zin[0][125] ), .B(n40864), .Z(n30998) );
  IV U43689 ( .A(n40862), .Z(n40864) );
  XOR U43690 ( .A(n40862), .B(n30999), .Z(n40863) );
  XNOR U43691 ( .A(n40865), .B(n40866), .Z(n30999) );
  ANDN U43692 ( .B(\modmult_1/xin[1023] ), .A(n40867), .Z(n40865) );
  IV U43693 ( .A(n40866), .Z(n40867) );
  XNOR U43694 ( .A(m[126]), .B(n40868), .Z(n40866) );
  NAND U43695 ( .A(n40869), .B(mul_pow), .Z(n40868) );
  XOR U43696 ( .A(m[126]), .B(c[126]), .Z(n40869) );
  XOR U43697 ( .A(n40870), .B(n40871), .Z(n40862) );
  ANDN U43698 ( .B(n40872), .A(n30996), .Z(n40870) );
  XNOR U43699 ( .A(\modmult_1/zin[0][124] ), .B(n40873), .Z(n30996) );
  IV U43700 ( .A(n40871), .Z(n40873) );
  XOR U43701 ( .A(n40871), .B(n30997), .Z(n40872) );
  XNOR U43702 ( .A(n40874), .B(n40875), .Z(n30997) );
  ANDN U43703 ( .B(\modmult_1/xin[1023] ), .A(n40876), .Z(n40874) );
  IV U43704 ( .A(n40875), .Z(n40876) );
  XNOR U43705 ( .A(m[125]), .B(n40877), .Z(n40875) );
  NAND U43706 ( .A(n40878), .B(mul_pow), .Z(n40877) );
  XOR U43707 ( .A(m[125]), .B(c[125]), .Z(n40878) );
  XOR U43708 ( .A(n40879), .B(n40880), .Z(n40871) );
  ANDN U43709 ( .B(n40881), .A(n30994), .Z(n40879) );
  XNOR U43710 ( .A(\modmult_1/zin[0][123] ), .B(n40882), .Z(n30994) );
  IV U43711 ( .A(n40880), .Z(n40882) );
  XOR U43712 ( .A(n40880), .B(n30995), .Z(n40881) );
  XNOR U43713 ( .A(n40883), .B(n40884), .Z(n30995) );
  ANDN U43714 ( .B(\modmult_1/xin[1023] ), .A(n40885), .Z(n40883) );
  IV U43715 ( .A(n40884), .Z(n40885) );
  XNOR U43716 ( .A(m[124]), .B(n40886), .Z(n40884) );
  NAND U43717 ( .A(n40887), .B(mul_pow), .Z(n40886) );
  XOR U43718 ( .A(m[124]), .B(c[124]), .Z(n40887) );
  XOR U43719 ( .A(n40888), .B(n40889), .Z(n40880) );
  ANDN U43720 ( .B(n40890), .A(n30992), .Z(n40888) );
  XNOR U43721 ( .A(\modmult_1/zin[0][122] ), .B(n40891), .Z(n30992) );
  IV U43722 ( .A(n40889), .Z(n40891) );
  XOR U43723 ( .A(n40889), .B(n30993), .Z(n40890) );
  XNOR U43724 ( .A(n40892), .B(n40893), .Z(n30993) );
  ANDN U43725 ( .B(\modmult_1/xin[1023] ), .A(n40894), .Z(n40892) );
  IV U43726 ( .A(n40893), .Z(n40894) );
  XNOR U43727 ( .A(m[123]), .B(n40895), .Z(n40893) );
  NAND U43728 ( .A(n40896), .B(mul_pow), .Z(n40895) );
  XOR U43729 ( .A(m[123]), .B(c[123]), .Z(n40896) );
  XOR U43730 ( .A(n40897), .B(n40898), .Z(n40889) );
  ANDN U43731 ( .B(n40899), .A(n30990), .Z(n40897) );
  XNOR U43732 ( .A(\modmult_1/zin[0][121] ), .B(n40900), .Z(n30990) );
  IV U43733 ( .A(n40898), .Z(n40900) );
  XOR U43734 ( .A(n40898), .B(n30991), .Z(n40899) );
  XNOR U43735 ( .A(n40901), .B(n40902), .Z(n30991) );
  ANDN U43736 ( .B(\modmult_1/xin[1023] ), .A(n40903), .Z(n40901) );
  IV U43737 ( .A(n40902), .Z(n40903) );
  XNOR U43738 ( .A(m[122]), .B(n40904), .Z(n40902) );
  NAND U43739 ( .A(n40905), .B(mul_pow), .Z(n40904) );
  XOR U43740 ( .A(m[122]), .B(c[122]), .Z(n40905) );
  XOR U43741 ( .A(n40906), .B(n40907), .Z(n40898) );
  ANDN U43742 ( .B(n40908), .A(n30988), .Z(n40906) );
  XNOR U43743 ( .A(\modmult_1/zin[0][120] ), .B(n40909), .Z(n30988) );
  IV U43744 ( .A(n40907), .Z(n40909) );
  XOR U43745 ( .A(n40907), .B(n30989), .Z(n40908) );
  XNOR U43746 ( .A(n40910), .B(n40911), .Z(n30989) );
  ANDN U43747 ( .B(\modmult_1/xin[1023] ), .A(n40912), .Z(n40910) );
  IV U43748 ( .A(n40911), .Z(n40912) );
  XNOR U43749 ( .A(m[121]), .B(n40913), .Z(n40911) );
  NAND U43750 ( .A(n40914), .B(mul_pow), .Z(n40913) );
  XOR U43751 ( .A(m[121]), .B(c[121]), .Z(n40914) );
  XOR U43752 ( .A(n40915), .B(n40916), .Z(n40907) );
  ANDN U43753 ( .B(n40917), .A(n30986), .Z(n40915) );
  XNOR U43754 ( .A(\modmult_1/zin[0][119] ), .B(n40918), .Z(n30986) );
  IV U43755 ( .A(n40916), .Z(n40918) );
  XOR U43756 ( .A(n40916), .B(n30987), .Z(n40917) );
  XNOR U43757 ( .A(n40919), .B(n40920), .Z(n30987) );
  ANDN U43758 ( .B(\modmult_1/xin[1023] ), .A(n40921), .Z(n40919) );
  IV U43759 ( .A(n40920), .Z(n40921) );
  XNOR U43760 ( .A(m[120]), .B(n40922), .Z(n40920) );
  NAND U43761 ( .A(n40923), .B(mul_pow), .Z(n40922) );
  XOR U43762 ( .A(m[120]), .B(c[120]), .Z(n40923) );
  XOR U43763 ( .A(n40924), .B(n40925), .Z(n40916) );
  ANDN U43764 ( .B(n40926), .A(n30984), .Z(n40924) );
  XNOR U43765 ( .A(\modmult_1/zin[0][118] ), .B(n40927), .Z(n30984) );
  IV U43766 ( .A(n40925), .Z(n40927) );
  XOR U43767 ( .A(n40925), .B(n30985), .Z(n40926) );
  XNOR U43768 ( .A(n40928), .B(n40929), .Z(n30985) );
  ANDN U43769 ( .B(\modmult_1/xin[1023] ), .A(n40930), .Z(n40928) );
  IV U43770 ( .A(n40929), .Z(n40930) );
  XNOR U43771 ( .A(m[119]), .B(n40931), .Z(n40929) );
  NAND U43772 ( .A(n40932), .B(mul_pow), .Z(n40931) );
  XOR U43773 ( .A(m[119]), .B(c[119]), .Z(n40932) );
  XOR U43774 ( .A(n40933), .B(n40934), .Z(n40925) );
  ANDN U43775 ( .B(n40935), .A(n30982), .Z(n40933) );
  XNOR U43776 ( .A(\modmult_1/zin[0][117] ), .B(n40936), .Z(n30982) );
  IV U43777 ( .A(n40934), .Z(n40936) );
  XOR U43778 ( .A(n40934), .B(n30983), .Z(n40935) );
  XNOR U43779 ( .A(n40937), .B(n40938), .Z(n30983) );
  ANDN U43780 ( .B(\modmult_1/xin[1023] ), .A(n40939), .Z(n40937) );
  IV U43781 ( .A(n40938), .Z(n40939) );
  XNOR U43782 ( .A(m[118]), .B(n40940), .Z(n40938) );
  NAND U43783 ( .A(n40941), .B(mul_pow), .Z(n40940) );
  XOR U43784 ( .A(m[118]), .B(c[118]), .Z(n40941) );
  XOR U43785 ( .A(n40942), .B(n40943), .Z(n40934) );
  ANDN U43786 ( .B(n40944), .A(n30980), .Z(n40942) );
  XNOR U43787 ( .A(\modmult_1/zin[0][116] ), .B(n40945), .Z(n30980) );
  IV U43788 ( .A(n40943), .Z(n40945) );
  XOR U43789 ( .A(n40943), .B(n30981), .Z(n40944) );
  XNOR U43790 ( .A(n40946), .B(n40947), .Z(n30981) );
  ANDN U43791 ( .B(\modmult_1/xin[1023] ), .A(n40948), .Z(n40946) );
  IV U43792 ( .A(n40947), .Z(n40948) );
  XNOR U43793 ( .A(m[117]), .B(n40949), .Z(n40947) );
  NAND U43794 ( .A(n40950), .B(mul_pow), .Z(n40949) );
  XOR U43795 ( .A(m[117]), .B(c[117]), .Z(n40950) );
  XOR U43796 ( .A(n40951), .B(n40952), .Z(n40943) );
  ANDN U43797 ( .B(n40953), .A(n30978), .Z(n40951) );
  XNOR U43798 ( .A(\modmult_1/zin[0][115] ), .B(n40954), .Z(n30978) );
  IV U43799 ( .A(n40952), .Z(n40954) );
  XOR U43800 ( .A(n40952), .B(n30979), .Z(n40953) );
  XNOR U43801 ( .A(n40955), .B(n40956), .Z(n30979) );
  ANDN U43802 ( .B(\modmult_1/xin[1023] ), .A(n40957), .Z(n40955) );
  IV U43803 ( .A(n40956), .Z(n40957) );
  XNOR U43804 ( .A(m[116]), .B(n40958), .Z(n40956) );
  NAND U43805 ( .A(n40959), .B(mul_pow), .Z(n40958) );
  XOR U43806 ( .A(m[116]), .B(c[116]), .Z(n40959) );
  XOR U43807 ( .A(n40960), .B(n40961), .Z(n40952) );
  ANDN U43808 ( .B(n40962), .A(n30976), .Z(n40960) );
  XNOR U43809 ( .A(\modmult_1/zin[0][114] ), .B(n40963), .Z(n30976) );
  IV U43810 ( .A(n40961), .Z(n40963) );
  XOR U43811 ( .A(n40961), .B(n30977), .Z(n40962) );
  XNOR U43812 ( .A(n40964), .B(n40965), .Z(n30977) );
  ANDN U43813 ( .B(\modmult_1/xin[1023] ), .A(n40966), .Z(n40964) );
  IV U43814 ( .A(n40965), .Z(n40966) );
  XNOR U43815 ( .A(m[115]), .B(n40967), .Z(n40965) );
  NAND U43816 ( .A(n40968), .B(mul_pow), .Z(n40967) );
  XOR U43817 ( .A(m[115]), .B(c[115]), .Z(n40968) );
  XOR U43818 ( .A(n40969), .B(n40970), .Z(n40961) );
  ANDN U43819 ( .B(n40971), .A(n30974), .Z(n40969) );
  XNOR U43820 ( .A(\modmult_1/zin[0][113] ), .B(n40972), .Z(n30974) );
  IV U43821 ( .A(n40970), .Z(n40972) );
  XOR U43822 ( .A(n40970), .B(n30975), .Z(n40971) );
  XNOR U43823 ( .A(n40973), .B(n40974), .Z(n30975) );
  ANDN U43824 ( .B(\modmult_1/xin[1023] ), .A(n40975), .Z(n40973) );
  IV U43825 ( .A(n40974), .Z(n40975) );
  XNOR U43826 ( .A(m[114]), .B(n40976), .Z(n40974) );
  NAND U43827 ( .A(n40977), .B(mul_pow), .Z(n40976) );
  XOR U43828 ( .A(m[114]), .B(c[114]), .Z(n40977) );
  XOR U43829 ( .A(n40978), .B(n40979), .Z(n40970) );
  ANDN U43830 ( .B(n40980), .A(n30972), .Z(n40978) );
  XNOR U43831 ( .A(\modmult_1/zin[0][112] ), .B(n40981), .Z(n30972) );
  IV U43832 ( .A(n40979), .Z(n40981) );
  XOR U43833 ( .A(n40979), .B(n30973), .Z(n40980) );
  XNOR U43834 ( .A(n40982), .B(n40983), .Z(n30973) );
  ANDN U43835 ( .B(\modmult_1/xin[1023] ), .A(n40984), .Z(n40982) );
  IV U43836 ( .A(n40983), .Z(n40984) );
  XNOR U43837 ( .A(m[113]), .B(n40985), .Z(n40983) );
  NAND U43838 ( .A(n40986), .B(mul_pow), .Z(n40985) );
  XOR U43839 ( .A(m[113]), .B(c[113]), .Z(n40986) );
  XOR U43840 ( .A(n40987), .B(n40988), .Z(n40979) );
  ANDN U43841 ( .B(n40989), .A(n30970), .Z(n40987) );
  XNOR U43842 ( .A(\modmult_1/zin[0][111] ), .B(n40990), .Z(n30970) );
  IV U43843 ( .A(n40988), .Z(n40990) );
  XOR U43844 ( .A(n40988), .B(n30971), .Z(n40989) );
  XNOR U43845 ( .A(n40991), .B(n40992), .Z(n30971) );
  ANDN U43846 ( .B(\modmult_1/xin[1023] ), .A(n40993), .Z(n40991) );
  IV U43847 ( .A(n40992), .Z(n40993) );
  XNOR U43848 ( .A(m[112]), .B(n40994), .Z(n40992) );
  NAND U43849 ( .A(n40995), .B(mul_pow), .Z(n40994) );
  XOR U43850 ( .A(m[112]), .B(c[112]), .Z(n40995) );
  XOR U43851 ( .A(n40996), .B(n40997), .Z(n40988) );
  ANDN U43852 ( .B(n40998), .A(n30968), .Z(n40996) );
  XNOR U43853 ( .A(\modmult_1/zin[0][110] ), .B(n40999), .Z(n30968) );
  IV U43854 ( .A(n40997), .Z(n40999) );
  XOR U43855 ( .A(n40997), .B(n30969), .Z(n40998) );
  XNOR U43856 ( .A(n41000), .B(n41001), .Z(n30969) );
  ANDN U43857 ( .B(\modmult_1/xin[1023] ), .A(n41002), .Z(n41000) );
  IV U43858 ( .A(n41001), .Z(n41002) );
  XNOR U43859 ( .A(m[111]), .B(n41003), .Z(n41001) );
  NAND U43860 ( .A(n41004), .B(mul_pow), .Z(n41003) );
  XOR U43861 ( .A(m[111]), .B(c[111]), .Z(n41004) );
  XOR U43862 ( .A(n41005), .B(n41006), .Z(n40997) );
  ANDN U43863 ( .B(n41007), .A(n30966), .Z(n41005) );
  XNOR U43864 ( .A(\modmult_1/zin[0][109] ), .B(n41008), .Z(n30966) );
  IV U43865 ( .A(n41006), .Z(n41008) );
  XOR U43866 ( .A(n41006), .B(n30967), .Z(n41007) );
  XNOR U43867 ( .A(n41009), .B(n41010), .Z(n30967) );
  ANDN U43868 ( .B(\modmult_1/xin[1023] ), .A(n41011), .Z(n41009) );
  IV U43869 ( .A(n41010), .Z(n41011) );
  XNOR U43870 ( .A(m[110]), .B(n41012), .Z(n41010) );
  NAND U43871 ( .A(n41013), .B(mul_pow), .Z(n41012) );
  XOR U43872 ( .A(m[110]), .B(c[110]), .Z(n41013) );
  XOR U43873 ( .A(n41014), .B(n41015), .Z(n41006) );
  ANDN U43874 ( .B(n41016), .A(n30964), .Z(n41014) );
  XNOR U43875 ( .A(\modmult_1/zin[0][108] ), .B(n41017), .Z(n30964) );
  IV U43876 ( .A(n41015), .Z(n41017) );
  XOR U43877 ( .A(n41015), .B(n30965), .Z(n41016) );
  XNOR U43878 ( .A(n41018), .B(n41019), .Z(n30965) );
  ANDN U43879 ( .B(\modmult_1/xin[1023] ), .A(n41020), .Z(n41018) );
  IV U43880 ( .A(n41019), .Z(n41020) );
  XNOR U43881 ( .A(m[109]), .B(n41021), .Z(n41019) );
  NAND U43882 ( .A(n41022), .B(mul_pow), .Z(n41021) );
  XOR U43883 ( .A(m[109]), .B(c[109]), .Z(n41022) );
  XOR U43884 ( .A(n41023), .B(n41024), .Z(n41015) );
  ANDN U43885 ( .B(n41025), .A(n30962), .Z(n41023) );
  XNOR U43886 ( .A(\modmult_1/zin[0][107] ), .B(n41026), .Z(n30962) );
  IV U43887 ( .A(n41024), .Z(n41026) );
  XOR U43888 ( .A(n41024), .B(n30963), .Z(n41025) );
  XNOR U43889 ( .A(n41027), .B(n41028), .Z(n30963) );
  ANDN U43890 ( .B(\modmult_1/xin[1023] ), .A(n41029), .Z(n41027) );
  IV U43891 ( .A(n41028), .Z(n41029) );
  XNOR U43892 ( .A(m[108]), .B(n41030), .Z(n41028) );
  NAND U43893 ( .A(n41031), .B(mul_pow), .Z(n41030) );
  XOR U43894 ( .A(m[108]), .B(c[108]), .Z(n41031) );
  XOR U43895 ( .A(n41032), .B(n41033), .Z(n41024) );
  ANDN U43896 ( .B(n41034), .A(n30960), .Z(n41032) );
  XNOR U43897 ( .A(\modmult_1/zin[0][106] ), .B(n41035), .Z(n30960) );
  IV U43898 ( .A(n41033), .Z(n41035) );
  XOR U43899 ( .A(n41033), .B(n30961), .Z(n41034) );
  XNOR U43900 ( .A(n41036), .B(n41037), .Z(n30961) );
  ANDN U43901 ( .B(\modmult_1/xin[1023] ), .A(n41038), .Z(n41036) );
  IV U43902 ( .A(n41037), .Z(n41038) );
  XNOR U43903 ( .A(m[107]), .B(n41039), .Z(n41037) );
  NAND U43904 ( .A(n41040), .B(mul_pow), .Z(n41039) );
  XOR U43905 ( .A(m[107]), .B(c[107]), .Z(n41040) );
  XOR U43906 ( .A(n41041), .B(n41042), .Z(n41033) );
  ANDN U43907 ( .B(n41043), .A(n30958), .Z(n41041) );
  XNOR U43908 ( .A(\modmult_1/zin[0][105] ), .B(n41044), .Z(n30958) );
  IV U43909 ( .A(n41042), .Z(n41044) );
  XOR U43910 ( .A(n41042), .B(n30959), .Z(n41043) );
  XNOR U43911 ( .A(n41045), .B(n41046), .Z(n30959) );
  ANDN U43912 ( .B(\modmult_1/xin[1023] ), .A(n41047), .Z(n41045) );
  IV U43913 ( .A(n41046), .Z(n41047) );
  XNOR U43914 ( .A(m[106]), .B(n41048), .Z(n41046) );
  NAND U43915 ( .A(n41049), .B(mul_pow), .Z(n41048) );
  XOR U43916 ( .A(m[106]), .B(c[106]), .Z(n41049) );
  XOR U43917 ( .A(n41050), .B(n41051), .Z(n41042) );
  ANDN U43918 ( .B(n41052), .A(n30956), .Z(n41050) );
  XNOR U43919 ( .A(\modmult_1/zin[0][104] ), .B(n41053), .Z(n30956) );
  IV U43920 ( .A(n41051), .Z(n41053) );
  XOR U43921 ( .A(n41051), .B(n30957), .Z(n41052) );
  XNOR U43922 ( .A(n41054), .B(n41055), .Z(n30957) );
  ANDN U43923 ( .B(\modmult_1/xin[1023] ), .A(n41056), .Z(n41054) );
  IV U43924 ( .A(n41055), .Z(n41056) );
  XNOR U43925 ( .A(m[105]), .B(n41057), .Z(n41055) );
  NAND U43926 ( .A(n41058), .B(mul_pow), .Z(n41057) );
  XOR U43927 ( .A(m[105]), .B(c[105]), .Z(n41058) );
  XOR U43928 ( .A(n41059), .B(n41060), .Z(n41051) );
  ANDN U43929 ( .B(n41061), .A(n30954), .Z(n41059) );
  XNOR U43930 ( .A(\modmult_1/zin[0][103] ), .B(n41062), .Z(n30954) );
  IV U43931 ( .A(n41060), .Z(n41062) );
  XOR U43932 ( .A(n41060), .B(n30955), .Z(n41061) );
  XNOR U43933 ( .A(n41063), .B(n41064), .Z(n30955) );
  ANDN U43934 ( .B(\modmult_1/xin[1023] ), .A(n41065), .Z(n41063) );
  IV U43935 ( .A(n41064), .Z(n41065) );
  XNOR U43936 ( .A(m[104]), .B(n41066), .Z(n41064) );
  NAND U43937 ( .A(n41067), .B(mul_pow), .Z(n41066) );
  XOR U43938 ( .A(m[104]), .B(c[104]), .Z(n41067) );
  XOR U43939 ( .A(n41068), .B(n41069), .Z(n41060) );
  ANDN U43940 ( .B(n41070), .A(n30952), .Z(n41068) );
  XNOR U43941 ( .A(\modmult_1/zin[0][102] ), .B(n41071), .Z(n30952) );
  IV U43942 ( .A(n41069), .Z(n41071) );
  XOR U43943 ( .A(n41069), .B(n30953), .Z(n41070) );
  XNOR U43944 ( .A(n41072), .B(n41073), .Z(n30953) );
  ANDN U43945 ( .B(\modmult_1/xin[1023] ), .A(n41074), .Z(n41072) );
  IV U43946 ( .A(n41073), .Z(n41074) );
  XNOR U43947 ( .A(m[103]), .B(n41075), .Z(n41073) );
  NAND U43948 ( .A(n41076), .B(mul_pow), .Z(n41075) );
  XOR U43949 ( .A(m[103]), .B(c[103]), .Z(n41076) );
  XOR U43950 ( .A(n41077), .B(n41078), .Z(n41069) );
  ANDN U43951 ( .B(n41079), .A(n30950), .Z(n41077) );
  XNOR U43952 ( .A(\modmult_1/zin[0][101] ), .B(n41080), .Z(n30950) );
  IV U43953 ( .A(n41078), .Z(n41080) );
  XOR U43954 ( .A(n41078), .B(n30951), .Z(n41079) );
  XNOR U43955 ( .A(n41081), .B(n41082), .Z(n30951) );
  ANDN U43956 ( .B(\modmult_1/xin[1023] ), .A(n41083), .Z(n41081) );
  IV U43957 ( .A(n41082), .Z(n41083) );
  XNOR U43958 ( .A(m[102]), .B(n41084), .Z(n41082) );
  NAND U43959 ( .A(n41085), .B(mul_pow), .Z(n41084) );
  XOR U43960 ( .A(m[102]), .B(c[102]), .Z(n41085) );
  XOR U43961 ( .A(n41086), .B(n41087), .Z(n41078) );
  ANDN U43962 ( .B(n41088), .A(n30948), .Z(n41086) );
  XNOR U43963 ( .A(\modmult_1/zin[0][100] ), .B(n41089), .Z(n30948) );
  IV U43964 ( .A(n41087), .Z(n41089) );
  XOR U43965 ( .A(n41087), .B(n30949), .Z(n41088) );
  XNOR U43966 ( .A(n41090), .B(n41091), .Z(n30949) );
  ANDN U43967 ( .B(\modmult_1/xin[1023] ), .A(n41092), .Z(n41090) );
  IV U43968 ( .A(n41091), .Z(n41092) );
  XNOR U43969 ( .A(m[101]), .B(n41093), .Z(n41091) );
  NAND U43970 ( .A(n41094), .B(mul_pow), .Z(n41093) );
  XOR U43971 ( .A(m[101]), .B(c[101]), .Z(n41094) );
  XOR U43972 ( .A(n41095), .B(n41096), .Z(n41087) );
  ANDN U43973 ( .B(n41097), .A(n30946), .Z(n41095) );
  XNOR U43974 ( .A(\modmult_1/zin[0][99] ), .B(n41098), .Z(n30946) );
  IV U43975 ( .A(n41096), .Z(n41098) );
  XOR U43976 ( .A(n41096), .B(n30947), .Z(n41097) );
  XNOR U43977 ( .A(n41099), .B(n41100), .Z(n30947) );
  ANDN U43978 ( .B(\modmult_1/xin[1023] ), .A(n41101), .Z(n41099) );
  IV U43979 ( .A(n41100), .Z(n41101) );
  XNOR U43980 ( .A(m[100]), .B(n41102), .Z(n41100) );
  NAND U43981 ( .A(n41103), .B(mul_pow), .Z(n41102) );
  XOR U43982 ( .A(m[100]), .B(c[100]), .Z(n41103) );
  XOR U43983 ( .A(n41104), .B(n41105), .Z(n41096) );
  ANDN U43984 ( .B(n41106), .A(n30944), .Z(n41104) );
  XNOR U43985 ( .A(\modmult_1/zin[0][98] ), .B(n41107), .Z(n30944) );
  IV U43986 ( .A(n41105), .Z(n41107) );
  XOR U43987 ( .A(n41105), .B(n30945), .Z(n41106) );
  XNOR U43988 ( .A(n41108), .B(n41109), .Z(n30945) );
  ANDN U43989 ( .B(\modmult_1/xin[1023] ), .A(n41110), .Z(n41108) );
  IV U43990 ( .A(n41109), .Z(n41110) );
  XNOR U43991 ( .A(m[99]), .B(n41111), .Z(n41109) );
  NAND U43992 ( .A(n41112), .B(mul_pow), .Z(n41111) );
  XOR U43993 ( .A(m[99]), .B(c[99]), .Z(n41112) );
  XOR U43994 ( .A(n41113), .B(n41114), .Z(n41105) );
  ANDN U43995 ( .B(n41115), .A(n30942), .Z(n41113) );
  XNOR U43996 ( .A(\modmult_1/zin[0][97] ), .B(n41116), .Z(n30942) );
  IV U43997 ( .A(n41114), .Z(n41116) );
  XOR U43998 ( .A(n41114), .B(n30943), .Z(n41115) );
  XNOR U43999 ( .A(n41117), .B(n41118), .Z(n30943) );
  ANDN U44000 ( .B(\modmult_1/xin[1023] ), .A(n41119), .Z(n41117) );
  IV U44001 ( .A(n41118), .Z(n41119) );
  XNOR U44002 ( .A(m[98]), .B(n41120), .Z(n41118) );
  NAND U44003 ( .A(n41121), .B(mul_pow), .Z(n41120) );
  XOR U44004 ( .A(m[98]), .B(c[98]), .Z(n41121) );
  XOR U44005 ( .A(n41122), .B(n41123), .Z(n41114) );
  ANDN U44006 ( .B(n41124), .A(n30940), .Z(n41122) );
  XNOR U44007 ( .A(\modmult_1/zin[0][96] ), .B(n41125), .Z(n30940) );
  IV U44008 ( .A(n41123), .Z(n41125) );
  XOR U44009 ( .A(n41123), .B(n30941), .Z(n41124) );
  XNOR U44010 ( .A(n41126), .B(n41127), .Z(n30941) );
  ANDN U44011 ( .B(\modmult_1/xin[1023] ), .A(n41128), .Z(n41126) );
  IV U44012 ( .A(n41127), .Z(n41128) );
  XNOR U44013 ( .A(m[97]), .B(n41129), .Z(n41127) );
  NAND U44014 ( .A(n41130), .B(mul_pow), .Z(n41129) );
  XOR U44015 ( .A(m[97]), .B(c[97]), .Z(n41130) );
  XOR U44016 ( .A(n41131), .B(n41132), .Z(n41123) );
  ANDN U44017 ( .B(n41133), .A(n30938), .Z(n41131) );
  XNOR U44018 ( .A(\modmult_1/zin[0][95] ), .B(n41134), .Z(n30938) );
  IV U44019 ( .A(n41132), .Z(n41134) );
  XOR U44020 ( .A(n41132), .B(n30939), .Z(n41133) );
  XNOR U44021 ( .A(n41135), .B(n41136), .Z(n30939) );
  ANDN U44022 ( .B(\modmult_1/xin[1023] ), .A(n41137), .Z(n41135) );
  IV U44023 ( .A(n41136), .Z(n41137) );
  XNOR U44024 ( .A(m[96]), .B(n41138), .Z(n41136) );
  NAND U44025 ( .A(n41139), .B(mul_pow), .Z(n41138) );
  XOR U44026 ( .A(m[96]), .B(c[96]), .Z(n41139) );
  XOR U44027 ( .A(n41140), .B(n41141), .Z(n41132) );
  ANDN U44028 ( .B(n41142), .A(n30936), .Z(n41140) );
  XNOR U44029 ( .A(\modmult_1/zin[0][94] ), .B(n41143), .Z(n30936) );
  IV U44030 ( .A(n41141), .Z(n41143) );
  XOR U44031 ( .A(n41141), .B(n30937), .Z(n41142) );
  XNOR U44032 ( .A(n41144), .B(n41145), .Z(n30937) );
  ANDN U44033 ( .B(\modmult_1/xin[1023] ), .A(n41146), .Z(n41144) );
  IV U44034 ( .A(n41145), .Z(n41146) );
  XNOR U44035 ( .A(m[95]), .B(n41147), .Z(n41145) );
  NAND U44036 ( .A(n41148), .B(mul_pow), .Z(n41147) );
  XOR U44037 ( .A(m[95]), .B(c[95]), .Z(n41148) );
  XOR U44038 ( .A(n41149), .B(n41150), .Z(n41141) );
  ANDN U44039 ( .B(n41151), .A(n30934), .Z(n41149) );
  XNOR U44040 ( .A(\modmult_1/zin[0][93] ), .B(n41152), .Z(n30934) );
  IV U44041 ( .A(n41150), .Z(n41152) );
  XOR U44042 ( .A(n41150), .B(n30935), .Z(n41151) );
  XNOR U44043 ( .A(n41153), .B(n41154), .Z(n30935) );
  ANDN U44044 ( .B(\modmult_1/xin[1023] ), .A(n41155), .Z(n41153) );
  IV U44045 ( .A(n41154), .Z(n41155) );
  XNOR U44046 ( .A(m[94]), .B(n41156), .Z(n41154) );
  NAND U44047 ( .A(n41157), .B(mul_pow), .Z(n41156) );
  XOR U44048 ( .A(m[94]), .B(c[94]), .Z(n41157) );
  XOR U44049 ( .A(n41158), .B(n41159), .Z(n41150) );
  ANDN U44050 ( .B(n41160), .A(n30932), .Z(n41158) );
  XNOR U44051 ( .A(\modmult_1/zin[0][92] ), .B(n41161), .Z(n30932) );
  IV U44052 ( .A(n41159), .Z(n41161) );
  XOR U44053 ( .A(n41159), .B(n30933), .Z(n41160) );
  XNOR U44054 ( .A(n41162), .B(n41163), .Z(n30933) );
  ANDN U44055 ( .B(\modmult_1/xin[1023] ), .A(n41164), .Z(n41162) );
  IV U44056 ( .A(n41163), .Z(n41164) );
  XNOR U44057 ( .A(m[93]), .B(n41165), .Z(n41163) );
  NAND U44058 ( .A(n41166), .B(mul_pow), .Z(n41165) );
  XOR U44059 ( .A(m[93]), .B(c[93]), .Z(n41166) );
  XOR U44060 ( .A(n41167), .B(n41168), .Z(n41159) );
  ANDN U44061 ( .B(n41169), .A(n30930), .Z(n41167) );
  XNOR U44062 ( .A(\modmult_1/zin[0][91] ), .B(n41170), .Z(n30930) );
  IV U44063 ( .A(n41168), .Z(n41170) );
  XOR U44064 ( .A(n41168), .B(n30931), .Z(n41169) );
  XNOR U44065 ( .A(n41171), .B(n41172), .Z(n30931) );
  ANDN U44066 ( .B(\modmult_1/xin[1023] ), .A(n41173), .Z(n41171) );
  IV U44067 ( .A(n41172), .Z(n41173) );
  XNOR U44068 ( .A(m[92]), .B(n41174), .Z(n41172) );
  NAND U44069 ( .A(n41175), .B(mul_pow), .Z(n41174) );
  XOR U44070 ( .A(m[92]), .B(c[92]), .Z(n41175) );
  XOR U44071 ( .A(n41176), .B(n41177), .Z(n41168) );
  ANDN U44072 ( .B(n41178), .A(n30928), .Z(n41176) );
  XNOR U44073 ( .A(\modmult_1/zin[0][90] ), .B(n41179), .Z(n30928) );
  IV U44074 ( .A(n41177), .Z(n41179) );
  XOR U44075 ( .A(n41177), .B(n30929), .Z(n41178) );
  XNOR U44076 ( .A(n41180), .B(n41181), .Z(n30929) );
  ANDN U44077 ( .B(\modmult_1/xin[1023] ), .A(n41182), .Z(n41180) );
  IV U44078 ( .A(n41181), .Z(n41182) );
  XNOR U44079 ( .A(m[91]), .B(n41183), .Z(n41181) );
  NAND U44080 ( .A(n41184), .B(mul_pow), .Z(n41183) );
  XOR U44081 ( .A(m[91]), .B(c[91]), .Z(n41184) );
  XOR U44082 ( .A(n41185), .B(n41186), .Z(n41177) );
  ANDN U44083 ( .B(n41187), .A(n30926), .Z(n41185) );
  XNOR U44084 ( .A(\modmult_1/zin[0][89] ), .B(n41188), .Z(n30926) );
  IV U44085 ( .A(n41186), .Z(n41188) );
  XOR U44086 ( .A(n41186), .B(n30927), .Z(n41187) );
  XNOR U44087 ( .A(n41189), .B(n41190), .Z(n30927) );
  ANDN U44088 ( .B(\modmult_1/xin[1023] ), .A(n41191), .Z(n41189) );
  IV U44089 ( .A(n41190), .Z(n41191) );
  XNOR U44090 ( .A(m[90]), .B(n41192), .Z(n41190) );
  NAND U44091 ( .A(n41193), .B(mul_pow), .Z(n41192) );
  XOR U44092 ( .A(m[90]), .B(c[90]), .Z(n41193) );
  XOR U44093 ( .A(n41194), .B(n41195), .Z(n41186) );
  ANDN U44094 ( .B(n41196), .A(n30924), .Z(n41194) );
  XNOR U44095 ( .A(\modmult_1/zin[0][88] ), .B(n41197), .Z(n30924) );
  IV U44096 ( .A(n41195), .Z(n41197) );
  XOR U44097 ( .A(n41195), .B(n30925), .Z(n41196) );
  XNOR U44098 ( .A(n41198), .B(n41199), .Z(n30925) );
  ANDN U44099 ( .B(\modmult_1/xin[1023] ), .A(n41200), .Z(n41198) );
  IV U44100 ( .A(n41199), .Z(n41200) );
  XNOR U44101 ( .A(m[89]), .B(n41201), .Z(n41199) );
  NAND U44102 ( .A(n41202), .B(mul_pow), .Z(n41201) );
  XOR U44103 ( .A(m[89]), .B(c[89]), .Z(n41202) );
  XOR U44104 ( .A(n41203), .B(n41204), .Z(n41195) );
  ANDN U44105 ( .B(n41205), .A(n30922), .Z(n41203) );
  XNOR U44106 ( .A(\modmult_1/zin[0][87] ), .B(n41206), .Z(n30922) );
  IV U44107 ( .A(n41204), .Z(n41206) );
  XOR U44108 ( .A(n41204), .B(n30923), .Z(n41205) );
  XNOR U44109 ( .A(n41207), .B(n41208), .Z(n30923) );
  ANDN U44110 ( .B(\modmult_1/xin[1023] ), .A(n41209), .Z(n41207) );
  IV U44111 ( .A(n41208), .Z(n41209) );
  XNOR U44112 ( .A(m[88]), .B(n41210), .Z(n41208) );
  NAND U44113 ( .A(n41211), .B(mul_pow), .Z(n41210) );
  XOR U44114 ( .A(m[88]), .B(c[88]), .Z(n41211) );
  XOR U44115 ( .A(n41212), .B(n41213), .Z(n41204) );
  ANDN U44116 ( .B(n41214), .A(n30920), .Z(n41212) );
  XNOR U44117 ( .A(\modmult_1/zin[0][86] ), .B(n41215), .Z(n30920) );
  IV U44118 ( .A(n41213), .Z(n41215) );
  XOR U44119 ( .A(n41213), .B(n30921), .Z(n41214) );
  XNOR U44120 ( .A(n41216), .B(n41217), .Z(n30921) );
  ANDN U44121 ( .B(\modmult_1/xin[1023] ), .A(n41218), .Z(n41216) );
  IV U44122 ( .A(n41217), .Z(n41218) );
  XNOR U44123 ( .A(m[87]), .B(n41219), .Z(n41217) );
  NAND U44124 ( .A(n41220), .B(mul_pow), .Z(n41219) );
  XOR U44125 ( .A(m[87]), .B(c[87]), .Z(n41220) );
  XOR U44126 ( .A(n41221), .B(n41222), .Z(n41213) );
  ANDN U44127 ( .B(n41223), .A(n30918), .Z(n41221) );
  XNOR U44128 ( .A(\modmult_1/zin[0][85] ), .B(n41224), .Z(n30918) );
  IV U44129 ( .A(n41222), .Z(n41224) );
  XOR U44130 ( .A(n41222), .B(n30919), .Z(n41223) );
  XNOR U44131 ( .A(n41225), .B(n41226), .Z(n30919) );
  ANDN U44132 ( .B(\modmult_1/xin[1023] ), .A(n41227), .Z(n41225) );
  IV U44133 ( .A(n41226), .Z(n41227) );
  XNOR U44134 ( .A(m[86]), .B(n41228), .Z(n41226) );
  NAND U44135 ( .A(n41229), .B(mul_pow), .Z(n41228) );
  XOR U44136 ( .A(m[86]), .B(c[86]), .Z(n41229) );
  XOR U44137 ( .A(n41230), .B(n41231), .Z(n41222) );
  ANDN U44138 ( .B(n41232), .A(n30916), .Z(n41230) );
  XNOR U44139 ( .A(\modmult_1/zin[0][84] ), .B(n41233), .Z(n30916) );
  IV U44140 ( .A(n41231), .Z(n41233) );
  XOR U44141 ( .A(n41231), .B(n30917), .Z(n41232) );
  XNOR U44142 ( .A(n41234), .B(n41235), .Z(n30917) );
  ANDN U44143 ( .B(\modmult_1/xin[1023] ), .A(n41236), .Z(n41234) );
  IV U44144 ( .A(n41235), .Z(n41236) );
  XNOR U44145 ( .A(m[85]), .B(n41237), .Z(n41235) );
  NAND U44146 ( .A(n41238), .B(mul_pow), .Z(n41237) );
  XOR U44147 ( .A(m[85]), .B(c[85]), .Z(n41238) );
  XOR U44148 ( .A(n41239), .B(n41240), .Z(n41231) );
  ANDN U44149 ( .B(n41241), .A(n30914), .Z(n41239) );
  XNOR U44150 ( .A(\modmult_1/zin[0][83] ), .B(n41242), .Z(n30914) );
  IV U44151 ( .A(n41240), .Z(n41242) );
  XOR U44152 ( .A(n41240), .B(n30915), .Z(n41241) );
  XNOR U44153 ( .A(n41243), .B(n41244), .Z(n30915) );
  ANDN U44154 ( .B(\modmult_1/xin[1023] ), .A(n41245), .Z(n41243) );
  IV U44155 ( .A(n41244), .Z(n41245) );
  XNOR U44156 ( .A(m[84]), .B(n41246), .Z(n41244) );
  NAND U44157 ( .A(n41247), .B(mul_pow), .Z(n41246) );
  XOR U44158 ( .A(m[84]), .B(c[84]), .Z(n41247) );
  XOR U44159 ( .A(n41248), .B(n41249), .Z(n41240) );
  ANDN U44160 ( .B(n41250), .A(n30912), .Z(n41248) );
  XNOR U44161 ( .A(\modmult_1/zin[0][82] ), .B(n41251), .Z(n30912) );
  IV U44162 ( .A(n41249), .Z(n41251) );
  XOR U44163 ( .A(n41249), .B(n30913), .Z(n41250) );
  XNOR U44164 ( .A(n41252), .B(n41253), .Z(n30913) );
  ANDN U44165 ( .B(\modmult_1/xin[1023] ), .A(n41254), .Z(n41252) );
  IV U44166 ( .A(n41253), .Z(n41254) );
  XNOR U44167 ( .A(m[83]), .B(n41255), .Z(n41253) );
  NAND U44168 ( .A(n41256), .B(mul_pow), .Z(n41255) );
  XOR U44169 ( .A(m[83]), .B(c[83]), .Z(n41256) );
  XOR U44170 ( .A(n41257), .B(n41258), .Z(n41249) );
  ANDN U44171 ( .B(n41259), .A(n30910), .Z(n41257) );
  XNOR U44172 ( .A(\modmult_1/zin[0][81] ), .B(n41260), .Z(n30910) );
  IV U44173 ( .A(n41258), .Z(n41260) );
  XOR U44174 ( .A(n41258), .B(n30911), .Z(n41259) );
  XNOR U44175 ( .A(n41261), .B(n41262), .Z(n30911) );
  ANDN U44176 ( .B(\modmult_1/xin[1023] ), .A(n41263), .Z(n41261) );
  IV U44177 ( .A(n41262), .Z(n41263) );
  XNOR U44178 ( .A(m[82]), .B(n41264), .Z(n41262) );
  NAND U44179 ( .A(n41265), .B(mul_pow), .Z(n41264) );
  XOR U44180 ( .A(m[82]), .B(c[82]), .Z(n41265) );
  XOR U44181 ( .A(n41266), .B(n41267), .Z(n41258) );
  ANDN U44182 ( .B(n41268), .A(n30908), .Z(n41266) );
  XNOR U44183 ( .A(\modmult_1/zin[0][80] ), .B(n41269), .Z(n30908) );
  IV U44184 ( .A(n41267), .Z(n41269) );
  XOR U44185 ( .A(n41267), .B(n30909), .Z(n41268) );
  XNOR U44186 ( .A(n41270), .B(n41271), .Z(n30909) );
  ANDN U44187 ( .B(\modmult_1/xin[1023] ), .A(n41272), .Z(n41270) );
  IV U44188 ( .A(n41271), .Z(n41272) );
  XNOR U44189 ( .A(m[81]), .B(n41273), .Z(n41271) );
  NAND U44190 ( .A(n41274), .B(mul_pow), .Z(n41273) );
  XOR U44191 ( .A(m[81]), .B(c[81]), .Z(n41274) );
  XOR U44192 ( .A(n41275), .B(n41276), .Z(n41267) );
  ANDN U44193 ( .B(n41277), .A(n30906), .Z(n41275) );
  XNOR U44194 ( .A(\modmult_1/zin[0][79] ), .B(n41278), .Z(n30906) );
  IV U44195 ( .A(n41276), .Z(n41278) );
  XOR U44196 ( .A(n41276), .B(n30907), .Z(n41277) );
  XNOR U44197 ( .A(n41279), .B(n41280), .Z(n30907) );
  ANDN U44198 ( .B(\modmult_1/xin[1023] ), .A(n41281), .Z(n41279) );
  IV U44199 ( .A(n41280), .Z(n41281) );
  XNOR U44200 ( .A(m[80]), .B(n41282), .Z(n41280) );
  NAND U44201 ( .A(n41283), .B(mul_pow), .Z(n41282) );
  XOR U44202 ( .A(m[80]), .B(c[80]), .Z(n41283) );
  XOR U44203 ( .A(n41284), .B(n41285), .Z(n41276) );
  ANDN U44204 ( .B(n41286), .A(n30904), .Z(n41284) );
  XNOR U44205 ( .A(\modmult_1/zin[0][78] ), .B(n41287), .Z(n30904) );
  IV U44206 ( .A(n41285), .Z(n41287) );
  XOR U44207 ( .A(n41285), .B(n30905), .Z(n41286) );
  XNOR U44208 ( .A(n41288), .B(n41289), .Z(n30905) );
  ANDN U44209 ( .B(\modmult_1/xin[1023] ), .A(n41290), .Z(n41288) );
  IV U44210 ( .A(n41289), .Z(n41290) );
  XNOR U44211 ( .A(m[79]), .B(n41291), .Z(n41289) );
  NAND U44212 ( .A(n41292), .B(mul_pow), .Z(n41291) );
  XOR U44213 ( .A(m[79]), .B(c[79]), .Z(n41292) );
  XOR U44214 ( .A(n41293), .B(n41294), .Z(n41285) );
  ANDN U44215 ( .B(n41295), .A(n30902), .Z(n41293) );
  XNOR U44216 ( .A(\modmult_1/zin[0][77] ), .B(n41296), .Z(n30902) );
  IV U44217 ( .A(n41294), .Z(n41296) );
  XOR U44218 ( .A(n41294), .B(n30903), .Z(n41295) );
  XNOR U44219 ( .A(n41297), .B(n41298), .Z(n30903) );
  ANDN U44220 ( .B(\modmult_1/xin[1023] ), .A(n41299), .Z(n41297) );
  IV U44221 ( .A(n41298), .Z(n41299) );
  XNOR U44222 ( .A(m[78]), .B(n41300), .Z(n41298) );
  NAND U44223 ( .A(n41301), .B(mul_pow), .Z(n41300) );
  XOR U44224 ( .A(m[78]), .B(c[78]), .Z(n41301) );
  XOR U44225 ( .A(n41302), .B(n41303), .Z(n41294) );
  ANDN U44226 ( .B(n41304), .A(n30900), .Z(n41302) );
  XNOR U44227 ( .A(\modmult_1/zin[0][76] ), .B(n41305), .Z(n30900) );
  IV U44228 ( .A(n41303), .Z(n41305) );
  XOR U44229 ( .A(n41303), .B(n30901), .Z(n41304) );
  XNOR U44230 ( .A(n41306), .B(n41307), .Z(n30901) );
  ANDN U44231 ( .B(\modmult_1/xin[1023] ), .A(n41308), .Z(n41306) );
  IV U44232 ( .A(n41307), .Z(n41308) );
  XNOR U44233 ( .A(m[77]), .B(n41309), .Z(n41307) );
  NAND U44234 ( .A(n41310), .B(mul_pow), .Z(n41309) );
  XOR U44235 ( .A(m[77]), .B(c[77]), .Z(n41310) );
  XOR U44236 ( .A(n41311), .B(n41312), .Z(n41303) );
  ANDN U44237 ( .B(n41313), .A(n30898), .Z(n41311) );
  XNOR U44238 ( .A(\modmult_1/zin[0][75] ), .B(n41314), .Z(n30898) );
  IV U44239 ( .A(n41312), .Z(n41314) );
  XOR U44240 ( .A(n41312), .B(n30899), .Z(n41313) );
  XNOR U44241 ( .A(n41315), .B(n41316), .Z(n30899) );
  ANDN U44242 ( .B(\modmult_1/xin[1023] ), .A(n41317), .Z(n41315) );
  IV U44243 ( .A(n41316), .Z(n41317) );
  XNOR U44244 ( .A(m[76]), .B(n41318), .Z(n41316) );
  NAND U44245 ( .A(n41319), .B(mul_pow), .Z(n41318) );
  XOR U44246 ( .A(m[76]), .B(c[76]), .Z(n41319) );
  XOR U44247 ( .A(n41320), .B(n41321), .Z(n41312) );
  ANDN U44248 ( .B(n41322), .A(n30896), .Z(n41320) );
  XNOR U44249 ( .A(\modmult_1/zin[0][74] ), .B(n41323), .Z(n30896) );
  IV U44250 ( .A(n41321), .Z(n41323) );
  XOR U44251 ( .A(n41321), .B(n30897), .Z(n41322) );
  XNOR U44252 ( .A(n41324), .B(n41325), .Z(n30897) );
  ANDN U44253 ( .B(\modmult_1/xin[1023] ), .A(n41326), .Z(n41324) );
  IV U44254 ( .A(n41325), .Z(n41326) );
  XNOR U44255 ( .A(m[75]), .B(n41327), .Z(n41325) );
  NAND U44256 ( .A(n41328), .B(mul_pow), .Z(n41327) );
  XOR U44257 ( .A(m[75]), .B(c[75]), .Z(n41328) );
  XOR U44258 ( .A(n41329), .B(n41330), .Z(n41321) );
  ANDN U44259 ( .B(n41331), .A(n30894), .Z(n41329) );
  XNOR U44260 ( .A(\modmult_1/zin[0][73] ), .B(n41332), .Z(n30894) );
  IV U44261 ( .A(n41330), .Z(n41332) );
  XOR U44262 ( .A(n41330), .B(n30895), .Z(n41331) );
  XNOR U44263 ( .A(n41333), .B(n41334), .Z(n30895) );
  ANDN U44264 ( .B(\modmult_1/xin[1023] ), .A(n41335), .Z(n41333) );
  IV U44265 ( .A(n41334), .Z(n41335) );
  XNOR U44266 ( .A(m[74]), .B(n41336), .Z(n41334) );
  NAND U44267 ( .A(n41337), .B(mul_pow), .Z(n41336) );
  XOR U44268 ( .A(m[74]), .B(c[74]), .Z(n41337) );
  XOR U44269 ( .A(n41338), .B(n41339), .Z(n41330) );
  ANDN U44270 ( .B(n41340), .A(n30892), .Z(n41338) );
  XNOR U44271 ( .A(\modmult_1/zin[0][72] ), .B(n41341), .Z(n30892) );
  IV U44272 ( .A(n41339), .Z(n41341) );
  XOR U44273 ( .A(n41339), .B(n30893), .Z(n41340) );
  XNOR U44274 ( .A(n41342), .B(n41343), .Z(n30893) );
  ANDN U44275 ( .B(\modmult_1/xin[1023] ), .A(n41344), .Z(n41342) );
  IV U44276 ( .A(n41343), .Z(n41344) );
  XNOR U44277 ( .A(m[73]), .B(n41345), .Z(n41343) );
  NAND U44278 ( .A(n41346), .B(mul_pow), .Z(n41345) );
  XOR U44279 ( .A(m[73]), .B(c[73]), .Z(n41346) );
  XOR U44280 ( .A(n41347), .B(n41348), .Z(n41339) );
  ANDN U44281 ( .B(n41349), .A(n30890), .Z(n41347) );
  XNOR U44282 ( .A(\modmult_1/zin[0][71] ), .B(n41350), .Z(n30890) );
  IV U44283 ( .A(n41348), .Z(n41350) );
  XOR U44284 ( .A(n41348), .B(n30891), .Z(n41349) );
  XNOR U44285 ( .A(n41351), .B(n41352), .Z(n30891) );
  ANDN U44286 ( .B(\modmult_1/xin[1023] ), .A(n41353), .Z(n41351) );
  IV U44287 ( .A(n41352), .Z(n41353) );
  XNOR U44288 ( .A(m[72]), .B(n41354), .Z(n41352) );
  NAND U44289 ( .A(n41355), .B(mul_pow), .Z(n41354) );
  XOR U44290 ( .A(m[72]), .B(c[72]), .Z(n41355) );
  XOR U44291 ( .A(n41356), .B(n41357), .Z(n41348) );
  ANDN U44292 ( .B(n41358), .A(n30888), .Z(n41356) );
  XNOR U44293 ( .A(\modmult_1/zin[0][70] ), .B(n41359), .Z(n30888) );
  IV U44294 ( .A(n41357), .Z(n41359) );
  XOR U44295 ( .A(n41357), .B(n30889), .Z(n41358) );
  XNOR U44296 ( .A(n41360), .B(n41361), .Z(n30889) );
  ANDN U44297 ( .B(\modmult_1/xin[1023] ), .A(n41362), .Z(n41360) );
  IV U44298 ( .A(n41361), .Z(n41362) );
  XNOR U44299 ( .A(m[71]), .B(n41363), .Z(n41361) );
  NAND U44300 ( .A(n41364), .B(mul_pow), .Z(n41363) );
  XOR U44301 ( .A(m[71]), .B(c[71]), .Z(n41364) );
  XOR U44302 ( .A(n41365), .B(n41366), .Z(n41357) );
  ANDN U44303 ( .B(n41367), .A(n30886), .Z(n41365) );
  XNOR U44304 ( .A(\modmult_1/zin[0][69] ), .B(n41368), .Z(n30886) );
  IV U44305 ( .A(n41366), .Z(n41368) );
  XOR U44306 ( .A(n41366), .B(n30887), .Z(n41367) );
  XNOR U44307 ( .A(n41369), .B(n41370), .Z(n30887) );
  ANDN U44308 ( .B(\modmult_1/xin[1023] ), .A(n41371), .Z(n41369) );
  IV U44309 ( .A(n41370), .Z(n41371) );
  XNOR U44310 ( .A(m[70]), .B(n41372), .Z(n41370) );
  NAND U44311 ( .A(n41373), .B(mul_pow), .Z(n41372) );
  XOR U44312 ( .A(m[70]), .B(c[70]), .Z(n41373) );
  XOR U44313 ( .A(n41374), .B(n41375), .Z(n41366) );
  ANDN U44314 ( .B(n41376), .A(n30884), .Z(n41374) );
  XNOR U44315 ( .A(\modmult_1/zin[0][68] ), .B(n41377), .Z(n30884) );
  IV U44316 ( .A(n41375), .Z(n41377) );
  XOR U44317 ( .A(n41375), .B(n30885), .Z(n41376) );
  XNOR U44318 ( .A(n41378), .B(n41379), .Z(n30885) );
  ANDN U44319 ( .B(\modmult_1/xin[1023] ), .A(n41380), .Z(n41378) );
  IV U44320 ( .A(n41379), .Z(n41380) );
  XNOR U44321 ( .A(m[69]), .B(n41381), .Z(n41379) );
  NAND U44322 ( .A(n41382), .B(mul_pow), .Z(n41381) );
  XOR U44323 ( .A(m[69]), .B(c[69]), .Z(n41382) );
  XOR U44324 ( .A(n41383), .B(n41384), .Z(n41375) );
  ANDN U44325 ( .B(n41385), .A(n30882), .Z(n41383) );
  XNOR U44326 ( .A(\modmult_1/zin[0][67] ), .B(n41386), .Z(n30882) );
  IV U44327 ( .A(n41384), .Z(n41386) );
  XOR U44328 ( .A(n41384), .B(n30883), .Z(n41385) );
  XNOR U44329 ( .A(n41387), .B(n41388), .Z(n30883) );
  ANDN U44330 ( .B(\modmult_1/xin[1023] ), .A(n41389), .Z(n41387) );
  IV U44331 ( .A(n41388), .Z(n41389) );
  XNOR U44332 ( .A(m[68]), .B(n41390), .Z(n41388) );
  NAND U44333 ( .A(n41391), .B(mul_pow), .Z(n41390) );
  XOR U44334 ( .A(m[68]), .B(c[68]), .Z(n41391) );
  XOR U44335 ( .A(n41392), .B(n41393), .Z(n41384) );
  ANDN U44336 ( .B(n41394), .A(n30880), .Z(n41392) );
  XNOR U44337 ( .A(\modmult_1/zin[0][66] ), .B(n41395), .Z(n30880) );
  IV U44338 ( .A(n41393), .Z(n41395) );
  XOR U44339 ( .A(n41393), .B(n30881), .Z(n41394) );
  XNOR U44340 ( .A(n41396), .B(n41397), .Z(n30881) );
  ANDN U44341 ( .B(\modmult_1/xin[1023] ), .A(n41398), .Z(n41396) );
  IV U44342 ( .A(n41397), .Z(n41398) );
  XNOR U44343 ( .A(m[67]), .B(n41399), .Z(n41397) );
  NAND U44344 ( .A(n41400), .B(mul_pow), .Z(n41399) );
  XOR U44345 ( .A(m[67]), .B(c[67]), .Z(n41400) );
  XOR U44346 ( .A(n41401), .B(n41402), .Z(n41393) );
  ANDN U44347 ( .B(n41403), .A(n30878), .Z(n41401) );
  XNOR U44348 ( .A(\modmult_1/zin[0][65] ), .B(n41404), .Z(n30878) );
  IV U44349 ( .A(n41402), .Z(n41404) );
  XOR U44350 ( .A(n41402), .B(n30879), .Z(n41403) );
  XNOR U44351 ( .A(n41405), .B(n41406), .Z(n30879) );
  ANDN U44352 ( .B(\modmult_1/xin[1023] ), .A(n41407), .Z(n41405) );
  IV U44353 ( .A(n41406), .Z(n41407) );
  XNOR U44354 ( .A(m[66]), .B(n41408), .Z(n41406) );
  NAND U44355 ( .A(n41409), .B(mul_pow), .Z(n41408) );
  XOR U44356 ( .A(m[66]), .B(c[66]), .Z(n41409) );
  XOR U44357 ( .A(n41410), .B(n41411), .Z(n41402) );
  ANDN U44358 ( .B(n41412), .A(n30876), .Z(n41410) );
  XNOR U44359 ( .A(\modmult_1/zin[0][64] ), .B(n41413), .Z(n30876) );
  IV U44360 ( .A(n41411), .Z(n41413) );
  XOR U44361 ( .A(n41411), .B(n30877), .Z(n41412) );
  XNOR U44362 ( .A(n41414), .B(n41415), .Z(n30877) );
  ANDN U44363 ( .B(\modmult_1/xin[1023] ), .A(n41416), .Z(n41414) );
  IV U44364 ( .A(n41415), .Z(n41416) );
  XNOR U44365 ( .A(m[65]), .B(n41417), .Z(n41415) );
  NAND U44366 ( .A(n41418), .B(mul_pow), .Z(n41417) );
  XOR U44367 ( .A(m[65]), .B(c[65]), .Z(n41418) );
  XOR U44368 ( .A(n41419), .B(n41420), .Z(n41411) );
  ANDN U44369 ( .B(n41421), .A(n30874), .Z(n41419) );
  XNOR U44370 ( .A(\modmult_1/zin[0][63] ), .B(n41422), .Z(n30874) );
  IV U44371 ( .A(n41420), .Z(n41422) );
  XOR U44372 ( .A(n41420), .B(n30875), .Z(n41421) );
  XNOR U44373 ( .A(n41423), .B(n41424), .Z(n30875) );
  ANDN U44374 ( .B(\modmult_1/xin[1023] ), .A(n41425), .Z(n41423) );
  IV U44375 ( .A(n41424), .Z(n41425) );
  XNOR U44376 ( .A(m[64]), .B(n41426), .Z(n41424) );
  NAND U44377 ( .A(n41427), .B(mul_pow), .Z(n41426) );
  XOR U44378 ( .A(m[64]), .B(c[64]), .Z(n41427) );
  XOR U44379 ( .A(n41428), .B(n41429), .Z(n41420) );
  ANDN U44380 ( .B(n41430), .A(n30872), .Z(n41428) );
  XNOR U44381 ( .A(\modmult_1/zin[0][62] ), .B(n41431), .Z(n30872) );
  IV U44382 ( .A(n41429), .Z(n41431) );
  XOR U44383 ( .A(n41429), .B(n30873), .Z(n41430) );
  XNOR U44384 ( .A(n41432), .B(n41433), .Z(n30873) );
  ANDN U44385 ( .B(\modmult_1/xin[1023] ), .A(n41434), .Z(n41432) );
  IV U44386 ( .A(n41433), .Z(n41434) );
  XNOR U44387 ( .A(m[63]), .B(n41435), .Z(n41433) );
  NAND U44388 ( .A(n41436), .B(mul_pow), .Z(n41435) );
  XOR U44389 ( .A(m[63]), .B(c[63]), .Z(n41436) );
  XOR U44390 ( .A(n41437), .B(n41438), .Z(n41429) );
  ANDN U44391 ( .B(n41439), .A(n30870), .Z(n41437) );
  XNOR U44392 ( .A(\modmult_1/zin[0][61] ), .B(n41440), .Z(n30870) );
  IV U44393 ( .A(n41438), .Z(n41440) );
  XOR U44394 ( .A(n41438), .B(n30871), .Z(n41439) );
  XNOR U44395 ( .A(n41441), .B(n41442), .Z(n30871) );
  ANDN U44396 ( .B(\modmult_1/xin[1023] ), .A(n41443), .Z(n41441) );
  IV U44397 ( .A(n41442), .Z(n41443) );
  XNOR U44398 ( .A(m[62]), .B(n41444), .Z(n41442) );
  NAND U44399 ( .A(n41445), .B(mul_pow), .Z(n41444) );
  XOR U44400 ( .A(m[62]), .B(c[62]), .Z(n41445) );
  XOR U44401 ( .A(n41446), .B(n41447), .Z(n41438) );
  ANDN U44402 ( .B(n41448), .A(n30868), .Z(n41446) );
  XNOR U44403 ( .A(\modmult_1/zin[0][60] ), .B(n41449), .Z(n30868) );
  IV U44404 ( .A(n41447), .Z(n41449) );
  XOR U44405 ( .A(n41447), .B(n30869), .Z(n41448) );
  XNOR U44406 ( .A(n41450), .B(n41451), .Z(n30869) );
  ANDN U44407 ( .B(\modmult_1/xin[1023] ), .A(n41452), .Z(n41450) );
  IV U44408 ( .A(n41451), .Z(n41452) );
  XNOR U44409 ( .A(m[61]), .B(n41453), .Z(n41451) );
  NAND U44410 ( .A(n41454), .B(mul_pow), .Z(n41453) );
  XOR U44411 ( .A(m[61]), .B(c[61]), .Z(n41454) );
  XOR U44412 ( .A(n41455), .B(n41456), .Z(n41447) );
  ANDN U44413 ( .B(n41457), .A(n30866), .Z(n41455) );
  XNOR U44414 ( .A(\modmult_1/zin[0][59] ), .B(n41458), .Z(n30866) );
  IV U44415 ( .A(n41456), .Z(n41458) );
  XOR U44416 ( .A(n41456), .B(n30867), .Z(n41457) );
  XNOR U44417 ( .A(n41459), .B(n41460), .Z(n30867) );
  ANDN U44418 ( .B(\modmult_1/xin[1023] ), .A(n41461), .Z(n41459) );
  IV U44419 ( .A(n41460), .Z(n41461) );
  XNOR U44420 ( .A(m[60]), .B(n41462), .Z(n41460) );
  NAND U44421 ( .A(n41463), .B(mul_pow), .Z(n41462) );
  XOR U44422 ( .A(m[60]), .B(c[60]), .Z(n41463) );
  XOR U44423 ( .A(n41464), .B(n41465), .Z(n41456) );
  ANDN U44424 ( .B(n41466), .A(n30864), .Z(n41464) );
  XNOR U44425 ( .A(\modmult_1/zin[0][58] ), .B(n41467), .Z(n30864) );
  IV U44426 ( .A(n41465), .Z(n41467) );
  XOR U44427 ( .A(n41465), .B(n30865), .Z(n41466) );
  XNOR U44428 ( .A(n41468), .B(n41469), .Z(n30865) );
  ANDN U44429 ( .B(\modmult_1/xin[1023] ), .A(n41470), .Z(n41468) );
  IV U44430 ( .A(n41469), .Z(n41470) );
  XNOR U44431 ( .A(m[59]), .B(n41471), .Z(n41469) );
  NAND U44432 ( .A(n41472), .B(mul_pow), .Z(n41471) );
  XOR U44433 ( .A(m[59]), .B(c[59]), .Z(n41472) );
  XOR U44434 ( .A(n41473), .B(n41474), .Z(n41465) );
  ANDN U44435 ( .B(n41475), .A(n30862), .Z(n41473) );
  XNOR U44436 ( .A(\modmult_1/zin[0][57] ), .B(n41476), .Z(n30862) );
  IV U44437 ( .A(n41474), .Z(n41476) );
  XOR U44438 ( .A(n41474), .B(n30863), .Z(n41475) );
  XNOR U44439 ( .A(n41477), .B(n41478), .Z(n30863) );
  ANDN U44440 ( .B(\modmult_1/xin[1023] ), .A(n41479), .Z(n41477) );
  IV U44441 ( .A(n41478), .Z(n41479) );
  XNOR U44442 ( .A(m[58]), .B(n41480), .Z(n41478) );
  NAND U44443 ( .A(n41481), .B(mul_pow), .Z(n41480) );
  XOR U44444 ( .A(m[58]), .B(c[58]), .Z(n41481) );
  XOR U44445 ( .A(n41482), .B(n41483), .Z(n41474) );
  ANDN U44446 ( .B(n41484), .A(n30860), .Z(n41482) );
  XNOR U44447 ( .A(\modmult_1/zin[0][56] ), .B(n41485), .Z(n30860) );
  IV U44448 ( .A(n41483), .Z(n41485) );
  XOR U44449 ( .A(n41483), .B(n30861), .Z(n41484) );
  XNOR U44450 ( .A(n41486), .B(n41487), .Z(n30861) );
  ANDN U44451 ( .B(\modmult_1/xin[1023] ), .A(n41488), .Z(n41486) );
  IV U44452 ( .A(n41487), .Z(n41488) );
  XNOR U44453 ( .A(m[57]), .B(n41489), .Z(n41487) );
  NAND U44454 ( .A(n41490), .B(mul_pow), .Z(n41489) );
  XOR U44455 ( .A(m[57]), .B(c[57]), .Z(n41490) );
  XOR U44456 ( .A(n41491), .B(n41492), .Z(n41483) );
  ANDN U44457 ( .B(n41493), .A(n30858), .Z(n41491) );
  XNOR U44458 ( .A(\modmult_1/zin[0][55] ), .B(n41494), .Z(n30858) );
  IV U44459 ( .A(n41492), .Z(n41494) );
  XOR U44460 ( .A(n41492), .B(n30859), .Z(n41493) );
  XNOR U44461 ( .A(n41495), .B(n41496), .Z(n30859) );
  ANDN U44462 ( .B(\modmult_1/xin[1023] ), .A(n41497), .Z(n41495) );
  IV U44463 ( .A(n41496), .Z(n41497) );
  XNOR U44464 ( .A(m[56]), .B(n41498), .Z(n41496) );
  NAND U44465 ( .A(n41499), .B(mul_pow), .Z(n41498) );
  XOR U44466 ( .A(m[56]), .B(c[56]), .Z(n41499) );
  XOR U44467 ( .A(n41500), .B(n41501), .Z(n41492) );
  ANDN U44468 ( .B(n41502), .A(n30856), .Z(n41500) );
  XNOR U44469 ( .A(\modmult_1/zin[0][54] ), .B(n41503), .Z(n30856) );
  IV U44470 ( .A(n41501), .Z(n41503) );
  XOR U44471 ( .A(n41501), .B(n30857), .Z(n41502) );
  XNOR U44472 ( .A(n41504), .B(n41505), .Z(n30857) );
  ANDN U44473 ( .B(\modmult_1/xin[1023] ), .A(n41506), .Z(n41504) );
  IV U44474 ( .A(n41505), .Z(n41506) );
  XNOR U44475 ( .A(m[55]), .B(n41507), .Z(n41505) );
  NAND U44476 ( .A(n41508), .B(mul_pow), .Z(n41507) );
  XOR U44477 ( .A(m[55]), .B(c[55]), .Z(n41508) );
  XOR U44478 ( .A(n41509), .B(n41510), .Z(n41501) );
  ANDN U44479 ( .B(n41511), .A(n30854), .Z(n41509) );
  XNOR U44480 ( .A(\modmult_1/zin[0][53] ), .B(n41512), .Z(n30854) );
  IV U44481 ( .A(n41510), .Z(n41512) );
  XOR U44482 ( .A(n41510), .B(n30855), .Z(n41511) );
  XNOR U44483 ( .A(n41513), .B(n41514), .Z(n30855) );
  ANDN U44484 ( .B(\modmult_1/xin[1023] ), .A(n41515), .Z(n41513) );
  IV U44485 ( .A(n41514), .Z(n41515) );
  XNOR U44486 ( .A(m[54]), .B(n41516), .Z(n41514) );
  NAND U44487 ( .A(n41517), .B(mul_pow), .Z(n41516) );
  XOR U44488 ( .A(m[54]), .B(c[54]), .Z(n41517) );
  XOR U44489 ( .A(n41518), .B(n41519), .Z(n41510) );
  ANDN U44490 ( .B(n41520), .A(n30852), .Z(n41518) );
  XNOR U44491 ( .A(\modmult_1/zin[0][52] ), .B(n41521), .Z(n30852) );
  IV U44492 ( .A(n41519), .Z(n41521) );
  XOR U44493 ( .A(n41519), .B(n30853), .Z(n41520) );
  XNOR U44494 ( .A(n41522), .B(n41523), .Z(n30853) );
  ANDN U44495 ( .B(\modmult_1/xin[1023] ), .A(n41524), .Z(n41522) );
  IV U44496 ( .A(n41523), .Z(n41524) );
  XNOR U44497 ( .A(m[53]), .B(n41525), .Z(n41523) );
  NAND U44498 ( .A(n41526), .B(mul_pow), .Z(n41525) );
  XOR U44499 ( .A(m[53]), .B(c[53]), .Z(n41526) );
  XOR U44500 ( .A(n41527), .B(n41528), .Z(n41519) );
  ANDN U44501 ( .B(n41529), .A(n30850), .Z(n41527) );
  XNOR U44502 ( .A(\modmult_1/zin[0][51] ), .B(n41530), .Z(n30850) );
  IV U44503 ( .A(n41528), .Z(n41530) );
  XOR U44504 ( .A(n41528), .B(n30851), .Z(n41529) );
  XNOR U44505 ( .A(n41531), .B(n41532), .Z(n30851) );
  ANDN U44506 ( .B(\modmult_1/xin[1023] ), .A(n41533), .Z(n41531) );
  IV U44507 ( .A(n41532), .Z(n41533) );
  XNOR U44508 ( .A(m[52]), .B(n41534), .Z(n41532) );
  NAND U44509 ( .A(n41535), .B(mul_pow), .Z(n41534) );
  XOR U44510 ( .A(m[52]), .B(c[52]), .Z(n41535) );
  XOR U44511 ( .A(n41536), .B(n41537), .Z(n41528) );
  ANDN U44512 ( .B(n41538), .A(n30848), .Z(n41536) );
  XNOR U44513 ( .A(\modmult_1/zin[0][50] ), .B(n41539), .Z(n30848) );
  IV U44514 ( .A(n41537), .Z(n41539) );
  XOR U44515 ( .A(n41537), .B(n30849), .Z(n41538) );
  XNOR U44516 ( .A(n41540), .B(n41541), .Z(n30849) );
  ANDN U44517 ( .B(\modmult_1/xin[1023] ), .A(n41542), .Z(n41540) );
  IV U44518 ( .A(n41541), .Z(n41542) );
  XNOR U44519 ( .A(m[51]), .B(n41543), .Z(n41541) );
  NAND U44520 ( .A(n41544), .B(mul_pow), .Z(n41543) );
  XOR U44521 ( .A(m[51]), .B(c[51]), .Z(n41544) );
  XOR U44522 ( .A(n41545), .B(n41546), .Z(n41537) );
  ANDN U44523 ( .B(n41547), .A(n30846), .Z(n41545) );
  XNOR U44524 ( .A(\modmult_1/zin[0][49] ), .B(n41548), .Z(n30846) );
  IV U44525 ( .A(n41546), .Z(n41548) );
  XOR U44526 ( .A(n41546), .B(n30847), .Z(n41547) );
  XNOR U44527 ( .A(n41549), .B(n41550), .Z(n30847) );
  ANDN U44528 ( .B(\modmult_1/xin[1023] ), .A(n41551), .Z(n41549) );
  IV U44529 ( .A(n41550), .Z(n41551) );
  XNOR U44530 ( .A(m[50]), .B(n41552), .Z(n41550) );
  NAND U44531 ( .A(n41553), .B(mul_pow), .Z(n41552) );
  XOR U44532 ( .A(m[50]), .B(c[50]), .Z(n41553) );
  XOR U44533 ( .A(n41554), .B(n41555), .Z(n41546) );
  ANDN U44534 ( .B(n41556), .A(n30844), .Z(n41554) );
  XNOR U44535 ( .A(\modmult_1/zin[0][48] ), .B(n41557), .Z(n30844) );
  IV U44536 ( .A(n41555), .Z(n41557) );
  XOR U44537 ( .A(n41555), .B(n30845), .Z(n41556) );
  XNOR U44538 ( .A(n41558), .B(n41559), .Z(n30845) );
  ANDN U44539 ( .B(\modmult_1/xin[1023] ), .A(n41560), .Z(n41558) );
  IV U44540 ( .A(n41559), .Z(n41560) );
  XNOR U44541 ( .A(m[49]), .B(n41561), .Z(n41559) );
  NAND U44542 ( .A(n41562), .B(mul_pow), .Z(n41561) );
  XOR U44543 ( .A(m[49]), .B(c[49]), .Z(n41562) );
  XOR U44544 ( .A(n41563), .B(n41564), .Z(n41555) );
  ANDN U44545 ( .B(n41565), .A(n30842), .Z(n41563) );
  XNOR U44546 ( .A(\modmult_1/zin[0][47] ), .B(n41566), .Z(n30842) );
  IV U44547 ( .A(n41564), .Z(n41566) );
  XOR U44548 ( .A(n41564), .B(n30843), .Z(n41565) );
  XNOR U44549 ( .A(n41567), .B(n41568), .Z(n30843) );
  ANDN U44550 ( .B(\modmult_1/xin[1023] ), .A(n41569), .Z(n41567) );
  IV U44551 ( .A(n41568), .Z(n41569) );
  XNOR U44552 ( .A(m[48]), .B(n41570), .Z(n41568) );
  NAND U44553 ( .A(n41571), .B(mul_pow), .Z(n41570) );
  XOR U44554 ( .A(m[48]), .B(c[48]), .Z(n41571) );
  XOR U44555 ( .A(n41572), .B(n41573), .Z(n41564) );
  ANDN U44556 ( .B(n41574), .A(n30840), .Z(n41572) );
  XNOR U44557 ( .A(\modmult_1/zin[0][46] ), .B(n41575), .Z(n30840) );
  IV U44558 ( .A(n41573), .Z(n41575) );
  XOR U44559 ( .A(n41573), .B(n30841), .Z(n41574) );
  XNOR U44560 ( .A(n41576), .B(n41577), .Z(n30841) );
  ANDN U44561 ( .B(\modmult_1/xin[1023] ), .A(n41578), .Z(n41576) );
  IV U44562 ( .A(n41577), .Z(n41578) );
  XNOR U44563 ( .A(m[47]), .B(n41579), .Z(n41577) );
  NAND U44564 ( .A(n41580), .B(mul_pow), .Z(n41579) );
  XOR U44565 ( .A(m[47]), .B(c[47]), .Z(n41580) );
  XOR U44566 ( .A(n41581), .B(n41582), .Z(n41573) );
  ANDN U44567 ( .B(n41583), .A(n30838), .Z(n41581) );
  XNOR U44568 ( .A(\modmult_1/zin[0][45] ), .B(n41584), .Z(n30838) );
  IV U44569 ( .A(n41582), .Z(n41584) );
  XOR U44570 ( .A(n41582), .B(n30839), .Z(n41583) );
  XNOR U44571 ( .A(n41585), .B(n41586), .Z(n30839) );
  ANDN U44572 ( .B(\modmult_1/xin[1023] ), .A(n41587), .Z(n41585) );
  IV U44573 ( .A(n41586), .Z(n41587) );
  XNOR U44574 ( .A(m[46]), .B(n41588), .Z(n41586) );
  NAND U44575 ( .A(n41589), .B(mul_pow), .Z(n41588) );
  XOR U44576 ( .A(m[46]), .B(c[46]), .Z(n41589) );
  XOR U44577 ( .A(n41590), .B(n41591), .Z(n41582) );
  ANDN U44578 ( .B(n41592), .A(n30836), .Z(n41590) );
  XNOR U44579 ( .A(\modmult_1/zin[0][44] ), .B(n41593), .Z(n30836) );
  IV U44580 ( .A(n41591), .Z(n41593) );
  XOR U44581 ( .A(n41591), .B(n30837), .Z(n41592) );
  XNOR U44582 ( .A(n41594), .B(n41595), .Z(n30837) );
  ANDN U44583 ( .B(\modmult_1/xin[1023] ), .A(n41596), .Z(n41594) );
  IV U44584 ( .A(n41595), .Z(n41596) );
  XNOR U44585 ( .A(m[45]), .B(n41597), .Z(n41595) );
  NAND U44586 ( .A(n41598), .B(mul_pow), .Z(n41597) );
  XOR U44587 ( .A(m[45]), .B(c[45]), .Z(n41598) );
  XOR U44588 ( .A(n41599), .B(n41600), .Z(n41591) );
  ANDN U44589 ( .B(n41601), .A(n30834), .Z(n41599) );
  XNOR U44590 ( .A(\modmult_1/zin[0][43] ), .B(n41602), .Z(n30834) );
  IV U44591 ( .A(n41600), .Z(n41602) );
  XOR U44592 ( .A(n41600), .B(n30835), .Z(n41601) );
  XNOR U44593 ( .A(n41603), .B(n41604), .Z(n30835) );
  ANDN U44594 ( .B(\modmult_1/xin[1023] ), .A(n41605), .Z(n41603) );
  IV U44595 ( .A(n41604), .Z(n41605) );
  XNOR U44596 ( .A(m[44]), .B(n41606), .Z(n41604) );
  NAND U44597 ( .A(n41607), .B(mul_pow), .Z(n41606) );
  XOR U44598 ( .A(m[44]), .B(c[44]), .Z(n41607) );
  XOR U44599 ( .A(n41608), .B(n41609), .Z(n41600) );
  ANDN U44600 ( .B(n41610), .A(n30832), .Z(n41608) );
  XNOR U44601 ( .A(\modmult_1/zin[0][42] ), .B(n41611), .Z(n30832) );
  IV U44602 ( .A(n41609), .Z(n41611) );
  XOR U44603 ( .A(n41609), .B(n30833), .Z(n41610) );
  XNOR U44604 ( .A(n41612), .B(n41613), .Z(n30833) );
  ANDN U44605 ( .B(\modmult_1/xin[1023] ), .A(n41614), .Z(n41612) );
  IV U44606 ( .A(n41613), .Z(n41614) );
  XNOR U44607 ( .A(m[43]), .B(n41615), .Z(n41613) );
  NAND U44608 ( .A(n41616), .B(mul_pow), .Z(n41615) );
  XOR U44609 ( .A(m[43]), .B(c[43]), .Z(n41616) );
  XOR U44610 ( .A(n41617), .B(n41618), .Z(n41609) );
  ANDN U44611 ( .B(n41619), .A(n30830), .Z(n41617) );
  XNOR U44612 ( .A(\modmult_1/zin[0][41] ), .B(n41620), .Z(n30830) );
  IV U44613 ( .A(n41618), .Z(n41620) );
  XOR U44614 ( .A(n41618), .B(n30831), .Z(n41619) );
  XNOR U44615 ( .A(n41621), .B(n41622), .Z(n30831) );
  ANDN U44616 ( .B(\modmult_1/xin[1023] ), .A(n41623), .Z(n41621) );
  IV U44617 ( .A(n41622), .Z(n41623) );
  XNOR U44618 ( .A(m[42]), .B(n41624), .Z(n41622) );
  NAND U44619 ( .A(n41625), .B(mul_pow), .Z(n41624) );
  XOR U44620 ( .A(m[42]), .B(c[42]), .Z(n41625) );
  XOR U44621 ( .A(n41626), .B(n41627), .Z(n41618) );
  ANDN U44622 ( .B(n41628), .A(n30828), .Z(n41626) );
  XNOR U44623 ( .A(\modmult_1/zin[0][40] ), .B(n41629), .Z(n30828) );
  IV U44624 ( .A(n41627), .Z(n41629) );
  XOR U44625 ( .A(n41627), .B(n30829), .Z(n41628) );
  XNOR U44626 ( .A(n41630), .B(n41631), .Z(n30829) );
  ANDN U44627 ( .B(\modmult_1/xin[1023] ), .A(n41632), .Z(n41630) );
  IV U44628 ( .A(n41631), .Z(n41632) );
  XNOR U44629 ( .A(m[41]), .B(n41633), .Z(n41631) );
  NAND U44630 ( .A(n41634), .B(mul_pow), .Z(n41633) );
  XOR U44631 ( .A(m[41]), .B(c[41]), .Z(n41634) );
  XOR U44632 ( .A(n41635), .B(n41636), .Z(n41627) );
  ANDN U44633 ( .B(n41637), .A(n30826), .Z(n41635) );
  XNOR U44634 ( .A(\modmult_1/zin[0][39] ), .B(n41638), .Z(n30826) );
  IV U44635 ( .A(n41636), .Z(n41638) );
  XOR U44636 ( .A(n41636), .B(n30827), .Z(n41637) );
  XNOR U44637 ( .A(n41639), .B(n41640), .Z(n30827) );
  ANDN U44638 ( .B(\modmult_1/xin[1023] ), .A(n41641), .Z(n41639) );
  IV U44639 ( .A(n41640), .Z(n41641) );
  XNOR U44640 ( .A(m[40]), .B(n41642), .Z(n41640) );
  NAND U44641 ( .A(n41643), .B(mul_pow), .Z(n41642) );
  XOR U44642 ( .A(m[40]), .B(c[40]), .Z(n41643) );
  XOR U44643 ( .A(n41644), .B(n41645), .Z(n41636) );
  ANDN U44644 ( .B(n41646), .A(n30824), .Z(n41644) );
  XNOR U44645 ( .A(\modmult_1/zin[0][38] ), .B(n41647), .Z(n30824) );
  IV U44646 ( .A(n41645), .Z(n41647) );
  XOR U44647 ( .A(n41645), .B(n30825), .Z(n41646) );
  XNOR U44648 ( .A(n41648), .B(n41649), .Z(n30825) );
  ANDN U44649 ( .B(\modmult_1/xin[1023] ), .A(n41650), .Z(n41648) );
  IV U44650 ( .A(n41649), .Z(n41650) );
  XNOR U44651 ( .A(m[39]), .B(n41651), .Z(n41649) );
  NAND U44652 ( .A(n41652), .B(mul_pow), .Z(n41651) );
  XOR U44653 ( .A(m[39]), .B(c[39]), .Z(n41652) );
  XOR U44654 ( .A(n41653), .B(n41654), .Z(n41645) );
  ANDN U44655 ( .B(n41655), .A(n30822), .Z(n41653) );
  XNOR U44656 ( .A(\modmult_1/zin[0][37] ), .B(n41656), .Z(n30822) );
  IV U44657 ( .A(n41654), .Z(n41656) );
  XOR U44658 ( .A(n41654), .B(n30823), .Z(n41655) );
  XNOR U44659 ( .A(n41657), .B(n41658), .Z(n30823) );
  ANDN U44660 ( .B(\modmult_1/xin[1023] ), .A(n41659), .Z(n41657) );
  IV U44661 ( .A(n41658), .Z(n41659) );
  XNOR U44662 ( .A(m[38]), .B(n41660), .Z(n41658) );
  NAND U44663 ( .A(n41661), .B(mul_pow), .Z(n41660) );
  XOR U44664 ( .A(m[38]), .B(c[38]), .Z(n41661) );
  XOR U44665 ( .A(n41662), .B(n41663), .Z(n41654) );
  ANDN U44666 ( .B(n41664), .A(n30820), .Z(n41662) );
  XNOR U44667 ( .A(\modmult_1/zin[0][36] ), .B(n41665), .Z(n30820) );
  IV U44668 ( .A(n41663), .Z(n41665) );
  XOR U44669 ( .A(n41663), .B(n30821), .Z(n41664) );
  XNOR U44670 ( .A(n41666), .B(n41667), .Z(n30821) );
  ANDN U44671 ( .B(\modmult_1/xin[1023] ), .A(n41668), .Z(n41666) );
  IV U44672 ( .A(n41667), .Z(n41668) );
  XNOR U44673 ( .A(m[37]), .B(n41669), .Z(n41667) );
  NAND U44674 ( .A(n41670), .B(mul_pow), .Z(n41669) );
  XOR U44675 ( .A(m[37]), .B(c[37]), .Z(n41670) );
  XOR U44676 ( .A(n41671), .B(n41672), .Z(n41663) );
  ANDN U44677 ( .B(n41673), .A(n30818), .Z(n41671) );
  XNOR U44678 ( .A(\modmult_1/zin[0][35] ), .B(n41674), .Z(n30818) );
  IV U44679 ( .A(n41672), .Z(n41674) );
  XOR U44680 ( .A(n41672), .B(n30819), .Z(n41673) );
  XNOR U44681 ( .A(n41675), .B(n41676), .Z(n30819) );
  ANDN U44682 ( .B(\modmult_1/xin[1023] ), .A(n41677), .Z(n41675) );
  IV U44683 ( .A(n41676), .Z(n41677) );
  XNOR U44684 ( .A(m[36]), .B(n41678), .Z(n41676) );
  NAND U44685 ( .A(n41679), .B(mul_pow), .Z(n41678) );
  XOR U44686 ( .A(m[36]), .B(c[36]), .Z(n41679) );
  XOR U44687 ( .A(n41680), .B(n41681), .Z(n41672) );
  ANDN U44688 ( .B(n41682), .A(n30816), .Z(n41680) );
  XNOR U44689 ( .A(\modmult_1/zin[0][34] ), .B(n41683), .Z(n30816) );
  IV U44690 ( .A(n41681), .Z(n41683) );
  XOR U44691 ( .A(n41681), .B(n30817), .Z(n41682) );
  XNOR U44692 ( .A(n41684), .B(n41685), .Z(n30817) );
  ANDN U44693 ( .B(\modmult_1/xin[1023] ), .A(n41686), .Z(n41684) );
  IV U44694 ( .A(n41685), .Z(n41686) );
  XNOR U44695 ( .A(m[35]), .B(n41687), .Z(n41685) );
  NAND U44696 ( .A(n41688), .B(mul_pow), .Z(n41687) );
  XOR U44697 ( .A(m[35]), .B(c[35]), .Z(n41688) );
  XOR U44698 ( .A(n41689), .B(n41690), .Z(n41681) );
  ANDN U44699 ( .B(n41691), .A(n30814), .Z(n41689) );
  XNOR U44700 ( .A(\modmult_1/zin[0][33] ), .B(n41692), .Z(n30814) );
  IV U44701 ( .A(n41690), .Z(n41692) );
  XOR U44702 ( .A(n41690), .B(n30815), .Z(n41691) );
  XNOR U44703 ( .A(n41693), .B(n41694), .Z(n30815) );
  ANDN U44704 ( .B(\modmult_1/xin[1023] ), .A(n41695), .Z(n41693) );
  IV U44705 ( .A(n41694), .Z(n41695) );
  XNOR U44706 ( .A(m[34]), .B(n41696), .Z(n41694) );
  NAND U44707 ( .A(n41697), .B(mul_pow), .Z(n41696) );
  XOR U44708 ( .A(m[34]), .B(c[34]), .Z(n41697) );
  XOR U44709 ( .A(n41698), .B(n41699), .Z(n41690) );
  ANDN U44710 ( .B(n41700), .A(n30812), .Z(n41698) );
  XNOR U44711 ( .A(\modmult_1/zin[0][32] ), .B(n41701), .Z(n30812) );
  IV U44712 ( .A(n41699), .Z(n41701) );
  XOR U44713 ( .A(n41699), .B(n30813), .Z(n41700) );
  XNOR U44714 ( .A(n41702), .B(n41703), .Z(n30813) );
  ANDN U44715 ( .B(\modmult_1/xin[1023] ), .A(n41704), .Z(n41702) );
  IV U44716 ( .A(n41703), .Z(n41704) );
  XNOR U44717 ( .A(m[33]), .B(n41705), .Z(n41703) );
  NAND U44718 ( .A(n41706), .B(mul_pow), .Z(n41705) );
  XOR U44719 ( .A(m[33]), .B(c[33]), .Z(n41706) );
  XOR U44720 ( .A(n41707), .B(n41708), .Z(n41699) );
  ANDN U44721 ( .B(n41709), .A(n30810), .Z(n41707) );
  XNOR U44722 ( .A(\modmult_1/zin[0][31] ), .B(n41710), .Z(n30810) );
  IV U44723 ( .A(n41708), .Z(n41710) );
  XOR U44724 ( .A(n41708), .B(n30811), .Z(n41709) );
  XNOR U44725 ( .A(n41711), .B(n41712), .Z(n30811) );
  ANDN U44726 ( .B(\modmult_1/xin[1023] ), .A(n41713), .Z(n41711) );
  IV U44727 ( .A(n41712), .Z(n41713) );
  XNOR U44728 ( .A(m[32]), .B(n41714), .Z(n41712) );
  NAND U44729 ( .A(n41715), .B(mul_pow), .Z(n41714) );
  XOR U44730 ( .A(m[32]), .B(c[32]), .Z(n41715) );
  XOR U44731 ( .A(n41716), .B(n41717), .Z(n41708) );
  ANDN U44732 ( .B(n41718), .A(n30808), .Z(n41716) );
  XNOR U44733 ( .A(\modmult_1/zin[0][30] ), .B(n41719), .Z(n30808) );
  IV U44734 ( .A(n41717), .Z(n41719) );
  XOR U44735 ( .A(n41717), .B(n30809), .Z(n41718) );
  XNOR U44736 ( .A(n41720), .B(n41721), .Z(n30809) );
  ANDN U44737 ( .B(\modmult_1/xin[1023] ), .A(n41722), .Z(n41720) );
  IV U44738 ( .A(n41721), .Z(n41722) );
  XNOR U44739 ( .A(m[31]), .B(n41723), .Z(n41721) );
  NAND U44740 ( .A(n41724), .B(mul_pow), .Z(n41723) );
  XOR U44741 ( .A(m[31]), .B(c[31]), .Z(n41724) );
  XOR U44742 ( .A(n41725), .B(n41726), .Z(n41717) );
  ANDN U44743 ( .B(n41727), .A(n30806), .Z(n41725) );
  XNOR U44744 ( .A(\modmult_1/zin[0][29] ), .B(n41728), .Z(n30806) );
  IV U44745 ( .A(n41726), .Z(n41728) );
  XOR U44746 ( .A(n41726), .B(n30807), .Z(n41727) );
  XNOR U44747 ( .A(n41729), .B(n41730), .Z(n30807) );
  ANDN U44748 ( .B(\modmult_1/xin[1023] ), .A(n41731), .Z(n41729) );
  IV U44749 ( .A(n41730), .Z(n41731) );
  XNOR U44750 ( .A(m[30]), .B(n41732), .Z(n41730) );
  NAND U44751 ( .A(n41733), .B(mul_pow), .Z(n41732) );
  XOR U44752 ( .A(m[30]), .B(c[30]), .Z(n41733) );
  XOR U44753 ( .A(n41734), .B(n41735), .Z(n41726) );
  ANDN U44754 ( .B(n41736), .A(n30804), .Z(n41734) );
  XNOR U44755 ( .A(\modmult_1/zin[0][28] ), .B(n41737), .Z(n30804) );
  IV U44756 ( .A(n41735), .Z(n41737) );
  XOR U44757 ( .A(n41735), .B(n30805), .Z(n41736) );
  XNOR U44758 ( .A(n41738), .B(n41739), .Z(n30805) );
  ANDN U44759 ( .B(\modmult_1/xin[1023] ), .A(n41740), .Z(n41738) );
  IV U44760 ( .A(n41739), .Z(n41740) );
  XNOR U44761 ( .A(m[29]), .B(n41741), .Z(n41739) );
  NAND U44762 ( .A(n41742), .B(mul_pow), .Z(n41741) );
  XOR U44763 ( .A(m[29]), .B(c[29]), .Z(n41742) );
  XOR U44764 ( .A(n41743), .B(n41744), .Z(n41735) );
  ANDN U44765 ( .B(n41745), .A(n30802), .Z(n41743) );
  XNOR U44766 ( .A(\modmult_1/zin[0][27] ), .B(n41746), .Z(n30802) );
  IV U44767 ( .A(n41744), .Z(n41746) );
  XOR U44768 ( .A(n41744), .B(n30803), .Z(n41745) );
  XNOR U44769 ( .A(n41747), .B(n41748), .Z(n30803) );
  ANDN U44770 ( .B(\modmult_1/xin[1023] ), .A(n41749), .Z(n41747) );
  IV U44771 ( .A(n41748), .Z(n41749) );
  XNOR U44772 ( .A(m[28]), .B(n41750), .Z(n41748) );
  NAND U44773 ( .A(n41751), .B(mul_pow), .Z(n41750) );
  XOR U44774 ( .A(m[28]), .B(c[28]), .Z(n41751) );
  XOR U44775 ( .A(n41752), .B(n41753), .Z(n41744) );
  ANDN U44776 ( .B(n41754), .A(n30800), .Z(n41752) );
  XNOR U44777 ( .A(\modmult_1/zin[0][26] ), .B(n41755), .Z(n30800) );
  IV U44778 ( .A(n41753), .Z(n41755) );
  XOR U44779 ( .A(n41753), .B(n30801), .Z(n41754) );
  XNOR U44780 ( .A(n41756), .B(n41757), .Z(n30801) );
  ANDN U44781 ( .B(\modmult_1/xin[1023] ), .A(n41758), .Z(n41756) );
  IV U44782 ( .A(n41757), .Z(n41758) );
  XNOR U44783 ( .A(m[27]), .B(n41759), .Z(n41757) );
  NAND U44784 ( .A(n41760), .B(mul_pow), .Z(n41759) );
  XOR U44785 ( .A(m[27]), .B(c[27]), .Z(n41760) );
  XOR U44786 ( .A(n41761), .B(n41762), .Z(n41753) );
  ANDN U44787 ( .B(n41763), .A(n30798), .Z(n41761) );
  XNOR U44788 ( .A(\modmult_1/zin[0][25] ), .B(n41764), .Z(n30798) );
  IV U44789 ( .A(n41762), .Z(n41764) );
  XOR U44790 ( .A(n41762), .B(n30799), .Z(n41763) );
  XNOR U44791 ( .A(n41765), .B(n41766), .Z(n30799) );
  ANDN U44792 ( .B(\modmult_1/xin[1023] ), .A(n41767), .Z(n41765) );
  IV U44793 ( .A(n41766), .Z(n41767) );
  XNOR U44794 ( .A(m[26]), .B(n41768), .Z(n41766) );
  NAND U44795 ( .A(n41769), .B(mul_pow), .Z(n41768) );
  XOR U44796 ( .A(m[26]), .B(c[26]), .Z(n41769) );
  XOR U44797 ( .A(n41770), .B(n41771), .Z(n41762) );
  ANDN U44798 ( .B(n41772), .A(n30796), .Z(n41770) );
  XNOR U44799 ( .A(\modmult_1/zin[0][24] ), .B(n41773), .Z(n30796) );
  IV U44800 ( .A(n41771), .Z(n41773) );
  XOR U44801 ( .A(n41771), .B(n30797), .Z(n41772) );
  XNOR U44802 ( .A(n41774), .B(n41775), .Z(n30797) );
  ANDN U44803 ( .B(\modmult_1/xin[1023] ), .A(n41776), .Z(n41774) );
  IV U44804 ( .A(n41775), .Z(n41776) );
  XNOR U44805 ( .A(m[25]), .B(n41777), .Z(n41775) );
  NAND U44806 ( .A(n41778), .B(mul_pow), .Z(n41777) );
  XOR U44807 ( .A(m[25]), .B(c[25]), .Z(n41778) );
  XOR U44808 ( .A(n41779), .B(n41780), .Z(n41771) );
  ANDN U44809 ( .B(n41781), .A(n30794), .Z(n41779) );
  XNOR U44810 ( .A(\modmult_1/zin[0][23] ), .B(n41782), .Z(n30794) );
  IV U44811 ( .A(n41780), .Z(n41782) );
  XOR U44812 ( .A(n41780), .B(n30795), .Z(n41781) );
  XNOR U44813 ( .A(n41783), .B(n41784), .Z(n30795) );
  ANDN U44814 ( .B(\modmult_1/xin[1023] ), .A(n41785), .Z(n41783) );
  IV U44815 ( .A(n41784), .Z(n41785) );
  XNOR U44816 ( .A(m[24]), .B(n41786), .Z(n41784) );
  NAND U44817 ( .A(n41787), .B(mul_pow), .Z(n41786) );
  XOR U44818 ( .A(m[24]), .B(c[24]), .Z(n41787) );
  XOR U44819 ( .A(n41788), .B(n41789), .Z(n41780) );
  ANDN U44820 ( .B(n41790), .A(n30792), .Z(n41788) );
  XNOR U44821 ( .A(\modmult_1/zin[0][22] ), .B(n41791), .Z(n30792) );
  IV U44822 ( .A(n41789), .Z(n41791) );
  XOR U44823 ( .A(n41789), .B(n30793), .Z(n41790) );
  XNOR U44824 ( .A(n41792), .B(n41793), .Z(n30793) );
  ANDN U44825 ( .B(\modmult_1/xin[1023] ), .A(n41794), .Z(n41792) );
  IV U44826 ( .A(n41793), .Z(n41794) );
  XNOR U44827 ( .A(m[23]), .B(n41795), .Z(n41793) );
  NAND U44828 ( .A(n41796), .B(mul_pow), .Z(n41795) );
  XOR U44829 ( .A(m[23]), .B(c[23]), .Z(n41796) );
  XOR U44830 ( .A(n41797), .B(n41798), .Z(n41789) );
  ANDN U44831 ( .B(n41799), .A(n30790), .Z(n41797) );
  XNOR U44832 ( .A(\modmult_1/zin[0][21] ), .B(n41800), .Z(n30790) );
  IV U44833 ( .A(n41798), .Z(n41800) );
  XOR U44834 ( .A(n41798), .B(n30791), .Z(n41799) );
  XNOR U44835 ( .A(n41801), .B(n41802), .Z(n30791) );
  ANDN U44836 ( .B(\modmult_1/xin[1023] ), .A(n41803), .Z(n41801) );
  IV U44837 ( .A(n41802), .Z(n41803) );
  XNOR U44838 ( .A(m[22]), .B(n41804), .Z(n41802) );
  NAND U44839 ( .A(n41805), .B(mul_pow), .Z(n41804) );
  XOR U44840 ( .A(m[22]), .B(c[22]), .Z(n41805) );
  XOR U44841 ( .A(n41806), .B(n41807), .Z(n41798) );
  ANDN U44842 ( .B(n41808), .A(n30788), .Z(n41806) );
  XNOR U44843 ( .A(\modmult_1/zin[0][20] ), .B(n41809), .Z(n30788) );
  IV U44844 ( .A(n41807), .Z(n41809) );
  XOR U44845 ( .A(n41807), .B(n30789), .Z(n41808) );
  XNOR U44846 ( .A(n41810), .B(n41811), .Z(n30789) );
  ANDN U44847 ( .B(\modmult_1/xin[1023] ), .A(n41812), .Z(n41810) );
  IV U44848 ( .A(n41811), .Z(n41812) );
  XNOR U44849 ( .A(m[21]), .B(n41813), .Z(n41811) );
  NAND U44850 ( .A(n41814), .B(mul_pow), .Z(n41813) );
  XOR U44851 ( .A(m[21]), .B(c[21]), .Z(n41814) );
  XOR U44852 ( .A(n41815), .B(n41816), .Z(n41807) );
  ANDN U44853 ( .B(n41817), .A(n30786), .Z(n41815) );
  XNOR U44854 ( .A(\modmult_1/zin[0][19] ), .B(n41818), .Z(n30786) );
  IV U44855 ( .A(n41816), .Z(n41818) );
  XOR U44856 ( .A(n41816), .B(n30787), .Z(n41817) );
  XNOR U44857 ( .A(n41819), .B(n41820), .Z(n30787) );
  ANDN U44858 ( .B(\modmult_1/xin[1023] ), .A(n41821), .Z(n41819) );
  IV U44859 ( .A(n41820), .Z(n41821) );
  XNOR U44860 ( .A(m[20]), .B(n41822), .Z(n41820) );
  NAND U44861 ( .A(n41823), .B(mul_pow), .Z(n41822) );
  XOR U44862 ( .A(m[20]), .B(c[20]), .Z(n41823) );
  XOR U44863 ( .A(n41824), .B(n41825), .Z(n41816) );
  ANDN U44864 ( .B(n41826), .A(n30784), .Z(n41824) );
  XNOR U44865 ( .A(\modmult_1/zin[0][18] ), .B(n41827), .Z(n30784) );
  IV U44866 ( .A(n41825), .Z(n41827) );
  XOR U44867 ( .A(n41825), .B(n30785), .Z(n41826) );
  XNOR U44868 ( .A(n41828), .B(n41829), .Z(n30785) );
  ANDN U44869 ( .B(\modmult_1/xin[1023] ), .A(n41830), .Z(n41828) );
  IV U44870 ( .A(n41829), .Z(n41830) );
  XNOR U44871 ( .A(m[19]), .B(n41831), .Z(n41829) );
  NAND U44872 ( .A(n41832), .B(mul_pow), .Z(n41831) );
  XOR U44873 ( .A(m[19]), .B(c[19]), .Z(n41832) );
  XOR U44874 ( .A(n41833), .B(n41834), .Z(n41825) );
  ANDN U44875 ( .B(n41835), .A(n30782), .Z(n41833) );
  XNOR U44876 ( .A(\modmult_1/zin[0][17] ), .B(n41836), .Z(n30782) );
  IV U44877 ( .A(n41834), .Z(n41836) );
  XOR U44878 ( .A(n41834), .B(n30783), .Z(n41835) );
  XNOR U44879 ( .A(n41837), .B(n41838), .Z(n30783) );
  ANDN U44880 ( .B(\modmult_1/xin[1023] ), .A(n41839), .Z(n41837) );
  IV U44881 ( .A(n41838), .Z(n41839) );
  XNOR U44882 ( .A(m[18]), .B(n41840), .Z(n41838) );
  NAND U44883 ( .A(n41841), .B(mul_pow), .Z(n41840) );
  XOR U44884 ( .A(m[18]), .B(c[18]), .Z(n41841) );
  XOR U44885 ( .A(n41842), .B(n41843), .Z(n41834) );
  ANDN U44886 ( .B(n41844), .A(n30780), .Z(n41842) );
  XNOR U44887 ( .A(\modmult_1/zin[0][16] ), .B(n41845), .Z(n30780) );
  IV U44888 ( .A(n41843), .Z(n41845) );
  XOR U44889 ( .A(n41843), .B(n30781), .Z(n41844) );
  XNOR U44890 ( .A(n41846), .B(n41847), .Z(n30781) );
  ANDN U44891 ( .B(\modmult_1/xin[1023] ), .A(n41848), .Z(n41846) );
  IV U44892 ( .A(n41847), .Z(n41848) );
  XNOR U44893 ( .A(m[17]), .B(n41849), .Z(n41847) );
  NAND U44894 ( .A(n41850), .B(mul_pow), .Z(n41849) );
  XOR U44895 ( .A(m[17]), .B(c[17]), .Z(n41850) );
  XOR U44896 ( .A(n41851), .B(n41852), .Z(n41843) );
  ANDN U44897 ( .B(n41853), .A(n30778), .Z(n41851) );
  XNOR U44898 ( .A(\modmult_1/zin[0][15] ), .B(n41854), .Z(n30778) );
  IV U44899 ( .A(n41852), .Z(n41854) );
  XOR U44900 ( .A(n41852), .B(n30779), .Z(n41853) );
  XNOR U44901 ( .A(n41855), .B(n41856), .Z(n30779) );
  ANDN U44902 ( .B(\modmult_1/xin[1023] ), .A(n41857), .Z(n41855) );
  IV U44903 ( .A(n41856), .Z(n41857) );
  XNOR U44904 ( .A(m[16]), .B(n41858), .Z(n41856) );
  NAND U44905 ( .A(n41859), .B(mul_pow), .Z(n41858) );
  XOR U44906 ( .A(m[16]), .B(c[16]), .Z(n41859) );
  XOR U44907 ( .A(n41860), .B(n41861), .Z(n41852) );
  ANDN U44908 ( .B(n41862), .A(n30776), .Z(n41860) );
  XNOR U44909 ( .A(\modmult_1/zin[0][14] ), .B(n41863), .Z(n30776) );
  IV U44910 ( .A(n41861), .Z(n41863) );
  XOR U44911 ( .A(n41861), .B(n30777), .Z(n41862) );
  XNOR U44912 ( .A(n41864), .B(n41865), .Z(n30777) );
  ANDN U44913 ( .B(\modmult_1/xin[1023] ), .A(n41866), .Z(n41864) );
  IV U44914 ( .A(n41865), .Z(n41866) );
  XNOR U44915 ( .A(m[15]), .B(n41867), .Z(n41865) );
  NAND U44916 ( .A(n41868), .B(mul_pow), .Z(n41867) );
  XOR U44917 ( .A(m[15]), .B(c[15]), .Z(n41868) );
  XOR U44918 ( .A(n41869), .B(n41870), .Z(n41861) );
  ANDN U44919 ( .B(n41871), .A(n30774), .Z(n41869) );
  XNOR U44920 ( .A(\modmult_1/zin[0][13] ), .B(n41872), .Z(n30774) );
  IV U44921 ( .A(n41870), .Z(n41872) );
  XOR U44922 ( .A(n41870), .B(n30775), .Z(n41871) );
  XNOR U44923 ( .A(n41873), .B(n41874), .Z(n30775) );
  ANDN U44924 ( .B(\modmult_1/xin[1023] ), .A(n41875), .Z(n41873) );
  IV U44925 ( .A(n41874), .Z(n41875) );
  XNOR U44926 ( .A(m[14]), .B(n41876), .Z(n41874) );
  NAND U44927 ( .A(n41877), .B(mul_pow), .Z(n41876) );
  XOR U44928 ( .A(m[14]), .B(c[14]), .Z(n41877) );
  XOR U44929 ( .A(n41878), .B(n41879), .Z(n41870) );
  ANDN U44930 ( .B(n41880), .A(n30772), .Z(n41878) );
  XNOR U44931 ( .A(\modmult_1/zin[0][12] ), .B(n41881), .Z(n30772) );
  IV U44932 ( .A(n41879), .Z(n41881) );
  XOR U44933 ( .A(n41879), .B(n30773), .Z(n41880) );
  XNOR U44934 ( .A(n41882), .B(n41883), .Z(n30773) );
  ANDN U44935 ( .B(\modmult_1/xin[1023] ), .A(n41884), .Z(n41882) );
  IV U44936 ( .A(n41883), .Z(n41884) );
  XNOR U44937 ( .A(m[13]), .B(n41885), .Z(n41883) );
  NAND U44938 ( .A(n41886), .B(mul_pow), .Z(n41885) );
  XOR U44939 ( .A(m[13]), .B(c[13]), .Z(n41886) );
  XOR U44940 ( .A(n41887), .B(n41888), .Z(n41879) );
  ANDN U44941 ( .B(n41889), .A(n30770), .Z(n41887) );
  XNOR U44942 ( .A(\modmult_1/zin[0][11] ), .B(n41890), .Z(n30770) );
  IV U44943 ( .A(n41888), .Z(n41890) );
  XOR U44944 ( .A(n41888), .B(n30771), .Z(n41889) );
  XNOR U44945 ( .A(n41891), .B(n41892), .Z(n30771) );
  ANDN U44946 ( .B(\modmult_1/xin[1023] ), .A(n41893), .Z(n41891) );
  IV U44947 ( .A(n41892), .Z(n41893) );
  XNOR U44948 ( .A(m[12]), .B(n41894), .Z(n41892) );
  NAND U44949 ( .A(n41895), .B(mul_pow), .Z(n41894) );
  XOR U44950 ( .A(m[12]), .B(c[12]), .Z(n41895) );
  XOR U44951 ( .A(n41896), .B(n41897), .Z(n41888) );
  ANDN U44952 ( .B(n41898), .A(n30768), .Z(n41896) );
  XNOR U44953 ( .A(\modmult_1/zin[0][10] ), .B(n41899), .Z(n30768) );
  IV U44954 ( .A(n41897), .Z(n41899) );
  XOR U44955 ( .A(n41897), .B(n30769), .Z(n41898) );
  XNOR U44956 ( .A(n41900), .B(n41901), .Z(n30769) );
  ANDN U44957 ( .B(\modmult_1/xin[1023] ), .A(n41902), .Z(n41900) );
  IV U44958 ( .A(n41901), .Z(n41902) );
  XNOR U44959 ( .A(m[11]), .B(n41903), .Z(n41901) );
  NAND U44960 ( .A(n41904), .B(mul_pow), .Z(n41903) );
  XOR U44961 ( .A(m[11]), .B(c[11]), .Z(n41904) );
  XOR U44962 ( .A(n41905), .B(n41906), .Z(n41897) );
  ANDN U44963 ( .B(n41907), .A(n30766), .Z(n41905) );
  XNOR U44964 ( .A(\modmult_1/zin[0][9] ), .B(n41908), .Z(n30766) );
  IV U44965 ( .A(n41906), .Z(n41908) );
  XOR U44966 ( .A(n41906), .B(n30767), .Z(n41907) );
  XNOR U44967 ( .A(n41909), .B(n41910), .Z(n30767) );
  ANDN U44968 ( .B(\modmult_1/xin[1023] ), .A(n41911), .Z(n41909) );
  IV U44969 ( .A(n41910), .Z(n41911) );
  XNOR U44970 ( .A(m[10]), .B(n41912), .Z(n41910) );
  NAND U44971 ( .A(n41913), .B(mul_pow), .Z(n41912) );
  XOR U44972 ( .A(m[10]), .B(c[10]), .Z(n41913) );
  XOR U44973 ( .A(n41914), .B(n41915), .Z(n41906) );
  ANDN U44974 ( .B(n41916), .A(n30764), .Z(n41914) );
  XNOR U44975 ( .A(\modmult_1/zin[0][8] ), .B(n41917), .Z(n30764) );
  IV U44976 ( .A(n41915), .Z(n41917) );
  XOR U44977 ( .A(n41915), .B(n30765), .Z(n41916) );
  XNOR U44978 ( .A(n41918), .B(n41919), .Z(n30765) );
  ANDN U44979 ( .B(\modmult_1/xin[1023] ), .A(n41920), .Z(n41918) );
  IV U44980 ( .A(n41919), .Z(n41920) );
  XNOR U44981 ( .A(m[9]), .B(n41921), .Z(n41919) );
  NAND U44982 ( .A(n41922), .B(mul_pow), .Z(n41921) );
  XOR U44983 ( .A(m[9]), .B(c[9]), .Z(n41922) );
  XOR U44984 ( .A(n41923), .B(n41924), .Z(n41915) );
  ANDN U44985 ( .B(n41925), .A(n30762), .Z(n41923) );
  XNOR U44986 ( .A(\modmult_1/zin[0][7] ), .B(n41926), .Z(n30762) );
  IV U44987 ( .A(n41924), .Z(n41926) );
  XOR U44988 ( .A(n41924), .B(n30763), .Z(n41925) );
  XNOR U44989 ( .A(n41927), .B(n41928), .Z(n30763) );
  ANDN U44990 ( .B(\modmult_1/xin[1023] ), .A(n41929), .Z(n41927) );
  IV U44991 ( .A(n41928), .Z(n41929) );
  XNOR U44992 ( .A(m[8]), .B(n41930), .Z(n41928) );
  NAND U44993 ( .A(n41931), .B(mul_pow), .Z(n41930) );
  XOR U44994 ( .A(m[8]), .B(c[8]), .Z(n41931) );
  XOR U44995 ( .A(n41932), .B(n41933), .Z(n41924) );
  ANDN U44996 ( .B(n41934), .A(n30760), .Z(n41932) );
  XNOR U44997 ( .A(\modmult_1/zin[0][6] ), .B(n41935), .Z(n30760) );
  IV U44998 ( .A(n41933), .Z(n41935) );
  XOR U44999 ( .A(n41933), .B(n30761), .Z(n41934) );
  XNOR U45000 ( .A(n41936), .B(n41937), .Z(n30761) );
  ANDN U45001 ( .B(\modmult_1/xin[1023] ), .A(n41938), .Z(n41936) );
  IV U45002 ( .A(n41937), .Z(n41938) );
  XNOR U45003 ( .A(m[7]), .B(n41939), .Z(n41937) );
  NAND U45004 ( .A(n41940), .B(mul_pow), .Z(n41939) );
  XOR U45005 ( .A(m[7]), .B(c[7]), .Z(n41940) );
  XOR U45006 ( .A(n41941), .B(n41942), .Z(n41933) );
  ANDN U45007 ( .B(n41943), .A(n30758), .Z(n41941) );
  XNOR U45008 ( .A(\modmult_1/zin[0][5] ), .B(n41944), .Z(n30758) );
  IV U45009 ( .A(n41942), .Z(n41944) );
  XOR U45010 ( .A(n41942), .B(n30759), .Z(n41943) );
  XNOR U45011 ( .A(n41945), .B(n41946), .Z(n30759) );
  ANDN U45012 ( .B(\modmult_1/xin[1023] ), .A(n41947), .Z(n41945) );
  IV U45013 ( .A(n41946), .Z(n41947) );
  XNOR U45014 ( .A(m[6]), .B(n41948), .Z(n41946) );
  NAND U45015 ( .A(n41949), .B(mul_pow), .Z(n41948) );
  XOR U45016 ( .A(m[6]), .B(c[6]), .Z(n41949) );
  XOR U45017 ( .A(n41950), .B(n41951), .Z(n41942) );
  ANDN U45018 ( .B(n41952), .A(n30756), .Z(n41950) );
  XNOR U45019 ( .A(\modmult_1/zin[0][4] ), .B(n41953), .Z(n30756) );
  IV U45020 ( .A(n41951), .Z(n41953) );
  XOR U45021 ( .A(n41951), .B(n30757), .Z(n41952) );
  XNOR U45022 ( .A(n41954), .B(n41955), .Z(n30757) );
  ANDN U45023 ( .B(\modmult_1/xin[1023] ), .A(n41956), .Z(n41954) );
  IV U45024 ( .A(n41955), .Z(n41956) );
  XNOR U45025 ( .A(m[5]), .B(n41957), .Z(n41955) );
  NAND U45026 ( .A(n41958), .B(mul_pow), .Z(n41957) );
  XOR U45027 ( .A(m[5]), .B(c[5]), .Z(n41958) );
  XOR U45028 ( .A(n41959), .B(n41960), .Z(n41951) );
  ANDN U45029 ( .B(n41961), .A(n30754), .Z(n41959) );
  XNOR U45030 ( .A(\modmult_1/zin[0][3] ), .B(n41962), .Z(n30754) );
  IV U45031 ( .A(n41960), .Z(n41962) );
  XOR U45032 ( .A(n41960), .B(n30755), .Z(n41961) );
  XNOR U45033 ( .A(n41963), .B(n41964), .Z(n30755) );
  ANDN U45034 ( .B(\modmult_1/xin[1023] ), .A(n41965), .Z(n41963) );
  IV U45035 ( .A(n41964), .Z(n41965) );
  XNOR U45036 ( .A(m[4]), .B(n41966), .Z(n41964) );
  NAND U45037 ( .A(n41967), .B(mul_pow), .Z(n41966) );
  XOR U45038 ( .A(m[4]), .B(c[4]), .Z(n41967) );
  XOR U45039 ( .A(n41968), .B(n41969), .Z(n41960) );
  ANDN U45040 ( .B(n41970), .A(n30752), .Z(n41968) );
  XOR U45041 ( .A(\modmult_1/zin[0][2] ), .B(n41969), .Z(n30752) );
  XOR U45042 ( .A(n41969), .B(n30753), .Z(n41970) );
  XNOR U45043 ( .A(n41971), .B(n41972), .Z(n30753) );
  ANDN U45044 ( .B(\modmult_1/xin[1023] ), .A(n41973), .Z(n41971) );
  IV U45045 ( .A(n41972), .Z(n41973) );
  XNOR U45046 ( .A(m[3]), .B(n41974), .Z(n41972) );
  NAND U45047 ( .A(n41975), .B(mul_pow), .Z(n41974) );
  XOR U45048 ( .A(m[3]), .B(c[3]), .Z(n41975) );
  XNOR U45049 ( .A(n41976), .B(n41977), .Z(n41969) );
  NAND U45050 ( .A(n41978), .B(n30750), .Z(n41977) );
  XOR U45051 ( .A(\modmult_1/zin[0][1] ), .B(n41979), .Z(n30750) );
  IV U45052 ( .A(n41976), .Z(n41979) );
  XOR U45053 ( .A(n41976), .B(n30751), .Z(n41978) );
  XNOR U45054 ( .A(n41980), .B(n41981), .Z(n30751) );
  ANDN U45055 ( .B(\modmult_1/xin[1023] ), .A(n41982), .Z(n41980) );
  IV U45056 ( .A(n41981), .Z(n41982) );
  XNOR U45057 ( .A(m[2]), .B(n41983), .Z(n41981) );
  NAND U45058 ( .A(n41984), .B(mul_pow), .Z(n41983) );
  XOR U45059 ( .A(m[2]), .B(c[2]), .Z(n41984) );
  NANDN U45060 ( .A(n30744), .B(\modmult_1/zin[0][0] ), .Z(n41976) );
  XNOR U45061 ( .A(n41985), .B(n41986), .Z(n30744) );
  ANDN U45062 ( .B(\modmult_1/xin[1023] ), .A(n41987), .Z(n41985) );
  IV U45063 ( .A(n41986), .Z(n41987) );
  XNOR U45064 ( .A(m[1]), .B(n41988), .Z(n41986) );
  NAND U45065 ( .A(n41989), .B(mul_pow), .Z(n41988) );
  XOR U45066 ( .A(m[1]), .B(c[1]), .Z(n41989) );
  NAND U45067 ( .A(n41990), .B(n41991), .Z(n3090) );
  NANDN U45068 ( .A(mul_pow), .B(first_one), .Z(n41991) );
  NAND U45069 ( .A(first_one), .B(ein[1023]), .Z(n41990) );
endmodule

