
module matrixMult_N_M_0_N3_M32 ( clk, rst, x, y, o );
  input [287:0] x;
  input [287:0] y;
  output [287:0] o;
  input clk, rst;
  wire   \oijt[2][2][1][31] , \oijt[2][2][1][30] , \oijt[2][2][1][29] ,
         \oijt[2][2][1][28] , \oijt[2][2][1][27] , \oijt[2][2][1][26] ,
         \oijt[2][2][1][25] , \oijt[2][2][1][24] , \oijt[2][2][1][23] ,
         \oijt[2][2][1][22] , \oijt[2][2][1][21] , \oijt[2][2][1][20] ,
         \oijt[2][2][1][19] , \oijt[2][2][1][18] , \oijt[2][2][1][17] ,
         \oijt[2][2][1][16] , \oijt[2][2][1][15] , \oijt[2][2][1][14] ,
         \oijt[2][2][1][13] , \oijt[2][2][1][12] , \oijt[2][2][1][11] ,
         \oijt[2][2][1][10] , \oijt[2][2][1][9] , \oijt[2][2][1][8] ,
         \oijt[2][2][1][7] , \oijt[2][2][1][6] , \oijt[2][2][1][5] ,
         \oijt[2][2][1][4] , \oijt[2][2][1][3] , \oijt[2][2][1][2] ,
         \oijt[2][2][1][1] , \oijt[2][2][0][31] , \oijt[2][2][0][30] ,
         \oijt[2][2][0][29] , \oijt[2][2][0][28] , \oijt[2][2][0][27] ,
         \oijt[2][2][0][26] , \oijt[2][2][0][25] , \oijt[2][2][0][24] ,
         \oijt[2][2][0][23] , \oijt[2][2][0][22] , \oijt[2][2][0][21] ,
         \oijt[2][2][0][20] , \oijt[2][2][0][19] , \oijt[2][2][0][18] ,
         \oijt[2][2][0][17] , \oijt[2][2][0][16] , \oijt[2][2][0][15] ,
         \oijt[2][2][0][14] , \oijt[2][2][0][13] , \oijt[2][2][0][12] ,
         \oijt[2][2][0][11] , \oijt[2][2][0][10] , \oijt[2][2][0][9] ,
         \oijt[2][2][0][8] , \oijt[2][2][0][7] , \oijt[2][2][0][6] ,
         \oijt[2][2][0][5] , \oijt[2][2][0][4] , \oijt[2][2][0][3] ,
         \oijt[2][2][0][2] , \oijt[2][2][0][1] , \oijt[2][1][1][31] ,
         \oijt[2][1][1][30] , \oijt[2][1][1][29] , \oijt[2][1][1][28] ,
         \oijt[2][1][1][27] , \oijt[2][1][1][26] , \oijt[2][1][1][25] ,
         \oijt[2][1][1][24] , \oijt[2][1][1][23] , \oijt[2][1][1][22] ,
         \oijt[2][1][1][21] , \oijt[2][1][1][20] , \oijt[2][1][1][19] ,
         \oijt[2][1][1][18] , \oijt[2][1][1][17] , \oijt[2][1][1][16] ,
         \oijt[2][1][1][15] , \oijt[2][1][1][14] , \oijt[2][1][1][13] ,
         \oijt[2][1][1][12] , \oijt[2][1][1][11] , \oijt[2][1][1][10] ,
         \oijt[2][1][1][9] , \oijt[2][1][1][8] , \oijt[2][1][1][7] ,
         \oijt[2][1][1][6] , \oijt[2][1][1][5] , \oijt[2][1][1][4] ,
         \oijt[2][1][1][3] , \oijt[2][1][1][2] , \oijt[2][1][1][1] ,
         \oijt[2][1][0][31] , \oijt[2][1][0][30] , \oijt[2][1][0][29] ,
         \oijt[2][1][0][28] , \oijt[2][1][0][27] , \oijt[2][1][0][26] ,
         \oijt[2][1][0][25] , \oijt[2][1][0][24] , \oijt[2][1][0][23] ,
         \oijt[2][1][0][22] , \oijt[2][1][0][21] , \oijt[2][1][0][20] ,
         \oijt[2][1][0][19] , \oijt[2][1][0][18] , \oijt[2][1][0][17] ,
         \oijt[2][1][0][16] , \oijt[2][1][0][15] , \oijt[2][1][0][14] ,
         \oijt[2][1][0][13] , \oijt[2][1][0][12] , \oijt[2][1][0][11] ,
         \oijt[2][1][0][10] , \oijt[2][1][0][9] , \oijt[2][1][0][8] ,
         \oijt[2][1][0][7] , \oijt[2][1][0][6] , \oijt[2][1][0][5] ,
         \oijt[2][1][0][4] , \oijt[2][1][0][3] , \oijt[2][1][0][2] ,
         \oijt[2][1][0][1] , \oijt[2][0][1][31] , \oijt[2][0][1][30] ,
         \oijt[2][0][1][29] , \oijt[2][0][1][28] , \oijt[2][0][1][27] ,
         \oijt[2][0][1][26] , \oijt[2][0][1][25] , \oijt[2][0][1][24] ,
         \oijt[2][0][1][23] , \oijt[2][0][1][22] , \oijt[2][0][1][21] ,
         \oijt[2][0][1][20] , \oijt[2][0][1][19] , \oijt[2][0][1][18] ,
         \oijt[2][0][1][17] , \oijt[2][0][1][16] , \oijt[2][0][1][15] ,
         \oijt[2][0][1][14] , \oijt[2][0][1][13] , \oijt[2][0][1][12] ,
         \oijt[2][0][1][11] , \oijt[2][0][1][10] , \oijt[2][0][1][9] ,
         \oijt[2][0][1][8] , \oijt[2][0][1][7] , \oijt[2][0][1][6] ,
         \oijt[2][0][1][5] , \oijt[2][0][1][4] , \oijt[2][0][1][3] ,
         \oijt[2][0][1][2] , \oijt[2][0][1][1] , \oijt[2][0][0][31] ,
         \oijt[2][0][0][30] , \oijt[2][0][0][29] , \oijt[2][0][0][28] ,
         \oijt[2][0][0][27] , \oijt[2][0][0][26] , \oijt[2][0][0][25] ,
         \oijt[2][0][0][24] , \oijt[2][0][0][23] , \oijt[2][0][0][22] ,
         \oijt[2][0][0][21] , \oijt[2][0][0][20] , \oijt[2][0][0][19] ,
         \oijt[2][0][0][18] , \oijt[2][0][0][17] , \oijt[2][0][0][16] ,
         \oijt[2][0][0][15] , \oijt[2][0][0][14] , \oijt[2][0][0][13] ,
         \oijt[2][0][0][12] , \oijt[2][0][0][11] , \oijt[2][0][0][10] ,
         \oijt[2][0][0][9] , \oijt[2][0][0][8] , \oijt[2][0][0][7] ,
         \oijt[2][0][0][6] , \oijt[2][0][0][5] , \oijt[2][0][0][4] ,
         \oijt[2][0][0][3] , \oijt[2][0][0][2] , \oijt[2][0][0][1] ,
         \oijt[1][2][1][31] , \oijt[1][2][1][30] , \oijt[1][2][1][29] ,
         \oijt[1][2][1][28] , \oijt[1][2][1][27] , \oijt[1][2][1][26] ,
         \oijt[1][2][1][25] , \oijt[1][2][1][24] , \oijt[1][2][1][23] ,
         \oijt[1][2][1][22] , \oijt[1][2][1][21] , \oijt[1][2][1][20] ,
         \oijt[1][2][1][19] , \oijt[1][2][1][18] , \oijt[1][2][1][17] ,
         \oijt[1][2][1][16] , \oijt[1][2][1][15] , \oijt[1][2][1][14] ,
         \oijt[1][2][1][13] , \oijt[1][2][1][12] , \oijt[1][2][1][11] ,
         \oijt[1][2][1][10] , \oijt[1][2][1][9] , \oijt[1][2][1][8] ,
         \oijt[1][2][1][7] , \oijt[1][2][1][6] , \oijt[1][2][1][5] ,
         \oijt[1][2][1][4] , \oijt[1][2][1][3] , \oijt[1][2][1][2] ,
         \oijt[1][2][1][1] , \oijt[1][2][0][31] , \oijt[1][2][0][30] ,
         \oijt[1][2][0][29] , \oijt[1][2][0][28] , \oijt[1][2][0][27] ,
         \oijt[1][2][0][26] , \oijt[1][2][0][25] , \oijt[1][2][0][24] ,
         \oijt[1][2][0][23] , \oijt[1][2][0][22] , \oijt[1][2][0][21] ,
         \oijt[1][2][0][20] , \oijt[1][2][0][19] , \oijt[1][2][0][18] ,
         \oijt[1][2][0][17] , \oijt[1][2][0][16] , \oijt[1][2][0][15] ,
         \oijt[1][2][0][14] , \oijt[1][2][0][13] , \oijt[1][2][0][12] ,
         \oijt[1][2][0][11] , \oijt[1][2][0][10] , \oijt[1][2][0][9] ,
         \oijt[1][2][0][8] , \oijt[1][2][0][7] , \oijt[1][2][0][6] ,
         \oijt[1][2][0][5] , \oijt[1][2][0][4] , \oijt[1][2][0][3] ,
         \oijt[1][2][0][2] , \oijt[1][2][0][1] , \oijt[1][1][1][31] ,
         \oijt[1][1][1][30] , \oijt[1][1][1][29] , \oijt[1][1][1][28] ,
         \oijt[1][1][1][27] , \oijt[1][1][1][26] , \oijt[1][1][1][25] ,
         \oijt[1][1][1][24] , \oijt[1][1][1][23] , \oijt[1][1][1][22] ,
         \oijt[1][1][1][21] , \oijt[1][1][1][20] , \oijt[1][1][1][19] ,
         \oijt[1][1][1][18] , \oijt[1][1][1][17] , \oijt[1][1][1][16] ,
         \oijt[1][1][1][15] , \oijt[1][1][1][14] , \oijt[1][1][1][13] ,
         \oijt[1][1][1][12] , \oijt[1][1][1][11] , \oijt[1][1][1][10] ,
         \oijt[1][1][1][9] , \oijt[1][1][1][8] , \oijt[1][1][1][7] ,
         \oijt[1][1][1][6] , \oijt[1][1][1][5] , \oijt[1][1][1][4] ,
         \oijt[1][1][1][3] , \oijt[1][1][1][2] , \oijt[1][1][1][1] ,
         \oijt[1][1][0][31] , \oijt[1][1][0][30] , \oijt[1][1][0][29] ,
         \oijt[1][1][0][28] , \oijt[1][1][0][27] , \oijt[1][1][0][26] ,
         \oijt[1][1][0][25] , \oijt[1][1][0][24] , \oijt[1][1][0][23] ,
         \oijt[1][1][0][22] , \oijt[1][1][0][21] , \oijt[1][1][0][20] ,
         \oijt[1][1][0][19] , \oijt[1][1][0][18] , \oijt[1][1][0][17] ,
         \oijt[1][1][0][16] , \oijt[1][1][0][15] , \oijt[1][1][0][14] ,
         \oijt[1][1][0][13] , \oijt[1][1][0][12] , \oijt[1][1][0][11] ,
         \oijt[1][1][0][10] , \oijt[1][1][0][9] , \oijt[1][1][0][8] ,
         \oijt[1][1][0][7] , \oijt[1][1][0][6] , \oijt[1][1][0][5] ,
         \oijt[1][1][0][4] , \oijt[1][1][0][3] , \oijt[1][1][0][2] ,
         \oijt[1][1][0][1] , \oijt[1][0][1][31] , \oijt[1][0][1][30] ,
         \oijt[1][0][1][29] , \oijt[1][0][1][28] , \oijt[1][0][1][27] ,
         \oijt[1][0][1][26] , \oijt[1][0][1][25] , \oijt[1][0][1][24] ,
         \oijt[1][0][1][23] , \oijt[1][0][1][22] , \oijt[1][0][1][21] ,
         \oijt[1][0][1][20] , \oijt[1][0][1][19] , \oijt[1][0][1][18] ,
         \oijt[1][0][1][17] , \oijt[1][0][1][16] , \oijt[1][0][1][15] ,
         \oijt[1][0][1][14] , \oijt[1][0][1][13] , \oijt[1][0][1][12] ,
         \oijt[1][0][1][11] , \oijt[1][0][1][10] , \oijt[1][0][1][9] ,
         \oijt[1][0][1][8] , \oijt[1][0][1][7] , \oijt[1][0][1][6] ,
         \oijt[1][0][1][5] , \oijt[1][0][1][4] , \oijt[1][0][1][3] ,
         \oijt[1][0][1][2] , \oijt[1][0][1][1] , \oijt[1][0][0][31] ,
         \oijt[1][0][0][30] , \oijt[1][0][0][29] , \oijt[1][0][0][28] ,
         \oijt[1][0][0][27] , \oijt[1][0][0][26] , \oijt[1][0][0][25] ,
         \oijt[1][0][0][24] , \oijt[1][0][0][23] , \oijt[1][0][0][22] ,
         \oijt[1][0][0][21] , \oijt[1][0][0][20] , \oijt[1][0][0][19] ,
         \oijt[1][0][0][18] , \oijt[1][0][0][17] , \oijt[1][0][0][16] ,
         \oijt[1][0][0][15] , \oijt[1][0][0][14] , \oijt[1][0][0][13] ,
         \oijt[1][0][0][12] , \oijt[1][0][0][11] , \oijt[1][0][0][10] ,
         \oijt[1][0][0][9] , \oijt[1][0][0][8] , \oijt[1][0][0][7] ,
         \oijt[1][0][0][6] , \oijt[1][0][0][5] , \oijt[1][0][0][4] ,
         \oijt[1][0][0][3] , \oijt[1][0][0][2] , \oijt[1][0][0][1] ,
         \oijt[0][2][1][31] , \oijt[0][2][1][30] , \oijt[0][2][1][29] ,
         \oijt[0][2][1][28] , \oijt[0][2][1][27] , \oijt[0][2][1][26] ,
         \oijt[0][2][1][25] , \oijt[0][2][1][24] , \oijt[0][2][1][23] ,
         \oijt[0][2][1][22] , \oijt[0][2][1][21] , \oijt[0][2][1][20] ,
         \oijt[0][2][1][19] , \oijt[0][2][1][18] , \oijt[0][2][1][17] ,
         \oijt[0][2][1][16] , \oijt[0][2][1][15] , \oijt[0][2][1][14] ,
         \oijt[0][2][1][13] , \oijt[0][2][1][12] , \oijt[0][2][1][11] ,
         \oijt[0][2][1][10] , \oijt[0][2][1][9] , \oijt[0][2][1][8] ,
         \oijt[0][2][1][7] , \oijt[0][2][1][6] , \oijt[0][2][1][5] ,
         \oijt[0][2][1][4] , \oijt[0][2][1][3] , \oijt[0][2][1][2] ,
         \oijt[0][2][1][1] , \oijt[0][2][0][31] , \oijt[0][2][0][30] ,
         \oijt[0][2][0][29] , \oijt[0][2][0][28] , \oijt[0][2][0][27] ,
         \oijt[0][2][0][26] , \oijt[0][2][0][25] , \oijt[0][2][0][24] ,
         \oijt[0][2][0][23] , \oijt[0][2][0][22] , \oijt[0][2][0][21] ,
         \oijt[0][2][0][20] , \oijt[0][2][0][19] , \oijt[0][2][0][18] ,
         \oijt[0][2][0][17] , \oijt[0][2][0][16] , \oijt[0][2][0][15] ,
         \oijt[0][2][0][14] , \oijt[0][2][0][13] , \oijt[0][2][0][12] ,
         \oijt[0][2][0][11] , \oijt[0][2][0][10] , \oijt[0][2][0][9] ,
         \oijt[0][2][0][8] , \oijt[0][2][0][7] , \oijt[0][2][0][6] ,
         \oijt[0][2][0][5] , \oijt[0][2][0][4] , \oijt[0][2][0][3] ,
         \oijt[0][2][0][2] , \oijt[0][2][0][1] , \oijt[0][1][1][31] ,
         \oijt[0][1][1][30] , \oijt[0][1][1][29] , \oijt[0][1][1][28] ,
         \oijt[0][1][1][27] , \oijt[0][1][1][26] , \oijt[0][1][1][25] ,
         \oijt[0][1][1][24] , \oijt[0][1][1][23] , \oijt[0][1][1][22] ,
         \oijt[0][1][1][21] , \oijt[0][1][1][20] , \oijt[0][1][1][19] ,
         \oijt[0][1][1][18] , \oijt[0][1][1][17] , \oijt[0][1][1][16] ,
         \oijt[0][1][1][15] , \oijt[0][1][1][14] , \oijt[0][1][1][13] ,
         \oijt[0][1][1][12] , \oijt[0][1][1][11] , \oijt[0][1][1][10] ,
         \oijt[0][1][1][9] , \oijt[0][1][1][8] , \oijt[0][1][1][7] ,
         \oijt[0][1][1][6] , \oijt[0][1][1][5] , \oijt[0][1][1][4] ,
         \oijt[0][1][1][3] , \oijt[0][1][1][2] , \oijt[0][1][1][1] ,
         \oijt[0][1][0][31] , \oijt[0][1][0][30] , \oijt[0][1][0][29] ,
         \oijt[0][1][0][28] , \oijt[0][1][0][27] , \oijt[0][1][0][26] ,
         \oijt[0][1][0][25] , \oijt[0][1][0][24] , \oijt[0][1][0][23] ,
         \oijt[0][1][0][22] , \oijt[0][1][0][21] , \oijt[0][1][0][20] ,
         \oijt[0][1][0][19] , \oijt[0][1][0][18] , \oijt[0][1][0][17] ,
         \oijt[0][1][0][16] , \oijt[0][1][0][15] , \oijt[0][1][0][14] ,
         \oijt[0][1][0][13] , \oijt[0][1][0][12] , \oijt[0][1][0][11] ,
         \oijt[0][1][0][10] , \oijt[0][1][0][9] , \oijt[0][1][0][8] ,
         \oijt[0][1][0][7] , \oijt[0][1][0][6] , \oijt[0][1][0][5] ,
         \oijt[0][1][0][4] , \oijt[0][1][0][3] , \oijt[0][1][0][2] ,
         \oijt[0][1][0][1] , \oijt[0][0][1][31] , \oijt[0][0][1][30] ,
         \oijt[0][0][1][29] , \oijt[0][0][1][28] , \oijt[0][0][1][27] ,
         \oijt[0][0][1][26] , \oijt[0][0][1][25] , \oijt[0][0][1][24] ,
         \oijt[0][0][1][23] , \oijt[0][0][1][22] , \oijt[0][0][1][21] ,
         \oijt[0][0][1][20] , \oijt[0][0][1][19] , \oijt[0][0][1][18] ,
         \oijt[0][0][1][17] , \oijt[0][0][1][16] , \oijt[0][0][1][15] ,
         \oijt[0][0][1][14] , \oijt[0][0][1][13] , \oijt[0][0][1][12] ,
         \oijt[0][0][1][11] , \oijt[0][0][1][10] , \oijt[0][0][1][9] ,
         \oijt[0][0][1][8] , \oijt[0][0][1][7] , \oijt[0][0][1][6] ,
         \oijt[0][0][1][5] , \oijt[0][0][1][4] , \oijt[0][0][1][3] ,
         \oijt[0][0][1][2] , \oijt[0][0][1][1] , \oijt[0][0][0][31] ,
         \oijt[0][0][0][30] , \oijt[0][0][0][29] , \oijt[0][0][0][28] ,
         \oijt[0][0][0][27] , \oijt[0][0][0][26] , \oijt[0][0][0][25] ,
         \oijt[0][0][0][24] , \oijt[0][0][0][23] , \oijt[0][0][0][22] ,
         \oijt[0][0][0][21] , \oijt[0][0][0][20] , \oijt[0][0][0][19] ,
         \oijt[0][0][0][18] , \oijt[0][0][0][17] , \oijt[0][0][0][16] ,
         \oijt[0][0][0][15] , \oijt[0][0][0][14] , \oijt[0][0][0][13] ,
         \oijt[0][0][0][12] , \oijt[0][0][0][11] , \oijt[0][0][0][10] ,
         \oijt[0][0][0][9] , \oijt[0][0][0][8] , \oijt[0][0][0][7] ,
         \oijt[0][0][0][6] , \oijt[0][0][0][5] , \oijt[0][0][0][4] ,
         \oijt[0][0][0][3] , \oijt[0][0][0][2] , \oijt[0][0][0][1] ,
         \_0_net_[31] , \_0_net_[30] , \_0_net_[29] , \_0_net_[28] ,
         \_0_net_[27] , \_0_net_[26] , \_0_net_[25] , \_0_net_[24] ,
         \_0_net_[23] , \_0_net_[22] , \_0_net_[21] , \_0_net_[20] ,
         \_0_net_[19] , \_0_net_[18] , \_0_net_[17] , \_0_net_[16] ,
         \_0_net_[15] , \_0_net_[14] , \_0_net_[13] , \_0_net_[12] ,
         \_0_net_[11] , \_0_net_[10] , \_0_net_[9] , \_0_net_[8] ,
         \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] , \_0_net_[3] ,
         \_0_net_[2] , \_0_net_[1] , \_4_net_[31] , \_4_net_[30] ,
         \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] ,
         \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] ,
         \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] ,
         \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] ,
         \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] ,
         \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] ,
         \_4_net_[4] , \_4_net_[3] , \_4_net_[2] , \_4_net_[1] , \_8_net_[31] ,
         \_8_net_[30] , \_8_net_[29] , \_8_net_[28] , \_8_net_[27] ,
         \_8_net_[26] , \_8_net_[25] , \_8_net_[24] , \_8_net_[23] ,
         \_8_net_[22] , \_8_net_[21] , \_8_net_[20] , \_8_net_[19] ,
         \_8_net_[18] , \_8_net_[17] , \_8_net_[16] , \_8_net_[15] ,
         \_8_net_[14] , \_8_net_[13] , \_8_net_[12] , \_8_net_[11] ,
         \_8_net_[10] , \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] ,
         \_8_net_[5] , \_8_net_[4] , \_8_net_[3] , \_8_net_[2] , \_8_net_[1] ,
         \_12_net_[31] , \_12_net_[30] , \_12_net_[29] , \_12_net_[28] ,
         \_12_net_[27] , \_12_net_[26] , \_12_net_[25] , \_12_net_[24] ,
         \_12_net_[23] , \_12_net_[22] , \_12_net_[21] , \_12_net_[20] ,
         \_12_net_[19] , \_12_net_[18] , \_12_net_[17] , \_12_net_[16] ,
         \_12_net_[15] , \_12_net_[14] , \_12_net_[13] , \_12_net_[12] ,
         \_12_net_[11] , \_12_net_[10] , \_12_net_[9] , \_12_net_[8] ,
         \_12_net_[7] , \_12_net_[6] , \_12_net_[5] , \_12_net_[4] ,
         \_12_net_[3] , \_12_net_[2] , \_12_net_[1] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_16_net_[8] , \_16_net_[7] ,
         \_16_net_[6] , \_16_net_[5] , \_16_net_[4] , \_16_net_[3] ,
         \_16_net_[2] , \_16_net_[1] , \_20_net_[31] , \_20_net_[30] ,
         \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] ,
         \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] ,
         \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] ,
         \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] ,
         \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , \_20_net_[10] ,
         \_20_net_[9] , \_20_net_[8] , \_20_net_[7] , \_20_net_[6] ,
         \_20_net_[5] , \_20_net_[4] , \_20_net_[3] , \_20_net_[2] ,
         \_20_net_[1] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_24_net_[12] , \_24_net_[11] , \_24_net_[10] , \_24_net_[9] ,
         \_24_net_[8] , \_24_net_[7] , \_24_net_[6] , \_24_net_[5] ,
         \_24_net_[4] , \_24_net_[3] , \_24_net_[2] , \_24_net_[1] ,
         \_28_net_[31] , \_28_net_[30] , \_28_net_[29] , \_28_net_[28] ,
         \_28_net_[27] , \_28_net_[26] , \_28_net_[25] , \_28_net_[24] ,
         \_28_net_[23] , \_28_net_[22] , \_28_net_[21] , \_28_net_[20] ,
         \_28_net_[19] , \_28_net_[18] , \_28_net_[17] , \_28_net_[16] ,
         \_28_net_[15] , \_28_net_[14] , \_28_net_[13] , \_28_net_[12] ,
         \_28_net_[11] , \_28_net_[10] , \_28_net_[9] , \_28_net_[8] ,
         \_28_net_[7] , \_28_net_[6] , \_28_net_[5] , \_28_net_[4] ,
         \_28_net_[3] , \_28_net_[2] , \_28_net_[1] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_32_net_[16] , \_32_net_[15] ,
         \_32_net_[14] , \_32_net_[13] , \_32_net_[12] , \_32_net_[11] ,
         \_32_net_[10] , \_32_net_[9] , \_32_net_[8] , \_32_net_[7] ,
         \_32_net_[6] , \_32_net_[5] , \_32_net_[4] , \_32_net_[3] ,
         \_32_net_[2] , \_32_net_[1] , \_36_net_[31] , \_36_net_[30] ,
         \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] ,
         \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] ,
         \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , \_36_net_[18] ,
         \_36_net_[17] , \_36_net_[16] , \_36_net_[15] , \_36_net_[14] ,
         \_36_net_[13] , \_36_net_[12] , \_36_net_[11] , \_36_net_[10] ,
         \_36_net_[9] , \_36_net_[8] , \_36_net_[7] , \_36_net_[6] ,
         \_36_net_[5] , \_36_net_[4] , \_36_net_[3] , \_36_net_[2] ,
         \_36_net_[1] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_40_net_[20] , \_40_net_[19] , \_40_net_[18] , \_40_net_[17] ,
         \_40_net_[16] , \_40_net_[15] , \_40_net_[14] , \_40_net_[13] ,
         \_40_net_[12] , \_40_net_[11] , \_40_net_[10] , \_40_net_[9] ,
         \_40_net_[8] , \_40_net_[7] , \_40_net_[6] , \_40_net_[5] ,
         \_40_net_[4] , \_40_net_[3] , \_40_net_[2] , \_40_net_[1] ,
         \_44_net_[31] , \_44_net_[30] , \_44_net_[29] , \_44_net_[28] ,
         \_44_net_[27] , \_44_net_[26] , \_44_net_[25] , \_44_net_[24] ,
         \_44_net_[23] , \_44_net_[22] , \_44_net_[21] , \_44_net_[20] ,
         \_44_net_[19] , \_44_net_[18] , \_44_net_[17] , \_44_net_[16] ,
         \_44_net_[15] , \_44_net_[14] , \_44_net_[13] , \_44_net_[12] ,
         \_44_net_[11] , \_44_net_[10] , \_44_net_[9] , \_44_net_[8] ,
         \_44_net_[7] , \_44_net_[6] , \_44_net_[5] , \_44_net_[4] ,
         \_44_net_[3] , \_44_net_[2] , \_44_net_[1] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_48_net_[24] , \_48_net_[23] ,
         \_48_net_[22] , \_48_net_[21] , \_48_net_[20] , \_48_net_[19] ,
         \_48_net_[18] , \_48_net_[17] , \_48_net_[16] , \_48_net_[15] ,
         \_48_net_[14] , \_48_net_[13] , \_48_net_[12] , \_48_net_[11] ,
         \_48_net_[10] , \_48_net_[9] , \_48_net_[8] , \_48_net_[7] ,
         \_48_net_[6] , \_48_net_[5] , \_48_net_[4] , \_48_net_[3] ,
         \_48_net_[2] , \_48_net_[1] , \_52_net_[31] , \_52_net_[30] ,
         \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , \_52_net_[26] ,
         \_52_net_[25] , \_52_net_[24] , \_52_net_[23] , \_52_net_[22] ,
         \_52_net_[21] , \_52_net_[20] , \_52_net_[19] , \_52_net_[18] ,
         \_52_net_[17] , \_52_net_[16] , \_52_net_[15] , \_52_net_[14] ,
         \_52_net_[13] , \_52_net_[12] , \_52_net_[11] , \_52_net_[10] ,
         \_52_net_[9] , \_52_net_[8] , \_52_net_[7] , \_52_net_[6] ,
         \_52_net_[5] , \_52_net_[4] , \_52_net_[3] , \_52_net_[2] ,
         \_52_net_[1] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_56_net_[28] , \_56_net_[27] , \_56_net_[26] , \_56_net_[25] ,
         \_56_net_[24] , \_56_net_[23] , \_56_net_[22] , \_56_net_[21] ,
         \_56_net_[20] , \_56_net_[19] , \_56_net_[18] , \_56_net_[17] ,
         \_56_net_[16] , \_56_net_[15] , \_56_net_[14] , \_56_net_[13] ,
         \_56_net_[12] , \_56_net_[11] , \_56_net_[10] , \_56_net_[9] ,
         \_56_net_[8] , \_56_net_[7] , \_56_net_[6] , \_56_net_[5] ,
         \_56_net_[4] , \_56_net_[3] , \_56_net_[2] , \_56_net_[1] ,
         \_60_net_[31] , \_60_net_[30] , \_60_net_[29] , \_60_net_[28] ,
         \_60_net_[27] , \_60_net_[26] , \_60_net_[25] , \_60_net_[24] ,
         \_60_net_[23] , \_60_net_[22] , \_60_net_[21] , \_60_net_[20] ,
         \_60_net_[19] , \_60_net_[18] , \_60_net_[17] , \_60_net_[16] ,
         \_60_net_[15] , \_60_net_[14] , \_60_net_[13] , \_60_net_[12] ,
         \_60_net_[11] , \_60_net_[10] , \_60_net_[9] , \_60_net_[8] ,
         \_60_net_[7] , \_60_net_[6] , \_60_net_[5] , \_60_net_[4] ,
         \_60_net_[3] , \_60_net_[2] , \_60_net_[1] , \_64_net_[31] ,
         \_64_net_[30] , \_64_net_[29] , \_64_net_[28] , \_64_net_[27] ,
         \_64_net_[26] , \_64_net_[25] , \_64_net_[24] , \_64_net_[23] ,
         \_64_net_[22] , \_64_net_[21] , \_64_net_[20] , \_64_net_[19] ,
         \_64_net_[18] , \_64_net_[17] , \_64_net_[16] , \_64_net_[15] ,
         \_64_net_[14] , \_64_net_[13] , \_64_net_[12] , \_64_net_[11] ,
         \_64_net_[10] , \_64_net_[9] , \_64_net_[8] , \_64_net_[7] ,
         \_64_net_[6] , \_64_net_[5] , \_64_net_[4] , \_64_net_[3] ,
         \_64_net_[2] , \_64_net_[1] , \_68_net_[31] , \_68_net_[30] ,
         \_68_net_[29] , \_68_net_[28] , \_68_net_[27] , \_68_net_[26] ,
         \_68_net_[25] , \_68_net_[24] , \_68_net_[23] , \_68_net_[22] ,
         \_68_net_[21] , \_68_net_[20] , \_68_net_[19] , \_68_net_[18] ,
         \_68_net_[17] , \_68_net_[16] , \_68_net_[15] , \_68_net_[14] ,
         \_68_net_[13] , \_68_net_[12] , \_68_net_[11] , \_68_net_[10] ,
         \_68_net_[9] , \_68_net_[8] , \_68_net_[7] , \_68_net_[6] ,
         \_68_net_[5] , \_68_net_[4] , \_68_net_[3] , \_68_net_[2] ,
         \_68_net_[1] , \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[1] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[31] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[30] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[29] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[28] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[27] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[26] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[25] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[24] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[23] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[22] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[21] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[20] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[19] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[18] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[17] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[16] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[15] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[14] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[13] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[12] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[11] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[10] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[9] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[8] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[7] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[6] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[5] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[4] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[3] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[2] ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[1] ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ,
         \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ;

  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][2][1][31] ), .Z(o[287]) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_68_net_[31] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][2][1][30] ), .Z(o[286]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][2][1][30] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_68_net_[30] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][2][1][29] ), .Z(o[285]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][2][1][29] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_68_net_[29] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][2][1][28] ), .Z(o[284]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][2][1][28] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_68_net_[28] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][2][1][27] ), .Z(o[283]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][2][1][27] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_68_net_[27] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][2][1][26] ), .Z(o[282]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][2][1][26] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_68_net_[26] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][2][1][25] ), .Z(o[281]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][2][1][25] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_68_net_[25] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][2][1][24] ), .Z(o[280]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][2][1][24] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_68_net_[24] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][2][1][23] ), .Z(o[279]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][2][1][23] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_68_net_[23] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][2][1][22] ), .Z(o[278]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][2][1][22] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_68_net_[22] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][2][1][21] ), .Z(o[277]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][2][1][21] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_68_net_[21] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][2][1][20] ), .Z(o[276]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][2][1][20] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_68_net_[20] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][2][1][19] ), .Z(o[275]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][2][1][19] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_68_net_[19] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][2][1][18] ), .Z(o[274]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][2][1][18] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_68_net_[18] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][2][1][17] ), .Z(o[273]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][2][1][17] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_68_net_[17] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][2][1][16] ), .Z(o[272]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][2][1][16] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_68_net_[16] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][2][1][15] ), .Z(o[271]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][2][1][15] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_68_net_[15] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][2][1][14] ), .Z(o[270]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][2][1][14] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_68_net_[14] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][2][1][13] ), .Z(o[269]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][2][1][13] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_68_net_[13] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][2][1][12] ), .Z(o[268]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][2][1][12] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_68_net_[12] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][2][1][11] ), .Z(o[267]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][2][1][11] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_68_net_[11] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][2][1][10] ), .Z(o[266]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][2][1][10] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_68_net_[10] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][2][1][9] ), .Z(o[265]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][2][1][9] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_68_net_[9] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][2][1][8] ), .Z(o[264]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][2][1][8] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_68_net_[8] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][2][1][7] ), .Z(o[263]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][2][1][7] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_68_net_[7] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][2][1][6] ), .Z(o[262]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][2][1][6] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_68_net_[6] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][2][1][5] ), .Z(o[261]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][2][1][5] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_68_net_[5] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][2][1][4] ), .Z(o[260]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][2][1][4] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_68_net_[4] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][2][1][3] ), .Z(o[259]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][2][1][3] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_68_net_[3] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][2][1][2] ), .Z(o[258]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][2][1][2] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_68_net_[2] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][2][1][1] ), .Z(o[257]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][2][1][1] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_68_net_[1] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[256]) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][2][0][31] ), .Z(\oijt[2][2][1][31] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_64_net_[31] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][2][0][30] ), .Z(\oijt[2][2][1][30] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][2][0][30] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_64_net_[30] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][2][0][29] ), .Z(\oijt[2][2][1][29] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][2][0][29] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_64_net_[29] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][2][0][28] ), .Z(\oijt[2][2][1][28] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][2][0][28] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_64_net_[28] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][2][0][27] ), .Z(\oijt[2][2][1][27] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][2][0][27] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_64_net_[27] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][2][0][26] ), .Z(\oijt[2][2][1][26] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][2][0][26] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_64_net_[26] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][2][0][25] ), .Z(\oijt[2][2][1][25] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][2][0][25] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_64_net_[25] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][2][0][24] ), .Z(\oijt[2][2][1][24] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][2][0][24] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_64_net_[24] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][2][0][23] ), .Z(\oijt[2][2][1][23] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][2][0][23] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_64_net_[23] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][2][0][22] ), .Z(\oijt[2][2][1][22] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][2][0][22] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_64_net_[22] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][2][0][21] ), .Z(\oijt[2][2][1][21] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][2][0][21] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_64_net_[21] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][2][0][20] ), .Z(\oijt[2][2][1][20] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][2][0][20] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_64_net_[20] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][2][0][19] ), .Z(\oijt[2][2][1][19] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][2][0][19] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_64_net_[19] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][2][0][18] ), .Z(\oijt[2][2][1][18] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][2][0][18] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_64_net_[18] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][2][0][17] ), .Z(\oijt[2][2][1][17] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][2][0][17] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_64_net_[17] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][2][0][16] ), .Z(\oijt[2][2][1][16] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][2][0][16] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_64_net_[16] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][2][0][15] ), .Z(\oijt[2][2][1][15] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][2][0][15] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_64_net_[15] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][2][0][14] ), .Z(\oijt[2][2][1][14] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][2][0][14] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_64_net_[14] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][2][0][13] ), .Z(\oijt[2][2][1][13] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][2][0][13] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_64_net_[13] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][2][0][12] ), .Z(\oijt[2][2][1][12] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][2][0][12] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_64_net_[12] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][2][0][11] ), .Z(\oijt[2][2][1][11] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][2][0][11] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_64_net_[11] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][2][0][10] ), .Z(\oijt[2][2][1][10] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][2][0][10] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_64_net_[10] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][2][0][9] ), .Z(\oijt[2][2][1][9] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][2][0][9] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_64_net_[9] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][2][0][8] ), .Z(\oijt[2][2][1][8] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][2][0][8] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_64_net_[8] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][2][0][7] ), .Z(\oijt[2][2][1][7] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][2][0][7] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_64_net_[7] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][2][0][6] ), .Z(\oijt[2][2][1][6] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][2][0][6] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_64_net_[6] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][2][0][5] ), .Z(\oijt[2][2][1][5] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][2][0][5] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_64_net_[5] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][2][0][4] ), .Z(\oijt[2][2][1][4] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][2][0][4] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_64_net_[4] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][2][0][3] ), .Z(\oijt[2][2][1][3] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][2][0][3] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_64_net_[3] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][2][0][2] ), .Z(\oijt[2][2][1][2] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][2][0][2] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_64_net_[2] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][2][0][1] ), .Z(\oijt[2][2][1][1] ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][2][0][1] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_64_net_[1] ), .B(\MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][1][1][31] ), .Z(o[255]) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_60_net_[31] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][1][1][30] ), .Z(o[254]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][1][1][30] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_60_net_[30] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][1][1][29] ), .Z(o[253]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][1][1][29] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_60_net_[29] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][1][1][28] ), .Z(o[252]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][1][1][28] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_60_net_[28] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][1][1][27] ), .Z(o[251]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][1][1][27] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_60_net_[27] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][1][1][26] ), .Z(o[250]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][1][1][26] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_60_net_[26] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][1][1][25] ), .Z(o[249]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][1][1][25] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_60_net_[25] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][1][1][24] ), .Z(o[248]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][1][1][24] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_60_net_[24] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][1][1][23] ), .Z(o[247]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][1][1][23] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_60_net_[23] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][1][1][22] ), .Z(o[246]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][1][1][22] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_60_net_[22] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][1][1][21] ), .Z(o[245]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][1][1][21] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_60_net_[21] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][1][1][20] ), .Z(o[244]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][1][1][20] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_60_net_[20] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][1][1][19] ), .Z(o[243]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][1][1][19] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_60_net_[19] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][1][1][18] ), .Z(o[242]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][1][1][18] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_60_net_[18] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][1][1][17] ), .Z(o[241]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][1][1][17] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_60_net_[17] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][1][1][16] ), .Z(o[240]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][1][1][16] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_60_net_[16] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][1][1][15] ), .Z(o[239]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][1][1][15] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_60_net_[15] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][1][1][14] ), .Z(o[238]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][1][1][14] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_60_net_[14] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][1][1][13] ), .Z(o[237]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][1][1][13] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_60_net_[13] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][1][1][12] ), .Z(o[236]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][1][1][12] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_60_net_[12] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][1][1][11] ), .Z(o[235]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][1][1][11] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_60_net_[11] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][1][1][10] ), .Z(o[234]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][1][1][10] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_60_net_[10] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][1][1][9] ), .Z(o[233]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][1][1][9] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_60_net_[9] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][1][1][8] ), .Z(o[232]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][1][1][8] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_60_net_[8] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][1][1][7] ), .Z(o[231]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][1][1][7] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_60_net_[7] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][1][1][6] ), .Z(o[230]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][1][1][6] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_60_net_[6] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][1][1][5] ), .Z(o[229]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][1][1][5] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_60_net_[5] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][1][1][4] ), .Z(o[228]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][1][1][4] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_60_net_[4] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][1][1][3] ), .Z(o[227]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][1][1][3] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_60_net_[3] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][1][1][2] ), .Z(o[226]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][1][1][2] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_60_net_[2] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][1][1][1] ), .Z(o[225]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][1][1][1] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_60_net_[1] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[224]) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][1][0][31] ), .Z(\oijt[2][1][1][31] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_56_net_[31] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][1][0][30] ), .Z(\oijt[2][1][1][30] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][1][0][30] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_56_net_[30] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][1][0][29] ), .Z(\oijt[2][1][1][29] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][1][0][29] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_56_net_[29] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][1][0][28] ), .Z(\oijt[2][1][1][28] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][1][0][28] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_56_net_[28] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][1][0][27] ), .Z(\oijt[2][1][1][27] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][1][0][27] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_56_net_[27] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][1][0][26] ), .Z(\oijt[2][1][1][26] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][1][0][26] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_56_net_[26] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][1][0][25] ), .Z(\oijt[2][1][1][25] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][1][0][25] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_56_net_[25] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][1][0][24] ), .Z(\oijt[2][1][1][24] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][1][0][24] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_56_net_[24] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][1][0][23] ), .Z(\oijt[2][1][1][23] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][1][0][23] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_56_net_[23] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][1][0][22] ), .Z(\oijt[2][1][1][22] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][1][0][22] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_56_net_[22] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][1][0][21] ), .Z(\oijt[2][1][1][21] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][1][0][21] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_56_net_[21] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][1][0][20] ), .Z(\oijt[2][1][1][20] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][1][0][20] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_56_net_[20] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][1][0][19] ), .Z(\oijt[2][1][1][19] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][1][0][19] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_56_net_[19] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][1][0][18] ), .Z(\oijt[2][1][1][18] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][1][0][18] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_56_net_[18] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][1][0][17] ), .Z(\oijt[2][1][1][17] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][1][0][17] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_56_net_[17] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][1][0][16] ), .Z(\oijt[2][1][1][16] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][1][0][16] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_56_net_[16] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][1][0][15] ), .Z(\oijt[2][1][1][15] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][1][0][15] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_56_net_[15] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][1][0][14] ), .Z(\oijt[2][1][1][14] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][1][0][14] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_56_net_[14] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][1][0][13] ), .Z(\oijt[2][1][1][13] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][1][0][13] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_56_net_[13] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][1][0][12] ), .Z(\oijt[2][1][1][12] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][1][0][12] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_56_net_[12] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][1][0][11] ), .Z(\oijt[2][1][1][11] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][1][0][11] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_56_net_[11] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][1][0][10] ), .Z(\oijt[2][1][1][10] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][1][0][10] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_56_net_[10] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][1][0][9] ), .Z(\oijt[2][1][1][9] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][1][0][9] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_56_net_[9] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][1][0][8] ), .Z(\oijt[2][1][1][8] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][1][0][8] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_56_net_[8] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][1][0][7] ), .Z(\oijt[2][1][1][7] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][1][0][7] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_56_net_[7] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][1][0][6] ), .Z(\oijt[2][1][1][6] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][1][0][6] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_56_net_[6] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][1][0][5] ), .Z(\oijt[2][1][1][5] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][1][0][5] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_56_net_[5] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][1][0][4] ), .Z(\oijt[2][1][1][4] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][1][0][4] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_56_net_[4] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][1][0][3] ), .Z(\oijt[2][1][1][3] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][1][0][3] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_56_net_[3] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][1][0][2] ), .Z(\oijt[2][1][1][2] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][1][0][2] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_56_net_[2] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][1][0][1] ), .Z(\oijt[2][1][1][1] ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][1][0][1] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_56_net_[1] ), .B(\MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][0][1][31] ), .Z(o[223]) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_52_net_[31] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][0][1][30] ), .Z(o[222]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][0][1][30] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_52_net_[30] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][0][1][29] ), .Z(o[221]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][0][1][29] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_52_net_[29] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][0][1][28] ), .Z(o[220]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][0][1][28] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_52_net_[28] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][0][1][27] ), .Z(o[219]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][0][1][27] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_52_net_[27] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][0][1][26] ), .Z(o[218]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][0][1][26] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_52_net_[26] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][0][1][25] ), .Z(o[217]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][0][1][25] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_52_net_[25] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][0][1][24] ), .Z(o[216]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][0][1][24] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_52_net_[24] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][0][1][23] ), .Z(o[215]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][0][1][23] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_52_net_[23] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][0][1][22] ), .Z(o[214]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][0][1][22] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_52_net_[22] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][0][1][21] ), .Z(o[213]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][0][1][21] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_52_net_[21] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][0][1][20] ), .Z(o[212]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][0][1][20] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_52_net_[20] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][0][1][19] ), .Z(o[211]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][0][1][19] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_52_net_[19] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][0][1][18] ), .Z(o[210]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][0][1][18] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_52_net_[18] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][0][1][17] ), .Z(o[209]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][0][1][17] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_52_net_[17] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][0][1][16] ), .Z(o[208]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][0][1][16] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_52_net_[16] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][0][1][15] ), .Z(o[207]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][0][1][15] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_52_net_[15] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][0][1][14] ), .Z(o[206]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][0][1][14] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_52_net_[14] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][0][1][13] ), .Z(o[205]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][0][1][13] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_52_net_[13] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][0][1][12] ), .Z(o[204]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][0][1][12] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_52_net_[12] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][0][1][11] ), .Z(o[203]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][0][1][11] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_52_net_[11] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][0][1][10] ), .Z(o[202]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][0][1][10] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_52_net_[10] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][0][1][9] ), .Z(o[201]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][0][1][9] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_52_net_[9] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][0][1][8] ), .Z(o[200]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][0][1][8] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_52_net_[8] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][0][1][7] ), .Z(o[199]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][0][1][7] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_52_net_[7] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][0][1][6] ), .Z(o[198]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][0][1][6] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_52_net_[6] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][0][1][5] ), .Z(o[197]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][0][1][5] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_52_net_[5] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][0][1][4] ), .Z(o[196]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][0][1][4] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_52_net_[4] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][0][1][3] ), .Z(o[195]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][0][1][3] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_52_net_[3] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][0][1][2] ), .Z(o[194]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][0][1][2] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_52_net_[2] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][0][1][1] ), .Z(o[193]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][0][1][1] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_52_net_[1] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[192]) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[2][0][0][31] ), .Z(\oijt[2][0][1][31] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_48_net_[31] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[2][0][0][30] ), .Z(\oijt[2][0][1][30] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[2][0][0][30] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_48_net_[30] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[2][0][0][29] ), .Z(\oijt[2][0][1][29] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[2][0][0][29] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_48_net_[29] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[2][0][0][28] ), .Z(\oijt[2][0][1][28] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[2][0][0][28] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_48_net_[28] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[2][0][0][27] ), .Z(\oijt[2][0][1][27] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[2][0][0][27] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_48_net_[27] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[2][0][0][26] ), .Z(\oijt[2][0][1][26] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[2][0][0][26] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_48_net_[26] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[2][0][0][25] ), .Z(\oijt[2][0][1][25] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[2][0][0][25] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_48_net_[25] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[2][0][0][24] ), .Z(\oijt[2][0][1][24] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[2][0][0][24] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_48_net_[24] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[2][0][0][23] ), .Z(\oijt[2][0][1][23] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[2][0][0][23] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_48_net_[23] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[2][0][0][22] ), .Z(\oijt[2][0][1][22] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[2][0][0][22] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_48_net_[22] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[2][0][0][21] ), .Z(\oijt[2][0][1][21] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[2][0][0][21] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_48_net_[21] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[2][0][0][20] ), .Z(\oijt[2][0][1][20] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[2][0][0][20] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_48_net_[20] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[2][0][0][19] ), .Z(\oijt[2][0][1][19] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[2][0][0][19] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_48_net_[19] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[2][0][0][18] ), .Z(\oijt[2][0][1][18] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[2][0][0][18] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_48_net_[18] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[2][0][0][17] ), .Z(\oijt[2][0][1][17] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[2][0][0][17] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_48_net_[17] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[2][0][0][16] ), .Z(\oijt[2][0][1][16] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[2][0][0][16] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_48_net_[16] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[2][0][0][15] ), .Z(\oijt[2][0][1][15] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[2][0][0][15] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_48_net_[15] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[2][0][0][14] ), .Z(\oijt[2][0][1][14] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[2][0][0][14] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_48_net_[14] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[2][0][0][13] ), .Z(\oijt[2][0][1][13] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[2][0][0][13] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_48_net_[13] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[2][0][0][12] ), .Z(\oijt[2][0][1][12] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[2][0][0][12] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_48_net_[12] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[2][0][0][11] ), .Z(\oijt[2][0][1][11] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[2][0][0][11] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_48_net_[11] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[2][0][0][10] ), .Z(\oijt[2][0][1][10] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[2][0][0][10] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_48_net_[10] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[2][0][0][9] ), .Z(\oijt[2][0][1][9] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[2][0][0][9] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_48_net_[9] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[2][0][0][8] ), .Z(\oijt[2][0][1][8] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[2][0][0][8] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_48_net_[8] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[2][0][0][7] ), .Z(\oijt[2][0][1][7] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[2][0][0][7] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_48_net_[7] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[2][0][0][6] ), .Z(\oijt[2][0][1][6] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[2][0][0][6] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_48_net_[6] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[2][0][0][5] ), .Z(\oijt[2][0][1][5] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[2][0][0][5] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_48_net_[5] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[2][0][0][4] ), .Z(\oijt[2][0][1][4] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[2][0][0][4] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_48_net_[4] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[2][0][0][3] ), .Z(\oijt[2][0][1][3] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[2][0][0][3] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_48_net_[3] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[2][0][0][2] ), .Z(\oijt[2][0][1][2] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[2][0][0][2] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_48_net_[2] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[2][0][0][1] ), .Z(\oijt[2][0][1][1] ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[2][0][0][1] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_48_net_[1] ), .B(\MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][2][1][31] ), .Z(o[191]) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_44_net_[31] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][2][1][30] ), .Z(o[190]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][2][1][30] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_44_net_[30] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][2][1][29] ), .Z(o[189]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][2][1][29] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_44_net_[29] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][2][1][28] ), .Z(o[188]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][2][1][28] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_44_net_[28] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][2][1][27] ), .Z(o[187]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][2][1][27] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_44_net_[27] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][2][1][26] ), .Z(o[186]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][2][1][26] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_44_net_[26] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][2][1][25] ), .Z(o[185]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][2][1][25] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_44_net_[25] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][2][1][24] ), .Z(o[184]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][2][1][24] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_44_net_[24] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][2][1][23] ), .Z(o[183]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][2][1][23] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_44_net_[23] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][2][1][22] ), .Z(o[182]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][2][1][22] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_44_net_[22] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][2][1][21] ), .Z(o[181]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][2][1][21] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_44_net_[21] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][2][1][20] ), .Z(o[180]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][2][1][20] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_44_net_[20] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][2][1][19] ), .Z(o[179]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][2][1][19] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_44_net_[19] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][2][1][18] ), .Z(o[178]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][2][1][18] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_44_net_[18] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][2][1][17] ), .Z(o[177]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][2][1][17] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_44_net_[17] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][2][1][16] ), .Z(o[176]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][2][1][16] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_44_net_[16] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][2][1][15] ), .Z(o[175]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][2][1][15] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_44_net_[15] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][2][1][14] ), .Z(o[174]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][2][1][14] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_44_net_[14] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][2][1][13] ), .Z(o[173]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][2][1][13] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_44_net_[13] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][2][1][12] ), .Z(o[172]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][2][1][12] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_44_net_[12] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][2][1][11] ), .Z(o[171]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][2][1][11] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_44_net_[11] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][2][1][10] ), .Z(o[170]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][2][1][10] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_44_net_[10] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][2][1][9] ), .Z(o[169]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][2][1][9] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_44_net_[9] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][2][1][8] ), .Z(o[168]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][2][1][8] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_44_net_[8] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][2][1][7] ), .Z(o[167]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][2][1][7] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_44_net_[7] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][2][1][6] ), .Z(o[166]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][2][1][6] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_44_net_[6] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][2][1][5] ), .Z(o[165]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][2][1][5] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_44_net_[5] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][2][1][4] ), .Z(o[164]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][2][1][4] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_44_net_[4] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][2][1][3] ), .Z(o[163]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][2][1][3] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_44_net_[3] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][2][1][2] ), .Z(o[162]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][2][1][2] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_44_net_[2] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][2][1][1] ), .Z(o[161]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][2][1][1] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_44_net_[1] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[160]) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][2][0][31] ), .Z(\oijt[1][2][1][31] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_40_net_[31] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][2][0][30] ), .Z(\oijt[1][2][1][30] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][2][0][30] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_40_net_[30] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][2][0][29] ), .Z(\oijt[1][2][1][29] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][2][0][29] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_40_net_[29] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][2][0][28] ), .Z(\oijt[1][2][1][28] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][2][0][28] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_40_net_[28] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][2][0][27] ), .Z(\oijt[1][2][1][27] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][2][0][27] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_40_net_[27] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][2][0][26] ), .Z(\oijt[1][2][1][26] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][2][0][26] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_40_net_[26] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][2][0][25] ), .Z(\oijt[1][2][1][25] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][2][0][25] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_40_net_[25] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][2][0][24] ), .Z(\oijt[1][2][1][24] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][2][0][24] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_40_net_[24] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][2][0][23] ), .Z(\oijt[1][2][1][23] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][2][0][23] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_40_net_[23] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][2][0][22] ), .Z(\oijt[1][2][1][22] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][2][0][22] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_40_net_[22] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][2][0][21] ), .Z(\oijt[1][2][1][21] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][2][0][21] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_40_net_[21] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][2][0][20] ), .Z(\oijt[1][2][1][20] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][2][0][20] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_40_net_[20] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][2][0][19] ), .Z(\oijt[1][2][1][19] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][2][0][19] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_40_net_[19] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][2][0][18] ), .Z(\oijt[1][2][1][18] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][2][0][18] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_40_net_[18] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][2][0][17] ), .Z(\oijt[1][2][1][17] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][2][0][17] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_40_net_[17] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][2][0][16] ), .Z(\oijt[1][2][1][16] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][2][0][16] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_40_net_[16] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][2][0][15] ), .Z(\oijt[1][2][1][15] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][2][0][15] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_40_net_[15] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][2][0][14] ), .Z(\oijt[1][2][1][14] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][2][0][14] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_40_net_[14] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][2][0][13] ), .Z(\oijt[1][2][1][13] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][2][0][13] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_40_net_[13] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][2][0][12] ), .Z(\oijt[1][2][1][12] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][2][0][12] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_40_net_[12] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][2][0][11] ), .Z(\oijt[1][2][1][11] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][2][0][11] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_40_net_[11] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][2][0][10] ), .Z(\oijt[1][2][1][10] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][2][0][10] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_40_net_[10] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][2][0][9] ), .Z(\oijt[1][2][1][9] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][2][0][9] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_40_net_[9] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][2][0][8] ), .Z(\oijt[1][2][1][8] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][2][0][8] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_40_net_[8] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][2][0][7] ), .Z(\oijt[1][2][1][7] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][2][0][7] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_40_net_[7] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][2][0][6] ), .Z(\oijt[1][2][1][6] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][2][0][6] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_40_net_[6] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][2][0][5] ), .Z(\oijt[1][2][1][5] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][2][0][5] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_40_net_[5] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][2][0][4] ), .Z(\oijt[1][2][1][4] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][2][0][4] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_40_net_[4] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][2][0][3] ), .Z(\oijt[1][2][1][3] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][2][0][3] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_40_net_[3] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][2][0][2] ), .Z(\oijt[1][2][1][2] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][2][0][2] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_40_net_[2] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][2][0][1] ), .Z(\oijt[1][2][1][1] ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][2][0][1] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_40_net_[1] ), .B(\MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][1][1][31] ), .Z(o[159]) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_36_net_[31] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][1][1][30] ), .Z(o[158]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][1][1][30] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_36_net_[30] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][1][1][29] ), .Z(o[157]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][1][1][29] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_36_net_[29] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][1][1][28] ), .Z(o[156]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][1][1][28] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_36_net_[28] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][1][1][27] ), .Z(o[155]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][1][1][27] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_36_net_[27] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][1][1][26] ), .Z(o[154]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][1][1][26] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_36_net_[26] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][1][1][25] ), .Z(o[153]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][1][1][25] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_36_net_[25] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][1][1][24] ), .Z(o[152]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][1][1][24] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_36_net_[24] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][1][1][23] ), .Z(o[151]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][1][1][23] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_36_net_[23] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][1][1][22] ), .Z(o[150]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][1][1][22] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_36_net_[22] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][1][1][21] ), .Z(o[149]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][1][1][21] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_36_net_[21] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][1][1][20] ), .Z(o[148]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][1][1][20] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_36_net_[20] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][1][1][19] ), .Z(o[147]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][1][1][19] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_36_net_[19] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][1][1][18] ), .Z(o[146]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][1][1][18] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_36_net_[18] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][1][1][17] ), .Z(o[145]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][1][1][17] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_36_net_[17] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][1][1][16] ), .Z(o[144]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][1][1][16] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_36_net_[16] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][1][1][15] ), .Z(o[143]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][1][1][15] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_36_net_[15] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][1][1][14] ), .Z(o[142]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][1][1][14] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_36_net_[14] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][1][1][13] ), .Z(o[141]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][1][1][13] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_36_net_[13] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][1][1][12] ), .Z(o[140]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][1][1][12] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_36_net_[12] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][1][1][11] ), .Z(o[139]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][1][1][11] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_36_net_[11] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][1][1][10] ), .Z(o[138]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][1][1][10] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_36_net_[10] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][1][1][9] ), .Z(o[137]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][1][1][9] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_36_net_[9] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][1][1][8] ), .Z(o[136]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][1][1][8] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_36_net_[8] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][1][1][7] ), .Z(o[135]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][1][1][7] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_36_net_[7] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][1][1][6] ), .Z(o[134]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][1][1][6] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_36_net_[6] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][1][1][5] ), .Z(o[133]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][1][1][5] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_36_net_[5] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][1][1][4] ), .Z(o[132]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][1][1][4] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_36_net_[4] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][1][1][3] ), .Z(o[131]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][1][1][3] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_36_net_[3] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][1][1][2] ), .Z(o[130]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][1][1][2] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_36_net_[2] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][1][1][1] ), .Z(o[129]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][1][1][1] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_36_net_[1] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[128]) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][1][0][31] ), .Z(\oijt[1][1][1][31] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_32_net_[31] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][1][0][30] ), .Z(\oijt[1][1][1][30] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][1][0][30] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_32_net_[30] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][1][0][29] ), .Z(\oijt[1][1][1][29] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][1][0][29] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_32_net_[29] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][1][0][28] ), .Z(\oijt[1][1][1][28] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][1][0][28] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_32_net_[28] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][1][0][27] ), .Z(\oijt[1][1][1][27] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][1][0][27] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_32_net_[27] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][1][0][26] ), .Z(\oijt[1][1][1][26] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][1][0][26] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_32_net_[26] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][1][0][25] ), .Z(\oijt[1][1][1][25] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][1][0][25] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_32_net_[25] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][1][0][24] ), .Z(\oijt[1][1][1][24] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][1][0][24] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_32_net_[24] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][1][0][23] ), .Z(\oijt[1][1][1][23] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][1][0][23] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_32_net_[23] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][1][0][22] ), .Z(\oijt[1][1][1][22] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][1][0][22] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_32_net_[22] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][1][0][21] ), .Z(\oijt[1][1][1][21] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][1][0][21] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_32_net_[21] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][1][0][20] ), .Z(\oijt[1][1][1][20] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][1][0][20] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_32_net_[20] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][1][0][19] ), .Z(\oijt[1][1][1][19] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][1][0][19] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_32_net_[19] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][1][0][18] ), .Z(\oijt[1][1][1][18] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][1][0][18] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_32_net_[18] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][1][0][17] ), .Z(\oijt[1][1][1][17] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][1][0][17] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_32_net_[17] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][1][0][16] ), .Z(\oijt[1][1][1][16] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][1][0][16] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_32_net_[16] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][1][0][15] ), .Z(\oijt[1][1][1][15] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][1][0][15] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_32_net_[15] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][1][0][14] ), .Z(\oijt[1][1][1][14] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][1][0][14] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_32_net_[14] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][1][0][13] ), .Z(\oijt[1][1][1][13] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][1][0][13] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_32_net_[13] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][1][0][12] ), .Z(\oijt[1][1][1][12] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][1][0][12] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_32_net_[12] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][1][0][11] ), .Z(\oijt[1][1][1][11] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][1][0][11] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_32_net_[11] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][1][0][10] ), .Z(\oijt[1][1][1][10] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][1][0][10] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_32_net_[10] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][1][0][9] ), .Z(\oijt[1][1][1][9] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][1][0][9] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_32_net_[9] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][1][0][8] ), .Z(\oijt[1][1][1][8] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][1][0][8] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_32_net_[8] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][1][0][7] ), .Z(\oijt[1][1][1][7] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][1][0][7] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_32_net_[7] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][1][0][6] ), .Z(\oijt[1][1][1][6] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][1][0][6] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_32_net_[6] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][1][0][5] ), .Z(\oijt[1][1][1][5] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][1][0][5] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_32_net_[5] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][1][0][4] ), .Z(\oijt[1][1][1][4] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][1][0][4] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_32_net_[4] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][1][0][3] ), .Z(\oijt[1][1][1][3] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][1][0][3] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_32_net_[3] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][1][0][2] ), .Z(\oijt[1][1][1][2] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][1][0][2] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_32_net_[2] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][1][0][1] ), .Z(\oijt[1][1][1][1] ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][1][0][1] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_32_net_[1] ), .B(\MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][0][1][31] ), .Z(o[127]) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_28_net_[31] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][0][1][30] ), .Z(o[126]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][0][1][30] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_28_net_[30] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][0][1][29] ), .Z(o[125]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][0][1][29] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_28_net_[29] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][0][1][28] ), .Z(o[124]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][0][1][28] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_28_net_[28] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][0][1][27] ), .Z(o[123]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][0][1][27] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_28_net_[27] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][0][1][26] ), .Z(o[122]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][0][1][26] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_28_net_[26] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][0][1][25] ), .Z(o[121]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][0][1][25] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_28_net_[25] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][0][1][24] ), .Z(o[120]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][0][1][24] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_28_net_[24] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][0][1][23] ), .Z(o[119]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][0][1][23] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_28_net_[23] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][0][1][22] ), .Z(o[118]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][0][1][22] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_28_net_[22] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][0][1][21] ), .Z(o[117]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][0][1][21] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_28_net_[21] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][0][1][20] ), .Z(o[116]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][0][1][20] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_28_net_[20] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][0][1][19] ), .Z(o[115]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][0][1][19] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_28_net_[19] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][0][1][18] ), .Z(o[114]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][0][1][18] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_28_net_[18] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][0][1][17] ), .Z(o[113]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][0][1][17] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_28_net_[17] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][0][1][16] ), .Z(o[112]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][0][1][16] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_28_net_[16] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][0][1][15] ), .Z(o[111]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][0][1][15] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_28_net_[15] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][0][1][14] ), .Z(o[110]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][0][1][14] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_28_net_[14] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][0][1][13] ), .Z(o[109]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][0][1][13] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_28_net_[13] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][0][1][12] ), .Z(o[108]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][0][1][12] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_28_net_[12] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][0][1][11] ), .Z(o[107]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][0][1][11] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_28_net_[11] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][0][1][10] ), .Z(o[106]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][0][1][10] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_28_net_[10] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][0][1][9] ), .Z(o[105]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][0][1][9] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_28_net_[9] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][0][1][8] ), .Z(o[104]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][0][1][8] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_28_net_[8] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][0][1][7] ), .Z(o[103]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][0][1][7] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_28_net_[7] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][0][1][6] ), .Z(o[102]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][0][1][6] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_28_net_[6] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][0][1][5] ), .Z(o[101]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][0][1][5] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_28_net_[5] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][0][1][4] ), .Z(o[100]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][0][1][4] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_28_net_[4] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][0][1][3] ), .Z(o[99]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][0][1][3] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_28_net_[3] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][0][1][2] ), .Z(o[98]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][0][1][2] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_28_net_[2] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][0][1][1] ), .Z(o[97]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][0][1][1] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_28_net_[1] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[96]) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[1][0][0][31] ), .Z(\oijt[1][0][1][31] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_24_net_[31] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[1][0][0][30] ), .Z(\oijt[1][0][1][30] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[1][0][0][30] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_24_net_[30] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[1][0][0][29] ), .Z(\oijt[1][0][1][29] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[1][0][0][29] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_24_net_[29] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[1][0][0][28] ), .Z(\oijt[1][0][1][28] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[1][0][0][28] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_24_net_[28] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[1][0][0][27] ), .Z(\oijt[1][0][1][27] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[1][0][0][27] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_24_net_[27] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[1][0][0][26] ), .Z(\oijt[1][0][1][26] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[1][0][0][26] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_24_net_[26] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[1][0][0][25] ), .Z(\oijt[1][0][1][25] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[1][0][0][25] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_24_net_[25] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[1][0][0][24] ), .Z(\oijt[1][0][1][24] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[1][0][0][24] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_24_net_[24] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[1][0][0][23] ), .Z(\oijt[1][0][1][23] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[1][0][0][23] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_24_net_[23] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[1][0][0][22] ), .Z(\oijt[1][0][1][22] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[1][0][0][22] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_24_net_[22] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[1][0][0][21] ), .Z(\oijt[1][0][1][21] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[1][0][0][21] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_24_net_[21] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[1][0][0][20] ), .Z(\oijt[1][0][1][20] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[1][0][0][20] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_24_net_[20] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[1][0][0][19] ), .Z(\oijt[1][0][1][19] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[1][0][0][19] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_24_net_[19] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[1][0][0][18] ), .Z(\oijt[1][0][1][18] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[1][0][0][18] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_24_net_[18] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[1][0][0][17] ), .Z(\oijt[1][0][1][17] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[1][0][0][17] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_24_net_[17] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[1][0][0][16] ), .Z(\oijt[1][0][1][16] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[1][0][0][16] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_24_net_[16] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[1][0][0][15] ), .Z(\oijt[1][0][1][15] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[1][0][0][15] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_24_net_[15] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[1][0][0][14] ), .Z(\oijt[1][0][1][14] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[1][0][0][14] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_24_net_[14] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[1][0][0][13] ), .Z(\oijt[1][0][1][13] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[1][0][0][13] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_24_net_[13] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[1][0][0][12] ), .Z(\oijt[1][0][1][12] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[1][0][0][12] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_24_net_[12] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[1][0][0][11] ), .Z(\oijt[1][0][1][11] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[1][0][0][11] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_24_net_[11] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[1][0][0][10] ), .Z(\oijt[1][0][1][10] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[1][0][0][10] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_24_net_[10] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[1][0][0][9] ), .Z(\oijt[1][0][1][9] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[1][0][0][9] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_24_net_[9] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[1][0][0][8] ), .Z(\oijt[1][0][1][8] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[1][0][0][8] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_24_net_[8] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[1][0][0][7] ), .Z(\oijt[1][0][1][7] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[1][0][0][7] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_24_net_[7] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[1][0][0][6] ), .Z(\oijt[1][0][1][6] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[1][0][0][6] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_24_net_[6] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[1][0][0][5] ), .Z(\oijt[1][0][1][5] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[1][0][0][5] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_24_net_[5] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[1][0][0][4] ), .Z(\oijt[1][0][1][4] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[1][0][0][4] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_24_net_[4] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[1][0][0][3] ), .Z(\oijt[1][0][1][3] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[1][0][0][3] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_24_net_[3] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[1][0][0][2] ), .Z(\oijt[1][0][1][2] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[1][0][0][2] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_24_net_[2] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[1][0][0][1] ), .Z(\oijt[1][0][1][1] ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[1][0][0][1] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_24_net_[1] ), .B(\MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][2][1][31] ), .Z(o[95]) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_20_net_[31] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][2][1][30] ), .Z(o[94]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][2][1][30] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_20_net_[30] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][2][1][29] ), .Z(o[93]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][2][1][29] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_20_net_[29] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][2][1][28] ), .Z(o[92]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][2][1][28] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_20_net_[28] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][2][1][27] ), .Z(o[91]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][2][1][27] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_20_net_[27] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][2][1][26] ), .Z(o[90]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][2][1][26] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_20_net_[26] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][2][1][25] ), .Z(o[89]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][2][1][25] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_20_net_[25] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][2][1][24] ), .Z(o[88]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][2][1][24] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_20_net_[24] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][2][1][23] ), .Z(o[87]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][2][1][23] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_20_net_[23] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][2][1][22] ), .Z(o[86]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][2][1][22] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_20_net_[22] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][2][1][21] ), .Z(o[85]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][2][1][21] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_20_net_[21] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][2][1][20] ), .Z(o[84]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][2][1][20] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_20_net_[20] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][2][1][19] ), .Z(o[83]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][2][1][19] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_20_net_[19] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][2][1][18] ), .Z(o[82]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][2][1][18] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_20_net_[18] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][2][1][17] ), .Z(o[81]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][2][1][17] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_20_net_[17] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][2][1][16] ), .Z(o[80]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][2][1][16] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_20_net_[16] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][2][1][15] ), .Z(o[79]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][2][1][15] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_20_net_[15] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][2][1][14] ), .Z(o[78]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][2][1][14] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_20_net_[14] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][2][1][13] ), .Z(o[77]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][2][1][13] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_20_net_[13] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][2][1][12] ), .Z(o[76]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][2][1][12] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_20_net_[12] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][2][1][11] ), .Z(o[75]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][2][1][11] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_20_net_[11] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][2][1][10] ), .Z(o[74]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][2][1][10] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_20_net_[10] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][2][1][9] ), .Z(o[73]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][2][1][9] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_20_net_[9] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][2][1][8] ), .Z(o[72]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][2][1][8] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_20_net_[8] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][2][1][7] ), .Z(o[71]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][2][1][7] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_20_net_[7] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][2][1][6] ), .Z(o[70]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][2][1][6] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_20_net_[6] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][2][1][5] ), .Z(o[69]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][2][1][5] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_20_net_[5] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][2][1][4] ), .Z(o[68]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][2][1][4] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_20_net_[4] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][2][1][3] ), .Z(o[67]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][2][1][3] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_20_net_[3] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][2][1][2] ), .Z(o[66]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][2][1][2] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_20_net_[2] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][2][1][1] ), .Z(o[65]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][2][1][1] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_20_net_[1] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[64]) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][2][0][31] ), .Z(\oijt[0][2][1][31] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_16_net_[31] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][2][0][30] ), .Z(\oijt[0][2][1][30] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][2][0][30] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_16_net_[30] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][2][0][29] ), .Z(\oijt[0][2][1][29] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][2][0][29] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_16_net_[29] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][2][0][28] ), .Z(\oijt[0][2][1][28] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][2][0][28] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_16_net_[28] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][2][0][27] ), .Z(\oijt[0][2][1][27] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][2][0][27] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_16_net_[27] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][2][0][26] ), .Z(\oijt[0][2][1][26] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][2][0][26] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_16_net_[26] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][2][0][25] ), .Z(\oijt[0][2][1][25] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][2][0][25] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_16_net_[25] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][2][0][24] ), .Z(\oijt[0][2][1][24] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][2][0][24] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_16_net_[24] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][2][0][23] ), .Z(\oijt[0][2][1][23] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][2][0][23] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_16_net_[23] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][2][0][22] ), .Z(\oijt[0][2][1][22] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][2][0][22] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_16_net_[22] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][2][0][21] ), .Z(\oijt[0][2][1][21] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][2][0][21] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_16_net_[21] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][2][0][20] ), .Z(\oijt[0][2][1][20] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][2][0][20] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_16_net_[20] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][2][0][19] ), .Z(\oijt[0][2][1][19] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][2][0][19] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_16_net_[19] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][2][0][18] ), .Z(\oijt[0][2][1][18] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][2][0][18] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_16_net_[18] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][2][0][17] ), .Z(\oijt[0][2][1][17] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][2][0][17] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_16_net_[17] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][2][0][16] ), .Z(\oijt[0][2][1][16] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][2][0][16] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_16_net_[16] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][2][0][15] ), .Z(\oijt[0][2][1][15] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][2][0][15] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_16_net_[15] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][2][0][14] ), .Z(\oijt[0][2][1][14] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][2][0][14] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_16_net_[14] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][2][0][13] ), .Z(\oijt[0][2][1][13] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][2][0][13] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_16_net_[13] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][2][0][12] ), .Z(\oijt[0][2][1][12] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][2][0][12] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_16_net_[12] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][2][0][11] ), .Z(\oijt[0][2][1][11] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][2][0][11] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_16_net_[11] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][2][0][10] ), .Z(\oijt[0][2][1][10] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][2][0][10] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_16_net_[10] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][2][0][9] ), .Z(\oijt[0][2][1][9] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][2][0][9] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(
        \_16_net_[9] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][2][0][8] ), .Z(\oijt[0][2][1][8] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][2][0][8] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(
        \_16_net_[8] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][2][0][7] ), .Z(\oijt[0][2][1][7] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][2][0][7] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(
        \_16_net_[7] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][2][0][6] ), .Z(\oijt[0][2][1][6] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][2][0][6] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(
        \_16_net_[6] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][2][0][5] ), .Z(\oijt[0][2][1][5] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][2][0][5] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(
        \_16_net_[5] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][2][0][4] ), .Z(\oijt[0][2][1][4] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][2][0][4] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(
        \_16_net_[4] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][2][0][3] ), .Z(\oijt[0][2][1][3] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][2][0][3] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(
        \_16_net_[3] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][2][0][2] ), .Z(\oijt[0][2][1][2] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][2][0][2] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(
        \_16_net_[2] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][2][0][1] ), .Z(\oijt[0][2][1][1] ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][2][0][1] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(
        \_16_net_[1] ), .B(\MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][1][1][31] ), .Z(o[63]) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_12_net_[31] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][1][1][30] ), .Z(o[62]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][1][1][30] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_12_net_[30] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][1][1][29] ), .Z(o[61]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][1][1][29] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_12_net_[29] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][1][1][28] ), .Z(o[60]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][1][1][28] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_12_net_[28] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][1][1][27] ), .Z(o[59]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][1][1][27] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_12_net_[27] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][1][1][26] ), .Z(o[58]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][1][1][26] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_12_net_[26] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][1][1][25] ), .Z(o[57]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][1][1][25] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_12_net_[25] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][1][1][24] ), .Z(o[56]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][1][1][24] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_12_net_[24] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][1][1][23] ), .Z(o[55]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][1][1][23] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_12_net_[23] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][1][1][22] ), .Z(o[54]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][1][1][22] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_12_net_[22] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][1][1][21] ), .Z(o[53]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][1][1][21] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_12_net_[21] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][1][1][20] ), .Z(o[52]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][1][1][20] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_12_net_[20] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][1][1][19] ), .Z(o[51]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][1][1][19] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_12_net_[19] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][1][1][18] ), .Z(o[50]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][1][1][18] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_12_net_[18] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][1][1][17] ), .Z(o[49]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][1][1][17] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_12_net_[17] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][1][1][16] ), .Z(o[48]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][1][1][16] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_12_net_[16] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][1][1][15] ), .Z(o[47]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][1][1][15] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_12_net_[15] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][1][1][14] ), .Z(o[46]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][1][1][14] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_12_net_[14] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][1][1][13] ), .Z(o[45]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][1][1][13] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_12_net_[13] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][1][1][12] ), .Z(o[44]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][1][1][12] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_12_net_[12] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][1][1][11] ), .Z(o[43]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][1][1][11] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_12_net_[11] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][1][1][10] ), .Z(o[42]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][1][1][10] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_12_net_[10] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][1][1][9] ), .Z(o[41]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][1][1][9] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(
        \_12_net_[9] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][1][1][8] ), .Z(o[40]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][1][1][8] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(
        \_12_net_[8] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][1][1][7] ), .Z(o[39]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][1][1][7] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(
        \_12_net_[7] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][1][1][6] ), .Z(o[38]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][1][1][6] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(
        \_12_net_[6] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][1][1][5] ), .Z(o[37]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][1][1][5] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(
        \_12_net_[5] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][1][1][4] ), .Z(o[36]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][1][1][4] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(
        \_12_net_[4] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][1][1][3] ), .Z(o[35]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][1][1][3] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(
        \_12_net_[3] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][1][1][2] ), .Z(o[34]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][1][1][2] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(
        \_12_net_[2] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][1][1][1] ), .Z(o[33]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][1][1][1] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(
        \_12_net_[1] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[32]) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][1][0][31] ), .Z(\oijt[0][1][1][31] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_8_net_[31] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][1][0][30] ), .Z(\oijt[0][1][1][30] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][1][0][30] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_8_net_[30] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][1][0][29] ), .Z(\oijt[0][1][1][29] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][1][0][29] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_8_net_[29] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][1][0][28] ), .Z(\oijt[0][1][1][28] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][1][0][28] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_8_net_[28] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][1][0][27] ), .Z(\oijt[0][1][1][27] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][1][0][27] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_8_net_[27] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][1][0][26] ), .Z(\oijt[0][1][1][26] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][1][0][26] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_8_net_[26] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][1][0][25] ), .Z(\oijt[0][1][1][25] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][1][0][25] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_8_net_[25] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][1][0][24] ), .Z(\oijt[0][1][1][24] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][1][0][24] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_8_net_[24] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][1][0][23] ), .Z(\oijt[0][1][1][23] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][1][0][23] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_8_net_[23] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][1][0][22] ), .Z(\oijt[0][1][1][22] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][1][0][22] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_8_net_[22] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][1][0][21] ), .Z(\oijt[0][1][1][21] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][1][0][21] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_8_net_[21] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][1][0][20] ), .Z(\oijt[0][1][1][20] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][1][0][20] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_8_net_[20] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][1][0][19] ), .Z(\oijt[0][1][1][19] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][1][0][19] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_8_net_[19] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][1][0][18] ), .Z(\oijt[0][1][1][18] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][1][0][18] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_8_net_[18] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][1][0][17] ), .Z(\oijt[0][1][1][17] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][1][0][17] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_8_net_[17] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][1][0][16] ), .Z(\oijt[0][1][1][16] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][1][0][16] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_8_net_[16] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][1][0][15] ), .Z(\oijt[0][1][1][15] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][1][0][15] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_8_net_[15] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][1][0][14] ), .Z(\oijt[0][1][1][14] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][1][0][14] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_8_net_[14] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][1][0][13] ), .Z(\oijt[0][1][1][13] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][1][0][13] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_8_net_[13] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][1][0][12] ), .Z(\oijt[0][1][1][12] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][1][0][12] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_8_net_[12] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][1][0][11] ), .Z(\oijt[0][1][1][11] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][1][0][11] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_8_net_[11] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][1][0][10] ), .Z(\oijt[0][1][1][10] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][1][0][10] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_8_net_[10] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][1][0][9] ), .Z(\oijt[0][1][1][9] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][1][0][9] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(\_8_net_[9] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][1][0][8] ), .Z(\oijt[0][1][1][8] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][1][0][8] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(\_8_net_[8] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][1][0][7] ), .Z(\oijt[0][1][1][7] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][1][0][7] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(\_8_net_[7] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][1][0][6] ), .Z(\oijt[0][1][1][6] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][1][0][6] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(\_8_net_[6] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][1][0][5] ), .Z(\oijt[0][1][1][5] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][1][0][5] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(\_8_net_[5] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][1][0][4] ), .Z(\oijt[0][1][1][4] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][1][0][4] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(\_8_net_[4] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][1][0][3] ), .Z(\oijt[0][1][1][3] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][1][0][3] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(\_8_net_[3] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][1][0][2] ), .Z(\oijt[0][1][1][2] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][1][0][2] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(\_8_net_[2] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][1][0][1] ), .Z(\oijt[0][1][1][1] ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][1][0][1] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(\_8_net_[1] ), .B(\MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n2 ) );
  AND \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][0][1][31] ), .Z(o[31]) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/U1  ( .A(
        \_4_net_[31] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][0][1][30] ), .Z(o[30]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][0][1][30] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/U1  ( .A(
        \_4_net_[30] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][0][1][29] ), .Z(o[29]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][0][1][29] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/U1  ( .A(
        \_4_net_[29] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][0][1][28] ), .Z(o[28]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][0][1][28] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/U1  ( .A(
        \_4_net_[28] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][0][1][27] ), .Z(o[27]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][0][1][27] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/U1  ( .A(
        \_4_net_[27] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][0][1][26] ), .Z(o[26]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][0][1][26] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/U1  ( .A(
        \_4_net_[26] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][0][1][25] ), .Z(o[25]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][0][1][25] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/U1  ( .A(
        \_4_net_[25] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][0][1][24] ), .Z(o[24]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][0][1][24] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/U1  ( .A(
        \_4_net_[24] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][0][1][23] ), .Z(o[23]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][0][1][23] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/U1  ( .A(
        \_4_net_[23] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][0][1][22] ), .Z(o[22]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][0][1][22] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/U1  ( .A(
        \_4_net_[22] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][0][1][21] ), .Z(o[21]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][0][1][21] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/U1  ( .A(
        \_4_net_[21] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][0][1][20] ), .Z(o[20]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][0][1][20] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/U1  ( .A(
        \_4_net_[20] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][0][1][19] ), .Z(o[19]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][0][1][19] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/U1  ( .A(
        \_4_net_[19] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][0][1][18] ), .Z(o[18]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][0][1][18] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/U1  ( .A(
        \_4_net_[18] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][0][1][17] ), .Z(o[17]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][0][1][17] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/U1  ( .A(
        \_4_net_[17] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][0][1][16] ), .Z(o[16]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][0][1][16] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/U1  ( .A(
        \_4_net_[16] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][0][1][15] ), .Z(o[15]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][0][1][15] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/U1  ( .A(
        \_4_net_[15] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][0][1][14] ), .Z(o[14]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][0][1][14] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/U1  ( .A(
        \_4_net_[14] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][0][1][13] ), .Z(o[13]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][0][1][13] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/U1  ( .A(
        \_4_net_[13] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][0][1][12] ), .Z(o[12]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][0][1][12] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/U1  ( .A(
        \_4_net_[12] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][0][1][11] ), .Z(o[11]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][0][1][11] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/U1  ( .A(
        \_4_net_[11] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][0][1][10] ), .Z(o[10]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][0][1][10] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/U1  ( .A(
        \_4_net_[10] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][0][1][9] ), .Z(o[9]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][0][1][9] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/U1  ( .A(\_4_net_[9] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][0][1][8] ), .Z(o[8]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][0][1][8] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/U1  ( .A(\_4_net_[8] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][0][1][7] ), .Z(o[7]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][0][1][7] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/U1  ( .A(\_4_net_[7] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][0][1][6] ), .Z(o[6]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][0][1][6] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/U1  ( .A(\_4_net_[6] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][0][1][5] ), .Z(o[5]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][0][1][5] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/U1  ( .A(\_4_net_[5] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][0][1][4] ), .Z(o[4]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][0][1][4] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/U1  ( .A(\_4_net_[4] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][0][1][3] ), .Z(o[3]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][0][1][3] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/U1  ( .A(\_4_net_[3] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][0][1][2] ), .Z(o[2]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][0][1][2] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/U1  ( .A(\_4_net_[2] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][0][1][1] ), .Z(o[1]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][0][1][1] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/U1  ( .A(\_4_net_[1] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[1].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(o[0]) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/c[1] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ), .B(
        \oijt[0][0][0][31] ), .Z(\oijt[0][0][1][31] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/U1  ( .A(
        \_0_net_[31] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[31] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[31].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[31] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \oijt[0][0][0][30] ), .Z(\oijt[0][0][1][30] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U2  ( .A(
        \oijt[0][0][0][30] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[30] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/U1  ( .A(
        \_0_net_[30] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[30] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[30].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[30] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \oijt[0][0][0][29] ), .Z(\oijt[0][0][1][29] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U2  ( .A(
        \oijt[0][0][0][29] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[29] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/U1  ( .A(
        \_0_net_[29] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[29] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[29].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[29] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \oijt[0][0][0][28] ), .Z(\oijt[0][0][1][28] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U2  ( .A(
        \oijt[0][0][0][28] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[28] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/U1  ( .A(
        \_0_net_[28] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[28] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[28].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[28] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \oijt[0][0][0][27] ), .Z(\oijt[0][0][1][27] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U2  ( .A(
        \oijt[0][0][0][27] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[27] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/U1  ( .A(
        \_0_net_[27] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[27] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[27].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[27] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \oijt[0][0][0][26] ), .Z(\oijt[0][0][1][26] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U2  ( .A(
        \oijt[0][0][0][26] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[26] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/U1  ( .A(
        \_0_net_[26] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[26] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[26].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[26] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \oijt[0][0][0][25] ), .Z(\oijt[0][0][1][25] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U2  ( .A(
        \oijt[0][0][0][25] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[25] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/U1  ( .A(
        \_0_net_[25] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[25] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[25].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[25] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \oijt[0][0][0][24] ), .Z(\oijt[0][0][1][24] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U2  ( .A(
        \oijt[0][0][0][24] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[24] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/U1  ( .A(
        \_0_net_[24] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[24] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[24].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[24] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \oijt[0][0][0][23] ), .Z(\oijt[0][0][1][23] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U2  ( .A(
        \oijt[0][0][0][23] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[23] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/U1  ( .A(
        \_0_net_[23] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[23] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[23].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[23] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \oijt[0][0][0][22] ), .Z(\oijt[0][0][1][22] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U2  ( .A(
        \oijt[0][0][0][22] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[22] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/U1  ( .A(
        \_0_net_[22] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[22] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[22].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[22] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \oijt[0][0][0][21] ), .Z(\oijt[0][0][1][21] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U2  ( .A(
        \oijt[0][0][0][21] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[21] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/U1  ( .A(
        \_0_net_[21] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[21] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[21].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[21] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \oijt[0][0][0][20] ), .Z(\oijt[0][0][1][20] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U2  ( .A(
        \oijt[0][0][0][20] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[20] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/U1  ( .A(
        \_0_net_[20] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[20] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[20].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[20] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \oijt[0][0][0][19] ), .Z(\oijt[0][0][1][19] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U2  ( .A(
        \oijt[0][0][0][19] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[19] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/U1  ( .A(
        \_0_net_[19] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[19] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[19].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[19] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \oijt[0][0][0][18] ), .Z(\oijt[0][0][1][18] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U2  ( .A(
        \oijt[0][0][0][18] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[18] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/U1  ( .A(
        \_0_net_[18] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[18] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[18].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[18] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \oijt[0][0][0][17] ), .Z(\oijt[0][0][1][17] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U2  ( .A(
        \oijt[0][0][0][17] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[17] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/U1  ( .A(
        \_0_net_[17] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[17] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[17].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[17] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \oijt[0][0][0][16] ), .Z(\oijt[0][0][1][16] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U2  ( .A(
        \oijt[0][0][0][16] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[16] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/U1  ( .A(
        \_0_net_[16] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[16] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[16].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[16] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \oijt[0][0][0][15] ), .Z(\oijt[0][0][1][15] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U2  ( .A(
        \oijt[0][0][0][15] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[15] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/U1  ( .A(
        \_0_net_[15] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[15] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[15].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[15] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \oijt[0][0][0][14] ), .Z(\oijt[0][0][1][14] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U2  ( .A(
        \oijt[0][0][0][14] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[14] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/U1  ( .A(
        \_0_net_[14] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[14] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[14].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[14] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \oijt[0][0][0][13] ), .Z(\oijt[0][0][1][13] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U2  ( .A(
        \oijt[0][0][0][13] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[13] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/U1  ( .A(
        \_0_net_[13] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[13] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[13].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[13] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \oijt[0][0][0][12] ), .Z(\oijt[0][0][1][12] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U2  ( .A(
        \oijt[0][0][0][12] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[12] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/U1  ( .A(
        \_0_net_[12] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[12] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[12].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[12] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \oijt[0][0][0][11] ), .Z(\oijt[0][0][1][11] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U2  ( .A(
        \oijt[0][0][0][11] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[11] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/U1  ( .A(
        \_0_net_[11] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[11] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[11].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[11] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \oijt[0][0][0][10] ), .Z(\oijt[0][0][1][10] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U2  ( .A(
        \oijt[0][0][0][10] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[10] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/U1  ( .A(
        \_0_net_[10] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[10] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[10].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[10] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \oijt[0][0][0][9] ), .Z(\oijt[0][0][1][9] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U2  ( .A(
        \oijt[0][0][0][9] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[9] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/U1  ( .A(\_0_net_[9] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[9] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[9].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[9] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \oijt[0][0][0][8] ), .Z(\oijt[0][0][1][8] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U2  ( .A(
        \oijt[0][0][0][8] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[8] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/U1  ( .A(\_0_net_[8] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[8] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[8].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[8] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \oijt[0][0][0][7] ), .Z(\oijt[0][0][1][7] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U2  ( .A(
        \oijt[0][0][0][7] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[7] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/U1  ( .A(\_0_net_[7] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[7] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[7].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[7] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \oijt[0][0][0][6] ), .Z(\oijt[0][0][1][6] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U2  ( .A(
        \oijt[0][0][0][6] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[6] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/U1  ( .A(\_0_net_[6] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[6] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[6].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[6] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \oijt[0][0][0][5] ), .Z(\oijt[0][0][1][5] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U2  ( .A(
        \oijt[0][0][0][5] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[5] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/U1  ( .A(\_0_net_[5] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[5] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[5].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[5] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \oijt[0][0][0][4] ), .Z(\oijt[0][0][1][4] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U2  ( .A(
        \oijt[0][0][0][4] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[4] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/U1  ( .A(\_0_net_[4] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[4] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[4].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[4] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \oijt[0][0][0][3] ), .Z(\oijt[0][0][1][3] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U2  ( .A(
        \oijt[0][0][0][3] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[3] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/U1  ( .A(\_0_net_[3] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[3] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[3].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[3] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \oijt[0][0][0][2] ), .Z(\oijt[0][0][1][2] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U2  ( .A(
        \oijt[0][0][0][2] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[2] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/U1  ( .A(\_0_net_[2] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[2] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[2].FA_/n1 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U5  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[2] ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U4  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \oijt[0][0][0][1] ), .Z(\oijt[0][0][1][1] ) );
  AND \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U3  ( .A(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ), .B(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n3 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U2  ( .A(
        \oijt[0][0][0][1] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[1] ), 
        .Z(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n2 ) );
  XOR \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/U1  ( .A(\_0_net_[1] ), .B(\MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/c[1] ), .Z(
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[1].FA_/n1 ) );
  MULT_UNS_OP mult_37 ( .A(x[31:0]), .B(y[31:0]), .Z({\oijt[0][0][0][31] , 
        \oijt[0][0][0][30] , \oijt[0][0][0][29] , \oijt[0][0][0][28] , 
        \oijt[0][0][0][27] , \oijt[0][0][0][26] , \oijt[0][0][0][25] , 
        \oijt[0][0][0][24] , \oijt[0][0][0][23] , \oijt[0][0][0][22] , 
        \oijt[0][0][0][21] , \oijt[0][0][0][20] , \oijt[0][0][0][19] , 
        \oijt[0][0][0][18] , \oijt[0][0][0][17] , \oijt[0][0][0][16] , 
        \oijt[0][0][0][15] , \oijt[0][0][0][14] , \oijt[0][0][0][13] , 
        \oijt[0][0][0][12] , \oijt[0][0][0][11] , \oijt[0][0][0][10] , 
        \oijt[0][0][0][9] , \oijt[0][0][0][8] , \oijt[0][0][0][7] , 
        \oijt[0][0][0][6] , \oijt[0][0][0][5] , \oijt[0][0][0][4] , 
        \oijt[0][0][0][3] , \oijt[0][0][0][2] , \oijt[0][0][0][1] , 
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G2_G1 ( .A(x[31:0]), .B(y[63:32]), .Z({
        \oijt[0][1][0][31] , \oijt[0][1][0][30] , \oijt[0][1][0][29] , 
        \oijt[0][1][0][28] , \oijt[0][1][0][27] , \oijt[0][1][0][26] , 
        \oijt[0][1][0][25] , \oijt[0][1][0][24] , \oijt[0][1][0][23] , 
        \oijt[0][1][0][22] , \oijt[0][1][0][21] , \oijt[0][1][0][20] , 
        \oijt[0][1][0][19] , \oijt[0][1][0][18] , \oijt[0][1][0][17] , 
        \oijt[0][1][0][16] , \oijt[0][1][0][15] , \oijt[0][1][0][14] , 
        \oijt[0][1][0][13] , \oijt[0][1][0][12] , \oijt[0][1][0][11] , 
        \oijt[0][1][0][10] , \oijt[0][1][0][9] , \oijt[0][1][0][8] , 
        \oijt[0][1][0][7] , \oijt[0][1][0][6] , \oijt[0][1][0][5] , 
        \oijt[0][1][0][4] , \oijt[0][1][0][3] , \oijt[0][1][0][2] , 
        \oijt[0][1][0][1] , 
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G3_G1 ( .A(x[31:0]), .B(y[95:64]), .Z({
        \oijt[0][2][0][31] , \oijt[0][2][0][30] , \oijt[0][2][0][29] , 
        \oijt[0][2][0][28] , \oijt[0][2][0][27] , \oijt[0][2][0][26] , 
        \oijt[0][2][0][25] , \oijt[0][2][0][24] , \oijt[0][2][0][23] , 
        \oijt[0][2][0][22] , \oijt[0][2][0][21] , \oijt[0][2][0][20] , 
        \oijt[0][2][0][19] , \oijt[0][2][0][18] , \oijt[0][2][0][17] , 
        \oijt[0][2][0][16] , \oijt[0][2][0][15] , \oijt[0][2][0][14] , 
        \oijt[0][2][0][13] , \oijt[0][2][0][12] , \oijt[0][2][0][11] , 
        \oijt[0][2][0][10] , \oijt[0][2][0][9] , \oijt[0][2][0][8] , 
        \oijt[0][2][0][7] , \oijt[0][2][0][6] , \oijt[0][2][0][5] , 
        \oijt[0][2][0][4] , \oijt[0][2][0][3] , \oijt[0][2][0][2] , 
        \oijt[0][2][0][1] , 
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G2 ( .A(x[127:96]), .B(y[31:0]), .Z({\oijt[1][0][0][31] , 
        \oijt[1][0][0][30] , \oijt[1][0][0][29] , \oijt[1][0][0][28] , 
        \oijt[1][0][0][27] , \oijt[1][0][0][26] , \oijt[1][0][0][25] , 
        \oijt[1][0][0][24] , \oijt[1][0][0][23] , \oijt[1][0][0][22] , 
        \oijt[1][0][0][21] , \oijt[1][0][0][20] , \oijt[1][0][0][19] , 
        \oijt[1][0][0][18] , \oijt[1][0][0][17] , \oijt[1][0][0][16] , 
        \oijt[1][0][0][15] , \oijt[1][0][0][14] , \oijt[1][0][0][13] , 
        \oijt[1][0][0][12] , \oijt[1][0][0][11] , \oijt[1][0][0][10] , 
        \oijt[1][0][0][9] , \oijt[1][0][0][8] , \oijt[1][0][0][7] , 
        \oijt[1][0][0][6] , \oijt[1][0][0][5] , \oijt[1][0][0][4] , 
        \oijt[1][0][0][3] , \oijt[1][0][0][2] , \oijt[1][0][0][1] , 
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G2_G2 ( .A(x[127:96]), .B(y[63:32]), .Z({
        \oijt[1][1][0][31] , \oijt[1][1][0][30] , \oijt[1][1][0][29] , 
        \oijt[1][1][0][28] , \oijt[1][1][0][27] , \oijt[1][1][0][26] , 
        \oijt[1][1][0][25] , \oijt[1][1][0][24] , \oijt[1][1][0][23] , 
        \oijt[1][1][0][22] , \oijt[1][1][0][21] , \oijt[1][1][0][20] , 
        \oijt[1][1][0][19] , \oijt[1][1][0][18] , \oijt[1][1][0][17] , 
        \oijt[1][1][0][16] , \oijt[1][1][0][15] , \oijt[1][1][0][14] , 
        \oijt[1][1][0][13] , \oijt[1][1][0][12] , \oijt[1][1][0][11] , 
        \oijt[1][1][0][10] , \oijt[1][1][0][9] , \oijt[1][1][0][8] , 
        \oijt[1][1][0][7] , \oijt[1][1][0][6] , \oijt[1][1][0][5] , 
        \oijt[1][1][0][4] , \oijt[1][1][0][3] , \oijt[1][1][0][2] , 
        \oijt[1][1][0][1] , 
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G3_G2 ( .A(x[127:96]), .B(y[95:64]), .Z({
        \oijt[1][2][0][31] , \oijt[1][2][0][30] , \oijt[1][2][0][29] , 
        \oijt[1][2][0][28] , \oijt[1][2][0][27] , \oijt[1][2][0][26] , 
        \oijt[1][2][0][25] , \oijt[1][2][0][24] , \oijt[1][2][0][23] , 
        \oijt[1][2][0][22] , \oijt[1][2][0][21] , \oijt[1][2][0][20] , 
        \oijt[1][2][0][19] , \oijt[1][2][0][18] , \oijt[1][2][0][17] , 
        \oijt[1][2][0][16] , \oijt[1][2][0][15] , \oijt[1][2][0][14] , 
        \oijt[1][2][0][13] , \oijt[1][2][0][12] , \oijt[1][2][0][11] , 
        \oijt[1][2][0][10] , \oijt[1][2][0][9] , \oijt[1][2][0][8] , 
        \oijt[1][2][0][7] , \oijt[1][2][0][6] , \oijt[1][2][0][5] , 
        \oijt[1][2][0][4] , \oijt[1][2][0][3] , \oijt[1][2][0][2] , 
        \oijt[1][2][0][1] , 
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G3 ( .A(x[223:192]), .B(y[31:0]), .Z({
        \oijt[2][0][0][31] , \oijt[2][0][0][30] , \oijt[2][0][0][29] , 
        \oijt[2][0][0][28] , \oijt[2][0][0][27] , \oijt[2][0][0][26] , 
        \oijt[2][0][0][25] , \oijt[2][0][0][24] , \oijt[2][0][0][23] , 
        \oijt[2][0][0][22] , \oijt[2][0][0][21] , \oijt[2][0][0][20] , 
        \oijt[2][0][0][19] , \oijt[2][0][0][18] , \oijt[2][0][0][17] , 
        \oijt[2][0][0][16] , \oijt[2][0][0][15] , \oijt[2][0][0][14] , 
        \oijt[2][0][0][13] , \oijt[2][0][0][12] , \oijt[2][0][0][11] , 
        \oijt[2][0][0][10] , \oijt[2][0][0][9] , \oijt[2][0][0][8] , 
        \oijt[2][0][0][7] , \oijt[2][0][0][6] , \oijt[2][0][0][5] , 
        \oijt[2][0][0][4] , \oijt[2][0][0][3] , \oijt[2][0][0][2] , 
        \oijt[2][0][0][1] , 
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G2_G3 ( .A(x[223:192]), .B(y[63:32]), .Z({
        \oijt[2][1][0][31] , \oijt[2][1][0][30] , \oijt[2][1][0][29] , 
        \oijt[2][1][0][28] , \oijt[2][1][0][27] , \oijt[2][1][0][26] , 
        \oijt[2][1][0][25] , \oijt[2][1][0][24] , \oijt[2][1][0][23] , 
        \oijt[2][1][0][22] , \oijt[2][1][0][21] , \oijt[2][1][0][20] , 
        \oijt[2][1][0][19] , \oijt[2][1][0][18] , \oijt[2][1][0][17] , 
        \oijt[2][1][0][16] , \oijt[2][1][0][15] , \oijt[2][1][0][14] , 
        \oijt[2][1][0][13] , \oijt[2][1][0][12] , \oijt[2][1][0][11] , 
        \oijt[2][1][0][10] , \oijt[2][1][0][9] , \oijt[2][1][0][8] , 
        \oijt[2][1][0][7] , \oijt[2][1][0][6] , \oijt[2][1][0][5] , 
        \oijt[2][1][0][4] , \oijt[2][1][0][3] , \oijt[2][1][0][2] , 
        \oijt[2][1][0][1] , 
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_37_G3_G3 ( .A(x[223:192]), .B(y[95:64]), .Z({
        \oijt[2][2][0][31] , \oijt[2][2][0][30] , \oijt[2][2][0][29] , 
        \oijt[2][2][0][28] , \oijt[2][2][0][27] , \oijt[2][2][0][26] , 
        \oijt[2][2][0][25] , \oijt[2][2][0][24] , \oijt[2][2][0][23] , 
        \oijt[2][2][0][22] , \oijt[2][2][0][21] , \oijt[2][2][0][20] , 
        \oijt[2][2][0][19] , \oijt[2][2][0][18] , \oijt[2][2][0][17] , 
        \oijt[2][2][0][16] , \oijt[2][2][0][15] , \oijt[2][2][0][14] , 
        \oijt[2][2][0][13] , \oijt[2][2][0][12] , \oijt[2][2][0][11] , 
        \oijt[2][2][0][10] , \oijt[2][2][0][9] , \oijt[2][2][0][8] , 
        \oijt[2][2][0][7] , \oijt[2][2][0][6] , \oijt[2][2][0][5] , 
        \oijt[2][2][0][4] , \oijt[2][2][0][3] , \oijt[2][2][0][2] , 
        \oijt[2][2][0][1] , 
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n2 }) );
  MULT_UNS_OP mult_55 ( .A(x[63:32]), .B(y[127:96]), .Z({\_0_net_[31] , 
        \_0_net_[30] , \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , 
        \_0_net_[26] , \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , 
        \_0_net_[22] , \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , 
        \_0_net_[18] , \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , 
        \_0_net_[14] , \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , 
        \_0_net_[10] , \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , 
        \_0_net_[5] , \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 
        \MUL_ROW[0].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G1_G1 ( .A(x[95:64]), .B(y[223:192]), .Z({
        \_4_net_[31] , \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , 
        \_4_net_[27] , \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , 
        \_4_net_[23] , \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , 
        \_4_net_[19] , \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , 
        \_4_net_[15] , \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , 
        \_4_net_[11] , \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , 
        \_4_net_[6] , \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_4_net_[2] , 
        \_4_net_[1] , \MUL_ROW[0].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 })
         );
  MULT_UNS_OP mult_55_G2_G1 ( .A(x[63:32]), .B(y[159:128]), .Z({\_8_net_[31] , 
        \_8_net_[30] , \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , 
        \_8_net_[26] , \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , 
        \_8_net_[22] , \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , 
        \_8_net_[18] , \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , 
        \_8_net_[14] , \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , 
        \_8_net_[10] , \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , 
        \_8_net_[5] , \_8_net_[4] , \_8_net_[3] , \_8_net_[2] , \_8_net_[1] , 
        \MUL_ROW[0].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G2_G1 ( .A(x[95:64]), .B(y[255:224]), .Z({
        \_12_net_[31] , \_12_net_[30] , \_12_net_[29] , \_12_net_[28] , 
        \_12_net_[27] , \_12_net_[26] , \_12_net_[25] , \_12_net_[24] , 
        \_12_net_[23] , \_12_net_[22] , \_12_net_[21] , \_12_net_[20] , 
        \_12_net_[19] , \_12_net_[18] , \_12_net_[17] , \_12_net_[16] , 
        \_12_net_[15] , \_12_net_[14] , \_12_net_[13] , \_12_net_[12] , 
        \_12_net_[11] , \_12_net_[10] , \_12_net_[9] , \_12_net_[8] , 
        \_12_net_[7] , \_12_net_[6] , \_12_net_[5] , \_12_net_[4] , 
        \_12_net_[3] , \_12_net_[2] , \_12_net_[1] , 
        \MUL_ROW[0].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G3_G1 ( .A(x[63:32]), .B(y[191:160]), .Z({\_16_net_[31] , 
        \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , 
        \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , 
        \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , 
        \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , 
        \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , 
        \_16_net_[10] , \_16_net_[9] , \_16_net_[8] , \_16_net_[7] , 
        \_16_net_[6] , \_16_net_[5] , \_16_net_[4] , \_16_net_[3] , 
        \_16_net_[2] , \_16_net_[1] , 
        \MUL_ROW[0].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G3_G1 ( .A(x[95:64]), .B(y[287:256]), .Z({
        \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] , 
        \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] , 
        \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] , 
        \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] , 
        \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] , 
        \_20_net_[11] , \_20_net_[10] , \_20_net_[9] , \_20_net_[8] , 
        \_20_net_[7] , \_20_net_[6] , \_20_net_[5] , \_20_net_[4] , 
        \_20_net_[3] , \_20_net_[2] , \_20_net_[1] , 
        \MUL_ROW[0].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2 ( .A(x[159:128]), .B(y[127:96]), .Z({\_24_net_[31] , 
        \_24_net_[30] , \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , 
        \_24_net_[26] , \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , 
        \_24_net_[22] , \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , 
        \_24_net_[18] , \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , 
        \_24_net_[14] , \_24_net_[13] , \_24_net_[12] , \_24_net_[11] , 
        \_24_net_[10] , \_24_net_[9] , \_24_net_[8] , \_24_net_[7] , 
        \_24_net_[6] , \_24_net_[5] , \_24_net_[4] , \_24_net_[3] , 
        \_24_net_[2] , \_24_net_[1] , 
        \MUL_ROW[1].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G1_G2 ( .A(x[191:160]), .B(y[223:192]), .Z({
        \_28_net_[31] , \_28_net_[30] , \_28_net_[29] , \_28_net_[28] , 
        \_28_net_[27] , \_28_net_[26] , \_28_net_[25] , \_28_net_[24] , 
        \_28_net_[23] , \_28_net_[22] , \_28_net_[21] , \_28_net_[20] , 
        \_28_net_[19] , \_28_net_[18] , \_28_net_[17] , \_28_net_[16] , 
        \_28_net_[15] , \_28_net_[14] , \_28_net_[13] , \_28_net_[12] , 
        \_28_net_[11] , \_28_net_[10] , \_28_net_[9] , \_28_net_[8] , 
        \_28_net_[7] , \_28_net_[6] , \_28_net_[5] , \_28_net_[4] , 
        \_28_net_[3] , \_28_net_[2] , \_28_net_[1] , 
        \MUL_ROW[1].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G2 ( .A(x[159:128]), .B(y[159:128]), .Z({
        \_32_net_[31] , \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , 
        \_32_net_[27] , \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , 
        \_32_net_[23] , \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , 
        \_32_net_[19] , \_32_net_[18] , \_32_net_[17] , \_32_net_[16] , 
        \_32_net_[15] , \_32_net_[14] , \_32_net_[13] , \_32_net_[12] , 
        \_32_net_[11] , \_32_net_[10] , \_32_net_[9] , \_32_net_[8] , 
        \_32_net_[7] , \_32_net_[6] , \_32_net_[5] , \_32_net_[4] , 
        \_32_net_[3] , \_32_net_[2] , \_32_net_[1] , 
        \MUL_ROW[1].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G2_G2 ( .A(x[191:160]), .B(y[255:224]), .Z({
        \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] , 
        \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] , 
        \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] , 
        \_36_net_[19] , \_36_net_[18] , \_36_net_[17] , \_36_net_[16] , 
        \_36_net_[15] , \_36_net_[14] , \_36_net_[13] , \_36_net_[12] , 
        \_36_net_[11] , \_36_net_[10] , \_36_net_[9] , \_36_net_[8] , 
        \_36_net_[7] , \_36_net_[6] , \_36_net_[5] , \_36_net_[4] , 
        \_36_net_[3] , \_36_net_[2] , \_36_net_[1] , 
        \MUL_ROW[1].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G3_G2 ( .A(x[159:128]), .B(y[191:160]), .Z({
        \_40_net_[31] , \_40_net_[30] , \_40_net_[29] , \_40_net_[28] , 
        \_40_net_[27] , \_40_net_[26] , \_40_net_[25] , \_40_net_[24] , 
        \_40_net_[23] , \_40_net_[22] , \_40_net_[21] , \_40_net_[20] , 
        \_40_net_[19] , \_40_net_[18] , \_40_net_[17] , \_40_net_[16] , 
        \_40_net_[15] , \_40_net_[14] , \_40_net_[13] , \_40_net_[12] , 
        \_40_net_[11] , \_40_net_[10] , \_40_net_[9] , \_40_net_[8] , 
        \_40_net_[7] , \_40_net_[6] , \_40_net_[5] , \_40_net_[4] , 
        \_40_net_[3] , \_40_net_[2] , \_40_net_[1] , 
        \MUL_ROW[1].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G3_G2 ( .A(x[191:160]), .B(y[287:256]), .Z({
        \_44_net_[31] , \_44_net_[30] , \_44_net_[29] , \_44_net_[28] , 
        \_44_net_[27] , \_44_net_[26] , \_44_net_[25] , \_44_net_[24] , 
        \_44_net_[23] , \_44_net_[22] , \_44_net_[21] , \_44_net_[20] , 
        \_44_net_[19] , \_44_net_[18] , \_44_net_[17] , \_44_net_[16] , 
        \_44_net_[15] , \_44_net_[14] , \_44_net_[13] , \_44_net_[12] , 
        \_44_net_[11] , \_44_net_[10] , \_44_net_[9] , \_44_net_[8] , 
        \_44_net_[7] , \_44_net_[6] , \_44_net_[5] , \_44_net_[4] , 
        \_44_net_[3] , \_44_net_[2] , \_44_net_[1] , 
        \MUL_ROW[1].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G3 ( .A(x[255:224]), .B(y[127:96]), .Z({\_48_net_[31] , 
        \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , 
        \_48_net_[26] , \_48_net_[25] , \_48_net_[24] , \_48_net_[23] , 
        \_48_net_[22] , \_48_net_[21] , \_48_net_[20] , \_48_net_[19] , 
        \_48_net_[18] , \_48_net_[17] , \_48_net_[16] , \_48_net_[15] , 
        \_48_net_[14] , \_48_net_[13] , \_48_net_[12] , \_48_net_[11] , 
        \_48_net_[10] , \_48_net_[9] , \_48_net_[8] , \_48_net_[7] , 
        \_48_net_[6] , \_48_net_[5] , \_48_net_[4] , \_48_net_[3] , 
        \_48_net_[2] , \_48_net_[1] , 
        \MUL_ROW[2].MUL_COL[0].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G1_G3 ( .A(x[287:256]), .B(y[223:192]), .Z({
        \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] , 
        \_52_net_[27] , \_52_net_[26] , \_52_net_[25] , \_52_net_[24] , 
        \_52_net_[23] , \_52_net_[22] , \_52_net_[21] , \_52_net_[20] , 
        \_52_net_[19] , \_52_net_[18] , \_52_net_[17] , \_52_net_[16] , 
        \_52_net_[15] , \_52_net_[14] , \_52_net_[13] , \_52_net_[12] , 
        \_52_net_[11] , \_52_net_[10] , \_52_net_[9] , \_52_net_[8] , 
        \_52_net_[7] , \_52_net_[6] , \_52_net_[5] , \_52_net_[4] , 
        \_52_net_[3] , \_52_net_[2] , \_52_net_[1] , 
        \MUL_ROW[2].MUL_COL[0].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G3 ( .A(x[255:224]), .B(y[159:128]), .Z({
        \_56_net_[31] , \_56_net_[30] , \_56_net_[29] , \_56_net_[28] , 
        \_56_net_[27] , \_56_net_[26] , \_56_net_[25] , \_56_net_[24] , 
        \_56_net_[23] , \_56_net_[22] , \_56_net_[21] , \_56_net_[20] , 
        \_56_net_[19] , \_56_net_[18] , \_56_net_[17] , \_56_net_[16] , 
        \_56_net_[15] , \_56_net_[14] , \_56_net_[13] , \_56_net_[12] , 
        \_56_net_[11] , \_56_net_[10] , \_56_net_[9] , \_56_net_[8] , 
        \_56_net_[7] , \_56_net_[6] , \_56_net_[5] , \_56_net_[4] , 
        \_56_net_[3] , \_56_net_[2] , \_56_net_[1] , 
        \MUL_ROW[2].MUL_COL[1].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G2_G3 ( .A(x[287:256]), .B(y[255:224]), .Z({
        \_60_net_[31] , \_60_net_[30] , \_60_net_[29] , \_60_net_[28] , 
        \_60_net_[27] , \_60_net_[26] , \_60_net_[25] , \_60_net_[24] , 
        \_60_net_[23] , \_60_net_[22] , \_60_net_[21] , \_60_net_[20] , 
        \_60_net_[19] , \_60_net_[18] , \_60_net_[17] , \_60_net_[16] , 
        \_60_net_[15] , \_60_net_[14] , \_60_net_[13] , \_60_net_[12] , 
        \_60_net_[11] , \_60_net_[10] , \_60_net_[9] , \_60_net_[8] , 
        \_60_net_[7] , \_60_net_[6] , \_60_net_[5] , \_60_net_[4] , 
        \_60_net_[3] , \_60_net_[2] , \_60_net_[1] , 
        \MUL_ROW[2].MUL_COL[1].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G3_G3 ( .A(x[255:224]), .B(y[191:160]), .Z({
        \_64_net_[31] , \_64_net_[30] , \_64_net_[29] , \_64_net_[28] , 
        \_64_net_[27] , \_64_net_[26] , \_64_net_[25] , \_64_net_[24] , 
        \_64_net_[23] , \_64_net_[22] , \_64_net_[21] , \_64_net_[20] , 
        \_64_net_[19] , \_64_net_[18] , \_64_net_[17] , \_64_net_[16] , 
        \_64_net_[15] , \_64_net_[14] , \_64_net_[13] , \_64_net_[12] , 
        \_64_net_[11] , \_64_net_[10] , \_64_net_[9] , \_64_net_[8] , 
        \_64_net_[7] , \_64_net_[6] , \_64_net_[5] , \_64_net_[4] , 
        \_64_net_[3] , \_64_net_[2] , \_64_net_[1] , 
        \MUL_ROW[2].MUL_COL[2].ADD_O[1].ADD_/FAINST[0].FA_/n1 }) );
  MULT_UNS_OP mult_55_G2_G3_G3 ( .A(x[287:256]), .B(y[287:256]), .Z({
        \_68_net_[31] , \_68_net_[30] , \_68_net_[29] , \_68_net_[28] , 
        \_68_net_[27] , \_68_net_[26] , \_68_net_[25] , \_68_net_[24] , 
        \_68_net_[23] , \_68_net_[22] , \_68_net_[21] , \_68_net_[20] , 
        \_68_net_[19] , \_68_net_[18] , \_68_net_[17] , \_68_net_[16] , 
        \_68_net_[15] , \_68_net_[14] , \_68_net_[13] , \_68_net_[12] , 
        \_68_net_[11] , \_68_net_[10] , \_68_net_[9] , \_68_net_[8] , 
        \_68_net_[7] , \_68_net_[6] , \_68_net_[5] , \_68_net_[4] , 
        \_68_net_[3] , \_68_net_[2] , \_68_net_[1] , 
        \MUL_ROW[2].MUL_COL[2].ADD_O[2].ADD_/FAINST[0].FA_/n1 }) );
endmodule

