
module compare_N16384_CC32 ( clk, rst, x, y, g, e );
  input [511:0] x;
  input [511:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  AND U10 ( .A(n2086), .B(n2087), .Z(n8) );
  NANDN U11 ( .A(n2085), .B(n2084), .Z(n9) );
  AND U12 ( .A(n8), .B(n9), .Z(n10) );
  OR U13 ( .A(n2088), .B(n10), .Z(n11) );
  NANDN U14 ( .A(n2089), .B(n11), .Z(n12) );
  ANDN U15 ( .B(n12), .A(n2090), .Z(n13) );
  ANDN U16 ( .B(n2091), .A(n13), .Z(n14) );
  NAND U17 ( .A(n14), .B(n2092), .Z(n15) );
  ANDN U18 ( .B(n15), .A(n2093), .Z(n16) );
  OR U19 ( .A(n2094), .B(n16), .Z(n17) );
  NANDN U20 ( .A(n2095), .B(n17), .Z(n18) );
  ANDN U21 ( .B(n18), .A(n2096), .Z(n19) );
  NOR U22 ( .A(n19), .B(n2098), .Z(n20) );
  NANDN U23 ( .A(n2097), .B(n20), .Z(n21) );
  NAND U24 ( .A(n21), .B(n2099), .Z(n22) );
  XNOR U25 ( .A(n22), .B(x[247]), .Z(n23) );
  NANDN U26 ( .A(y[247]), .B(n23), .Z(n24) );
  NANDN U27 ( .A(n22), .B(x[247]), .Z(n25) );
  AND U28 ( .A(n24), .B(n25), .Z(n2100) );
  NANDN U29 ( .A(y[256]), .B(x[256]), .Z(n26) );
  AND U30 ( .A(n1597), .B(n26), .Z(n27) );
  OR U31 ( .A(y[248]), .B(n2100), .Z(n28) );
  NAND U32 ( .A(n28), .B(n2103), .Z(n29) );
  AND U33 ( .A(n2104), .B(n29), .Z(n30) );
  OR U34 ( .A(n2105), .B(n30), .Z(n31) );
  NANDN U35 ( .A(n2106), .B(n31), .Z(n32) );
  ANDN U36 ( .B(n32), .A(n2107), .Z(n33) );
  OR U37 ( .A(n2108), .B(n33), .Z(n34) );
  NANDN U38 ( .A(n2109), .B(n34), .Z(n35) );
  ANDN U39 ( .B(n35), .A(n2110), .Z(n36) );
  NANDN U40 ( .A(x[256]), .B(y[256]), .Z(n37) );
  NANDN U41 ( .A(n36), .B(n27), .Z(n38) );
  NAND U42 ( .A(n38), .B(n37), .Z(n39) );
  NAND U43 ( .A(n39), .B(n1598), .Z(n40) );
  NANDN U44 ( .A(n2111), .B(n40), .Z(n41) );
  NANDN U45 ( .A(n2112), .B(n41), .Z(n42) );
  ANDN U46 ( .B(n42), .A(n2113), .Z(n2114) );
  ANDN U47 ( .B(n1991), .A(n1990), .Z(n43) );
  OR U48 ( .A(y[182]), .B(n43), .Z(n44) );
  XOR U49 ( .A(y[182]), .B(n43), .Z(n45) );
  NAND U50 ( .A(n45), .B(x[182]), .Z(n46) );
  NAND U51 ( .A(n44), .B(n46), .Z(n47) );
  AND U52 ( .A(n1992), .B(n47), .Z(n48) );
  OR U53 ( .A(n1993), .B(n48), .Z(n49) );
  NANDN U54 ( .A(n1994), .B(n49), .Z(n50) );
  ANDN U55 ( .B(n50), .A(n1995), .Z(n51) );
  OR U56 ( .A(n1996), .B(n51), .Z(n52) );
  NANDN U57 ( .A(n1997), .B(n52), .Z(n53) );
  ANDN U58 ( .B(n53), .A(n1998), .Z(n54) );
  OR U59 ( .A(n1999), .B(n54), .Z(n55) );
  NANDN U60 ( .A(n2000), .B(n55), .Z(n56) );
  ANDN U61 ( .B(n56), .A(n2001), .Z(n57) );
  OR U62 ( .A(n2002), .B(n57), .Z(n58) );
  NANDN U63 ( .A(n2003), .B(n58), .Z(n59) );
  NANDN U64 ( .A(n2004), .B(n59), .Z(n60) );
  NANDN U65 ( .A(n2005), .B(n60), .Z(n2006) );
  NANDN U66 ( .A(n2305), .B(n2304), .Z(n61) );
  AND U67 ( .A(n2306), .B(n61), .Z(n62) );
  NANDN U68 ( .A(x[346]), .B(y[346]), .Z(n63) );
  AND U69 ( .A(n62), .B(n63), .Z(n64) );
  ANDN U70 ( .B(n2309), .A(n2308), .Z(n65) );
  OR U71 ( .A(n2307), .B(n64), .Z(n66) );
  AND U72 ( .A(n65), .B(n66), .Z(n67) );
  NANDN U73 ( .A(y[349]), .B(x[349]), .Z(n68) );
  NANDN U74 ( .A(n67), .B(n68), .Z(n69) );
  ANDN U75 ( .B(n69), .A(n2310), .Z(n70) );
  AND U76 ( .A(n1587), .B(n1588), .Z(n71) );
  OR U77 ( .A(n2311), .B(n70), .Z(n72) );
  AND U78 ( .A(n71), .B(n72), .Z(n73) );
  OR U79 ( .A(n2312), .B(n73), .Z(n74) );
  NANDN U80 ( .A(n2313), .B(n74), .Z(n75) );
  NANDN U81 ( .A(n2314), .B(n75), .Z(n76) );
  NANDN U82 ( .A(n2315), .B(n76), .Z(n77) );
  NANDN U83 ( .A(n2316), .B(n77), .Z(n78) );
  ANDN U84 ( .B(n78), .A(n2317), .Z(n2318) );
  NANDN U85 ( .A(x[255]), .B(y[255]), .Z(n79) );
  NANDN U86 ( .A(x[254]), .B(y[254]), .Z(n80) );
  NAND U87 ( .A(n79), .B(n80), .Z(n2110) );
  ANDN U88 ( .B(y[384]), .A(x[384]), .Z(n1325) );
  NANDN U89 ( .A(n2549), .B(n2548), .Z(n81) );
  ANDN U90 ( .B(n81), .A(n2550), .Z(n82) );
  NANDN U91 ( .A(x[468]), .B(y[468]), .Z(n83) );
  ANDN U92 ( .B(n83), .A(n2551), .Z(n84) );
  XNOR U93 ( .A(x[468]), .B(y[468]), .Z(n85) );
  NAND U94 ( .A(n85), .B(n82), .Z(n86) );
  AND U95 ( .A(n84), .B(n86), .Z(n87) );
  OR U96 ( .A(n2552), .B(n87), .Z(n88) );
  NANDN U97 ( .A(n2553), .B(n88), .Z(n89) );
  ANDN U98 ( .B(n89), .A(n2554), .Z(n90) );
  OR U99 ( .A(n2555), .B(n90), .Z(n91) );
  NANDN U100 ( .A(n2556), .B(n91), .Z(n92) );
  ANDN U101 ( .B(n92), .A(n2557), .Z(n93) );
  OR U102 ( .A(n2558), .B(n93), .Z(n94) );
  NANDN U103 ( .A(n2559), .B(n94), .Z(n95) );
  ANDN U104 ( .B(n95), .A(n2560), .Z(n96) );
  OR U105 ( .A(n2561), .B(n96), .Z(n97) );
  NANDN U106 ( .A(n2562), .B(n97), .Z(n98) );
  AND U107 ( .A(n2563), .B(n98), .Z(n2565) );
  IV U108 ( .A(ebreg), .Z(e) );
  NANDN U109 ( .A(x[62]), .B(y[62]), .Z(n100) );
  NANDN U110 ( .A(x[63]), .B(y[63]), .Z(n99) );
  NAND U111 ( .A(n100), .B(n99), .Z(n1731) );
  NANDN U112 ( .A(x[58]), .B(y[58]), .Z(n102) );
  NANDN U113 ( .A(x[59]), .B(y[59]), .Z(n101) );
  NAND U114 ( .A(n102), .B(n101), .Z(n1724) );
  NANDN U115 ( .A(y[61]), .B(x[61]), .Z(n104) );
  NANDN U116 ( .A(y[62]), .B(x[62]), .Z(n103) );
  NAND U117 ( .A(n104), .B(n103), .Z(n1730) );
  NOR U118 ( .A(n1724), .B(n1730), .Z(n107) );
  NANDN U119 ( .A(y[65]), .B(x[65]), .Z(n106) );
  NANDN U120 ( .A(y[66]), .B(x[66]), .Z(n105) );
  NAND U121 ( .A(n106), .B(n105), .Z(n1738) );
  ANDN U122 ( .B(n107), .A(n1738), .Z(n108) );
  NANDN U123 ( .A(n1731), .B(n108), .Z(n144) );
  NANDN U124 ( .A(y[41]), .B(x[41]), .Z(n110) );
  NANDN U125 ( .A(y[42]), .B(x[42]), .Z(n109) );
  NAND U126 ( .A(n110), .B(n109), .Z(n1690) );
  NANDN U127 ( .A(x[30]), .B(y[30]), .Z(n112) );
  NANDN U128 ( .A(x[31]), .B(y[31]), .Z(n111) );
  NAND U129 ( .A(n112), .B(n111), .Z(n1667) );
  NANDN U130 ( .A(y[33]), .B(x[33]), .Z(n114) );
  NANDN U131 ( .A(y[34]), .B(x[34]), .Z(n113) );
  NAND U132 ( .A(n114), .B(n113), .Z(n1674) );
  NOR U133 ( .A(n1667), .B(n1674), .Z(n117) );
  NANDN U134 ( .A(x[42]), .B(y[42]), .Z(n116) );
  NANDN U135 ( .A(x[43]), .B(y[43]), .Z(n115) );
  NAND U136 ( .A(n116), .B(n115), .Z(n1691) );
  ANDN U137 ( .B(n117), .A(n1691), .Z(n118) );
  NANDN U138 ( .A(n1690), .B(n118), .Z(n130) );
  NANDN U139 ( .A(x[28]), .B(y[28]), .Z(n120) );
  NANDN U140 ( .A(x[29]), .B(y[29]), .Z(n119) );
  NAND U141 ( .A(n120), .B(n119), .Z(n1664) );
  NANDN U142 ( .A(x[22]), .B(y[22]), .Z(n122) );
  NANDN U143 ( .A(x[23]), .B(y[23]), .Z(n121) );
  NAND U144 ( .A(n122), .B(n121), .Z(n1652) );
  NANDN U145 ( .A(x[24]), .B(y[24]), .Z(n124) );
  NANDN U146 ( .A(x[25]), .B(y[25]), .Z(n123) );
  NAND U147 ( .A(n124), .B(n123), .Z(n1655) );
  NOR U148 ( .A(n1652), .B(n1655), .Z(n127) );
  NANDN U149 ( .A(x[36]), .B(y[36]), .Z(n126) );
  NANDN U150 ( .A(x[37]), .B(y[37]), .Z(n125) );
  NAND U151 ( .A(n126), .B(n125), .Z(n1679) );
  ANDN U152 ( .B(n127), .A(n1679), .Z(n128) );
  NANDN U153 ( .A(n1664), .B(n128), .Z(n129) );
  NOR U154 ( .A(n130), .B(n129), .Z(n142) );
  NANDN U155 ( .A(x[50]), .B(y[50]), .Z(n132) );
  NANDN U156 ( .A(x[51]), .B(y[51]), .Z(n131) );
  NAND U157 ( .A(n132), .B(n131), .Z(n1707) );
  NANDN U158 ( .A(y[51]), .B(x[51]), .Z(n134) );
  NANDN U159 ( .A(y[52]), .B(x[52]), .Z(n133) );
  NAND U160 ( .A(n134), .B(n133), .Z(n1710) );
  NANDN U161 ( .A(y[43]), .B(x[43]), .Z(n136) );
  NANDN U162 ( .A(y[44]), .B(x[44]), .Z(n135) );
  NAND U163 ( .A(n136), .B(n135), .Z(n1694) );
  NOR U164 ( .A(n1710), .B(n1694), .Z(n139) );
  NANDN U165 ( .A(y[57]), .B(x[57]), .Z(n138) );
  NANDN U166 ( .A(y[58]), .B(x[58]), .Z(n137) );
  NAND U167 ( .A(n138), .B(n137), .Z(n1722) );
  ANDN U168 ( .B(n139), .A(n1722), .Z(n140) );
  NANDN U169 ( .A(n1707), .B(n140), .Z(n141) );
  ANDN U170 ( .B(n142), .A(n141), .Z(n143) );
  NANDN U171 ( .A(n144), .B(n143), .Z(n476) );
  NANDN U172 ( .A(y[237]), .B(x[237]), .Z(n146) );
  NANDN U173 ( .A(y[238]), .B(x[238]), .Z(n145) );
  NAND U174 ( .A(n146), .B(n145), .Z(n2088) );
  NANDN U175 ( .A(y[285]), .B(x[285]), .Z(n148) );
  NANDN U176 ( .A(y[286]), .B(x[286]), .Z(n147) );
  NAND U177 ( .A(n148), .B(n147), .Z(n2167) );
  NANDN U178 ( .A(y[283]), .B(x[283]), .Z(n150) );
  NANDN U179 ( .A(y[284]), .B(x[284]), .Z(n149) );
  NAND U180 ( .A(n150), .B(n149), .Z(n2163) );
  NOR U181 ( .A(n2167), .B(n2163), .Z(n153) );
  NANDN U182 ( .A(y[147]), .B(x[147]), .Z(n152) );
  NANDN U183 ( .A(y[148]), .B(x[148]), .Z(n151) );
  NAND U184 ( .A(n152), .B(n151), .Z(n1921) );
  ANDN U185 ( .B(n153), .A(n1921), .Z(n154) );
  NANDN U186 ( .A(n2088), .B(n154), .Z(n236) );
  NANDN U187 ( .A(x[498]), .B(y[498]), .Z(n156) );
  NANDN U188 ( .A(x[499]), .B(y[499]), .Z(n155) );
  NAND U189 ( .A(n156), .B(n155), .Z(n2602) );
  ANDN U190 ( .B(x[264]), .A(y[264]), .Z(n1594) );
  NANDN U191 ( .A(y[263]), .B(x[263]), .Z(n158) );
  NANDN U192 ( .A(y[262]), .B(x[262]), .Z(n157) );
  AND U193 ( .A(n158), .B(n157), .Z(n159) );
  NANDN U194 ( .A(n1594), .B(n159), .Z(n2119) );
  NANDN U195 ( .A(y[499]), .B(x[499]), .Z(n161) );
  NANDN U196 ( .A(y[500]), .B(x[500]), .Z(n160) );
  NAND U197 ( .A(n161), .B(n160), .Z(n2605) );
  NOR U198 ( .A(n2119), .B(n2605), .Z(n173) );
  NANDN U199 ( .A(y[287]), .B(x[287]), .Z(n163) );
  NANDN U200 ( .A(y[288]), .B(x[288]), .Z(n162) );
  NAND U201 ( .A(n163), .B(n162), .Z(n2171) );
  NANDN U202 ( .A(x[344]), .B(y[344]), .Z(n165) );
  NANDN U203 ( .A(x[345]), .B(y[345]), .Z(n164) );
  NAND U204 ( .A(n165), .B(n164), .Z(n2303) );
  NANDN U205 ( .A(y[326]), .B(x[326]), .Z(n167) );
  NANDN U206 ( .A(y[327]), .B(x[327]), .Z(n166) );
  NAND U207 ( .A(n167), .B(n166), .Z(n2253) );
  NOR U208 ( .A(n2303), .B(n2253), .Z(n170) );
  NANDN U209 ( .A(x[284]), .B(y[284]), .Z(n169) );
  NANDN U210 ( .A(x[285]), .B(y[285]), .Z(n168) );
  NAND U211 ( .A(n169), .B(n168), .Z(n2165) );
  ANDN U212 ( .B(n170), .A(n2165), .Z(n171) );
  NANDN U213 ( .A(n2171), .B(n171), .Z(n172) );
  ANDN U214 ( .B(n173), .A(n172), .Z(n174) );
  NANDN U215 ( .A(n2602), .B(n174), .Z(n186) );
  NANDN U216 ( .A(x[3]), .B(y[3]), .Z(n176) );
  NANDN U217 ( .A(x[4]), .B(y[4]), .Z(n175) );
  NAND U218 ( .A(n176), .B(n175), .Z(n1610) );
  NANDN U219 ( .A(y[78]), .B(x[78]), .Z(n178) );
  NANDN U220 ( .A(y[79]), .B(x[79]), .Z(n177) );
  NAND U221 ( .A(n178), .B(n177), .Z(n1770) );
  NANDN U222 ( .A(x[1]), .B(y[1]), .Z(n180) );
  NANDN U223 ( .A(x[2]), .B(y[2]), .Z(n179) );
  NAND U224 ( .A(n180), .B(n179), .Z(n1604) );
  NOR U225 ( .A(n1770), .B(n1604), .Z(n183) );
  NANDN U226 ( .A(y[4]), .B(x[4]), .Z(n182) );
  NANDN U227 ( .A(y[5]), .B(x[5]), .Z(n181) );
  NAND U228 ( .A(n182), .B(n181), .Z(n1612) );
  ANDN U229 ( .B(n183), .A(n1612), .Z(n184) );
  NANDN U230 ( .A(n1610), .B(n184), .Z(n185) );
  NOR U231 ( .A(n186), .B(n185), .Z(n234) );
  NANDN U232 ( .A(y[23]), .B(x[23]), .Z(n188) );
  NANDN U233 ( .A(y[24]), .B(x[24]), .Z(n187) );
  NAND U234 ( .A(n188), .B(n187), .Z(n1654) );
  NANDN U235 ( .A(x[18]), .B(y[18]), .Z(n190) );
  NANDN U236 ( .A(x[19]), .B(y[19]), .Z(n189) );
  NAND U237 ( .A(n190), .B(n189), .Z(n1642) );
  NANDN U238 ( .A(y[19]), .B(x[19]), .Z(n192) );
  NANDN U239 ( .A(y[20]), .B(x[20]), .Z(n191) );
  NAND U240 ( .A(n192), .B(n191), .Z(n1644) );
  NOR U241 ( .A(n1642), .B(n1644), .Z(n195) );
  NANDN U242 ( .A(y[21]), .B(x[21]), .Z(n194) );
  NANDN U243 ( .A(y[22]), .B(x[22]), .Z(n193) );
  NAND U244 ( .A(n194), .B(n193), .Z(n1650) );
  ANDN U245 ( .B(n195), .A(n1650), .Z(n196) );
  NANDN U246 ( .A(n1654), .B(n196), .Z(n232) );
  NANDN U247 ( .A(y[11]), .B(x[11]), .Z(n198) );
  NANDN U248 ( .A(y[12]), .B(x[12]), .Z(n197) );
  NAND U249 ( .A(n198), .B(n197), .Z(n1628) );
  NANDN U250 ( .A(x[10]), .B(y[10]), .Z(n200) );
  NANDN U251 ( .A(x[11]), .B(y[11]), .Z(n199) );
  NAND U252 ( .A(n200), .B(n199), .Z(n1625) );
  NANDN U253 ( .A(y[13]), .B(x[13]), .Z(n202) );
  NANDN U254 ( .A(y[14]), .B(x[14]), .Z(n201) );
  NAND U255 ( .A(n202), .B(n201), .Z(n1632) );
  NOR U256 ( .A(n1625), .B(n1632), .Z(n205) );
  NANDN U257 ( .A(x[12]), .B(y[12]), .Z(n204) );
  NANDN U258 ( .A(x[13]), .B(y[13]), .Z(n203) );
  NAND U259 ( .A(n204), .B(n203), .Z(n1630) );
  ANDN U260 ( .B(n205), .A(n1630), .Z(n206) );
  NANDN U261 ( .A(n1628), .B(n206), .Z(n218) );
  NANDN U262 ( .A(y[6]), .B(x[6]), .Z(n208) );
  NANDN U263 ( .A(y[7]), .B(x[7]), .Z(n207) );
  NAND U264 ( .A(n208), .B(n207), .Z(n1616) );
  NANDN U265 ( .A(x[8]), .B(y[8]), .Z(n210) );
  NANDN U266 ( .A(x[9]), .B(y[9]), .Z(n209) );
  NAND U267 ( .A(n210), .B(n209), .Z(n1622) );
  NANDN U268 ( .A(x[5]), .B(y[5]), .Z(n212) );
  NANDN U269 ( .A(x[6]), .B(y[6]), .Z(n211) );
  NAND U270 ( .A(n212), .B(n211), .Z(n1613) );
  NOR U271 ( .A(n1622), .B(n1613), .Z(n215) );
  NANDN U272 ( .A(y[9]), .B(x[9]), .Z(n214) );
  NANDN U273 ( .A(y[10]), .B(x[10]), .Z(n213) );
  NAND U274 ( .A(n214), .B(n213), .Z(n1624) );
  ANDN U275 ( .B(n215), .A(n1624), .Z(n216) );
  NANDN U276 ( .A(n1616), .B(n216), .Z(n217) );
  NOR U277 ( .A(n218), .B(n217), .Z(n230) );
  NANDN U278 ( .A(x[16]), .B(y[16]), .Z(n220) );
  NANDN U279 ( .A(x[17]), .B(y[17]), .Z(n219) );
  NAND U280 ( .A(n220), .B(n219), .Z(n1637) );
  NANDN U281 ( .A(x[14]), .B(y[14]), .Z(n222) );
  NANDN U282 ( .A(x[15]), .B(y[15]), .Z(n221) );
  NAND U283 ( .A(n222), .B(n221), .Z(n1634) );
  NANDN U284 ( .A(y[15]), .B(x[15]), .Z(n224) );
  NANDN U285 ( .A(y[16]), .B(x[16]), .Z(n223) );
  NAND U286 ( .A(n224), .B(n223), .Z(n1636) );
  NOR U287 ( .A(n1634), .B(n1636), .Z(n227) );
  NANDN U288 ( .A(y[17]), .B(x[17]), .Z(n226) );
  NANDN U289 ( .A(y[18]), .B(x[18]), .Z(n225) );
  NAND U290 ( .A(n226), .B(n225), .Z(n1640) );
  ANDN U291 ( .B(n227), .A(n1640), .Z(n228) );
  NANDN U292 ( .A(n1637), .B(n228), .Z(n229) );
  ANDN U293 ( .B(n230), .A(n229), .Z(n231) );
  NANDN U294 ( .A(n232), .B(n231), .Z(n233) );
  ANDN U295 ( .B(n234), .A(n233), .Z(n235) );
  NANDN U296 ( .A(n236), .B(n235), .Z(n284) );
  NANDN U297 ( .A(y[101]), .B(x[101]), .Z(n238) );
  NANDN U298 ( .A(y[102]), .B(x[102]), .Z(n237) );
  NAND U299 ( .A(n238), .B(n237), .Z(n1820) );
  NANDN U300 ( .A(y[87]), .B(x[87]), .Z(n240) );
  NANDN U301 ( .A(y[88]), .B(x[88]), .Z(n239) );
  NAND U302 ( .A(n240), .B(n239), .Z(n1790) );
  NANDN U303 ( .A(x[100]), .B(y[100]), .Z(n242) );
  NANDN U304 ( .A(x[101]), .B(y[101]), .Z(n241) );
  NAND U305 ( .A(n242), .B(n241), .Z(n1818) );
  NOR U306 ( .A(n1790), .B(n1818), .Z(n245) );
  NANDN U307 ( .A(x[102]), .B(y[102]), .Z(n244) );
  NANDN U308 ( .A(x[103]), .B(y[103]), .Z(n243) );
  NAND U309 ( .A(n244), .B(n243), .Z(n1821) );
  ANDN U310 ( .B(n245), .A(n1821), .Z(n246) );
  NANDN U311 ( .A(n1820), .B(n246), .Z(n282) );
  NANDN U312 ( .A(x[82]), .B(y[82]), .Z(n248) );
  NANDN U313 ( .A(x[83]), .B(y[83]), .Z(n247) );
  NAND U314 ( .A(n248), .B(n247), .Z(n1779) );
  NANDN U315 ( .A(x[77]), .B(y[77]), .Z(n250) );
  NANDN U316 ( .A(x[76]), .B(y[76]), .Z(n249) );
  NAND U317 ( .A(n250), .B(n249), .Z(n1764) );
  NANDN U318 ( .A(x[80]), .B(y[80]), .Z(n252) );
  NANDN U319 ( .A(x[81]), .B(y[81]), .Z(n251) );
  NAND U320 ( .A(n252), .B(n251), .Z(n1776) );
  NOR U321 ( .A(n1764), .B(n1776), .Z(n255) );
  NANDN U322 ( .A(y[83]), .B(x[83]), .Z(n254) );
  NANDN U323 ( .A(y[84]), .B(x[84]), .Z(n253) );
  NAND U324 ( .A(n254), .B(n253), .Z(n1782) );
  ANDN U325 ( .B(n255), .A(n1782), .Z(n256) );
  NANDN U326 ( .A(n1779), .B(n256), .Z(n268) );
  NANDN U327 ( .A(y[71]), .B(x[71]), .Z(n258) );
  NANDN U328 ( .A(y[72]), .B(x[72]), .Z(n257) );
  NAND U329 ( .A(n258), .B(n257), .Z(n1752) );
  NANDN U330 ( .A(x[70]), .B(y[70]), .Z(n260) );
  NANDN U331 ( .A(x[71]), .B(y[71]), .Z(n259) );
  NAND U332 ( .A(n260), .B(n259), .Z(n1749) );
  NANDN U333 ( .A(x[74]), .B(y[74]), .Z(n262) );
  NANDN U334 ( .A(x[75]), .B(y[75]), .Z(n261) );
  NAND U335 ( .A(n262), .B(n261), .Z(n1758) );
  NOR U336 ( .A(n1749), .B(n1758), .Z(n265) );
  NANDN U337 ( .A(x[72]), .B(y[72]), .Z(n264) );
  NANDN U338 ( .A(x[73]), .B(y[73]), .Z(n263) );
  NAND U339 ( .A(n264), .B(n263), .Z(n1754) );
  ANDN U340 ( .B(n265), .A(n1754), .Z(n266) );
  NANDN U341 ( .A(n1752), .B(n266), .Z(n267) );
  NOR U342 ( .A(n268), .B(n267), .Z(n280) );
  NANDN U343 ( .A(x[90]), .B(y[90]), .Z(n270) );
  NANDN U344 ( .A(x[91]), .B(y[91]), .Z(n269) );
  NAND U345 ( .A(n270), .B(n269), .Z(n1797) );
  NANDN U346 ( .A(x[84]), .B(y[84]), .Z(n272) );
  NANDN U347 ( .A(x[85]), .B(y[85]), .Z(n271) );
  NAND U348 ( .A(n272), .B(n271), .Z(n1784) );
  NANDN U349 ( .A(y[85]), .B(x[85]), .Z(n274) );
  NANDN U350 ( .A(y[86]), .B(x[86]), .Z(n273) );
  NAND U351 ( .A(n274), .B(n273), .Z(n1786) );
  NOR U352 ( .A(n1784), .B(n1786), .Z(n277) );
  NANDN U353 ( .A(x[86]), .B(y[86]), .Z(n276) );
  NANDN U354 ( .A(x[87]), .B(y[87]), .Z(n275) );
  NAND U355 ( .A(n276), .B(n275), .Z(n1788) );
  ANDN U356 ( .B(n277), .A(n1788), .Z(n278) );
  NANDN U357 ( .A(n1797), .B(n278), .Z(n279) );
  ANDN U358 ( .B(n280), .A(n279), .Z(n281) );
  NANDN U359 ( .A(n282), .B(n281), .Z(n283) );
  NOR U360 ( .A(n284), .B(n283), .Z(n474) );
  NANDN U361 ( .A(y[305]), .B(x[305]), .Z(n286) );
  NANDN U362 ( .A(y[306]), .B(x[306]), .Z(n285) );
  NAND U363 ( .A(n286), .B(n285), .Z(n2209) );
  NANDN U364 ( .A(x[302]), .B(y[302]), .Z(n288) );
  NANDN U365 ( .A(x[303]), .B(y[303]), .Z(n287) );
  NAND U366 ( .A(n288), .B(n287), .Z(n2203) );
  NANDN U367 ( .A(x[304]), .B(y[304]), .Z(n290) );
  NANDN U368 ( .A(x[305]), .B(y[305]), .Z(n289) );
  NAND U369 ( .A(n290), .B(n289), .Z(n2207) );
  NOR U370 ( .A(n2203), .B(n2207), .Z(n293) );
  NANDN U371 ( .A(x[306]), .B(y[306]), .Z(n292) );
  NANDN U372 ( .A(x[307]), .B(y[307]), .Z(n291) );
  NAND U373 ( .A(n292), .B(n291), .Z(n2210) );
  ANDN U374 ( .B(n293), .A(n2210), .Z(n294) );
  NANDN U375 ( .A(n2209), .B(n294), .Z(n330) );
  NANDN U376 ( .A(y[291]), .B(x[291]), .Z(n296) );
  NANDN U377 ( .A(y[292]), .B(x[292]), .Z(n295) );
  NAND U378 ( .A(n296), .B(n295), .Z(n2181) );
  NANDN U379 ( .A(x[286]), .B(y[286]), .Z(n298) );
  NANDN U380 ( .A(x[287]), .B(y[287]), .Z(n297) );
  NAND U381 ( .A(n298), .B(n297), .Z(n2168) );
  NANDN U382 ( .A(y[289]), .B(x[289]), .Z(n300) );
  NANDN U383 ( .A(y[290]), .B(x[290]), .Z(n299) );
  NAND U384 ( .A(n300), .B(n299), .Z(n2175) );
  NOR U385 ( .A(n2168), .B(n2175), .Z(n303) );
  NANDN U386 ( .A(y[295]), .B(x[295]), .Z(n302) );
  NANDN U387 ( .A(y[296]), .B(x[296]), .Z(n301) );
  NAND U388 ( .A(n302), .B(n301), .Z(n2189) );
  ANDN U389 ( .B(n303), .A(n2189), .Z(n304) );
  NANDN U390 ( .A(n2181), .B(n304), .Z(n316) );
  NANDN U391 ( .A(y[277]), .B(x[277]), .Z(n306) );
  NANDN U392 ( .A(y[278]), .B(x[278]), .Z(n305) );
  NAND U393 ( .A(n306), .B(n305), .Z(n2149) );
  NANDN U394 ( .A(x[276]), .B(y[276]), .Z(n308) );
  NANDN U395 ( .A(x[277]), .B(y[277]), .Z(n307) );
  NAND U396 ( .A(n308), .B(n307), .Z(n2147) );
  NANDN U397 ( .A(y[281]), .B(x[281]), .Z(n310) );
  NANDN U398 ( .A(y[282]), .B(x[282]), .Z(n309) );
  NAND U399 ( .A(n310), .B(n309), .Z(n2157) );
  NOR U400 ( .A(n2147), .B(n2157), .Z(n313) );
  NANDN U401 ( .A(x[280]), .B(y[280]), .Z(n312) );
  NANDN U402 ( .A(x[281]), .B(y[281]), .Z(n311) );
  NAND U403 ( .A(n312), .B(n311), .Z(n2155) );
  ANDN U404 ( .B(n313), .A(n2155), .Z(n314) );
  NANDN U405 ( .A(n2149), .B(n314), .Z(n315) );
  NOR U406 ( .A(n316), .B(n315), .Z(n328) );
  NANDN U407 ( .A(y[303]), .B(x[303]), .Z(n318) );
  NANDN U408 ( .A(y[304]), .B(x[304]), .Z(n317) );
  NAND U409 ( .A(n318), .B(n317), .Z(n2205) );
  NANDN U410 ( .A(x[296]), .B(y[296]), .Z(n320) );
  NANDN U411 ( .A(x[297]), .B(y[297]), .Z(n319) );
  NAND U412 ( .A(n320), .B(n319), .Z(n2191) );
  NANDN U413 ( .A(x[298]), .B(y[298]), .Z(n322) );
  NANDN U414 ( .A(x[299]), .B(y[299]), .Z(n321) );
  NAND U415 ( .A(n322), .B(n321), .Z(n2195) );
  NOR U416 ( .A(n2191), .B(n2195), .Z(n325) );
  NANDN U417 ( .A(x[300]), .B(y[300]), .Z(n324) );
  NANDN U418 ( .A(x[301]), .B(y[301]), .Z(n323) );
  NAND U419 ( .A(n324), .B(n323), .Z(n2198) );
  ANDN U420 ( .B(n325), .A(n2198), .Z(n326) );
  NANDN U421 ( .A(n2205), .B(n326), .Z(n327) );
  ANDN U422 ( .B(n328), .A(n327), .Z(n329) );
  NANDN U423 ( .A(n330), .B(n329), .Z(n472) );
  NANDN U424 ( .A(x[228]), .B(y[228]), .Z(n332) );
  NANDN U425 ( .A(x[229]), .B(y[229]), .Z(n331) );
  NAND U426 ( .A(n332), .B(n331), .Z(n2071) );
  NANDN U427 ( .A(y[207]), .B(x[207]), .Z(n334) );
  NANDN U428 ( .A(y[208]), .B(x[208]), .Z(n333) );
  NAND U429 ( .A(n334), .B(n333), .Z(n2029) );
  NANDN U430 ( .A(y[215]), .B(x[215]), .Z(n336) );
  NANDN U431 ( .A(y[216]), .B(x[216]), .Z(n335) );
  NAND U432 ( .A(n336), .B(n335), .Z(n2045) );
  NOR U433 ( .A(n2029), .B(n2045), .Z(n339) );
  NANDN U434 ( .A(x[234]), .B(y[234]), .Z(n338) );
  NANDN U435 ( .A(x[235]), .B(y[235]), .Z(n337) );
  NAND U436 ( .A(n338), .B(n337), .Z(n2083) );
  ANDN U437 ( .B(n339), .A(n2083), .Z(n340) );
  NANDN U438 ( .A(n2071), .B(n340), .Z(n376) );
  NANDN U439 ( .A(x[204]), .B(y[204]), .Z(n342) );
  NANDN U440 ( .A(x[205]), .B(y[205]), .Z(n341) );
  NAND U441 ( .A(n342), .B(n341), .Z(n2023) );
  NANDN U442 ( .A(x[194]), .B(y[194]), .Z(n344) );
  NANDN U443 ( .A(x[195]), .B(y[195]), .Z(n343) );
  NAND U444 ( .A(n344), .B(n343), .Z(n2004) );
  NANDN U445 ( .A(x[198]), .B(y[198]), .Z(n346) );
  NANDN U446 ( .A(x[199]), .B(y[199]), .Z(n345) );
  NAND U447 ( .A(n346), .B(n345), .Z(n2011) );
  NOR U448 ( .A(n2004), .B(n2011), .Z(n349) );
  NANDN U449 ( .A(x[202]), .B(y[202]), .Z(n348) );
  NANDN U450 ( .A(x[203]), .B(y[203]), .Z(n347) );
  NAND U451 ( .A(n348), .B(n347), .Z(n2019) );
  ANDN U452 ( .B(n349), .A(n2019), .Z(n350) );
  NANDN U453 ( .A(n2023), .B(n350), .Z(n362) );
  NANDN U454 ( .A(y[187]), .B(x[187]), .Z(n352) );
  NANDN U455 ( .A(y[188]), .B(x[188]), .Z(n351) );
  NAND U456 ( .A(n352), .B(n351), .Z(n1997) );
  NANDN U457 ( .A(x[176]), .B(y[176]), .Z(n354) );
  NANDN U458 ( .A(x[177]), .B(y[177]), .Z(n353) );
  NAND U459 ( .A(n354), .B(n353), .Z(n1981) );
  NANDN U460 ( .A(x[180]), .B(y[180]), .Z(n356) );
  NANDN U461 ( .A(x[181]), .B(y[181]), .Z(n355) );
  NAND U462 ( .A(n356), .B(n355), .Z(n1989) );
  NOR U463 ( .A(n1981), .B(n1989), .Z(n359) );
  NANDN U464 ( .A(x[190]), .B(y[190]), .Z(n358) );
  NANDN U465 ( .A(x[191]), .B(y[191]), .Z(n357) );
  NAND U466 ( .A(n358), .B(n357), .Z(n2000) );
  ANDN U467 ( .B(n359), .A(n2000), .Z(n360) );
  NANDN U468 ( .A(n1997), .B(n360), .Z(n361) );
  NOR U469 ( .A(n362), .B(n361), .Z(n374) );
  NANDN U470 ( .A(x[206]), .B(y[206]), .Z(n364) );
  NANDN U471 ( .A(x[207]), .B(y[207]), .Z(n363) );
  NAND U472 ( .A(n364), .B(n363), .Z(n2026) );
  NANDN U473 ( .A(y[203]), .B(x[203]), .Z(n366) );
  NANDN U474 ( .A(y[204]), .B(x[204]), .Z(n365) );
  NAND U475 ( .A(n366), .B(n365), .Z(n2021) );
  NANDN U476 ( .A(y[205]), .B(x[205]), .Z(n368) );
  NANDN U477 ( .A(y[206]), .B(x[206]), .Z(n367) );
  NAND U478 ( .A(n368), .B(n367), .Z(n2025) );
  NOR U479 ( .A(n2021), .B(n2025), .Z(n371) );
  NANDN U480 ( .A(y[227]), .B(x[227]), .Z(n370) );
  NANDN U481 ( .A(y[228]), .B(x[228]), .Z(n369) );
  NAND U482 ( .A(n370), .B(n369), .Z(n2069) );
  ANDN U483 ( .B(n371), .A(n2069), .Z(n372) );
  NANDN U484 ( .A(n2026), .B(n372), .Z(n373) );
  ANDN U485 ( .B(n374), .A(n373), .Z(n375) );
  NANDN U486 ( .A(n376), .B(n375), .Z(n424) );
  NANDN U487 ( .A(y[167]), .B(x[167]), .Z(n378) );
  NANDN U488 ( .A(y[168]), .B(x[168]), .Z(n377) );
  NAND U489 ( .A(n378), .B(n377), .Z(n1963) );
  NANDN U490 ( .A(x[164]), .B(y[164]), .Z(n380) );
  NANDN U491 ( .A(x[165]), .B(y[165]), .Z(n379) );
  NAND U492 ( .A(n380), .B(n379), .Z(n1957) );
  NANDN U493 ( .A(x[174]), .B(y[174]), .Z(n382) );
  NANDN U494 ( .A(x[175]), .B(y[175]), .Z(n381) );
  NAND U495 ( .A(n382), .B(n381), .Z(n1977) );
  NOR U496 ( .A(n1957), .B(n1977), .Z(n385) );
  NANDN U497 ( .A(x[170]), .B(y[170]), .Z(n384) );
  NANDN U498 ( .A(x[171]), .B(y[171]), .Z(n383) );
  NAND U499 ( .A(n384), .B(n383), .Z(n1969) );
  ANDN U500 ( .B(n385), .A(n1969), .Z(n386) );
  NANDN U501 ( .A(n1963), .B(n386), .Z(n422) );
  NANDN U502 ( .A(x[126]), .B(y[126]), .Z(n388) );
  NANDN U503 ( .A(x[127]), .B(y[127]), .Z(n387) );
  NAND U504 ( .A(n388), .B(n387), .Z(n1869) );
  NANDN U505 ( .A(y[119]), .B(x[119]), .Z(n390) );
  NANDN U506 ( .A(y[120]), .B(x[120]), .Z(n389) );
  NAND U507 ( .A(n390), .B(n389), .Z(n1856) );
  NANDN U508 ( .A(x[120]), .B(y[120]), .Z(n392) );
  NANDN U509 ( .A(x[121]), .B(y[121]), .Z(n391) );
  NAND U510 ( .A(n392), .B(n391), .Z(n1857) );
  NOR U511 ( .A(n1856), .B(n1857), .Z(n395) );
  NANDN U512 ( .A(y[135]), .B(x[135]), .Z(n394) );
  NANDN U513 ( .A(y[136]), .B(x[136]), .Z(n393) );
  NAND U514 ( .A(n394), .B(n393), .Z(n1890) );
  ANDN U515 ( .B(n395), .A(n1890), .Z(n396) );
  NANDN U516 ( .A(n1869), .B(n396), .Z(n408) );
  NANDN U517 ( .A(x[112]), .B(y[112]), .Z(n398) );
  NANDN U518 ( .A(x[113]), .B(y[113]), .Z(n397) );
  NAND U519 ( .A(n398), .B(n397), .Z(n1842) );
  NANDN U520 ( .A(y[103]), .B(x[103]), .Z(n400) );
  NANDN U521 ( .A(y[104]), .B(x[104]), .Z(n399) );
  NAND U522 ( .A(n400), .B(n399), .Z(n1824) );
  NANDN U523 ( .A(y[107]), .B(x[107]), .Z(n402) );
  NANDN U524 ( .A(y[108]), .B(x[108]), .Z(n401) );
  NAND U525 ( .A(n402), .B(n401), .Z(n1832) );
  NOR U526 ( .A(n1824), .B(n1832), .Z(n405) );
  NANDN U527 ( .A(y[121]), .B(x[121]), .Z(n404) );
  NANDN U528 ( .A(y[122]), .B(x[122]), .Z(n403) );
  NAND U529 ( .A(n404), .B(n403), .Z(n1860) );
  ANDN U530 ( .B(n405), .A(n1860), .Z(n406) );
  NANDN U531 ( .A(n1842), .B(n406), .Z(n407) );
  NOR U532 ( .A(n408), .B(n407), .Z(n420) );
  NANDN U533 ( .A(x[148]), .B(y[148]), .Z(n410) );
  NANDN U534 ( .A(x[149]), .B(y[149]), .Z(n409) );
  NAND U535 ( .A(n410), .B(n409), .Z(n1923) );
  NANDN U536 ( .A(y[159]), .B(x[159]), .Z(n412) );
  NANDN U537 ( .A(y[160]), .B(x[160]), .Z(n411) );
  NAND U538 ( .A(n412), .B(n411), .Z(n1947) );
  NANDN U539 ( .A(x[136]), .B(y[136]), .Z(n414) );
  NANDN U540 ( .A(x[137]), .B(y[137]), .Z(n413) );
  NAND U541 ( .A(n414), .B(n413), .Z(n1892) );
  NOR U542 ( .A(n1947), .B(n1892), .Z(n417) );
  NANDN U543 ( .A(x[160]), .B(y[160]), .Z(n416) );
  NANDN U544 ( .A(x[161]), .B(y[161]), .Z(n415) );
  NAND U545 ( .A(n416), .B(n415), .Z(n1948) );
  ANDN U546 ( .B(n417), .A(n1948), .Z(n418) );
  NANDN U547 ( .A(n1923), .B(n418), .Z(n419) );
  ANDN U548 ( .B(n420), .A(n419), .Z(n421) );
  NANDN U549 ( .A(n422), .B(n421), .Z(n423) );
  NOR U550 ( .A(n424), .B(n423), .Z(n470) );
  NANDN U551 ( .A(x[270]), .B(y[270]), .Z(n426) );
  NANDN U552 ( .A(x[271]), .B(y[271]), .Z(n425) );
  NAND U553 ( .A(n426), .B(n425), .Z(n2135) );
  NANDN U554 ( .A(y[271]), .B(x[271]), .Z(n428) );
  NANDN U555 ( .A(y[272]), .B(x[272]), .Z(n427) );
  NAND U556 ( .A(n428), .B(n427), .Z(n2137) );
  NANDN U557 ( .A(y[269]), .B(x[269]), .Z(n430) );
  NANDN U558 ( .A(y[270]), .B(x[270]), .Z(n429) );
  NAND U559 ( .A(n430), .B(n429), .Z(n2133) );
  NOR U560 ( .A(n2137), .B(n2133), .Z(n433) );
  NANDN U561 ( .A(y[275]), .B(x[275]), .Z(n432) );
  NANDN U562 ( .A(y[276]), .B(x[276]), .Z(n431) );
  NAND U563 ( .A(n432), .B(n431), .Z(n2145) );
  ANDN U564 ( .B(n433), .A(n2145), .Z(n434) );
  NANDN U565 ( .A(n2135), .B(n434), .Z(n468) );
  NANDN U566 ( .A(y[258]), .B(x[258]), .Z(n436) );
  NANDN U567 ( .A(y[259]), .B(x[259]), .Z(n435) );
  NAND U568 ( .A(n436), .B(n435), .Z(n2112) );
  NANDN U569 ( .A(x[257]), .B(y[257]), .Z(n438) );
  NANDN U570 ( .A(x[258]), .B(y[258]), .Z(n437) );
  NAND U571 ( .A(n438), .B(n437), .Z(n2111) );
  NOR U572 ( .A(n2110), .B(n2111), .Z(n441) );
  NANDN U573 ( .A(x[259]), .B(y[259]), .Z(n440) );
  NANDN U574 ( .A(x[260]), .B(y[260]), .Z(n439) );
  NAND U575 ( .A(n440), .B(n439), .Z(n2113) );
  ANDN U576 ( .B(n441), .A(n2113), .Z(n442) );
  NANDN U577 ( .A(n2112), .B(n442), .Z(n454) );
  NANDN U578 ( .A(y[241]), .B(x[241]), .Z(n444) );
  NANDN U579 ( .A(y[242]), .B(x[242]), .Z(n443) );
  NAND U580 ( .A(n444), .B(n443), .Z(n2093) );
  NANDN U581 ( .A(y[249]), .B(x[249]), .Z(n446) );
  NANDN U582 ( .A(y[250]), .B(x[250]), .Z(n445) );
  NAND U583 ( .A(n446), .B(n445), .Z(n2105) );
  NANDN U584 ( .A(x[238]), .B(y[238]), .Z(n448) );
  NANDN U585 ( .A(x[239]), .B(y[239]), .Z(n447) );
  NAND U586 ( .A(n448), .B(n447), .Z(n2089) );
  NOR U587 ( .A(n2105), .B(n2089), .Z(n451) );
  NANDN U588 ( .A(x[252]), .B(y[252]), .Z(n450) );
  NANDN U589 ( .A(x[253]), .B(y[253]), .Z(n449) );
  NAND U590 ( .A(n450), .B(n449), .Z(n2108) );
  ANDN U591 ( .B(n451), .A(n2108), .Z(n452) );
  NANDN U592 ( .A(n2093), .B(n452), .Z(n453) );
  NOR U593 ( .A(n454), .B(n453), .Z(n466) );
  NANDN U594 ( .A(x[266]), .B(y[266]), .Z(n456) );
  NANDN U595 ( .A(x[267]), .B(y[267]), .Z(n455) );
  NAND U596 ( .A(n456), .B(n455), .Z(n2126) );
  NANDN U597 ( .A(y[260]), .B(x[260]), .Z(n458) );
  NANDN U598 ( .A(y[261]), .B(x[261]), .Z(n457) );
  NAND U599 ( .A(n458), .B(n457), .Z(n2115) );
  NANDN U600 ( .A(x[264]), .B(y[264]), .Z(n460) );
  NANDN U601 ( .A(x[265]), .B(y[265]), .Z(n459) );
  NAND U602 ( .A(n460), .B(n459), .Z(n2123) );
  NOR U603 ( .A(n2115), .B(n2123), .Z(n463) );
  NANDN U604 ( .A(x[268]), .B(y[268]), .Z(n462) );
  NANDN U605 ( .A(x[269]), .B(y[269]), .Z(n461) );
  NAND U606 ( .A(n462), .B(n461), .Z(n2131) );
  ANDN U607 ( .B(n463), .A(n2131), .Z(n464) );
  NANDN U608 ( .A(n2126), .B(n464), .Z(n465) );
  ANDN U609 ( .B(n466), .A(n465), .Z(n467) );
  NANDN U610 ( .A(n468), .B(n467), .Z(n469) );
  ANDN U611 ( .B(n470), .A(n469), .Z(n471) );
  NANDN U612 ( .A(n472), .B(n471), .Z(n473) );
  ANDN U613 ( .B(n474), .A(n473), .Z(n475) );
  NANDN U614 ( .A(n476), .B(n475), .Z(n668) );
  NANDN U615 ( .A(x[92]), .B(y[92]), .Z(n478) );
  NANDN U616 ( .A(x[93]), .B(y[93]), .Z(n477) );
  NAND U617 ( .A(n478), .B(n477), .Z(n1802) );
  NANDN U618 ( .A(y[89]), .B(x[89]), .Z(n480) );
  NANDN U619 ( .A(y[90]), .B(x[90]), .Z(n479) );
  NAND U620 ( .A(n480), .B(n479), .Z(n1796) );
  NANDN U621 ( .A(y[91]), .B(x[91]), .Z(n482) );
  NANDN U622 ( .A(y[92]), .B(x[92]), .Z(n481) );
  NAND U623 ( .A(n482), .B(n481), .Z(n1800) );
  NOR U624 ( .A(n1796), .B(n1800), .Z(n485) );
  NANDN U625 ( .A(x[94]), .B(y[94]), .Z(n484) );
  NANDN U626 ( .A(x[95]), .B(y[95]), .Z(n483) );
  NAND U627 ( .A(n484), .B(n483), .Z(n1806) );
  ANDN U628 ( .B(n485), .A(n1806), .Z(n486) );
  NANDN U629 ( .A(n1802), .B(n486), .Z(n522) );
  NANDN U630 ( .A(y[63]), .B(x[63]), .Z(n488) );
  NANDN U631 ( .A(y[64]), .B(x[64]), .Z(n487) );
  NAND U632 ( .A(n488), .B(n487), .Z(n1734) );
  NANDN U633 ( .A(x[56]), .B(y[56]), .Z(n490) );
  NANDN U634 ( .A(x[57]), .B(y[57]), .Z(n489) );
  NAND U635 ( .A(n490), .B(n489), .Z(n1719) );
  NANDN U636 ( .A(x[60]), .B(y[60]), .Z(n492) );
  NANDN U637 ( .A(x[61]), .B(y[61]), .Z(n491) );
  NAND U638 ( .A(n492), .B(n491), .Z(n1728) );
  NOR U639 ( .A(n1719), .B(n1728), .Z(n495) );
  NANDN U640 ( .A(x[68]), .B(y[68]), .Z(n494) );
  NANDN U641 ( .A(x[69]), .B(y[69]), .Z(n493) );
  NAND U642 ( .A(n494), .B(n493), .Z(n1746) );
  ANDN U643 ( .B(n495), .A(n1746), .Z(n496) );
  NANDN U644 ( .A(n1734), .B(n496), .Z(n508) );
  NANDN U645 ( .A(y[59]), .B(x[59]), .Z(n498) );
  NANDN U646 ( .A(y[60]), .B(x[60]), .Z(n497) );
  NAND U647 ( .A(n498), .B(n497), .Z(n1726) );
  NANDN U648 ( .A(x[52]), .B(y[52]), .Z(n500) );
  NANDN U649 ( .A(x[53]), .B(y[53]), .Z(n499) );
  NAND U650 ( .A(n500), .B(n499), .Z(n1712) );
  NANDN U651 ( .A(y[53]), .B(x[53]), .Z(n502) );
  NANDN U652 ( .A(y[54]), .B(x[54]), .Z(n501) );
  NAND U653 ( .A(n502), .B(n501), .Z(n1714) );
  NOR U654 ( .A(n1712), .B(n1714), .Z(n505) );
  NANDN U655 ( .A(y[55]), .B(x[55]), .Z(n504) );
  NANDN U656 ( .A(y[56]), .B(x[56]), .Z(n503) );
  NAND U657 ( .A(n504), .B(n503), .Z(n1718) );
  ANDN U658 ( .B(n505), .A(n1718), .Z(n506) );
  NANDN U659 ( .A(n1726), .B(n506), .Z(n507) );
  NOR U660 ( .A(n508), .B(n507), .Z(n520) );
  NANDN U661 ( .A(y[69]), .B(x[69]), .Z(n510) );
  NANDN U662 ( .A(y[70]), .B(x[70]), .Z(n509) );
  NAND U663 ( .A(n510), .B(n509), .Z(n1748) );
  NANDN U664 ( .A(x[64]), .B(y[64]), .Z(n512) );
  NANDN U665 ( .A(x[65]), .B(y[65]), .Z(n511) );
  NAND U666 ( .A(n512), .B(n511), .Z(n1736) );
  NANDN U667 ( .A(x[66]), .B(y[66]), .Z(n514) );
  NANDN U668 ( .A(x[67]), .B(y[67]), .Z(n513) );
  NAND U669 ( .A(n514), .B(n513), .Z(n1740) );
  NOR U670 ( .A(n1736), .B(n1740), .Z(n517) );
  NANDN U671 ( .A(y[73]), .B(x[73]), .Z(n516) );
  NANDN U672 ( .A(y[74]), .B(x[74]), .Z(n515) );
  NAND U673 ( .A(n516), .B(n515), .Z(n1756) );
  ANDN U674 ( .B(n517), .A(n1756), .Z(n518) );
  NANDN U675 ( .A(n1748), .B(n518), .Z(n519) );
  ANDN U676 ( .B(n520), .A(n519), .Z(n521) );
  NANDN U677 ( .A(n522), .B(n521), .Z(n666) );
  NANDN U678 ( .A(y[105]), .B(x[105]), .Z(n524) );
  NANDN U679 ( .A(y[106]), .B(x[106]), .Z(n523) );
  NAND U680 ( .A(n524), .B(n523), .Z(n1828) );
  NANDN U681 ( .A(y[157]), .B(x[157]), .Z(n526) );
  NANDN U682 ( .A(y[158]), .B(x[158]), .Z(n525) );
  NAND U683 ( .A(n526), .B(n525), .Z(n1943) );
  NANDN U684 ( .A(y[169]), .B(x[169]), .Z(n528) );
  NANDN U685 ( .A(y[170]), .B(x[170]), .Z(n527) );
  NAND U686 ( .A(n528), .B(n527), .Z(n1967) );
  NOR U687 ( .A(n1943), .B(n1967), .Z(n531) );
  NANDN U688 ( .A(y[93]), .B(x[93]), .Z(n530) );
  NANDN U689 ( .A(y[94]), .B(x[94]), .Z(n529) );
  NAND U690 ( .A(n530), .B(n529), .Z(n1804) );
  ANDN U691 ( .B(n531), .A(n1804), .Z(n532) );
  NANDN U692 ( .A(n1828), .B(n532), .Z(n568) );
  NANDN U693 ( .A(x[472]), .B(y[472]), .Z(n534) );
  NANDN U694 ( .A(x[473]), .B(y[473]), .Z(n533) );
  NAND U695 ( .A(n534), .B(n533), .Z(n2555) );
  NANDN U696 ( .A(y[0]), .B(x[0]), .Z(n536) );
  NANDN U697 ( .A(y[1]), .B(x[1]), .Z(n535) );
  AND U698 ( .A(n536), .B(n535), .Z(n1603) );
  NANDN U699 ( .A(x[510]), .B(y[510]), .Z(n538) );
  NANDN U700 ( .A(x[511]), .B(y[511]), .Z(n537) );
  NAND U701 ( .A(n538), .B(n537), .Z(n2631) );
  ANDN U702 ( .B(n1603), .A(n2631), .Z(n541) );
  NANDN U703 ( .A(x[412]), .B(y[412]), .Z(n540) );
  NANDN U704 ( .A(x[413]), .B(y[413]), .Z(n539) );
  NAND U705 ( .A(n540), .B(n539), .Z(n2433) );
  ANDN U706 ( .B(n541), .A(n2433), .Z(n542) );
  NANDN U707 ( .A(n2555), .B(n542), .Z(n554) );
  NANDN U708 ( .A(x[504]), .B(y[504]), .Z(n544) );
  NANDN U709 ( .A(x[505]), .B(y[505]), .Z(n543) );
  NAND U710 ( .A(n544), .B(n543), .Z(n2614) );
  NANDN U711 ( .A(x[502]), .B(y[502]), .Z(n546) );
  NANDN U712 ( .A(x[503]), .B(y[503]), .Z(n545) );
  NAND U713 ( .A(n546), .B(n545), .Z(n2611) );
  NANDN U714 ( .A(y[503]), .B(x[503]), .Z(n548) );
  NANDN U715 ( .A(y[504]), .B(x[504]), .Z(n547) );
  NAND U716 ( .A(n548), .B(n547), .Z(n2613) );
  NOR U717 ( .A(n2611), .B(n2613), .Z(n551) );
  NANDN U718 ( .A(x[508]), .B(y[508]), .Z(n550) );
  NANDN U719 ( .A(x[509]), .B(y[509]), .Z(n549) );
  NAND U720 ( .A(n550), .B(n549), .Z(n2625) );
  ANDN U721 ( .B(n551), .A(n2625), .Z(n552) );
  NANDN U722 ( .A(n2614), .B(n552), .Z(n553) );
  NOR U723 ( .A(n554), .B(n553), .Z(n566) );
  NANDN U724 ( .A(x[312]), .B(y[312]), .Z(n556) );
  NANDN U725 ( .A(x[313]), .B(y[313]), .Z(n555) );
  NAND U726 ( .A(n556), .B(n555), .Z(n2222) );
  NANDN U727 ( .A(x[420]), .B(y[420]), .Z(n558) );
  NANDN U728 ( .A(x[421]), .B(y[421]), .Z(n557) );
  NAND U729 ( .A(n558), .B(n557), .Z(n2450) );
  NANDN U730 ( .A(x[402]), .B(y[402]), .Z(n560) );
  NANDN U731 ( .A(x[403]), .B(y[403]), .Z(n559) );
  NAND U732 ( .A(n560), .B(n559), .Z(n2414) );
  NOR U733 ( .A(n2450), .B(n2414), .Z(n563) );
  NANDN U734 ( .A(y[225]), .B(x[225]), .Z(n562) );
  NANDN U735 ( .A(y[226]), .B(x[226]), .Z(n561) );
  NAND U736 ( .A(n562), .B(n561), .Z(n2065) );
  ANDN U737 ( .B(n563), .A(n2065), .Z(n564) );
  NANDN U738 ( .A(n2222), .B(n564), .Z(n565) );
  ANDN U739 ( .B(n566), .A(n565), .Z(n567) );
  NANDN U740 ( .A(n568), .B(n567), .Z(n616) );
  NANDN U741 ( .A(y[497]), .B(x[497]), .Z(n570) );
  NANDN U742 ( .A(y[498]), .B(x[498]), .Z(n569) );
  NAND U743 ( .A(n570), .B(n569), .Z(n2601) );
  NANDN U744 ( .A(x[496]), .B(y[496]), .Z(n572) );
  NANDN U745 ( .A(x[497]), .B(y[497]), .Z(n571) );
  NAND U746 ( .A(n572), .B(n571), .Z(n2599) );
  NANDN U747 ( .A(y[501]), .B(x[501]), .Z(n574) );
  NANDN U748 ( .A(y[502]), .B(x[502]), .Z(n573) );
  NAND U749 ( .A(n574), .B(n573), .Z(n2609) );
  NOR U750 ( .A(n2599), .B(n2609), .Z(n577) );
  NANDN U751 ( .A(x[500]), .B(y[500]), .Z(n576) );
  NANDN U752 ( .A(x[501]), .B(y[501]), .Z(n575) );
  NAND U753 ( .A(n576), .B(n575), .Z(n2607) );
  ANDN U754 ( .B(n577), .A(n2607), .Z(n578) );
  NANDN U755 ( .A(n2601), .B(n578), .Z(n614) );
  NANDN U756 ( .A(x[482]), .B(y[482]), .Z(n580) );
  NANDN U757 ( .A(x[483]), .B(y[483]), .Z(n579) );
  NAND U758 ( .A(n580), .B(n579), .Z(n2568) );
  NANDN U759 ( .A(y[483]), .B(x[483]), .Z(n582) );
  NANDN U760 ( .A(y[484]), .B(x[484]), .Z(n581) );
  NAND U761 ( .A(n582), .B(n581), .Z(n2571) );
  NANDN U762 ( .A(y[481]), .B(x[481]), .Z(n584) );
  NANDN U763 ( .A(y[482]), .B(x[482]), .Z(n583) );
  NAND U764 ( .A(n584), .B(n583), .Z(n2567) );
  NOR U765 ( .A(n2571), .B(n2567), .Z(n587) );
  NANDN U766 ( .A(y[487]), .B(x[487]), .Z(n586) );
  NANDN U767 ( .A(y[488]), .B(x[488]), .Z(n585) );
  NAND U768 ( .A(n586), .B(n585), .Z(n2579) );
  ANDN U769 ( .B(n587), .A(n2579), .Z(n588) );
  NANDN U770 ( .A(n2568), .B(n588), .Z(n600) );
  NANDN U771 ( .A(y[475]), .B(x[475]), .Z(n590) );
  NANDN U772 ( .A(y[476]), .B(x[476]), .Z(n589) );
  NAND U773 ( .A(n590), .B(n589), .Z(n2558) );
  NANDN U774 ( .A(x[466]), .B(y[466]), .Z(n592) );
  NANDN U775 ( .A(x[467]), .B(y[467]), .Z(n591) );
  NAND U776 ( .A(n592), .B(n591), .Z(n2549) );
  NANDN U777 ( .A(y[469]), .B(x[469]), .Z(n594) );
  NANDN U778 ( .A(y[470]), .B(x[470]), .Z(n593) );
  NAND U779 ( .A(n594), .B(n593), .Z(n2552) );
  NOR U780 ( .A(n2549), .B(n2552), .Z(n597) );
  NANDN U781 ( .A(y[477]), .B(x[477]), .Z(n596) );
  NANDN U782 ( .A(y[478]), .B(x[478]), .Z(n595) );
  NAND U783 ( .A(n596), .B(n595), .Z(n2560) );
  ANDN U784 ( .B(n597), .A(n2560), .Z(n598) );
  NANDN U785 ( .A(n2558), .B(n598), .Z(n599) );
  NOR U786 ( .A(n600), .B(n599), .Z(n612) );
  NANDN U787 ( .A(x[494]), .B(y[494]), .Z(n602) );
  NANDN U788 ( .A(x[495]), .B(y[495]), .Z(n601) );
  NAND U789 ( .A(n602), .B(n601), .Z(n2595) );
  NANDN U790 ( .A(y[489]), .B(x[489]), .Z(n604) );
  NANDN U791 ( .A(y[490]), .B(x[490]), .Z(n603) );
  NAND U792 ( .A(n604), .B(n603), .Z(n2583) );
  NANDN U793 ( .A(x[490]), .B(y[490]), .Z(n606) );
  NANDN U794 ( .A(x[491]), .B(y[491]), .Z(n605) );
  NAND U795 ( .A(n606), .B(n605), .Z(n2584) );
  NOR U796 ( .A(n2583), .B(n2584), .Z(n609) );
  NANDN U797 ( .A(y[495]), .B(x[495]), .Z(n608) );
  NANDN U798 ( .A(y[496]), .B(x[496]), .Z(n607) );
  NAND U799 ( .A(n608), .B(n607), .Z(n2597) );
  ANDN U800 ( .B(n609), .A(n2597), .Z(n610) );
  NANDN U801 ( .A(n2595), .B(n610), .Z(n611) );
  ANDN U802 ( .B(n612), .A(n611), .Z(n613) );
  NANDN U803 ( .A(n614), .B(n613), .Z(n615) );
  NOR U804 ( .A(n616), .B(n615), .Z(n664) );
  NANDN U805 ( .A(y[47]), .B(x[47]), .Z(n618) );
  NANDN U806 ( .A(y[48]), .B(x[48]), .Z(n617) );
  NAND U807 ( .A(n618), .B(n617), .Z(n1702) );
  NANDN U808 ( .A(x[46]), .B(y[46]), .Z(n620) );
  NANDN U809 ( .A(x[47]), .B(y[47]), .Z(n619) );
  NAND U810 ( .A(n620), .B(n619), .Z(n1700) );
  NANDN U811 ( .A(y[49]), .B(x[49]), .Z(n622) );
  NANDN U812 ( .A(y[50]), .B(x[50]), .Z(n621) );
  NAND U813 ( .A(n622), .B(n621), .Z(n1706) );
  NOR U814 ( .A(n1700), .B(n1706), .Z(n625) );
  NANDN U815 ( .A(x[48]), .B(y[48]), .Z(n624) );
  NANDN U816 ( .A(x[49]), .B(y[49]), .Z(n623) );
  NAND U817 ( .A(n624), .B(n623), .Z(n1704) );
  ANDN U818 ( .B(n625), .A(n1704), .Z(n626) );
  NANDN U819 ( .A(n1702), .B(n626), .Z(n662) );
  NANDN U820 ( .A(x[34]), .B(y[34]), .Z(n628) );
  NANDN U821 ( .A(x[35]), .B(y[35]), .Z(n627) );
  NAND U822 ( .A(n628), .B(n627), .Z(n1676) );
  NANDN U823 ( .A(y[35]), .B(x[35]), .Z(n630) );
  NANDN U824 ( .A(y[36]), .B(x[36]), .Z(n629) );
  NAND U825 ( .A(n630), .B(n629), .Z(n1678) );
  NANDN U826 ( .A(x[32]), .B(y[32]), .Z(n632) );
  NANDN U827 ( .A(x[33]), .B(y[33]), .Z(n631) );
  NAND U828 ( .A(n632), .B(n631), .Z(n1672) );
  NOR U829 ( .A(n1678), .B(n1672), .Z(n635) );
  NANDN U830 ( .A(y[37]), .B(x[37]), .Z(n634) );
  NANDN U831 ( .A(y[38]), .B(x[38]), .Z(n633) );
  NAND U832 ( .A(n634), .B(n633), .Z(n1682) );
  ANDN U833 ( .B(n635), .A(n1682), .Z(n636) );
  NANDN U834 ( .A(n1676), .B(n636), .Z(n648) );
  NANDN U835 ( .A(y[27]), .B(x[27]), .Z(n638) );
  NANDN U836 ( .A(y[28]), .B(x[28]), .Z(n637) );
  NAND U837 ( .A(n638), .B(n637), .Z(n1662) );
  NANDN U838 ( .A(x[26]), .B(y[26]), .Z(n640) );
  NANDN U839 ( .A(x[27]), .B(y[27]), .Z(n639) );
  NAND U840 ( .A(n640), .B(n639), .Z(n1660) );
  NANDN U841 ( .A(y[25]), .B(x[25]), .Z(n642) );
  NANDN U842 ( .A(y[26]), .B(x[26]), .Z(n641) );
  NAND U843 ( .A(n642), .B(n641), .Z(n1658) );
  NOR U844 ( .A(n1660), .B(n1658), .Z(n645) );
  NANDN U845 ( .A(y[29]), .B(x[29]), .Z(n644) );
  NANDN U846 ( .A(y[30]), .B(x[30]), .Z(n643) );
  NAND U847 ( .A(n644), .B(n643), .Z(n1666) );
  ANDN U848 ( .B(n645), .A(n1666), .Z(n646) );
  NANDN U849 ( .A(n1662), .B(n646), .Z(n647) );
  NOR U850 ( .A(n648), .B(n647), .Z(n660) );
  NANDN U851 ( .A(x[40]), .B(y[40]), .Z(n650) );
  NANDN U852 ( .A(x[41]), .B(y[41]), .Z(n649) );
  NAND U853 ( .A(n650), .B(n649), .Z(n1688) );
  NANDN U854 ( .A(x[38]), .B(y[38]), .Z(n652) );
  NANDN U855 ( .A(x[39]), .B(y[39]), .Z(n651) );
  NAND U856 ( .A(n652), .B(n651), .Z(n1684) );
  NANDN U857 ( .A(y[39]), .B(x[39]), .Z(n654) );
  NANDN U858 ( .A(y[40]), .B(x[40]), .Z(n653) );
  NAND U859 ( .A(n654), .B(n653), .Z(n1686) );
  NOR U860 ( .A(n1684), .B(n1686), .Z(n657) );
  NANDN U861 ( .A(y[45]), .B(x[45]), .Z(n656) );
  NANDN U862 ( .A(y[46]), .B(x[46]), .Z(n655) );
  NAND U863 ( .A(n656), .B(n655), .Z(n1698) );
  ANDN U864 ( .B(n657), .A(n1698), .Z(n658) );
  NANDN U865 ( .A(n1688), .B(n658), .Z(n659) );
  ANDN U866 ( .B(n660), .A(n659), .Z(n661) );
  NANDN U867 ( .A(n662), .B(n661), .Z(n663) );
  ANDN U868 ( .B(n664), .A(n663), .Z(n665) );
  NANDN U869 ( .A(n666), .B(n665), .Z(n667) );
  NOR U870 ( .A(n668), .B(n667), .Z(n1391) );
  NANDN U871 ( .A(x[485]), .B(y[485]), .Z(n1585) );
  ANDN U872 ( .B(x[510]), .A(y[510]), .Z(n2629) );
  ANDN U873 ( .B(x[493]), .A(y[493]), .Z(n2593) );
  NOR U874 ( .A(n2629), .B(n2593), .Z(n669) );
  AND U875 ( .A(n1585), .B(n669), .Z(n670) );
  NANDN U876 ( .A(x[481]), .B(y[481]), .Z(n2564) );
  NAND U877 ( .A(n670), .B(n2564), .Z(n687) );
  NANDN U878 ( .A(y[507]), .B(x[507]), .Z(n672) );
  NANDN U879 ( .A(y[508]), .B(x[508]), .Z(n671) );
  NAND U880 ( .A(n672), .B(n671), .Z(n2623) );
  NANDN U881 ( .A(x[492]), .B(y[492]), .Z(n674) );
  NANDN U882 ( .A(x[493]), .B(y[493]), .Z(n673) );
  NAND U883 ( .A(n674), .B(n673), .Z(n2589) );
  NOR U884 ( .A(n2623), .B(n2589), .Z(n685) );
  ANDN U885 ( .B(x[505]), .A(y[505]), .Z(n2616) );
  ANDN U886 ( .B(x[385]), .A(y[385]), .Z(n676) );
  IV U887 ( .A(y[436]), .Z(n2482) );
  NOR U888 ( .A(n2482), .B(x[436]), .Z(n675) );
  NOR U889 ( .A(n676), .B(n675), .Z(n678) );
  XNOR U890 ( .A(x[468]), .B(y[468]), .Z(n677) );
  NAND U891 ( .A(n678), .B(n677), .Z(n681) );
  NANDN U892 ( .A(x[506]), .B(y[506]), .Z(n680) );
  NANDN U893 ( .A(x[507]), .B(y[507]), .Z(n679) );
  NAND U894 ( .A(n680), .B(n679), .Z(n2620) );
  NOR U895 ( .A(n681), .B(n2620), .Z(n682) );
  ANDN U896 ( .B(x[511]), .A(y[511]), .Z(n2633) );
  ANDN U897 ( .B(n682), .A(n2633), .Z(n683) );
  NANDN U898 ( .A(n2616), .B(n683), .Z(n684) );
  ANDN U899 ( .B(n685), .A(n684), .Z(n686) );
  NANDN U900 ( .A(n687), .B(n686), .Z(n759) );
  NANDN U901 ( .A(y[451]), .B(x[451]), .Z(n689) );
  NANDN U902 ( .A(y[452]), .B(x[452]), .Z(n688) );
  NAND U903 ( .A(n689), .B(n688), .Z(n2517) );
  NANDN U904 ( .A(y[447]), .B(x[447]), .Z(n691) );
  NANDN U905 ( .A(y[448]), .B(x[448]), .Z(n690) );
  NAND U906 ( .A(n691), .B(n690), .Z(n2509) );
  NANDN U907 ( .A(y[449]), .B(x[449]), .Z(n693) );
  NANDN U908 ( .A(y[450]), .B(x[450]), .Z(n692) );
  NAND U909 ( .A(n693), .B(n692), .Z(n2513) );
  NOR U910 ( .A(n2509), .B(n2513), .Z(n696) );
  NANDN U911 ( .A(y[455]), .B(x[455]), .Z(n695) );
  NANDN U912 ( .A(y[456]), .B(x[456]), .Z(n694) );
  NAND U913 ( .A(n695), .B(n694), .Z(n2525) );
  ANDN U914 ( .B(n696), .A(n2525), .Z(n697) );
  NANDN U915 ( .A(n2517), .B(n697), .Z(n709) );
  NANDN U916 ( .A(y[437]), .B(x[437]), .Z(n699) );
  NANDN U917 ( .A(y[438]), .B(x[438]), .Z(n698) );
  NAND U918 ( .A(n699), .B(n698), .Z(n2489) );
  NANDN U919 ( .A(y[433]), .B(x[433]), .Z(n701) );
  NANDN U920 ( .A(y[434]), .B(x[434]), .Z(n700) );
  NAND U921 ( .A(n701), .B(n700), .Z(n2476) );
  NANDN U922 ( .A(y[445]), .B(x[445]), .Z(n703) );
  NANDN U923 ( .A(y[446]), .B(x[446]), .Z(n702) );
  NAND U924 ( .A(n703), .B(n702), .Z(n2505) );
  NOR U925 ( .A(n2476), .B(n2505), .Z(n706) );
  NANDN U926 ( .A(y[443]), .B(x[443]), .Z(n705) );
  NANDN U927 ( .A(y[444]), .B(x[444]), .Z(n704) );
  NAND U928 ( .A(n705), .B(n704), .Z(n2501) );
  ANDN U929 ( .B(n706), .A(n2501), .Z(n707) );
  NANDN U930 ( .A(n2489), .B(n707), .Z(n708) );
  NOR U931 ( .A(n709), .B(n708), .Z(n757) );
  NANDN U932 ( .A(x[488]), .B(y[488]), .Z(n711) );
  NANDN U933 ( .A(x[489]), .B(y[489]), .Z(n710) );
  NAND U934 ( .A(n711), .B(n710), .Z(n2581) );
  NANDN U935 ( .A(y[479]), .B(x[479]), .Z(n713) );
  NANDN U936 ( .A(y[480]), .B(x[480]), .Z(n712) );
  NAND U937 ( .A(n713), .B(n712), .Z(n2562) );
  NANDN U938 ( .A(y[485]), .B(x[485]), .Z(n715) );
  NANDN U939 ( .A(y[486]), .B(x[486]), .Z(n714) );
  NAND U940 ( .A(n715), .B(n714), .Z(n2575) );
  NOR U941 ( .A(n2562), .B(n2575), .Z(n718) );
  NANDN U942 ( .A(y[491]), .B(x[491]), .Z(n717) );
  NANDN U943 ( .A(y[492]), .B(x[492]), .Z(n716) );
  NAND U944 ( .A(n717), .B(n716), .Z(n2587) );
  ANDN U945 ( .B(n718), .A(n2587), .Z(n719) );
  NANDN U946 ( .A(n2581), .B(n719), .Z(n755) );
  NANDN U947 ( .A(y[471]), .B(x[471]), .Z(n721) );
  NANDN U948 ( .A(y[472]), .B(x[472]), .Z(n720) );
  NAND U949 ( .A(n721), .B(n720), .Z(n2554) );
  NANDN U950 ( .A(x[462]), .B(y[462]), .Z(n723) );
  NANDN U951 ( .A(x[463]), .B(y[463]), .Z(n722) );
  NAND U952 ( .A(n723), .B(n722), .Z(n2540) );
  NANDN U953 ( .A(x[470]), .B(y[470]), .Z(n725) );
  NANDN U954 ( .A(x[471]), .B(y[471]), .Z(n724) );
  NAND U955 ( .A(n725), .B(n724), .Z(n2553) );
  NOR U956 ( .A(n2540), .B(n2553), .Z(n728) );
  NANDN U957 ( .A(y[473]), .B(x[473]), .Z(n727) );
  NANDN U958 ( .A(y[474]), .B(x[474]), .Z(n726) );
  NAND U959 ( .A(n727), .B(n726), .Z(n2556) );
  ANDN U960 ( .B(n728), .A(n2556), .Z(n729) );
  NANDN U961 ( .A(n2554), .B(n729), .Z(n741) );
  NANDN U962 ( .A(y[463]), .B(x[463]), .Z(n731) );
  NANDN U963 ( .A(y[464]), .B(x[464]), .Z(n730) );
  NAND U964 ( .A(n731), .B(n730), .Z(n2543) );
  NANDN U965 ( .A(y[457]), .B(x[457]), .Z(n733) );
  NANDN U966 ( .A(y[458]), .B(x[458]), .Z(n732) );
  NAND U967 ( .A(n733), .B(n732), .Z(n2529) );
  NANDN U968 ( .A(y[459]), .B(x[459]), .Z(n735) );
  NANDN U969 ( .A(y[460]), .B(x[460]), .Z(n734) );
  NAND U970 ( .A(n735), .B(n734), .Z(n2533) );
  NOR U971 ( .A(n2529), .B(n2533), .Z(n738) );
  NANDN U972 ( .A(x[460]), .B(y[460]), .Z(n737) );
  NANDN U973 ( .A(x[461]), .B(y[461]), .Z(n736) );
  NAND U974 ( .A(n737), .B(n736), .Z(n2534) );
  ANDN U975 ( .B(n738), .A(n2534), .Z(n739) );
  NANDN U976 ( .A(n2543), .B(n739), .Z(n740) );
  NOR U977 ( .A(n741), .B(n740), .Z(n753) );
  NANDN U978 ( .A(x[478]), .B(y[478]), .Z(n743) );
  NANDN U979 ( .A(x[479]), .B(y[479]), .Z(n742) );
  NAND U980 ( .A(n743), .B(n742), .Z(n2561) );
  NANDN U981 ( .A(x[474]), .B(y[474]), .Z(n745) );
  NANDN U982 ( .A(x[475]), .B(y[475]), .Z(n744) );
  NAND U983 ( .A(n745), .B(n744), .Z(n2557) );
  NANDN U984 ( .A(x[476]), .B(y[476]), .Z(n747) );
  NANDN U985 ( .A(x[477]), .B(y[477]), .Z(n746) );
  NAND U986 ( .A(n747), .B(n746), .Z(n2559) );
  NOR U987 ( .A(n2557), .B(n2559), .Z(n750) );
  NANDN U988 ( .A(x[486]), .B(y[486]), .Z(n749) );
  NANDN U989 ( .A(x[487]), .B(y[487]), .Z(n748) );
  NAND U990 ( .A(n749), .B(n748), .Z(n2577) );
  ANDN U991 ( .B(n750), .A(n2577), .Z(n751) );
  NANDN U992 ( .A(n2561), .B(n751), .Z(n752) );
  ANDN U993 ( .B(n753), .A(n752), .Z(n754) );
  NANDN U994 ( .A(n755), .B(n754), .Z(n756) );
  ANDN U995 ( .B(n757), .A(n756), .Z(n758) );
  NANDN U996 ( .A(n759), .B(n758), .Z(n1389) );
  NANDN U997 ( .A(y[362]), .B(x[362]), .Z(n761) );
  NANDN U998 ( .A(y[363]), .B(x[363]), .Z(n760) );
  NAND U999 ( .A(n761), .B(n760), .Z(n2327) );
  NANDN U1000 ( .A(y[358]), .B(x[358]), .Z(n763) );
  NANDN U1001 ( .A(y[359]), .B(x[359]), .Z(n762) );
  NAND U1002 ( .A(n763), .B(n762), .Z(n2319) );
  NANDN U1003 ( .A(x[359]), .B(y[359]), .Z(n765) );
  NANDN U1004 ( .A(x[360]), .B(y[360]), .Z(n764) );
  NAND U1005 ( .A(n765), .B(n764), .Z(n2321) );
  NOR U1006 ( .A(n2319), .B(n2321), .Z(n768) );
  NANDN U1007 ( .A(x[363]), .B(y[363]), .Z(n767) );
  NANDN U1008 ( .A(x[364]), .B(y[364]), .Z(n766) );
  NAND U1009 ( .A(n767), .B(n766), .Z(n2328) );
  ANDN U1010 ( .B(n768), .A(n2328), .Z(n769) );
  NANDN U1011 ( .A(n2327), .B(n769), .Z(n805) );
  NANDN U1012 ( .A(y[352]), .B(x[352]), .Z(n771) );
  NANDN U1013 ( .A(y[353]), .B(x[353]), .Z(n770) );
  NAND U1014 ( .A(n771), .B(n770), .Z(n2312) );
  NANDN U1015 ( .A(x[336]), .B(y[336]), .Z(n773) );
  NANDN U1016 ( .A(x[337]), .B(y[337]), .Z(n772) );
  NAND U1017 ( .A(n773), .B(n772), .Z(n2280) );
  NANDN U1018 ( .A(y[343]), .B(x[343]), .Z(n775) );
  NANDN U1019 ( .A(y[344]), .B(x[344]), .Z(n774) );
  NAND U1020 ( .A(n775), .B(n774), .Z(n2301) );
  NOR U1021 ( .A(n2280), .B(n2301), .Z(n778) );
  NANDN U1022 ( .A(y[347]), .B(x[347]), .Z(n777) );
  NANDN U1023 ( .A(y[348]), .B(x[348]), .Z(n776) );
  NAND U1024 ( .A(n777), .B(n776), .Z(n2307) );
  ANDN U1025 ( .B(n778), .A(n2307), .Z(n779) );
  NANDN U1026 ( .A(n2312), .B(n779), .Z(n791) );
  NANDN U1027 ( .A(x[322]), .B(y[322]), .Z(n781) );
  NANDN U1028 ( .A(x[323]), .B(y[323]), .Z(n780) );
  NAND U1029 ( .A(n781), .B(n780), .Z(n2243) );
  NANDN U1030 ( .A(y[321]), .B(x[321]), .Z(n783) );
  NANDN U1031 ( .A(y[322]), .B(x[322]), .Z(n782) );
  NAND U1032 ( .A(n783), .B(n782), .Z(n2241) );
  NANDN U1033 ( .A(y[333]), .B(x[333]), .Z(n785) );
  NANDN U1034 ( .A(y[334]), .B(x[334]), .Z(n784) );
  NAND U1035 ( .A(n785), .B(n784), .Z(n2273) );
  NOR U1036 ( .A(n2241), .B(n2273), .Z(n788) );
  NANDN U1037 ( .A(y[324]), .B(x[324]), .Z(n787) );
  NANDN U1038 ( .A(y[325]), .B(x[325]), .Z(n786) );
  NAND U1039 ( .A(n787), .B(n786), .Z(n2249) );
  ANDN U1040 ( .B(n788), .A(n2249), .Z(n789) );
  NANDN U1041 ( .A(n2243), .B(n789), .Z(n790) );
  NOR U1042 ( .A(n791), .B(n790), .Z(n803) );
  NANDN U1043 ( .A(y[356]), .B(x[356]), .Z(n793) );
  NANDN U1044 ( .A(y[357]), .B(x[357]), .Z(n792) );
  NAND U1045 ( .A(n793), .B(n792), .Z(n2316) );
  NANDN U1046 ( .A(y[350]), .B(x[350]), .Z(n795) );
  NANDN U1047 ( .A(y[351]), .B(x[351]), .Z(n794) );
  NAND U1048 ( .A(n795), .B(n794), .Z(n2311) );
  NANDN U1049 ( .A(y[354]), .B(x[354]), .Z(n797) );
  NANDN U1050 ( .A(y[355]), .B(x[355]), .Z(n796) );
  NAND U1051 ( .A(n797), .B(n796), .Z(n2314) );
  NOR U1052 ( .A(n2311), .B(n2314), .Z(n800) );
  NANDN U1053 ( .A(y[360]), .B(x[360]), .Z(n799) );
  NANDN U1054 ( .A(y[361]), .B(x[361]), .Z(n798) );
  NAND U1055 ( .A(n799), .B(n798), .Z(n2323) );
  ANDN U1056 ( .B(n800), .A(n2323), .Z(n801) );
  NANDN U1057 ( .A(n2316), .B(n801), .Z(n802) );
  ANDN U1058 ( .B(n803), .A(n802), .Z(n804) );
  NANDN U1059 ( .A(n805), .B(n804), .Z(n949) );
  NANDN U1060 ( .A(y[265]), .B(x[265]), .Z(n807) );
  NANDN U1061 ( .A(y[266]), .B(x[266]), .Z(n806) );
  NAND U1062 ( .A(n807), .B(n806), .Z(n2125) );
  NANDN U1063 ( .A(x[244]), .B(y[244]), .Z(n809) );
  NANDN U1064 ( .A(x[245]), .B(y[245]), .Z(n808) );
  NAND U1065 ( .A(n809), .B(n808), .Z(n2096) );
  NANDN U1066 ( .A(x[250]), .B(y[250]), .Z(n811) );
  NANDN U1067 ( .A(x[251]), .B(y[251]), .Z(n810) );
  NAND U1068 ( .A(n811), .B(n810), .Z(n2106) );
  NOR U1069 ( .A(n2096), .B(n2106), .Z(n814) );
  NANDN U1070 ( .A(y[251]), .B(x[251]), .Z(n813) );
  NANDN U1071 ( .A(y[252]), .B(x[252]), .Z(n812) );
  NAND U1072 ( .A(n813), .B(n812), .Z(n2107) );
  ANDN U1073 ( .B(n814), .A(n2107), .Z(n815) );
  NANDN U1074 ( .A(n2125), .B(n815), .Z(n851) );
  NANDN U1075 ( .A(x[230]), .B(y[230]), .Z(n817) );
  NANDN U1076 ( .A(x[231]), .B(y[231]), .Z(n816) );
  NAND U1077 ( .A(n817), .B(n816), .Z(n2075) );
  NANDN U1078 ( .A(y[229]), .B(x[229]), .Z(n819) );
  NANDN U1079 ( .A(y[230]), .B(x[230]), .Z(n818) );
  NAND U1080 ( .A(n819), .B(n818), .Z(n2073) );
  NANDN U1081 ( .A(x[232]), .B(y[232]), .Z(n821) );
  NANDN U1082 ( .A(x[233]), .B(y[233]), .Z(n820) );
  NAND U1083 ( .A(n821), .B(n820), .Z(n2078) );
  NOR U1084 ( .A(n2073), .B(n2078), .Z(n824) );
  NANDN U1085 ( .A(y[231]), .B(x[231]), .Z(n823) );
  NANDN U1086 ( .A(y[232]), .B(x[232]), .Z(n822) );
  NAND U1087 ( .A(n823), .B(n822), .Z(n2077) );
  ANDN U1088 ( .B(n824), .A(n2077), .Z(n825) );
  NANDN U1089 ( .A(n2075), .B(n825), .Z(n837) );
  NANDN U1090 ( .A(y[223]), .B(x[223]), .Z(n827) );
  NANDN U1091 ( .A(y[224]), .B(x[224]), .Z(n826) );
  NAND U1092 ( .A(n827), .B(n826), .Z(n2061) );
  NANDN U1093 ( .A(x[224]), .B(y[224]), .Z(n829) );
  NANDN U1094 ( .A(x[225]), .B(y[225]), .Z(n828) );
  NAND U1095 ( .A(n829), .B(n828), .Z(n2063) );
  NANDN U1096 ( .A(x[222]), .B(y[222]), .Z(n831) );
  NANDN U1097 ( .A(x[223]), .B(y[223]), .Z(n830) );
  NAND U1098 ( .A(n831), .B(n830), .Z(n2059) );
  NOR U1099 ( .A(n2063), .B(n2059), .Z(n834) );
  NANDN U1100 ( .A(x[226]), .B(y[226]), .Z(n833) );
  NANDN U1101 ( .A(x[227]), .B(y[227]), .Z(n832) );
  NAND U1102 ( .A(n833), .B(n832), .Z(n2066) );
  ANDN U1103 ( .B(n834), .A(n2066), .Z(n835) );
  NANDN U1104 ( .A(n2061), .B(n835), .Z(n836) );
  NOR U1105 ( .A(n837), .B(n836), .Z(n849) );
  NANDN U1106 ( .A(x[242]), .B(y[242]), .Z(n839) );
  NANDN U1107 ( .A(x[243]), .B(y[243]), .Z(n838) );
  NAND U1108 ( .A(n839), .B(n838), .Z(n2094) );
  NANDN U1109 ( .A(y[233]), .B(x[233]), .Z(n841) );
  NANDN U1110 ( .A(y[234]), .B(x[234]), .Z(n840) );
  NAND U1111 ( .A(n841), .B(n840), .Z(n2081) );
  NANDN U1112 ( .A(y[235]), .B(x[235]), .Z(n843) );
  NANDN U1113 ( .A(y[236]), .B(x[236]), .Z(n842) );
  NAND U1114 ( .A(n843), .B(n842), .Z(n2085) );
  NOR U1115 ( .A(n2081), .B(n2085), .Z(n846) );
  NANDN U1116 ( .A(y[243]), .B(x[243]), .Z(n845) );
  NANDN U1117 ( .A(y[244]), .B(x[244]), .Z(n844) );
  NAND U1118 ( .A(n845), .B(n844), .Z(n2095) );
  ANDN U1119 ( .B(n846), .A(n2095), .Z(n847) );
  NANDN U1120 ( .A(n2094), .B(n847), .Z(n848) );
  ANDN U1121 ( .B(n849), .A(n848), .Z(n850) );
  NANDN U1122 ( .A(n851), .B(n850), .Z(n899) );
  NANDN U1123 ( .A(x[220]), .B(y[220]), .Z(n853) );
  NANDN U1124 ( .A(x[221]), .B(y[221]), .Z(n852) );
  NAND U1125 ( .A(n853), .B(n852), .Z(n2054) );
  NANDN U1126 ( .A(x[216]), .B(y[216]), .Z(n855) );
  NANDN U1127 ( .A(x[217]), .B(y[217]), .Z(n854) );
  NAND U1128 ( .A(n855), .B(n854), .Z(n2047) );
  NANDN U1129 ( .A(x[218]), .B(y[218]), .Z(n857) );
  NANDN U1130 ( .A(x[219]), .B(y[219]), .Z(n856) );
  NAND U1131 ( .A(n857), .B(n856), .Z(n2051) );
  NOR U1132 ( .A(n2047), .B(n2051), .Z(n860) );
  NANDN U1133 ( .A(y[221]), .B(x[221]), .Z(n859) );
  NANDN U1134 ( .A(y[222]), .B(x[222]), .Z(n858) );
  NAND U1135 ( .A(n859), .B(n858), .Z(n2057) );
  ANDN U1136 ( .B(n860), .A(n2057), .Z(n861) );
  NANDN U1137 ( .A(n2054), .B(n861), .Z(n897) );
  NANDN U1138 ( .A(x[210]), .B(y[210]), .Z(n863) );
  NANDN U1139 ( .A(x[211]), .B(y[211]), .Z(n862) );
  NAND U1140 ( .A(n863), .B(n862), .Z(n2035) );
  NANDN U1141 ( .A(x[200]), .B(y[200]), .Z(n865) );
  NANDN U1142 ( .A(x[201]), .B(y[201]), .Z(n864) );
  NAND U1143 ( .A(n865), .B(n864), .Z(n2014) );
  NANDN U1144 ( .A(y[209]), .B(x[209]), .Z(n867) );
  NANDN U1145 ( .A(y[210]), .B(x[210]), .Z(n866) );
  NAND U1146 ( .A(n867), .B(n866), .Z(n2033) );
  NOR U1147 ( .A(n2014), .B(n2033), .Z(n870) );
  NANDN U1148 ( .A(y[211]), .B(x[211]), .Z(n869) );
  NANDN U1149 ( .A(y[212]), .B(x[212]), .Z(n868) );
  NAND U1150 ( .A(n869), .B(n868), .Z(n2037) );
  ANDN U1151 ( .B(n870), .A(n2037), .Z(n871) );
  NANDN U1152 ( .A(n2035), .B(n871), .Z(n883) );
  NANDN U1153 ( .A(y[201]), .B(x[201]), .Z(n873) );
  NANDN U1154 ( .A(y[202]), .B(x[202]), .Z(n872) );
  NAND U1155 ( .A(n873), .B(n872), .Z(n2017) );
  NANDN U1156 ( .A(x[196]), .B(y[196]), .Z(n875) );
  NANDN U1157 ( .A(x[197]), .B(y[197]), .Z(n874) );
  NAND U1158 ( .A(n875), .B(n874), .Z(n2007) );
  NANDN U1159 ( .A(y[197]), .B(x[197]), .Z(n877) );
  NANDN U1160 ( .A(y[198]), .B(x[198]), .Z(n876) );
  NAND U1161 ( .A(n877), .B(n876), .Z(n2009) );
  NOR U1162 ( .A(n2007), .B(n2009), .Z(n880) );
  NANDN U1163 ( .A(y[199]), .B(x[199]), .Z(n879) );
  NANDN U1164 ( .A(y[200]), .B(x[200]), .Z(n878) );
  NAND U1165 ( .A(n879), .B(n878), .Z(n2013) );
  ANDN U1166 ( .B(n880), .A(n2013), .Z(n881) );
  NANDN U1167 ( .A(n2017), .B(n881), .Z(n882) );
  NOR U1168 ( .A(n883), .B(n882), .Z(n895) );
  NANDN U1169 ( .A(x[214]), .B(y[214]), .Z(n885) );
  NANDN U1170 ( .A(x[215]), .B(y[215]), .Z(n884) );
  NAND U1171 ( .A(n885), .B(n884), .Z(n2042) );
  NANDN U1172 ( .A(x[212]), .B(y[212]), .Z(n887) );
  NANDN U1173 ( .A(x[213]), .B(y[213]), .Z(n886) );
  NAND U1174 ( .A(n887), .B(n886), .Z(n2039) );
  NANDN U1175 ( .A(y[213]), .B(x[213]), .Z(n889) );
  NANDN U1176 ( .A(y[214]), .B(x[214]), .Z(n888) );
  NAND U1177 ( .A(n889), .B(n888), .Z(n2041) );
  NOR U1178 ( .A(n2039), .B(n2041), .Z(n892) );
  NANDN U1179 ( .A(y[219]), .B(x[219]), .Z(n891) );
  NANDN U1180 ( .A(y[220]), .B(x[220]), .Z(n890) );
  NAND U1181 ( .A(n891), .B(n890), .Z(n2053) );
  ANDN U1182 ( .B(n892), .A(n2053), .Z(n893) );
  NANDN U1183 ( .A(n2042), .B(n893), .Z(n894) );
  ANDN U1184 ( .B(n895), .A(n894), .Z(n896) );
  NANDN U1185 ( .A(n897), .B(n896), .Z(n898) );
  NOR U1186 ( .A(n899), .B(n898), .Z(n947) );
  NANDN U1187 ( .A(y[315]), .B(x[315]), .Z(n901) );
  NANDN U1188 ( .A(y[316]), .B(x[316]), .Z(n900) );
  NAND U1189 ( .A(n901), .B(n900), .Z(n2229) );
  NANDN U1190 ( .A(y[309]), .B(x[309]), .Z(n903) );
  NANDN U1191 ( .A(y[310]), .B(x[310]), .Z(n902) );
  NAND U1192 ( .A(n903), .B(n902), .Z(n2217) );
  NANDN U1193 ( .A(x[314]), .B(y[314]), .Z(n905) );
  NANDN U1194 ( .A(x[315]), .B(y[315]), .Z(n904) );
  NAND U1195 ( .A(n905), .B(n904), .Z(n2227) );
  NOR U1196 ( .A(n2217), .B(n2227), .Z(n908) );
  NANDN U1197 ( .A(x[318]), .B(y[318]), .Z(n907) );
  NANDN U1198 ( .A(x[319]), .B(y[319]), .Z(n906) );
  NAND U1199 ( .A(n907), .B(n906), .Z(n2234) );
  ANDN U1200 ( .B(n908), .A(n2234), .Z(n909) );
  NANDN U1201 ( .A(n2229), .B(n909), .Z(n945) );
  NANDN U1202 ( .A(x[292]), .B(y[292]), .Z(n911) );
  NANDN U1203 ( .A(x[293]), .B(y[293]), .Z(n910) );
  NAND U1204 ( .A(n911), .B(n910), .Z(n2183) );
  NANDN U1205 ( .A(y[273]), .B(x[273]), .Z(n913) );
  NANDN U1206 ( .A(y[274]), .B(x[274]), .Z(n912) );
  NAND U1207 ( .A(n913), .B(n912), .Z(n2141) );
  NANDN U1208 ( .A(x[278]), .B(y[278]), .Z(n915) );
  NANDN U1209 ( .A(x[279]), .B(y[279]), .Z(n914) );
  NAND U1210 ( .A(n915), .B(n914), .Z(n2150) );
  NOR U1211 ( .A(n2141), .B(n2150), .Z(n918) );
  NANDN U1212 ( .A(y[293]), .B(x[293]), .Z(n917) );
  NANDN U1213 ( .A(y[294]), .B(x[294]), .Z(n916) );
  NAND U1214 ( .A(n917), .B(n916), .Z(n2185) );
  ANDN U1215 ( .B(n918), .A(n2185), .Z(n919) );
  NANDN U1216 ( .A(n2183), .B(n919), .Z(n931) );
  NANDN U1217 ( .A(x[272]), .B(y[272]), .Z(n921) );
  NANDN U1218 ( .A(x[273]), .B(y[273]), .Z(n920) );
  NAND U1219 ( .A(n921), .B(n920), .Z(n2138) );
  NANDN U1220 ( .A(y[253]), .B(x[253]), .Z(n923) );
  NANDN U1221 ( .A(y[254]), .B(x[254]), .Z(n922) );
  NAND U1222 ( .A(n923), .B(n922), .Z(n2109) );
  NANDN U1223 ( .A(y[267]), .B(x[267]), .Z(n925) );
  NANDN U1224 ( .A(y[268]), .B(x[268]), .Z(n924) );
  NAND U1225 ( .A(n925), .B(n924), .Z(n2129) );
  NOR U1226 ( .A(n2109), .B(n2129), .Z(n928) );
  NANDN U1227 ( .A(y[279]), .B(x[279]), .Z(n927) );
  NANDN U1228 ( .A(y[280]), .B(x[280]), .Z(n926) );
  NAND U1229 ( .A(n927), .B(n926), .Z(n2153) );
  ANDN U1230 ( .B(n928), .A(n2153), .Z(n929) );
  NANDN U1231 ( .A(n2138), .B(n929), .Z(n930) );
  NOR U1232 ( .A(n931), .B(n930), .Z(n943) );
  NANDN U1233 ( .A(y[299]), .B(x[299]), .Z(n933) );
  NANDN U1234 ( .A(y[300]), .B(x[300]), .Z(n932) );
  NAND U1235 ( .A(n933), .B(n932), .Z(n2197) );
  NANDN U1236 ( .A(y[301]), .B(x[301]), .Z(n935) );
  NANDN U1237 ( .A(y[302]), .B(x[302]), .Z(n934) );
  NAND U1238 ( .A(n935), .B(n934), .Z(n2201) );
  NANDN U1239 ( .A(y[297]), .B(x[297]), .Z(n937) );
  NANDN U1240 ( .A(y[298]), .B(x[298]), .Z(n936) );
  NAND U1241 ( .A(n937), .B(n936), .Z(n2193) );
  NOR U1242 ( .A(n2201), .B(n2193), .Z(n940) );
  NANDN U1243 ( .A(y[307]), .B(x[307]), .Z(n939) );
  NANDN U1244 ( .A(y[308]), .B(x[308]), .Z(n938) );
  NAND U1245 ( .A(n939), .B(n938), .Z(n2213) );
  ANDN U1246 ( .B(n940), .A(n2213), .Z(n941) );
  NANDN U1247 ( .A(n2197), .B(n941), .Z(n942) );
  ANDN U1248 ( .B(n943), .A(n942), .Z(n944) );
  NANDN U1249 ( .A(n945), .B(n944), .Z(n946) );
  ANDN U1250 ( .B(n947), .A(n946), .Z(n948) );
  NANDN U1251 ( .A(n949), .B(n948), .Z(n1141) );
  NANDN U1252 ( .A(y[191]), .B(x[191]), .Z(n951) );
  NANDN U1253 ( .A(y[192]), .B(x[192]), .Z(n950) );
  NAND U1254 ( .A(n951), .B(n950), .Z(n2001) );
  NANDN U1255 ( .A(y[189]), .B(x[189]), .Z(n953) );
  NANDN U1256 ( .A(y[190]), .B(x[190]), .Z(n952) );
  NAND U1257 ( .A(n953), .B(n952), .Z(n1999) );
  NANDN U1258 ( .A(y[195]), .B(x[195]), .Z(n955) );
  NANDN U1259 ( .A(y[196]), .B(x[196]), .Z(n954) );
  NAND U1260 ( .A(n955), .B(n954), .Z(n2005) );
  NOR U1261 ( .A(n1999), .B(n2005), .Z(n958) );
  NANDN U1262 ( .A(y[193]), .B(x[193]), .Z(n957) );
  NANDN U1263 ( .A(y[194]), .B(x[194]), .Z(n956) );
  NAND U1264 ( .A(n957), .B(n956), .Z(n2003) );
  ANDN U1265 ( .B(n958), .A(n2003), .Z(n959) );
  NANDN U1266 ( .A(n2001), .B(n959), .Z(n995) );
  NANDN U1267 ( .A(y[179]), .B(x[179]), .Z(n961) );
  NANDN U1268 ( .A(y[180]), .B(x[180]), .Z(n960) );
  NAND U1269 ( .A(n961), .B(n960), .Z(n1987) );
  NANDN U1270 ( .A(y[177]), .B(x[177]), .Z(n963) );
  NANDN U1271 ( .A(y[178]), .B(x[178]), .Z(n962) );
  NAND U1272 ( .A(n963), .B(n962), .Z(n1983) );
  NANDN U1273 ( .A(x[178]), .B(y[178]), .Z(n965) );
  NANDN U1274 ( .A(x[179]), .B(y[179]), .Z(n964) );
  NAND U1275 ( .A(n965), .B(n964), .Z(n1984) );
  NOR U1276 ( .A(n1983), .B(n1984), .Z(n968) );
  NANDN U1277 ( .A(y[183]), .B(x[183]), .Z(n967) );
  NANDN U1278 ( .A(y[184]), .B(x[184]), .Z(n966) );
  NAND U1279 ( .A(n967), .B(n966), .Z(n1993) );
  ANDN U1280 ( .B(n968), .A(n1993), .Z(n969) );
  NANDN U1281 ( .A(n1987), .B(n969), .Z(n981) );
  NANDN U1282 ( .A(y[173]), .B(x[173]), .Z(n971) );
  NANDN U1283 ( .A(y[174]), .B(x[174]), .Z(n970) );
  NAND U1284 ( .A(n971), .B(n970), .Z(n1975) );
  NANDN U1285 ( .A(x[168]), .B(y[168]), .Z(n973) );
  NANDN U1286 ( .A(x[169]), .B(y[169]), .Z(n972) );
  NAND U1287 ( .A(n973), .B(n972), .Z(n1965) );
  NANDN U1288 ( .A(y[171]), .B(x[171]), .Z(n975) );
  NANDN U1289 ( .A(y[172]), .B(x[172]), .Z(n974) );
  NAND U1290 ( .A(n975), .B(n974), .Z(n1971) );
  NOR U1291 ( .A(n1965), .B(n1971), .Z(n978) );
  NANDN U1292 ( .A(y[175]), .B(x[175]), .Z(n977) );
  NANDN U1293 ( .A(y[176]), .B(x[176]), .Z(n976) );
  NAND U1294 ( .A(n977), .B(n976), .Z(n1979) );
  ANDN U1295 ( .B(n978), .A(n1979), .Z(n979) );
  NANDN U1296 ( .A(n1975), .B(n979), .Z(n980) );
  NOR U1297 ( .A(n981), .B(n980), .Z(n993) );
  NANDN U1298 ( .A(y[185]), .B(x[185]), .Z(n983) );
  NANDN U1299 ( .A(y[186]), .B(x[186]), .Z(n982) );
  NAND U1300 ( .A(n983), .B(n982), .Z(n1995) );
  NANDN U1301 ( .A(x[186]), .B(y[186]), .Z(n985) );
  NANDN U1302 ( .A(x[187]), .B(y[187]), .Z(n984) );
  NAND U1303 ( .A(n985), .B(n984), .Z(n1996) );
  NANDN U1304 ( .A(x[184]), .B(y[184]), .Z(n987) );
  NANDN U1305 ( .A(x[185]), .B(y[185]), .Z(n986) );
  NAND U1306 ( .A(n987), .B(n986), .Z(n1994) );
  NOR U1307 ( .A(n1996), .B(n1994), .Z(n990) );
  NANDN U1308 ( .A(x[188]), .B(y[188]), .Z(n989) );
  NANDN U1309 ( .A(x[189]), .B(y[189]), .Z(n988) );
  NAND U1310 ( .A(n989), .B(n988), .Z(n1998) );
  ANDN U1311 ( .B(n990), .A(n1998), .Z(n991) );
  NANDN U1312 ( .A(n1995), .B(n991), .Z(n992) );
  ANDN U1313 ( .B(n993), .A(n992), .Z(n994) );
  NANDN U1314 ( .A(n995), .B(n994), .Z(n1139) );
  NANDN U1315 ( .A(x[140]), .B(y[140]), .Z(n997) );
  NANDN U1316 ( .A(x[141]), .B(y[141]), .Z(n996) );
  NAND U1317 ( .A(n997), .B(n996), .Z(n1902) );
  NANDN U1318 ( .A(y[141]), .B(x[141]), .Z(n999) );
  NANDN U1319 ( .A(y[142]), .B(x[142]), .Z(n998) );
  NAND U1320 ( .A(n999), .B(n998), .Z(n1904) );
  NANDN U1321 ( .A(y[139]), .B(x[139]), .Z(n1001) );
  NANDN U1322 ( .A(y[140]), .B(x[140]), .Z(n1000) );
  NAND U1323 ( .A(n1001), .B(n1000), .Z(n1900) );
  NOR U1324 ( .A(n1904), .B(n1900), .Z(n1004) );
  NANDN U1325 ( .A(x[142]), .B(y[142]), .Z(n1003) );
  NANDN U1326 ( .A(x[143]), .B(y[143]), .Z(n1002) );
  NAND U1327 ( .A(n1003), .B(n1002), .Z(n1905) );
  ANDN U1328 ( .B(n1004), .A(n1905), .Z(n1005) );
  NANDN U1329 ( .A(n1902), .B(n1005), .Z(n1041) );
  NANDN U1330 ( .A(x[130]), .B(y[130]), .Z(n1007) );
  NANDN U1331 ( .A(x[131]), .B(y[131]), .Z(n1006) );
  NAND U1332 ( .A(n1007), .B(n1006), .Z(n1880) );
  NANDN U1333 ( .A(y[125]), .B(x[125]), .Z(n1009) );
  NANDN U1334 ( .A(y[126]), .B(x[126]), .Z(n1008) );
  NAND U1335 ( .A(n1009), .B(n1008), .Z(n1868) );
  NANDN U1336 ( .A(x[128]), .B(y[128]), .Z(n1011) );
  NANDN U1337 ( .A(x[129]), .B(y[129]), .Z(n1010) );
  NAND U1338 ( .A(n1011), .B(n1010), .Z(n1875) );
  NOR U1339 ( .A(n1868), .B(n1875), .Z(n1014) );
  NANDN U1340 ( .A(y[131]), .B(x[131]), .Z(n1013) );
  NANDN U1341 ( .A(y[132]), .B(x[132]), .Z(n1012) );
  NAND U1342 ( .A(n1013), .B(n1012), .Z(n1882) );
  ANDN U1343 ( .B(n1014), .A(n1882), .Z(n1015) );
  NANDN U1344 ( .A(n1880), .B(n1015), .Z(n1027) );
  NANDN U1345 ( .A(x[124]), .B(y[124]), .Z(n1017) );
  NANDN U1346 ( .A(x[125]), .B(y[125]), .Z(n1016) );
  NAND U1347 ( .A(n1017), .B(n1016), .Z(n1866) );
  NANDN U1348 ( .A(x[122]), .B(y[122]), .Z(n1019) );
  NANDN U1349 ( .A(x[123]), .B(y[123]), .Z(n1018) );
  NAND U1350 ( .A(n1019), .B(n1018), .Z(n1862) );
  NANDN U1351 ( .A(y[123]), .B(x[123]), .Z(n1021) );
  NANDN U1352 ( .A(y[124]), .B(x[124]), .Z(n1020) );
  NAND U1353 ( .A(n1021), .B(n1020), .Z(n1864) );
  NOR U1354 ( .A(n1862), .B(n1864), .Z(n1024) );
  NANDN U1355 ( .A(y[129]), .B(x[129]), .Z(n1023) );
  NANDN U1356 ( .A(y[130]), .B(x[130]), .Z(n1022) );
  NAND U1357 ( .A(n1023), .B(n1022), .Z(n1878) );
  ANDN U1358 ( .B(n1024), .A(n1878), .Z(n1025) );
  NANDN U1359 ( .A(n1866), .B(n1025), .Z(n1026) );
  NOR U1360 ( .A(n1027), .B(n1026), .Z(n1039) );
  NANDN U1361 ( .A(x[134]), .B(y[134]), .Z(n1029) );
  NANDN U1362 ( .A(x[135]), .B(y[135]), .Z(n1028) );
  NAND U1363 ( .A(n1029), .B(n1028), .Z(n1887) );
  NANDN U1364 ( .A(x[132]), .B(y[132]), .Z(n1031) );
  NANDN U1365 ( .A(x[133]), .B(y[133]), .Z(n1030) );
  NAND U1366 ( .A(n1031), .B(n1030), .Z(n1884) );
  NANDN U1367 ( .A(y[133]), .B(x[133]), .Z(n1033) );
  NANDN U1368 ( .A(y[134]), .B(x[134]), .Z(n1032) );
  NAND U1369 ( .A(n1033), .B(n1032), .Z(n1886) );
  NOR U1370 ( .A(n1884), .B(n1886), .Z(n1036) );
  NANDN U1371 ( .A(x[138]), .B(y[138]), .Z(n1035) );
  NANDN U1372 ( .A(x[139]), .B(y[139]), .Z(n1034) );
  NAND U1373 ( .A(n1035), .B(n1034), .Z(n1898) );
  ANDN U1374 ( .B(n1036), .A(n1898), .Z(n1037) );
  NANDN U1375 ( .A(n1887), .B(n1037), .Z(n1038) );
  ANDN U1376 ( .B(n1039), .A(n1038), .Z(n1040) );
  NANDN U1377 ( .A(n1041), .B(n1040), .Z(n1089) );
  NANDN U1378 ( .A(y[117]), .B(x[117]), .Z(n1043) );
  NANDN U1379 ( .A(y[118]), .B(x[118]), .Z(n1042) );
  NAND U1380 ( .A(n1043), .B(n1042), .Z(n1852) );
  NANDN U1381 ( .A(y[113]), .B(x[113]), .Z(n1045) );
  NANDN U1382 ( .A(y[114]), .B(x[114]), .Z(n1044) );
  NAND U1383 ( .A(n1045), .B(n1044), .Z(n1844) );
  NANDN U1384 ( .A(x[116]), .B(y[116]), .Z(n1047) );
  NANDN U1385 ( .A(x[117]), .B(y[117]), .Z(n1046) );
  NAND U1386 ( .A(n1047), .B(n1046), .Z(n1850) );
  NOR U1387 ( .A(n1844), .B(n1850), .Z(n1050) );
  NANDN U1388 ( .A(x[118]), .B(y[118]), .Z(n1049) );
  NANDN U1389 ( .A(x[119]), .B(y[119]), .Z(n1048) );
  NAND U1390 ( .A(n1049), .B(n1048), .Z(n1854) );
  ANDN U1391 ( .B(n1050), .A(n1854), .Z(n1051) );
  NANDN U1392 ( .A(n1852), .B(n1051), .Z(n1087) );
  NANDN U1393 ( .A(x[104]), .B(y[104]), .Z(n1053) );
  NANDN U1394 ( .A(x[105]), .B(y[105]), .Z(n1052) );
  NAND U1395 ( .A(n1053), .B(n1052), .Z(n1826) );
  NANDN U1396 ( .A(y[99]), .B(x[99]), .Z(n1055) );
  NANDN U1397 ( .A(y[100]), .B(x[100]), .Z(n1054) );
  NAND U1398 ( .A(n1055), .B(n1054), .Z(n1816) );
  NANDN U1399 ( .A(x[108]), .B(y[108]), .Z(n1057) );
  NANDN U1400 ( .A(x[109]), .B(y[109]), .Z(n1056) );
  NAND U1401 ( .A(n1057), .B(n1056), .Z(n1833) );
  NOR U1402 ( .A(n1816), .B(n1833), .Z(n1060) );
  NANDN U1403 ( .A(x[106]), .B(y[106]), .Z(n1059) );
  NANDN U1404 ( .A(x[107]), .B(y[107]), .Z(n1058) );
  NAND U1405 ( .A(n1059), .B(n1058), .Z(n1830) );
  ANDN U1406 ( .B(n1060), .A(n1830), .Z(n1061) );
  NANDN U1407 ( .A(n1826), .B(n1061), .Z(n1073) );
  NANDN U1408 ( .A(x[96]), .B(y[96]), .Z(n1063) );
  NANDN U1409 ( .A(x[97]), .B(y[97]), .Z(n1062) );
  NAND U1410 ( .A(n1063), .B(n1062), .Z(n1809) );
  NANDN U1411 ( .A(y[97]), .B(x[97]), .Z(n1065) );
  NANDN U1412 ( .A(y[98]), .B(x[98]), .Z(n1064) );
  NAND U1413 ( .A(n1065), .B(n1064), .Z(n1812) );
  NANDN U1414 ( .A(y[95]), .B(x[95]), .Z(n1067) );
  NANDN U1415 ( .A(y[96]), .B(x[96]), .Z(n1066) );
  NAND U1416 ( .A(n1067), .B(n1066), .Z(n1808) );
  NOR U1417 ( .A(n1812), .B(n1808), .Z(n1070) );
  NANDN U1418 ( .A(x[98]), .B(y[98]), .Z(n1069) );
  NANDN U1419 ( .A(x[99]), .B(y[99]), .Z(n1068) );
  NAND U1420 ( .A(n1069), .B(n1068), .Z(n1814) );
  ANDN U1421 ( .B(n1070), .A(n1814), .Z(n1071) );
  NANDN U1422 ( .A(n1809), .B(n1071), .Z(n1072) );
  NOR U1423 ( .A(n1073), .B(n1072), .Z(n1085) );
  NANDN U1424 ( .A(x[114]), .B(y[114]), .Z(n1075) );
  NANDN U1425 ( .A(x[115]), .B(y[115]), .Z(n1074) );
  NAND U1426 ( .A(n1075), .B(n1074), .Z(n1845) );
  NANDN U1427 ( .A(y[109]), .B(x[109]), .Z(n1077) );
  NANDN U1428 ( .A(y[110]), .B(x[110]), .Z(n1076) );
  NAND U1429 ( .A(n1077), .B(n1076), .Z(n1836) );
  NANDN U1430 ( .A(x[110]), .B(y[110]), .Z(n1079) );
  NANDN U1431 ( .A(x[111]), .B(y[111]), .Z(n1078) );
  NAND U1432 ( .A(n1079), .B(n1078), .Z(n1838) );
  NOR U1433 ( .A(n1836), .B(n1838), .Z(n1082) );
  NANDN U1434 ( .A(y[111]), .B(x[111]), .Z(n1081) );
  NANDN U1435 ( .A(y[112]), .B(x[112]), .Z(n1080) );
  NAND U1436 ( .A(n1081), .B(n1080), .Z(n1840) );
  ANDN U1437 ( .B(n1082), .A(n1840), .Z(n1083) );
  NANDN U1438 ( .A(n1845), .B(n1083), .Z(n1084) );
  ANDN U1439 ( .B(n1085), .A(n1084), .Z(n1086) );
  NANDN U1440 ( .A(n1087), .B(n1086), .Z(n1088) );
  NOR U1441 ( .A(n1089), .B(n1088), .Z(n1137) );
  NANDN U1442 ( .A(x[166]), .B(y[166]), .Z(n1091) );
  NANDN U1443 ( .A(x[167]), .B(y[167]), .Z(n1090) );
  NAND U1444 ( .A(n1091), .B(n1090), .Z(n1960) );
  NANDN U1445 ( .A(x[162]), .B(y[162]), .Z(n1093) );
  NANDN U1446 ( .A(x[163]), .B(y[163]), .Z(n1092) );
  NAND U1447 ( .A(n1093), .B(n1092), .Z(n1953) );
  NANDN U1448 ( .A(y[165]), .B(x[165]), .Z(n1095) );
  NANDN U1449 ( .A(y[166]), .B(x[166]), .Z(n1094) );
  NAND U1450 ( .A(n1095), .B(n1094), .Z(n1959) );
  NOR U1451 ( .A(n1953), .B(n1959), .Z(n1098) );
  NANDN U1452 ( .A(x[172]), .B(y[172]), .Z(n1097) );
  NANDN U1453 ( .A(x[173]), .B(y[173]), .Z(n1096) );
  NAND U1454 ( .A(n1097), .B(n1096), .Z(n1972) );
  ANDN U1455 ( .B(n1098), .A(n1972), .Z(n1099) );
  NANDN U1456 ( .A(n1960), .B(n1099), .Z(n1135) );
  NANDN U1457 ( .A(y[153]), .B(x[153]), .Z(n1101) );
  NANDN U1458 ( .A(y[154]), .B(x[154]), .Z(n1100) );
  NAND U1459 ( .A(n1101), .B(n1100), .Z(n1935) );
  NANDN U1460 ( .A(x[152]), .B(y[152]), .Z(n1103) );
  NANDN U1461 ( .A(x[153]), .B(y[153]), .Z(n1102) );
  NAND U1462 ( .A(n1103), .B(n1102), .Z(n1933) );
  NANDN U1463 ( .A(y[155]), .B(x[155]), .Z(n1105) );
  NANDN U1464 ( .A(y[156]), .B(x[156]), .Z(n1104) );
  NAND U1465 ( .A(n1105), .B(n1104), .Z(n1939) );
  NOR U1466 ( .A(n1933), .B(n1939), .Z(n1108) );
  NANDN U1467 ( .A(x[154]), .B(y[154]), .Z(n1107) );
  NANDN U1468 ( .A(x[155]), .B(y[155]), .Z(n1106) );
  NAND U1469 ( .A(n1107), .B(n1106), .Z(n1936) );
  ANDN U1470 ( .B(n1108), .A(n1936), .Z(n1109) );
  NANDN U1471 ( .A(n1935), .B(n1109), .Z(n1121) );
  NANDN U1472 ( .A(x[150]), .B(y[150]), .Z(n1111) );
  NANDN U1473 ( .A(x[151]), .B(y[151]), .Z(n1110) );
  NAND U1474 ( .A(n1111), .B(n1110), .Z(n1929) );
  NANDN U1475 ( .A(y[143]), .B(x[143]), .Z(n1113) );
  NANDN U1476 ( .A(y[144]), .B(x[144]), .Z(n1112) );
  NAND U1477 ( .A(n1113), .B(n1112), .Z(n1908) );
  NANDN U1478 ( .A(x[144]), .B(y[144]), .Z(n1115) );
  NANDN U1479 ( .A(x[145]), .B(y[145]), .Z(n1114) );
  NAND U1480 ( .A(n1115), .B(n1114), .Z(n1910) );
  NOR U1481 ( .A(n1908), .B(n1910), .Z(n1118) );
  NANDN U1482 ( .A(y[151]), .B(x[151]), .Z(n1117) );
  NANDN U1483 ( .A(y[152]), .B(x[152]), .Z(n1116) );
  NAND U1484 ( .A(n1117), .B(n1116), .Z(n1931) );
  ANDN U1485 ( .B(n1118), .A(n1931), .Z(n1119) );
  NANDN U1486 ( .A(n1929), .B(n1119), .Z(n1120) );
  NOR U1487 ( .A(n1121), .B(n1120), .Z(n1133) );
  NANDN U1488 ( .A(y[163]), .B(x[163]), .Z(n1123) );
  NANDN U1489 ( .A(y[164]), .B(x[164]), .Z(n1122) );
  NAND U1490 ( .A(n1123), .B(n1122), .Z(n1955) );
  NANDN U1491 ( .A(x[156]), .B(y[156]), .Z(n1125) );
  NANDN U1492 ( .A(x[157]), .B(y[157]), .Z(n1124) );
  NAND U1493 ( .A(n1125), .B(n1124), .Z(n1941) );
  NANDN U1494 ( .A(x[158]), .B(y[158]), .Z(n1127) );
  NANDN U1495 ( .A(x[159]), .B(y[159]), .Z(n1126) );
  NAND U1496 ( .A(n1127), .B(n1126), .Z(n1945) );
  NOR U1497 ( .A(n1941), .B(n1945), .Z(n1130) );
  NANDN U1498 ( .A(y[161]), .B(x[161]), .Z(n1129) );
  NANDN U1499 ( .A(y[162]), .B(x[162]), .Z(n1128) );
  NAND U1500 ( .A(n1129), .B(n1128), .Z(n1951) );
  ANDN U1501 ( .B(n1130), .A(n1951), .Z(n1131) );
  NANDN U1502 ( .A(n1955), .B(n1131), .Z(n1132) );
  ANDN U1503 ( .B(n1133), .A(n1132), .Z(n1134) );
  NANDN U1504 ( .A(n1135), .B(n1134), .Z(n1136) );
  ANDN U1505 ( .B(n1137), .A(n1136), .Z(n1138) );
  NANDN U1506 ( .A(n1139), .B(n1138), .Z(n1140) );
  NOR U1507 ( .A(n1141), .B(n1140), .Z(n1387) );
  ANDN U1508 ( .B(y[348]), .A(x[348]), .Z(n2308) );
  ANDN U1509 ( .B(y[350]), .A(x[350]), .Z(n2310) );
  NOR U1510 ( .A(n2308), .B(n2310), .Z(n1142) );
  NANDN U1511 ( .A(x[383]), .B(y[383]), .Z(n2368) );
  NAND U1512 ( .A(n1142), .B(n2368), .Z(n1145) );
  XNOR U1513 ( .A(x[346]), .B(y[346]), .Z(n1143) );
  NANDN U1514 ( .A(y[345]), .B(x[345]), .Z(n1589) );
  NAND U1515 ( .A(n1143), .B(n1589), .Z(n1144) );
  NOR U1516 ( .A(n1145), .B(n1144), .Z(n1146) );
  XNOR U1517 ( .A(x[349]), .B(y[349]), .Z(n2309) );
  NAND U1518 ( .A(n1146), .B(n2309), .Z(n1212) );
  ANDN U1519 ( .B(x[384]), .A(y[384]), .Z(n1151) );
  NANDN U1520 ( .A(x[351]), .B(y[351]), .Z(n1587) );
  ANDN U1521 ( .B(x[436]), .A(y[436]), .Z(n1148) );
  IV U1522 ( .A(y[385]), .Z(n2377) );
  NOR U1523 ( .A(n2377), .B(x[385]), .Z(n1147) );
  NOR U1524 ( .A(n1148), .B(n1147), .Z(n1149) );
  AND U1525 ( .A(n1587), .B(n1149), .Z(n1150) );
  NANDN U1526 ( .A(n1151), .B(n1150), .Z(n1155) );
  ANDN U1527 ( .B(x[342]), .A(y[342]), .Z(n2297) );
  NANDN U1528 ( .A(x[341]), .B(y[341]), .Z(n2295) );
  NANDN U1529 ( .A(x[347]), .B(y[347]), .Z(n2306) );
  ANDN U1530 ( .B(y[340]), .A(x[340]), .Z(n2291) );
  ANDN U1531 ( .B(n2306), .A(n2291), .Z(n1152) );
  AND U1532 ( .A(n2295), .B(n1152), .Z(n1153) );
  NANDN U1533 ( .A(n2297), .B(n1153), .Z(n1154) );
  NOR U1534 ( .A(n1155), .B(n1154), .Z(n1210) );
  NANDN U1535 ( .A(x[324]), .B(y[324]), .Z(n2247) );
  NANDN U1536 ( .A(x[288]), .B(y[288]), .Z(n1157) );
  NANDN U1537 ( .A(x[289]), .B(y[289]), .Z(n1156) );
  NAND U1538 ( .A(n1157), .B(n1156), .Z(n2173) );
  NANDN U1539 ( .A(x[326]), .B(y[326]), .Z(n1591) );
  NANDN U1540 ( .A(x[330]), .B(y[330]), .Z(n2263) );
  ANDN U1541 ( .B(x[328]), .A(y[328]), .Z(n2257) );
  ANDN U1542 ( .B(n2263), .A(n2257), .Z(n1158) );
  AND U1543 ( .A(n1591), .B(n1158), .Z(n1159) );
  NANDN U1544 ( .A(x[327]), .B(y[327]), .Z(n2254) );
  NAND U1545 ( .A(n1159), .B(n2254), .Z(n1160) );
  NOR U1546 ( .A(n2173), .B(n1160), .Z(n1161) );
  AND U1547 ( .A(n2247), .B(n1161), .Z(n1162) );
  NANDN U1548 ( .A(x[325]), .B(y[325]), .Z(n1592) );
  NAND U1549 ( .A(n1162), .B(n1592), .Z(n1208) );
  NANDN U1550 ( .A(x[338]), .B(y[338]), .Z(n2284) );
  ANDN U1551 ( .B(x[335]), .A(y[335]), .Z(n2277) );
  ANDN U1552 ( .B(n2284), .A(n2277), .Z(n1164) );
  XNOR U1553 ( .A(y[339]), .B(x[339]), .Z(n1163) );
  NAND U1554 ( .A(n1164), .B(n1163), .Z(n1168) );
  ANDN U1555 ( .B(x[329]), .A(y[329]), .Z(n2261) );
  NANDN U1556 ( .A(x[331]), .B(y[331]), .Z(n2266) );
  ANDN U1557 ( .B(x[332]), .A(y[332]), .Z(n2269) );
  ANDN U1558 ( .B(x[336]), .A(y[336]), .Z(n2276) );
  NOR U1559 ( .A(n2269), .B(n2276), .Z(n1165) );
  AND U1560 ( .A(n2266), .B(n1165), .Z(n1166) );
  NANDN U1561 ( .A(n2261), .B(n1166), .Z(n1167) );
  NOR U1562 ( .A(n1168), .B(n1167), .Z(n1206) );
  NANDN U1563 ( .A(x[183]), .B(y[183]), .Z(n1992) );
  ANDN U1564 ( .B(x[181]), .A(y[181]), .Z(n1990) );
  NANDN U1565 ( .A(x[236]), .B(y[236]), .Z(n2087) );
  ANDN U1566 ( .B(x[150]), .A(y[150]), .Z(n1927) );
  ANDN U1567 ( .B(n2087), .A(n1927), .Z(n1170) );
  IV U1568 ( .A(y[146]), .Z(n1914) );
  NOR U1569 ( .A(n1914), .B(x[146]), .Z(n1169) );
  ANDN U1570 ( .B(n1170), .A(n1169), .Z(n1171) );
  NANDN U1571 ( .A(n1990), .B(n1171), .Z(n1174) );
  NANDN U1572 ( .A(y[240]), .B(x[240]), .Z(n1173) );
  NANDN U1573 ( .A(y[239]), .B(x[239]), .Z(n1172) );
  NAND U1574 ( .A(n1173), .B(n1172), .Z(n2090) );
  NOR U1575 ( .A(n1174), .B(n2090), .Z(n1175) );
  AND U1576 ( .A(n1992), .B(n1175), .Z(n1176) );
  NANDN U1577 ( .A(x[241]), .B(y[241]), .Z(n2092) );
  NAND U1578 ( .A(n1176), .B(n2092), .Z(n1204) );
  ANDN U1579 ( .B(x[248]), .A(y[248]), .Z(n1179) );
  NANDN U1580 ( .A(x[249]), .B(y[249]), .Z(n2104) );
  NANDN U1581 ( .A(x[291]), .B(y[291]), .Z(n2178) );
  ANDN U1582 ( .B(y[282]), .A(x[282]), .Z(n2161) );
  ANDN U1583 ( .B(n2178), .A(n2161), .Z(n1177) );
  AND U1584 ( .A(n2104), .B(n1177), .Z(n1178) );
  NANDN U1585 ( .A(n1179), .B(n1178), .Z(n1183) );
  NANDN U1586 ( .A(x[246]), .B(y[246]), .Z(n2099) );
  ANDN U1587 ( .B(x[245]), .A(y[245]), .Z(n2098) );
  ANDN U1588 ( .B(n2099), .A(n2098), .Z(n1181) );
  XNOR U1589 ( .A(x[247]), .B(y[247]), .Z(n1180) );
  NAND U1590 ( .A(n1181), .B(n1180), .Z(n1182) );
  NOR U1591 ( .A(n1183), .B(n1182), .Z(n1202) );
  ANDN U1592 ( .B(x[146]), .A(y[146]), .Z(n1200) );
  NANDN U1593 ( .A(x[147]), .B(y[147]), .Z(n1919) );
  NANDN U1594 ( .A(x[263]), .B(y[263]), .Z(n1593) );
  ANDN U1595 ( .B(x[2]), .A(y[2]), .Z(n1605) );
  ANDN U1596 ( .B(n1593), .A(n1605), .Z(n1185) );
  NANDN U1597 ( .A(x[0]), .B(y[0]), .Z(n1184) );
  NAND U1598 ( .A(n1185), .B(n1184), .Z(n1194) );
  NANDN U1599 ( .A(x[7]), .B(y[7]), .Z(n1617) );
  NANDN U1600 ( .A(x[78]), .B(y[78]), .Z(n1768) );
  NANDN U1601 ( .A(x[88]), .B(y[88]), .Z(n1793) );
  ANDN U1602 ( .B(x[80]), .A(y[80]), .Z(n1774) );
  ANDN U1603 ( .B(n1793), .A(n1774), .Z(n1186) );
  AND U1604 ( .A(n1768), .B(n1186), .Z(n1187) );
  NANDN U1605 ( .A(x[79]), .B(y[79]), .Z(n1771) );
  NAND U1606 ( .A(n1187), .B(n1771), .Z(n1191) );
  ANDN U1607 ( .B(x[8]), .A(y[8]), .Z(n1620) );
  NANDN U1608 ( .A(x[21]), .B(y[21]), .Z(n1647) );
  ANDN U1609 ( .B(x[77]), .A(y[77]), .Z(n1766) );
  ANDN U1610 ( .B(x[75]), .A(y[75]), .Z(n1762) );
  NOR U1611 ( .A(n1766), .B(n1762), .Z(n1188) );
  AND U1612 ( .A(n1647), .B(n1188), .Z(n1189) );
  NANDN U1613 ( .A(n1620), .B(n1189), .Z(n1190) );
  NOR U1614 ( .A(n1191), .B(n1190), .Z(n1192) );
  AND U1615 ( .A(n1617), .B(n1192), .Z(n1193) );
  NANDN U1616 ( .A(n1194), .B(n1193), .Z(n1197) );
  NANDN U1617 ( .A(y[81]), .B(x[81]), .Z(n1196) );
  NANDN U1618 ( .A(y[82]), .B(x[82]), .Z(n1195) );
  NAND U1619 ( .A(n1196), .B(n1195), .Z(n1778) );
  NOR U1620 ( .A(n1197), .B(n1778), .Z(n1198) );
  AND U1621 ( .A(n1919), .B(n1198), .Z(n1199) );
  NANDN U1622 ( .A(n1200), .B(n1199), .Z(n1201) );
  ANDN U1623 ( .B(n1202), .A(n1201), .Z(n1203) );
  NANDN U1624 ( .A(n1204), .B(n1203), .Z(n1205) );
  ANDN U1625 ( .B(n1206), .A(n1205), .Z(n1207) );
  NANDN U1626 ( .A(n1208), .B(n1207), .Z(n1209) );
  ANDN U1627 ( .B(n1210), .A(n1209), .Z(n1211) );
  NANDN U1628 ( .A(n1212), .B(n1211), .Z(n1385) );
  NANDN U1629 ( .A(x[422]), .B(y[422]), .Z(n1214) );
  NANDN U1630 ( .A(x[423]), .B(y[423]), .Z(n1213) );
  NAND U1631 ( .A(n1214), .B(n1213), .Z(n2454) );
  NANDN U1632 ( .A(y[427]), .B(x[427]), .Z(n1216) );
  NANDN U1633 ( .A(y[428]), .B(x[428]), .Z(n1215) );
  NAND U1634 ( .A(n1216), .B(n1215), .Z(n2464) );
  NANDN U1635 ( .A(y[421]), .B(x[421]), .Z(n1218) );
  NANDN U1636 ( .A(y[422]), .B(x[422]), .Z(n1217) );
  NAND U1637 ( .A(n1218), .B(n1217), .Z(n2452) );
  NOR U1638 ( .A(n2464), .B(n2452), .Z(n1221) );
  NANDN U1639 ( .A(y[429]), .B(x[429]), .Z(n1220) );
  NANDN U1640 ( .A(y[430]), .B(x[430]), .Z(n1219) );
  NAND U1641 ( .A(n1220), .B(n1219), .Z(n2468) );
  ANDN U1642 ( .B(n1221), .A(n2468), .Z(n1222) );
  NANDN U1643 ( .A(n2454), .B(n1222), .Z(n1258) );
  NANDN U1644 ( .A(y[411]), .B(x[411]), .Z(n1224) );
  NANDN U1645 ( .A(y[412]), .B(x[412]), .Z(n1223) );
  NAND U1646 ( .A(n1224), .B(n1223), .Z(n2432) );
  NANDN U1647 ( .A(x[406]), .B(y[406]), .Z(n1226) );
  NANDN U1648 ( .A(x[407]), .B(y[407]), .Z(n1225) );
  NAND U1649 ( .A(n1226), .B(n1225), .Z(n2421) );
  NANDN U1650 ( .A(x[410]), .B(y[410]), .Z(n1228) );
  NANDN U1651 ( .A(x[411]), .B(y[411]), .Z(n1227) );
  NAND U1652 ( .A(n1228), .B(n1227), .Z(n2430) );
  NOR U1653 ( .A(n2421), .B(n2430), .Z(n1231) );
  NANDN U1654 ( .A(x[416]), .B(y[416]), .Z(n1230) );
  NANDN U1655 ( .A(x[417]), .B(y[417]), .Z(n1229) );
  NAND U1656 ( .A(n1230), .B(n1229), .Z(n2442) );
  ANDN U1657 ( .B(n1231), .A(n2442), .Z(n1232) );
  NANDN U1658 ( .A(n2432), .B(n1232), .Z(n1244) );
  NANDN U1659 ( .A(y[403]), .B(x[403]), .Z(n1234) );
  NANDN U1660 ( .A(y[404]), .B(x[404]), .Z(n1233) );
  NAND U1661 ( .A(n1234), .B(n1233), .Z(n2416) );
  NANDN U1662 ( .A(x[398]), .B(y[398]), .Z(n1236) );
  NANDN U1663 ( .A(x[399]), .B(y[399]), .Z(n1235) );
  NAND U1664 ( .A(n1236), .B(n1235), .Z(n2406) );
  NANDN U1665 ( .A(y[401]), .B(x[401]), .Z(n1238) );
  NANDN U1666 ( .A(y[402]), .B(x[402]), .Z(n1237) );
  NAND U1667 ( .A(n1238), .B(n1237), .Z(n2412) );
  NOR U1668 ( .A(n2406), .B(n2412), .Z(n1241) );
  NANDN U1669 ( .A(x[404]), .B(y[404]), .Z(n1240) );
  NANDN U1670 ( .A(x[405]), .B(y[405]), .Z(n1239) );
  NAND U1671 ( .A(n1240), .B(n1239), .Z(n2418) );
  ANDN U1672 ( .B(n1241), .A(n2418), .Z(n1242) );
  NANDN U1673 ( .A(n2416), .B(n1242), .Z(n1243) );
  NOR U1674 ( .A(n1244), .B(n1243), .Z(n1256) );
  NANDN U1675 ( .A(x[418]), .B(y[418]), .Z(n1246) );
  NANDN U1676 ( .A(x[419]), .B(y[419]), .Z(n1245) );
  NAND U1677 ( .A(n1246), .B(n1245), .Z(n2445) );
  NANDN U1678 ( .A(y[413]), .B(x[413]), .Z(n1248) );
  NANDN U1679 ( .A(y[414]), .B(x[414]), .Z(n1247) );
  NAND U1680 ( .A(n1248), .B(n1247), .Z(n2436) );
  NANDN U1681 ( .A(x[414]), .B(y[414]), .Z(n1250) );
  NANDN U1682 ( .A(x[415]), .B(y[415]), .Z(n1249) );
  NAND U1683 ( .A(n1250), .B(n1249), .Z(n2438) );
  NOR U1684 ( .A(n2436), .B(n2438), .Z(n1253) );
  NANDN U1685 ( .A(y[419]), .B(x[419]), .Z(n1252) );
  NANDN U1686 ( .A(y[420]), .B(x[420]), .Z(n1251) );
  NAND U1687 ( .A(n1252), .B(n1251), .Z(n2448) );
  ANDN U1688 ( .B(n1253), .A(n2448), .Z(n1254) );
  NANDN U1689 ( .A(n2445), .B(n1254), .Z(n1255) );
  ANDN U1690 ( .B(n1256), .A(n1255), .Z(n1257) );
  NANDN U1691 ( .A(n1258), .B(n1257), .Z(n1306) );
  NANDN U1692 ( .A(x[400]), .B(y[400]), .Z(n1260) );
  NANDN U1693 ( .A(x[401]), .B(y[401]), .Z(n1259) );
  NAND U1694 ( .A(n1260), .B(n1259), .Z(n2409) );
  NANDN U1695 ( .A(y[393]), .B(x[393]), .Z(n1262) );
  NANDN U1696 ( .A(y[394]), .B(x[394]), .Z(n1261) );
  NAND U1697 ( .A(n1262), .B(n1261), .Z(n2396) );
  NANDN U1698 ( .A(y[395]), .B(x[395]), .Z(n1264) );
  NANDN U1699 ( .A(y[396]), .B(x[396]), .Z(n1263) );
  NAND U1700 ( .A(n1264), .B(n1263), .Z(n2400) );
  NOR U1701 ( .A(n2396), .B(n2400), .Z(n1267) );
  NANDN U1702 ( .A(x[396]), .B(y[396]), .Z(n1266) );
  NANDN U1703 ( .A(x[397]), .B(y[397]), .Z(n1265) );
  NAND U1704 ( .A(n1266), .B(n1265), .Z(n2402) );
  ANDN U1705 ( .B(n1267), .A(n2402), .Z(n1268) );
  NANDN U1706 ( .A(n2409), .B(n1268), .Z(n1304) );
  NANDN U1707 ( .A(x[373]), .B(y[373]), .Z(n1270) );
  NANDN U1708 ( .A(x[374]), .B(y[374]), .Z(n1269) );
  NAND U1709 ( .A(n1270), .B(n1269), .Z(n2349) );
  NANDN U1710 ( .A(y[378]), .B(x[378]), .Z(n1272) );
  NANDN U1711 ( .A(y[379]), .B(x[379]), .Z(n1271) );
  NAND U1712 ( .A(n1272), .B(n1271), .Z(n2359) );
  NANDN U1713 ( .A(y[370]), .B(x[370]), .Z(n1274) );
  NANDN U1714 ( .A(y[371]), .B(x[371]), .Z(n1273) );
  NAND U1715 ( .A(n1274), .B(n1273), .Z(n2343) );
  NOR U1716 ( .A(n2359), .B(n2343), .Z(n1277) );
  NANDN U1717 ( .A(x[379]), .B(y[379]), .Z(n1276) );
  NANDN U1718 ( .A(x[380]), .B(y[380]), .Z(n1275) );
  NAND U1719 ( .A(n1276), .B(n1275), .Z(n2361) );
  ANDN U1720 ( .B(n1277), .A(n2361), .Z(n1278) );
  NANDN U1721 ( .A(n2349), .B(n1278), .Z(n1290) );
  NANDN U1722 ( .A(y[366]), .B(x[366]), .Z(n1280) );
  NANDN U1723 ( .A(y[367]), .B(x[367]), .Z(n1279) );
  NAND U1724 ( .A(n1280), .B(n1279), .Z(n2335) );
  NANDN U1725 ( .A(y[364]), .B(x[364]), .Z(n1282) );
  NANDN U1726 ( .A(y[365]), .B(x[365]), .Z(n1281) );
  NAND U1727 ( .A(n1282), .B(n1281), .Z(n2331) );
  NANDN U1728 ( .A(x[365]), .B(y[365]), .Z(n1284) );
  NANDN U1729 ( .A(x[366]), .B(y[366]), .Z(n1283) );
  NAND U1730 ( .A(n1284), .B(n1283), .Z(n2333) );
  NOR U1731 ( .A(n2331), .B(n2333), .Z(n1287) );
  NANDN U1732 ( .A(y[368]), .B(x[368]), .Z(n1286) );
  NANDN U1733 ( .A(y[369]), .B(x[369]), .Z(n1285) );
  NAND U1734 ( .A(n1286), .B(n1285), .Z(n2339) );
  ANDN U1735 ( .B(n1287), .A(n2339), .Z(n1288) );
  NANDN U1736 ( .A(n2335), .B(n1288), .Z(n1289) );
  NOR U1737 ( .A(n1290), .B(n1289), .Z(n1302) );
  NANDN U1738 ( .A(y[387]), .B(x[387]), .Z(n1292) );
  NANDN U1739 ( .A(y[388]), .B(x[388]), .Z(n1291) );
  NAND U1740 ( .A(n1292), .B(n1291), .Z(n2384) );
  NANDN U1741 ( .A(x[386]), .B(y[386]), .Z(n1294) );
  NANDN U1742 ( .A(x[387]), .B(y[387]), .Z(n1293) );
  NAND U1743 ( .A(n1294), .B(n1293), .Z(n2382) );
  NANDN U1744 ( .A(x[392]), .B(y[392]), .Z(n1296) );
  NANDN U1745 ( .A(x[393]), .B(y[393]), .Z(n1295) );
  NAND U1746 ( .A(n1296), .B(n1295), .Z(n2394) );
  NOR U1747 ( .A(n2382), .B(n2394), .Z(n1299) );
  NANDN U1748 ( .A(x[390]), .B(y[390]), .Z(n1298) );
  NANDN U1749 ( .A(x[391]), .B(y[391]), .Z(n1297) );
  NAND U1750 ( .A(n1298), .B(n1297), .Z(n2390) );
  ANDN U1751 ( .B(n1299), .A(n2390), .Z(n1300) );
  NANDN U1752 ( .A(n2384), .B(n1300), .Z(n1301) );
  ANDN U1753 ( .B(n1302), .A(n1301), .Z(n1303) );
  NANDN U1754 ( .A(n1304), .B(n1303), .Z(n1305) );
  NOR U1755 ( .A(n1306), .B(n1305), .Z(n1383) );
  NANDN U1756 ( .A(x[290]), .B(y[290]), .Z(n2176) );
  NANDN U1757 ( .A(x[261]), .B(y[261]), .Z(n1595) );
  NANDN U1758 ( .A(x[237]), .B(y[237]), .Z(n2086) );
  ANDN U1759 ( .B(x[246]), .A(y[246]), .Z(n2097) );
  IV U1760 ( .A(y[248]), .Z(n2101) );
  NOR U1761 ( .A(n2101), .B(x[248]), .Z(n1307) );
  NOR U1762 ( .A(n2097), .B(n1307), .Z(n1308) );
  AND U1763 ( .A(n2086), .B(n1308), .Z(n1309) );
  NANDN U1764 ( .A(x[262]), .B(y[262]), .Z(n1596) );
  NAND U1765 ( .A(n1309), .B(n1596), .Z(n1312) );
  NANDN U1766 ( .A(x[274]), .B(y[274]), .Z(n1311) );
  NANDN U1767 ( .A(x[275]), .B(y[275]), .Z(n1310) );
  NAND U1768 ( .A(n1311), .B(n1310), .Z(n2143) );
  NOR U1769 ( .A(n1312), .B(n2143), .Z(n1313) );
  AND U1770 ( .A(n1595), .B(n1313), .Z(n1314) );
  NANDN U1771 ( .A(x[283]), .B(y[283]), .Z(n2158) );
  NAND U1772 ( .A(n1314), .B(n2158), .Z(n1317) );
  NANDN U1773 ( .A(x[294]), .B(y[294]), .Z(n1316) );
  NANDN U1774 ( .A(x[295]), .B(y[295]), .Z(n1315) );
  NAND U1775 ( .A(n1316), .B(n1315), .Z(n2186) );
  NOR U1776 ( .A(n1317), .B(n2186), .Z(n1318) );
  AND U1777 ( .A(n2176), .B(n1318), .Z(n1319) );
  NANDN U1778 ( .A(x[352]), .B(y[352]), .Z(n1588) );
  NAND U1779 ( .A(n1319), .B(n1588), .Z(n1322) );
  NANDN U1780 ( .A(x[368]), .B(y[368]), .Z(n1321) );
  NANDN U1781 ( .A(x[367]), .B(y[367]), .Z(n1320) );
  NAND U1782 ( .A(n1321), .B(n1320), .Z(n2337) );
  NOR U1783 ( .A(n1322), .B(n2337), .Z(n1323) );
  ANDN U1784 ( .B(x[323]), .A(y[323]), .Z(n2245) );
  ANDN U1785 ( .B(n1323), .A(n2245), .Z(n1324) );
  NANDN U1786 ( .A(n1325), .B(n1324), .Z(n1381) );
  ANDN U1787 ( .B(x[509]), .A(y[509]), .Z(n2627) );
  NANDN U1788 ( .A(x[480]), .B(y[480]), .Z(n2563) );
  NANDN U1789 ( .A(y[506]), .B(x[506]), .Z(n2617) );
  ANDN U1790 ( .B(x[494]), .A(y[494]), .Z(n2591) );
  ANDN U1791 ( .B(n2617), .A(n2591), .Z(n1326) );
  AND U1792 ( .A(n2563), .B(n1326), .Z(n1327) );
  NANDN U1793 ( .A(n2627), .B(n1327), .Z(n1341) );
  ANDN U1794 ( .B(x[462]), .A(y[462]), .Z(n2536) );
  ANDN U1795 ( .B(x[386]), .A(y[386]), .Z(n2374) );
  NANDN U1796 ( .A(x[437]), .B(y[437]), .Z(n2487) );
  NANDN U1797 ( .A(x[394]), .B(y[394]), .Z(n1329) );
  NANDN U1798 ( .A(x[395]), .B(y[395]), .Z(n1328) );
  NAND U1799 ( .A(n1329), .B(n1328), .Z(n2397) );
  NANDN U1800 ( .A(x[484]), .B(y[484]), .Z(n1586) );
  ANDN U1801 ( .B(y[469]), .A(x[469]), .Z(n2551) );
  ANDN U1802 ( .B(n1586), .A(n2551), .Z(n1330) );
  ANDN U1803 ( .B(x[467]), .A(y[467]), .Z(n2550) );
  ANDN U1804 ( .B(n1330), .A(n2550), .Z(n1331) );
  NANDN U1805 ( .A(y[461]), .B(x[461]), .Z(n2537) );
  NAND U1806 ( .A(n1331), .B(n2537), .Z(n1332) );
  NOR U1807 ( .A(n2397), .B(n1332), .Z(n1333) );
  AND U1808 ( .A(n2487), .B(n1333), .Z(n1334) );
  NANDN U1809 ( .A(n2374), .B(n1334), .Z(n1337) );
  NANDN U1810 ( .A(x[450]), .B(y[450]), .Z(n1336) );
  NANDN U1811 ( .A(x[451]), .B(y[451]), .Z(n1335) );
  NAND U1812 ( .A(n1336), .B(n1335), .Z(n2515) );
  NOR U1813 ( .A(n1337), .B(n2515), .Z(n1338) );
  ANDN U1814 ( .B(x[435]), .A(y[435]), .Z(n2479) );
  ANDN U1815 ( .B(n1338), .A(n2479), .Z(n1339) );
  NANDN U1816 ( .A(n2536), .B(n1339), .Z(n1340) );
  NOR U1817 ( .A(n1341), .B(n1340), .Z(n1379) );
  ANDN U1818 ( .B(x[68]), .A(y[68]), .Z(n1741) );
  NANDN U1819 ( .A(x[45]), .B(y[45]), .Z(n1601) );
  ANDN U1820 ( .B(x[3]), .A(y[3]), .Z(n1608) );
  NANDN U1821 ( .A(x[44]), .B(y[44]), .Z(n1602) );
  NANDN U1822 ( .A(y[32]), .B(x[32]), .Z(n1343) );
  NANDN U1823 ( .A(y[31]), .B(x[31]), .Z(n1342) );
  NAND U1824 ( .A(n1343), .B(n1342), .Z(n1670) );
  ANDN U1825 ( .B(x[67]), .A(y[67]), .Z(n1744) );
  NANDN U1826 ( .A(x[89]), .B(y[89]), .Z(n1792) );
  ANDN U1827 ( .B(x[128]), .A(y[128]), .Z(n1871) );
  ANDN U1828 ( .B(n1792), .A(n1871), .Z(n1344) );
  ANDN U1829 ( .B(x[76]), .A(y[76]), .Z(n1759) );
  ANDN U1830 ( .B(n1344), .A(n1759), .Z(n1345) );
  NANDN U1831 ( .A(n1744), .B(n1345), .Z(n1346) );
  NOR U1832 ( .A(n1670), .B(n1346), .Z(n1347) );
  AND U1833 ( .A(n1602), .B(n1347), .Z(n1348) );
  NANDN U1834 ( .A(n1608), .B(n1348), .Z(n1351) );
  NANDN U1835 ( .A(x[55]), .B(y[55]), .Z(n1350) );
  NANDN U1836 ( .A(x[54]), .B(y[54]), .Z(n1349) );
  NAND U1837 ( .A(n1350), .B(n1349), .Z(n1716) );
  NOR U1838 ( .A(n1351), .B(n1716), .Z(n1352) );
  AND U1839 ( .A(n1601), .B(n1352), .Z(n1353) );
  NANDN U1840 ( .A(n1741), .B(n1353), .Z(n1377) );
  NANDN U1841 ( .A(x[20]), .B(y[20]), .Z(n1645) );
  XNOR U1842 ( .A(y[256]), .B(x[256]), .Z(n1355) );
  NANDN U1843 ( .A(y[257]), .B(x[257]), .Z(n1598) );
  NANDN U1844 ( .A(y[255]), .B(x[255]), .Z(n1597) );
  AND U1845 ( .A(n1598), .B(n1597), .Z(n1354) );
  NAND U1846 ( .A(n1355), .B(n1354), .Z(n1374) );
  NANDN U1847 ( .A(x[209]), .B(y[209]), .Z(n1600) );
  NANDN U1848 ( .A(x[193]), .B(y[193]), .Z(n1357) );
  NANDN U1849 ( .A(x[192]), .B(y[192]), .Z(n1356) );
  NAND U1850 ( .A(n1357), .B(n1356), .Z(n2002) );
  ANDN U1851 ( .B(y[208]), .A(x[208]), .Z(n1599) );
  OR U1852 ( .A(n2002), .B(n1599), .Z(n1360) );
  ANDN U1853 ( .B(x[137]), .A(y[137]), .Z(n1896) );
  ANDN U1854 ( .B(x[145]), .A(y[145]), .Z(n1911) );
  ANDN U1855 ( .B(x[149]), .A(y[149]), .Z(n1925) );
  NOR U1856 ( .A(n1911), .B(n1925), .Z(n1358) );
  NANDN U1857 ( .A(n1896), .B(n1358), .Z(n1359) );
  NOR U1858 ( .A(n1360), .B(n1359), .Z(n1362) );
  XNOR U1859 ( .A(x[182]), .B(y[182]), .Z(n1361) );
  NAND U1860 ( .A(n1362), .B(n1361), .Z(n1365) );
  NANDN U1861 ( .A(y[116]), .B(x[116]), .Z(n1364) );
  NANDN U1862 ( .A(y[115]), .B(x[115]), .Z(n1363) );
  NAND U1863 ( .A(n1364), .B(n1363), .Z(n1848) );
  NOR U1864 ( .A(n1365), .B(n1848), .Z(n1366) );
  ANDN U1865 ( .B(x[138]), .A(y[138]), .Z(n1894) );
  ANDN U1866 ( .B(n1366), .A(n1894), .Z(n1367) );
  NANDN U1867 ( .A(y[127]), .B(x[127]), .Z(n1872) );
  NAND U1868 ( .A(n1367), .B(n1872), .Z(n1370) );
  NANDN U1869 ( .A(y[217]), .B(x[217]), .Z(n1369) );
  NANDN U1870 ( .A(y[218]), .B(x[218]), .Z(n1368) );
  NAND U1871 ( .A(n1369), .B(n1368), .Z(n2049) );
  NOR U1872 ( .A(n1370), .B(n2049), .Z(n1371) );
  AND U1873 ( .A(n1600), .B(n1371), .Z(n1372) );
  NANDN U1874 ( .A(x[240]), .B(y[240]), .Z(n2091) );
  NAND U1875 ( .A(n1372), .B(n2091), .Z(n1373) );
  NOR U1876 ( .A(n1374), .B(n1373), .Z(n1375) );
  AND U1877 ( .A(n1645), .B(n1375), .Z(n1376) );
  NANDN U1878 ( .A(n1377), .B(n1376), .Z(n1378) );
  ANDN U1879 ( .B(n1379), .A(n1378), .Z(n1380) );
  NANDN U1880 ( .A(n1381), .B(n1380), .Z(n1382) );
  ANDN U1881 ( .B(n1383), .A(n1382), .Z(n1384) );
  NANDN U1882 ( .A(n1385), .B(n1384), .Z(n1386) );
  ANDN U1883 ( .B(n1387), .A(n1386), .Z(n1388) );
  NANDN U1884 ( .A(n1389), .B(n1388), .Z(n1390) );
  ANDN U1885 ( .B(n1391), .A(n1390), .Z(n1583) );
  NANDN U1886 ( .A(x[464]), .B(y[464]), .Z(n1393) );
  NANDN U1887 ( .A(x[465]), .B(y[465]), .Z(n1392) );
  NAND U1888 ( .A(n1393), .B(n1392), .Z(n2544) );
  NANDN U1889 ( .A(x[454]), .B(y[454]), .Z(n1395) );
  NANDN U1890 ( .A(x[455]), .B(y[455]), .Z(n1394) );
  NAND U1891 ( .A(n1395), .B(n1394), .Z(n2522) );
  NANDN U1892 ( .A(x[456]), .B(y[456]), .Z(n1397) );
  NANDN U1893 ( .A(x[457]), .B(y[457]), .Z(n1396) );
  NAND U1894 ( .A(n1397), .B(n1396), .Z(n2527) );
  NOR U1895 ( .A(n2522), .B(n2527), .Z(n1400) );
  NANDN U1896 ( .A(y[465]), .B(x[465]), .Z(n1399) );
  NANDN U1897 ( .A(y[466]), .B(x[466]), .Z(n1398) );
  NAND U1898 ( .A(n1399), .B(n1398), .Z(n2547) );
  ANDN U1899 ( .B(n1400), .A(n2547), .Z(n1401) );
  NANDN U1900 ( .A(n2544), .B(n1401), .Z(n1437) );
  NANDN U1901 ( .A(x[448]), .B(y[448]), .Z(n1403) );
  NANDN U1902 ( .A(x[449]), .B(y[449]), .Z(n1402) );
  NAND U1903 ( .A(n1403), .B(n1402), .Z(n2510) );
  NANDN U1904 ( .A(y[441]), .B(x[441]), .Z(n1405) );
  NANDN U1905 ( .A(y[442]), .B(x[442]), .Z(n1404) );
  NAND U1906 ( .A(n1405), .B(n1404), .Z(n2497) );
  NANDN U1907 ( .A(x[442]), .B(y[442]), .Z(n1407) );
  NANDN U1908 ( .A(x[443]), .B(y[443]), .Z(n1406) );
  NAND U1909 ( .A(n1407), .B(n1406), .Z(n2498) );
  NOR U1910 ( .A(n2497), .B(n2498), .Z(n1410) );
  NANDN U1911 ( .A(x[444]), .B(y[444]), .Z(n1409) );
  NANDN U1912 ( .A(x[445]), .B(y[445]), .Z(n1408) );
  NAND U1913 ( .A(n1409), .B(n1408), .Z(n2503) );
  ANDN U1914 ( .B(n1410), .A(n2503), .Z(n1411) );
  NANDN U1915 ( .A(n2510), .B(n1411), .Z(n1423) );
  NANDN U1916 ( .A(x[438]), .B(y[438]), .Z(n1413) );
  NANDN U1917 ( .A(x[439]), .B(y[439]), .Z(n1412) );
  NAND U1918 ( .A(n1413), .B(n1412), .Z(n2491) );
  NANDN U1919 ( .A(x[434]), .B(y[434]), .Z(n1415) );
  NANDN U1920 ( .A(x[435]), .B(y[435]), .Z(n1414) );
  NAND U1921 ( .A(n1415), .B(n1414), .Z(n2478) );
  NANDN U1922 ( .A(x[440]), .B(y[440]), .Z(n1417) );
  NANDN U1923 ( .A(x[441]), .B(y[441]), .Z(n1416) );
  NAND U1924 ( .A(n1417), .B(n1416), .Z(n2495) );
  NOR U1925 ( .A(n2478), .B(n2495), .Z(n1420) );
  NANDN U1926 ( .A(y[439]), .B(x[439]), .Z(n1419) );
  NANDN U1927 ( .A(y[440]), .B(x[440]), .Z(n1418) );
  NAND U1928 ( .A(n1419), .B(n1418), .Z(n2493) );
  ANDN U1929 ( .B(n1420), .A(n2493), .Z(n1421) );
  NANDN U1930 ( .A(n2491), .B(n1421), .Z(n1422) );
  NOR U1931 ( .A(n1423), .B(n1422), .Z(n1435) );
  NANDN U1932 ( .A(y[453]), .B(x[453]), .Z(n1425) );
  NANDN U1933 ( .A(y[454]), .B(x[454]), .Z(n1424) );
  NAND U1934 ( .A(n1425), .B(n1424), .Z(n2521) );
  NANDN U1935 ( .A(x[446]), .B(y[446]), .Z(n1427) );
  NANDN U1936 ( .A(x[447]), .B(y[447]), .Z(n1426) );
  NAND U1937 ( .A(n1427), .B(n1426), .Z(n2507) );
  NANDN U1938 ( .A(x[452]), .B(y[452]), .Z(n1429) );
  NANDN U1939 ( .A(x[453]), .B(y[453]), .Z(n1428) );
  NAND U1940 ( .A(n1429), .B(n1428), .Z(n2519) );
  NOR U1941 ( .A(n2507), .B(n2519), .Z(n1432) );
  NANDN U1942 ( .A(x[458]), .B(y[458]), .Z(n1431) );
  NANDN U1943 ( .A(x[459]), .B(y[459]), .Z(n1430) );
  NAND U1944 ( .A(n1431), .B(n1430), .Z(n2531) );
  ANDN U1945 ( .B(n1432), .A(n2531), .Z(n1433) );
  NANDN U1946 ( .A(n2521), .B(n1433), .Z(n1434) );
  ANDN U1947 ( .B(n1435), .A(n1434), .Z(n1436) );
  NANDN U1948 ( .A(n1437), .B(n1436), .Z(n1581) );
  NANDN U1949 ( .A(y[389]), .B(x[389]), .Z(n1439) );
  NANDN U1950 ( .A(y[390]), .B(x[390]), .Z(n1438) );
  NAND U1951 ( .A(n1439), .B(n1438), .Z(n2388) );
  NANDN U1952 ( .A(y[382]), .B(x[382]), .Z(n1441) );
  NANDN U1953 ( .A(y[383]), .B(x[383]), .Z(n1440) );
  NAND U1954 ( .A(n1441), .B(n1440), .Z(n2367) );
  NANDN U1955 ( .A(x[388]), .B(y[388]), .Z(n1443) );
  NANDN U1956 ( .A(x[389]), .B(y[389]), .Z(n1442) );
  NAND U1957 ( .A(n1443), .B(n1442), .Z(n2385) );
  NOR U1958 ( .A(n2367), .B(n2385), .Z(n1446) );
  NANDN U1959 ( .A(y[399]), .B(x[399]), .Z(n1445) );
  NANDN U1960 ( .A(y[400]), .B(x[400]), .Z(n1444) );
  NAND U1961 ( .A(n1445), .B(n1444), .Z(n2408) );
  ANDN U1962 ( .B(n1446), .A(n2408), .Z(n1447) );
  NANDN U1963 ( .A(n2388), .B(n1447), .Z(n1483) );
  NANDN U1964 ( .A(y[376]), .B(x[376]), .Z(n1449) );
  NANDN U1965 ( .A(y[377]), .B(x[377]), .Z(n1448) );
  NAND U1966 ( .A(n1449), .B(n1448), .Z(n2355) );
  NANDN U1967 ( .A(x[371]), .B(y[371]), .Z(n1451) );
  NANDN U1968 ( .A(x[372]), .B(y[372]), .Z(n1450) );
  NAND U1969 ( .A(n1451), .B(n1450), .Z(n2345) );
  NANDN U1970 ( .A(y[372]), .B(x[372]), .Z(n1453) );
  NANDN U1971 ( .A(y[373]), .B(x[373]), .Z(n1452) );
  NAND U1972 ( .A(n1453), .B(n1452), .Z(n2347) );
  NOR U1973 ( .A(n2345), .B(n2347), .Z(n1456) );
  NANDN U1974 ( .A(y[374]), .B(x[374]), .Z(n1455) );
  NANDN U1975 ( .A(y[375]), .B(x[375]), .Z(n1454) );
  NAND U1976 ( .A(n1455), .B(n1454), .Z(n2351) );
  ANDN U1977 ( .B(n1456), .A(n2351), .Z(n1457) );
  NANDN U1978 ( .A(n2355), .B(n1457), .Z(n1469) );
  NANDN U1979 ( .A(x[357]), .B(y[357]), .Z(n1459) );
  NANDN U1980 ( .A(x[358]), .B(y[358]), .Z(n1458) );
  NAND U1981 ( .A(n1459), .B(n1458), .Z(n2317) );
  NANDN U1982 ( .A(x[355]), .B(y[355]), .Z(n1461) );
  NANDN U1983 ( .A(x[356]), .B(y[356]), .Z(n1460) );
  NAND U1984 ( .A(n1461), .B(n1460), .Z(n2315) );
  NANDN U1985 ( .A(x[369]), .B(y[369]), .Z(n1463) );
  NANDN U1986 ( .A(x[370]), .B(y[370]), .Z(n1462) );
  NAND U1987 ( .A(n1463), .B(n1462), .Z(n2340) );
  NOR U1988 ( .A(n2315), .B(n2340), .Z(n1466) );
  NANDN U1989 ( .A(x[361]), .B(y[361]), .Z(n1465) );
  NANDN U1990 ( .A(x[362]), .B(y[362]), .Z(n1464) );
  NAND U1991 ( .A(n1465), .B(n1464), .Z(n2325) );
  ANDN U1992 ( .B(n1466), .A(n2325), .Z(n1467) );
  NANDN U1993 ( .A(n2317), .B(n1467), .Z(n1468) );
  NOR U1994 ( .A(n1469), .B(n1468), .Z(n1481) );
  NANDN U1995 ( .A(y[380]), .B(x[380]), .Z(n1471) );
  NANDN U1996 ( .A(y[381]), .B(x[381]), .Z(n1470) );
  NAND U1997 ( .A(n1471), .B(n1470), .Z(n2363) );
  NANDN U1998 ( .A(x[375]), .B(y[375]), .Z(n1473) );
  NANDN U1999 ( .A(x[376]), .B(y[376]), .Z(n1472) );
  NAND U2000 ( .A(n1473), .B(n1472), .Z(n2352) );
  NANDN U2001 ( .A(x[377]), .B(y[377]), .Z(n1475) );
  NANDN U2002 ( .A(x[378]), .B(y[378]), .Z(n1474) );
  NAND U2003 ( .A(n1475), .B(n1474), .Z(n2357) );
  NOR U2004 ( .A(n2352), .B(n2357), .Z(n1478) );
  NANDN U2005 ( .A(x[381]), .B(y[381]), .Z(n1477) );
  NANDN U2006 ( .A(x[382]), .B(y[382]), .Z(n1476) );
  NAND U2007 ( .A(n1477), .B(n1476), .Z(n2364) );
  ANDN U2008 ( .B(n1478), .A(n2364), .Z(n1479) );
  NANDN U2009 ( .A(n2363), .B(n1479), .Z(n1480) );
  ANDN U2010 ( .B(n1481), .A(n1480), .Z(n1482) );
  NANDN U2011 ( .A(n1483), .B(n1482), .Z(n1531) );
  NANDN U2012 ( .A(y[340]), .B(x[340]), .Z(n1485) );
  NANDN U2013 ( .A(y[341]), .B(x[341]), .Z(n1484) );
  NAND U2014 ( .A(n1485), .B(n1484), .Z(n2293) );
  NANDN U2015 ( .A(x[342]), .B(y[342]), .Z(n1487) );
  NANDN U2016 ( .A(x[343]), .B(y[343]), .Z(n1486) );
  NAND U2017 ( .A(n1487), .B(n1486), .Z(n2299) );
  NANDN U2018 ( .A(y[337]), .B(x[337]), .Z(n1489) );
  NANDN U2019 ( .A(y[338]), .B(x[338]), .Z(n1488) );
  NAND U2020 ( .A(n1489), .B(n1488), .Z(n2283) );
  NOR U2021 ( .A(n2299), .B(n2283), .Z(n1492) );
  NANDN U2022 ( .A(x[353]), .B(y[353]), .Z(n1491) );
  NANDN U2023 ( .A(x[354]), .B(y[354]), .Z(n1490) );
  NAND U2024 ( .A(n1491), .B(n1490), .Z(n2313) );
  ANDN U2025 ( .B(n1492), .A(n2313), .Z(n1493) );
  NANDN U2026 ( .A(n2293), .B(n1493), .Z(n1529) );
  NANDN U2027 ( .A(y[319]), .B(x[319]), .Z(n1495) );
  NANDN U2028 ( .A(y[320]), .B(x[320]), .Z(n1494) );
  NAND U2029 ( .A(n1495), .B(n1494), .Z(n2237) );
  NANDN U2030 ( .A(y[313]), .B(x[313]), .Z(n1497) );
  NANDN U2031 ( .A(y[314]), .B(x[314]), .Z(n1496) );
  NAND U2032 ( .A(n1497), .B(n1496), .Z(n2225) );
  NANDN U2033 ( .A(x[316]), .B(y[316]), .Z(n1499) );
  NANDN U2034 ( .A(x[317]), .B(y[317]), .Z(n1498) );
  NAND U2035 ( .A(n1499), .B(n1498), .Z(n2231) );
  NOR U2036 ( .A(n2225), .B(n2231), .Z(n1502) );
  NANDN U2037 ( .A(x[320]), .B(y[320]), .Z(n1501) );
  NANDN U2038 ( .A(x[321]), .B(y[321]), .Z(n1500) );
  NAND U2039 ( .A(n1501), .B(n1500), .Z(n2239) );
  ANDN U2040 ( .B(n1502), .A(n2239), .Z(n1503) );
  NANDN U2041 ( .A(n2237), .B(n1503), .Z(n1515) );
  NANDN U2042 ( .A(y[311]), .B(x[311]), .Z(n1505) );
  NANDN U2043 ( .A(y[312]), .B(x[312]), .Z(n1504) );
  NAND U2044 ( .A(n1505), .B(n1504), .Z(n2221) );
  NANDN U2045 ( .A(x[308]), .B(y[308]), .Z(n1507) );
  NANDN U2046 ( .A(x[309]), .B(y[309]), .Z(n1506) );
  NAND U2047 ( .A(n1507), .B(n1506), .Z(n2215) );
  NANDN U2048 ( .A(x[310]), .B(y[310]), .Z(n1509) );
  NANDN U2049 ( .A(x[311]), .B(y[311]), .Z(n1508) );
  NAND U2050 ( .A(n1509), .B(n1508), .Z(n2219) );
  NOR U2051 ( .A(n2215), .B(n2219), .Z(n1512) );
  NANDN U2052 ( .A(y[317]), .B(x[317]), .Z(n1511) );
  NANDN U2053 ( .A(y[318]), .B(x[318]), .Z(n1510) );
  NAND U2054 ( .A(n1511), .B(n1510), .Z(n2233) );
  ANDN U2055 ( .B(n1512), .A(n2233), .Z(n1513) );
  NANDN U2056 ( .A(n2221), .B(n1513), .Z(n1514) );
  NOR U2057 ( .A(n1515), .B(n1514), .Z(n1527) );
  NANDN U2058 ( .A(x[332]), .B(y[332]), .Z(n1517) );
  NANDN U2059 ( .A(x[333]), .B(y[333]), .Z(n1516) );
  NAND U2060 ( .A(n1517), .B(n1516), .Z(n2271) );
  NANDN U2061 ( .A(x[329]), .B(y[329]), .Z(n1519) );
  NANDN U2062 ( .A(x[328]), .B(y[328]), .Z(n1518) );
  NAND U2063 ( .A(n1519), .B(n1518), .Z(n2259) );
  NANDN U2064 ( .A(y[331]), .B(x[331]), .Z(n1521) );
  NANDN U2065 ( .A(y[330]), .B(x[330]), .Z(n1520) );
  NAND U2066 ( .A(n1521), .B(n1520), .Z(n2265) );
  NOR U2067 ( .A(n2259), .B(n2265), .Z(n1524) );
  NANDN U2068 ( .A(x[334]), .B(y[334]), .Z(n1523) );
  NANDN U2069 ( .A(x[335]), .B(y[335]), .Z(n1522) );
  NAND U2070 ( .A(n1523), .B(n1522), .Z(n2274) );
  ANDN U2071 ( .B(n1524), .A(n2274), .Z(n1525) );
  NANDN U2072 ( .A(n2271), .B(n1525), .Z(n1526) );
  ANDN U2073 ( .B(n1527), .A(n1526), .Z(n1528) );
  NANDN U2074 ( .A(n1529), .B(n1528), .Z(n1530) );
  NOR U2075 ( .A(n1531), .B(n1530), .Z(n1579) );
  NANDN U2076 ( .A(y[431]), .B(x[431]), .Z(n1533) );
  NANDN U2077 ( .A(y[432]), .B(x[432]), .Z(n1532) );
  NAND U2078 ( .A(n1533), .B(n1532), .Z(n2472) );
  NANDN U2079 ( .A(x[428]), .B(y[428]), .Z(n1535) );
  NANDN U2080 ( .A(x[429]), .B(y[429]), .Z(n1534) );
  NAND U2081 ( .A(n1535), .B(n1534), .Z(n2466) );
  NANDN U2082 ( .A(x[430]), .B(y[430]), .Z(n1537) );
  NANDN U2083 ( .A(x[431]), .B(y[431]), .Z(n1536) );
  NAND U2084 ( .A(n1537), .B(n1536), .Z(n2469) );
  NOR U2085 ( .A(n2466), .B(n2469), .Z(n1540) );
  NANDN U2086 ( .A(x[432]), .B(y[432]), .Z(n1539) );
  NANDN U2087 ( .A(x[433]), .B(y[433]), .Z(n1538) );
  NAND U2088 ( .A(n1539), .B(n1538), .Z(n2473) );
  ANDN U2089 ( .B(n1540), .A(n2473), .Z(n1541) );
  NANDN U2090 ( .A(n2472), .B(n1541), .Z(n1577) );
  NANDN U2091 ( .A(y[415]), .B(x[415]), .Z(n1543) );
  NANDN U2092 ( .A(y[416]), .B(x[416]), .Z(n1542) );
  NAND U2093 ( .A(n1543), .B(n1542), .Z(n2440) );
  NANDN U2094 ( .A(x[408]), .B(y[408]), .Z(n1545) );
  NANDN U2095 ( .A(x[409]), .B(y[409]), .Z(n1544) );
  NAND U2096 ( .A(n1545), .B(n1544), .Z(n2426) );
  NANDN U2097 ( .A(y[409]), .B(x[409]), .Z(n1547) );
  NANDN U2098 ( .A(y[410]), .B(x[410]), .Z(n1546) );
  NAND U2099 ( .A(n1547), .B(n1546), .Z(n2428) );
  NOR U2100 ( .A(n2426), .B(n2428), .Z(n1550) );
  NANDN U2101 ( .A(y[417]), .B(x[417]), .Z(n1549) );
  NANDN U2102 ( .A(y[418]), .B(x[418]), .Z(n1548) );
  NAND U2103 ( .A(n1549), .B(n1548), .Z(n2444) );
  ANDN U2104 ( .B(n1550), .A(n2444), .Z(n1551) );
  NANDN U2105 ( .A(n2440), .B(n1551), .Z(n1563) );
  NANDN U2106 ( .A(y[405]), .B(x[405]), .Z(n1553) );
  NANDN U2107 ( .A(y[406]), .B(x[406]), .Z(n1552) );
  NAND U2108 ( .A(n1553), .B(n1552), .Z(n2420) );
  NANDN U2109 ( .A(y[391]), .B(x[391]), .Z(n1555) );
  NANDN U2110 ( .A(y[392]), .B(x[392]), .Z(n1554) );
  NAND U2111 ( .A(n1555), .B(n1554), .Z(n2392) );
  NANDN U2112 ( .A(y[397]), .B(x[397]), .Z(n1557) );
  NANDN U2113 ( .A(y[398]), .B(x[398]), .Z(n1556) );
  NAND U2114 ( .A(n1557), .B(n1556), .Z(n2404) );
  NOR U2115 ( .A(n2392), .B(n2404), .Z(n1560) );
  NANDN U2116 ( .A(y[407]), .B(x[407]), .Z(n1559) );
  NANDN U2117 ( .A(y[408]), .B(x[408]), .Z(n1558) );
  NAND U2118 ( .A(n1559), .B(n1558), .Z(n2424) );
  ANDN U2119 ( .B(n1560), .A(n2424), .Z(n1561) );
  NANDN U2120 ( .A(n2420), .B(n1561), .Z(n1562) );
  NOR U2121 ( .A(n1563), .B(n1562), .Z(n1575) );
  NANDN U2122 ( .A(x[424]), .B(y[424]), .Z(n1565) );
  NANDN U2123 ( .A(x[425]), .B(y[425]), .Z(n1564) );
  NAND U2124 ( .A(n1565), .B(n1564), .Z(n2457) );
  NANDN U2125 ( .A(y[425]), .B(x[425]), .Z(n1567) );
  NANDN U2126 ( .A(y[426]), .B(x[426]), .Z(n1566) );
  NAND U2127 ( .A(n1567), .B(n1566), .Z(n2460) );
  NANDN U2128 ( .A(y[423]), .B(x[423]), .Z(n1569) );
  NANDN U2129 ( .A(y[424]), .B(x[424]), .Z(n1568) );
  NAND U2130 ( .A(n1569), .B(n1568), .Z(n2456) );
  NOR U2131 ( .A(n2460), .B(n2456), .Z(n1572) );
  NANDN U2132 ( .A(x[426]), .B(y[426]), .Z(n1571) );
  NANDN U2133 ( .A(x[427]), .B(y[427]), .Z(n1570) );
  NAND U2134 ( .A(n1571), .B(n1570), .Z(n2462) );
  ANDN U2135 ( .B(n1572), .A(n2462), .Z(n1573) );
  NANDN U2136 ( .A(n2457), .B(n1573), .Z(n1574) );
  ANDN U2137 ( .B(n1575), .A(n1574), .Z(n1576) );
  NANDN U2138 ( .A(n1577), .B(n1576), .Z(n1578) );
  ANDN U2139 ( .B(n1579), .A(n1578), .Z(n1580) );
  NANDN U2140 ( .A(n1581), .B(n1580), .Z(n1582) );
  ANDN U2141 ( .B(n1583), .A(n1582), .Z(n1584) );
  NANDN U2142 ( .A(ebreg), .B(n1584), .Z(n5) );
  OR U2143 ( .A(n1584), .B(ebreg), .Z(n2635) );
  AND U2144 ( .A(n1586), .B(n1585), .Z(n2573) );
  NANDN U2145 ( .A(y[346]), .B(x[346]), .Z(n1590) );
  NAND U2146 ( .A(n1590), .B(n1589), .Z(n2305) );
  ANDN U2147 ( .B(x[339]), .A(y[339]), .Z(n2289) );
  AND U2148 ( .A(n1592), .B(n1591), .Z(n2251) );
  OR U2149 ( .A(n1594), .B(n1593), .Z(n2121) );
  AND U2150 ( .A(n1596), .B(n1595), .Z(n2117) );
  ANDN U2151 ( .B(n1600), .A(n1599), .Z(n2031) );
  AND U2152 ( .A(n1602), .B(n1601), .Z(n1696) );
  OR U2153 ( .A(n1604), .B(n1603), .Z(n1606) );
  ANDN U2154 ( .B(n1606), .A(n1605), .Z(n1607) );
  NANDN U2155 ( .A(n1608), .B(n1607), .Z(n1609) );
  NANDN U2156 ( .A(n1610), .B(n1609), .Z(n1611) );
  NANDN U2157 ( .A(n1612), .B(n1611), .Z(n1614) );
  ANDN U2158 ( .B(n1614), .A(n1613), .Z(n1615) );
  OR U2159 ( .A(n1616), .B(n1615), .Z(n1618) );
  NAND U2160 ( .A(n1618), .B(n1617), .Z(n1619) );
  NANDN U2161 ( .A(n1620), .B(n1619), .Z(n1621) );
  NANDN U2162 ( .A(n1622), .B(n1621), .Z(n1623) );
  NANDN U2163 ( .A(n1624), .B(n1623), .Z(n1626) );
  ANDN U2164 ( .B(n1626), .A(n1625), .Z(n1627) );
  OR U2165 ( .A(n1628), .B(n1627), .Z(n1629) );
  NANDN U2166 ( .A(n1630), .B(n1629), .Z(n1631) );
  NANDN U2167 ( .A(n1632), .B(n1631), .Z(n1633) );
  NANDN U2168 ( .A(n1634), .B(n1633), .Z(n1635) );
  NANDN U2169 ( .A(n1636), .B(n1635), .Z(n1638) );
  ANDN U2170 ( .B(n1638), .A(n1637), .Z(n1639) );
  OR U2171 ( .A(n1640), .B(n1639), .Z(n1641) );
  NANDN U2172 ( .A(n1642), .B(n1641), .Z(n1643) );
  NANDN U2173 ( .A(n1644), .B(n1643), .Z(n1646) );
  AND U2174 ( .A(n1646), .B(n1645), .Z(n1648) );
  NAND U2175 ( .A(n1648), .B(n1647), .Z(n1649) );
  NANDN U2176 ( .A(n1650), .B(n1649), .Z(n1651) );
  NANDN U2177 ( .A(n1652), .B(n1651), .Z(n1653) );
  NANDN U2178 ( .A(n1654), .B(n1653), .Z(n1656) );
  ANDN U2179 ( .B(n1656), .A(n1655), .Z(n1657) );
  OR U2180 ( .A(n1658), .B(n1657), .Z(n1659) );
  NANDN U2181 ( .A(n1660), .B(n1659), .Z(n1661) );
  NANDN U2182 ( .A(n1662), .B(n1661), .Z(n1663) );
  NANDN U2183 ( .A(n1664), .B(n1663), .Z(n1665) );
  NANDN U2184 ( .A(n1666), .B(n1665), .Z(n1668) );
  ANDN U2185 ( .B(n1668), .A(n1667), .Z(n1669) );
  OR U2186 ( .A(n1670), .B(n1669), .Z(n1671) );
  NANDN U2187 ( .A(n1672), .B(n1671), .Z(n1673) );
  NANDN U2188 ( .A(n1674), .B(n1673), .Z(n1675) );
  NANDN U2189 ( .A(n1676), .B(n1675), .Z(n1677) );
  NANDN U2190 ( .A(n1678), .B(n1677), .Z(n1680) );
  ANDN U2191 ( .B(n1680), .A(n1679), .Z(n1681) );
  OR U2192 ( .A(n1682), .B(n1681), .Z(n1683) );
  NANDN U2193 ( .A(n1684), .B(n1683), .Z(n1685) );
  NANDN U2194 ( .A(n1686), .B(n1685), .Z(n1687) );
  NANDN U2195 ( .A(n1688), .B(n1687), .Z(n1689) );
  NANDN U2196 ( .A(n1690), .B(n1689), .Z(n1692) );
  ANDN U2197 ( .B(n1692), .A(n1691), .Z(n1693) );
  OR U2198 ( .A(n1694), .B(n1693), .Z(n1695) );
  AND U2199 ( .A(n1696), .B(n1695), .Z(n1697) );
  OR U2200 ( .A(n1698), .B(n1697), .Z(n1699) );
  NANDN U2201 ( .A(n1700), .B(n1699), .Z(n1701) );
  NANDN U2202 ( .A(n1702), .B(n1701), .Z(n1703) );
  NANDN U2203 ( .A(n1704), .B(n1703), .Z(n1705) );
  NANDN U2204 ( .A(n1706), .B(n1705), .Z(n1708) );
  ANDN U2205 ( .B(n1708), .A(n1707), .Z(n1709) );
  OR U2206 ( .A(n1710), .B(n1709), .Z(n1711) );
  NANDN U2207 ( .A(n1712), .B(n1711), .Z(n1713) );
  NANDN U2208 ( .A(n1714), .B(n1713), .Z(n1715) );
  NANDN U2209 ( .A(n1716), .B(n1715), .Z(n1717) );
  NANDN U2210 ( .A(n1718), .B(n1717), .Z(n1720) );
  ANDN U2211 ( .B(n1720), .A(n1719), .Z(n1721) );
  OR U2212 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U2213 ( .A(n1724), .B(n1723), .Z(n1725) );
  NANDN U2214 ( .A(n1726), .B(n1725), .Z(n1727) );
  NANDN U2215 ( .A(n1728), .B(n1727), .Z(n1729) );
  NANDN U2216 ( .A(n1730), .B(n1729), .Z(n1732) );
  ANDN U2217 ( .B(n1732), .A(n1731), .Z(n1733) );
  OR U2218 ( .A(n1734), .B(n1733), .Z(n1735) );
  NANDN U2219 ( .A(n1736), .B(n1735), .Z(n1737) );
  NANDN U2220 ( .A(n1738), .B(n1737), .Z(n1739) );
  NANDN U2221 ( .A(n1740), .B(n1739), .Z(n1742) );
  ANDN U2222 ( .B(n1742), .A(n1741), .Z(n1743) );
  NANDN U2223 ( .A(n1744), .B(n1743), .Z(n1745) );
  NANDN U2224 ( .A(n1746), .B(n1745), .Z(n1747) );
  NANDN U2225 ( .A(n1748), .B(n1747), .Z(n1750) );
  ANDN U2226 ( .B(n1750), .A(n1749), .Z(n1751) );
  OR U2227 ( .A(n1752), .B(n1751), .Z(n1753) );
  NANDN U2228 ( .A(n1754), .B(n1753), .Z(n1755) );
  NANDN U2229 ( .A(n1756), .B(n1755), .Z(n1757) );
  NANDN U2230 ( .A(n1758), .B(n1757), .Z(n1760) );
  ANDN U2231 ( .B(n1760), .A(n1759), .Z(n1761) );
  NANDN U2232 ( .A(n1762), .B(n1761), .Z(n1763) );
  NANDN U2233 ( .A(n1764), .B(n1763), .Z(n1765) );
  NANDN U2234 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U2235 ( .A(n1768), .B(n1767), .Z(n1769) );
  OR U2236 ( .A(n1770), .B(n1769), .Z(n1772) );
  NAND U2237 ( .A(n1772), .B(n1771), .Z(n1773) );
  NANDN U2238 ( .A(n1774), .B(n1773), .Z(n1775) );
  NANDN U2239 ( .A(n1776), .B(n1775), .Z(n1777) );
  NANDN U2240 ( .A(n1778), .B(n1777), .Z(n1780) );
  ANDN U2241 ( .B(n1780), .A(n1779), .Z(n1781) );
  OR U2242 ( .A(n1782), .B(n1781), .Z(n1783) );
  NANDN U2243 ( .A(n1784), .B(n1783), .Z(n1785) );
  NANDN U2244 ( .A(n1786), .B(n1785), .Z(n1787) );
  NANDN U2245 ( .A(n1788), .B(n1787), .Z(n1789) );
  NANDN U2246 ( .A(n1790), .B(n1789), .Z(n1791) );
  AND U2247 ( .A(n1792), .B(n1791), .Z(n1794) );
  NAND U2248 ( .A(n1794), .B(n1793), .Z(n1795) );
  NANDN U2249 ( .A(n1796), .B(n1795), .Z(n1798) );
  ANDN U2250 ( .B(n1798), .A(n1797), .Z(n1799) );
  OR U2251 ( .A(n1800), .B(n1799), .Z(n1801) );
  NANDN U2252 ( .A(n1802), .B(n1801), .Z(n1803) );
  NANDN U2253 ( .A(n1804), .B(n1803), .Z(n1805) );
  NANDN U2254 ( .A(n1806), .B(n1805), .Z(n1807) );
  NANDN U2255 ( .A(n1808), .B(n1807), .Z(n1810) );
  ANDN U2256 ( .B(n1810), .A(n1809), .Z(n1811) );
  OR U2257 ( .A(n1812), .B(n1811), .Z(n1813) );
  NANDN U2258 ( .A(n1814), .B(n1813), .Z(n1815) );
  NANDN U2259 ( .A(n1816), .B(n1815), .Z(n1817) );
  NANDN U2260 ( .A(n1818), .B(n1817), .Z(n1819) );
  NANDN U2261 ( .A(n1820), .B(n1819), .Z(n1822) );
  ANDN U2262 ( .B(n1822), .A(n1821), .Z(n1823) );
  OR U2263 ( .A(n1824), .B(n1823), .Z(n1825) );
  NANDN U2264 ( .A(n1826), .B(n1825), .Z(n1827) );
  NANDN U2265 ( .A(n1828), .B(n1827), .Z(n1829) );
  NANDN U2266 ( .A(n1830), .B(n1829), .Z(n1831) );
  NANDN U2267 ( .A(n1832), .B(n1831), .Z(n1834) );
  ANDN U2268 ( .B(n1834), .A(n1833), .Z(n1835) );
  OR U2269 ( .A(n1836), .B(n1835), .Z(n1837) );
  NANDN U2270 ( .A(n1838), .B(n1837), .Z(n1839) );
  NANDN U2271 ( .A(n1840), .B(n1839), .Z(n1841) );
  NANDN U2272 ( .A(n1842), .B(n1841), .Z(n1843) );
  NANDN U2273 ( .A(n1844), .B(n1843), .Z(n1846) );
  ANDN U2274 ( .B(n1846), .A(n1845), .Z(n1847) );
  OR U2275 ( .A(n1848), .B(n1847), .Z(n1849) );
  NANDN U2276 ( .A(n1850), .B(n1849), .Z(n1851) );
  NANDN U2277 ( .A(n1852), .B(n1851), .Z(n1853) );
  NANDN U2278 ( .A(n1854), .B(n1853), .Z(n1855) );
  NANDN U2279 ( .A(n1856), .B(n1855), .Z(n1858) );
  ANDN U2280 ( .B(n1858), .A(n1857), .Z(n1859) );
  OR U2281 ( .A(n1860), .B(n1859), .Z(n1861) );
  NANDN U2282 ( .A(n1862), .B(n1861), .Z(n1863) );
  NANDN U2283 ( .A(n1864), .B(n1863), .Z(n1865) );
  NANDN U2284 ( .A(n1866), .B(n1865), .Z(n1867) );
  NANDN U2285 ( .A(n1868), .B(n1867), .Z(n1870) );
  ANDN U2286 ( .B(n1870), .A(n1869), .Z(n1874) );
  ANDN U2287 ( .B(n1872), .A(n1871), .Z(n1873) );
  NANDN U2288 ( .A(n1874), .B(n1873), .Z(n1876) );
  ANDN U2289 ( .B(n1876), .A(n1875), .Z(n1877) );
  OR U2290 ( .A(n1878), .B(n1877), .Z(n1879) );
  NANDN U2291 ( .A(n1880), .B(n1879), .Z(n1881) );
  NANDN U2292 ( .A(n1882), .B(n1881), .Z(n1883) );
  NANDN U2293 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U2294 ( .A(n1886), .B(n1885), .Z(n1888) );
  ANDN U2295 ( .B(n1888), .A(n1887), .Z(n1889) );
  OR U2296 ( .A(n1890), .B(n1889), .Z(n1891) );
  NANDN U2297 ( .A(n1892), .B(n1891), .Z(n1893) );
  NANDN U2298 ( .A(n1894), .B(n1893), .Z(n1895) );
  OR U2299 ( .A(n1896), .B(n1895), .Z(n1897) );
  NANDN U2300 ( .A(n1898), .B(n1897), .Z(n1899) );
  NANDN U2301 ( .A(n1900), .B(n1899), .Z(n1901) );
  NANDN U2302 ( .A(n1902), .B(n1901), .Z(n1903) );
  NANDN U2303 ( .A(n1904), .B(n1903), .Z(n1906) );
  ANDN U2304 ( .B(n1906), .A(n1905), .Z(n1907) );
  OR U2305 ( .A(n1908), .B(n1907), .Z(n1909) );
  NANDN U2306 ( .A(n1910), .B(n1909), .Z(n1912) );
  ANDN U2307 ( .B(n1912), .A(n1911), .Z(n1913) );
  OR U2308 ( .A(n1913), .B(y[146]), .Z(n1917) );
  XNOR U2309 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2310 ( .A(n1915), .B(x[146]), .Z(n1916) );
  NAND U2311 ( .A(n1917), .B(n1916), .Z(n1918) );
  AND U2312 ( .A(n1919), .B(n1918), .Z(n1920) );
  OR U2313 ( .A(n1921), .B(n1920), .Z(n1922) );
  NANDN U2314 ( .A(n1923), .B(n1922), .Z(n1924) );
  NANDN U2315 ( .A(n1925), .B(n1924), .Z(n1926) );
  OR U2316 ( .A(n1927), .B(n1926), .Z(n1928) );
  NANDN U2317 ( .A(n1929), .B(n1928), .Z(n1930) );
  NANDN U2318 ( .A(n1931), .B(n1930), .Z(n1932) );
  NANDN U2319 ( .A(n1933), .B(n1932), .Z(n1934) );
  NANDN U2320 ( .A(n1935), .B(n1934), .Z(n1937) );
  ANDN U2321 ( .B(n1937), .A(n1936), .Z(n1938) );
  OR U2322 ( .A(n1939), .B(n1938), .Z(n1940) );
  NANDN U2323 ( .A(n1941), .B(n1940), .Z(n1942) );
  NANDN U2324 ( .A(n1943), .B(n1942), .Z(n1944) );
  NANDN U2325 ( .A(n1945), .B(n1944), .Z(n1946) );
  NANDN U2326 ( .A(n1947), .B(n1946), .Z(n1949) );
  ANDN U2327 ( .B(n1949), .A(n1948), .Z(n1950) );
  OR U2328 ( .A(n1951), .B(n1950), .Z(n1952) );
  NANDN U2329 ( .A(n1953), .B(n1952), .Z(n1954) );
  NANDN U2330 ( .A(n1955), .B(n1954), .Z(n1956) );
  NANDN U2331 ( .A(n1957), .B(n1956), .Z(n1958) );
  NANDN U2332 ( .A(n1959), .B(n1958), .Z(n1961) );
  ANDN U2333 ( .B(n1961), .A(n1960), .Z(n1962) );
  OR U2334 ( .A(n1963), .B(n1962), .Z(n1964) );
  NANDN U2335 ( .A(n1965), .B(n1964), .Z(n1966) );
  NANDN U2336 ( .A(n1967), .B(n1966), .Z(n1968) );
  NANDN U2337 ( .A(n1969), .B(n1968), .Z(n1970) );
  NANDN U2338 ( .A(n1971), .B(n1970), .Z(n1973) );
  ANDN U2339 ( .B(n1973), .A(n1972), .Z(n1974) );
  OR U2340 ( .A(n1975), .B(n1974), .Z(n1976) );
  NANDN U2341 ( .A(n1977), .B(n1976), .Z(n1978) );
  NANDN U2342 ( .A(n1979), .B(n1978), .Z(n1980) );
  NANDN U2343 ( .A(n1981), .B(n1980), .Z(n1982) );
  NANDN U2344 ( .A(n1983), .B(n1982), .Z(n1985) );
  ANDN U2345 ( .B(n1985), .A(n1984), .Z(n1986) );
  OR U2346 ( .A(n1987), .B(n1986), .Z(n1988) );
  NANDN U2347 ( .A(n1989), .B(n1988), .Z(n1991) );
  NANDN U2348 ( .A(n2007), .B(n2006), .Z(n2008) );
  NANDN U2349 ( .A(n2009), .B(n2008), .Z(n2010) );
  NANDN U2350 ( .A(n2011), .B(n2010), .Z(n2012) );
  NANDN U2351 ( .A(n2013), .B(n2012), .Z(n2015) );
  ANDN U2352 ( .B(n2015), .A(n2014), .Z(n2016) );
  OR U2353 ( .A(n2017), .B(n2016), .Z(n2018) );
  NANDN U2354 ( .A(n2019), .B(n2018), .Z(n2020) );
  NANDN U2355 ( .A(n2021), .B(n2020), .Z(n2022) );
  NANDN U2356 ( .A(n2023), .B(n2022), .Z(n2024) );
  NANDN U2357 ( .A(n2025), .B(n2024), .Z(n2027) );
  ANDN U2358 ( .B(n2027), .A(n2026), .Z(n2028) );
  OR U2359 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U2360 ( .A(n2031), .B(n2030), .Z(n2032) );
  OR U2361 ( .A(n2033), .B(n2032), .Z(n2034) );
  NANDN U2362 ( .A(n2035), .B(n2034), .Z(n2036) );
  NANDN U2363 ( .A(n2037), .B(n2036), .Z(n2038) );
  NANDN U2364 ( .A(n2039), .B(n2038), .Z(n2040) );
  NANDN U2365 ( .A(n2041), .B(n2040), .Z(n2043) );
  ANDN U2366 ( .B(n2043), .A(n2042), .Z(n2044) );
  OR U2367 ( .A(n2045), .B(n2044), .Z(n2046) );
  NANDN U2368 ( .A(n2047), .B(n2046), .Z(n2048) );
  NANDN U2369 ( .A(n2049), .B(n2048), .Z(n2050) );
  NANDN U2370 ( .A(n2051), .B(n2050), .Z(n2052) );
  NANDN U2371 ( .A(n2053), .B(n2052), .Z(n2055) );
  ANDN U2372 ( .B(n2055), .A(n2054), .Z(n2056) );
  OR U2373 ( .A(n2057), .B(n2056), .Z(n2058) );
  NANDN U2374 ( .A(n2059), .B(n2058), .Z(n2060) );
  NANDN U2375 ( .A(n2061), .B(n2060), .Z(n2062) );
  NANDN U2376 ( .A(n2063), .B(n2062), .Z(n2064) );
  NANDN U2377 ( .A(n2065), .B(n2064), .Z(n2067) );
  ANDN U2378 ( .B(n2067), .A(n2066), .Z(n2068) );
  OR U2379 ( .A(n2069), .B(n2068), .Z(n2070) );
  NANDN U2380 ( .A(n2071), .B(n2070), .Z(n2072) );
  NANDN U2381 ( .A(n2073), .B(n2072), .Z(n2074) );
  NANDN U2382 ( .A(n2075), .B(n2074), .Z(n2076) );
  NANDN U2383 ( .A(n2077), .B(n2076), .Z(n2079) );
  ANDN U2384 ( .B(n2079), .A(n2078), .Z(n2080) );
  OR U2385 ( .A(n2081), .B(n2080), .Z(n2082) );
  NANDN U2386 ( .A(n2083), .B(n2082), .Z(n2084) );
  XNOR U2387 ( .A(n2101), .B(n2100), .Z(n2102) );
  NAND U2388 ( .A(x[248]), .B(n2102), .Z(n2103) );
  OR U2389 ( .A(n2115), .B(n2114), .Z(n2116) );
  AND U2390 ( .A(n2117), .B(n2116), .Z(n2118) );
  OR U2391 ( .A(n2119), .B(n2118), .Z(n2120) );
  AND U2392 ( .A(n2121), .B(n2120), .Z(n2122) );
  NANDN U2393 ( .A(n2123), .B(n2122), .Z(n2124) );
  NANDN U2394 ( .A(n2125), .B(n2124), .Z(n2127) );
  ANDN U2395 ( .B(n2127), .A(n2126), .Z(n2128) );
  OR U2396 ( .A(n2129), .B(n2128), .Z(n2130) );
  NANDN U2397 ( .A(n2131), .B(n2130), .Z(n2132) );
  NANDN U2398 ( .A(n2133), .B(n2132), .Z(n2134) );
  NANDN U2399 ( .A(n2135), .B(n2134), .Z(n2136) );
  NANDN U2400 ( .A(n2137), .B(n2136), .Z(n2139) );
  ANDN U2401 ( .B(n2139), .A(n2138), .Z(n2140) );
  OR U2402 ( .A(n2141), .B(n2140), .Z(n2142) );
  NANDN U2403 ( .A(n2143), .B(n2142), .Z(n2144) );
  NANDN U2404 ( .A(n2145), .B(n2144), .Z(n2146) );
  NANDN U2405 ( .A(n2147), .B(n2146), .Z(n2148) );
  NANDN U2406 ( .A(n2149), .B(n2148), .Z(n2151) );
  ANDN U2407 ( .B(n2151), .A(n2150), .Z(n2152) );
  OR U2408 ( .A(n2153), .B(n2152), .Z(n2154) );
  NANDN U2409 ( .A(n2155), .B(n2154), .Z(n2156) );
  NANDN U2410 ( .A(n2157), .B(n2156), .Z(n2159) );
  AND U2411 ( .A(n2159), .B(n2158), .Z(n2160) );
  NANDN U2412 ( .A(n2161), .B(n2160), .Z(n2162) );
  NANDN U2413 ( .A(n2163), .B(n2162), .Z(n2164) );
  NANDN U2414 ( .A(n2165), .B(n2164), .Z(n2166) );
  NANDN U2415 ( .A(n2167), .B(n2166), .Z(n2169) );
  ANDN U2416 ( .B(n2169), .A(n2168), .Z(n2170) );
  OR U2417 ( .A(n2171), .B(n2170), .Z(n2172) );
  NANDN U2418 ( .A(n2173), .B(n2172), .Z(n2174) );
  NANDN U2419 ( .A(n2175), .B(n2174), .Z(n2177) );
  AND U2420 ( .A(n2177), .B(n2176), .Z(n2179) );
  NAND U2421 ( .A(n2179), .B(n2178), .Z(n2180) );
  NANDN U2422 ( .A(n2181), .B(n2180), .Z(n2182) );
  NANDN U2423 ( .A(n2183), .B(n2182), .Z(n2184) );
  NANDN U2424 ( .A(n2185), .B(n2184), .Z(n2187) );
  ANDN U2425 ( .B(n2187), .A(n2186), .Z(n2188) );
  OR U2426 ( .A(n2189), .B(n2188), .Z(n2190) );
  NANDN U2427 ( .A(n2191), .B(n2190), .Z(n2192) );
  NANDN U2428 ( .A(n2193), .B(n2192), .Z(n2194) );
  NANDN U2429 ( .A(n2195), .B(n2194), .Z(n2196) );
  NANDN U2430 ( .A(n2197), .B(n2196), .Z(n2199) );
  ANDN U2431 ( .B(n2199), .A(n2198), .Z(n2200) );
  OR U2432 ( .A(n2201), .B(n2200), .Z(n2202) );
  NANDN U2433 ( .A(n2203), .B(n2202), .Z(n2204) );
  NANDN U2434 ( .A(n2205), .B(n2204), .Z(n2206) );
  NANDN U2435 ( .A(n2207), .B(n2206), .Z(n2208) );
  NANDN U2436 ( .A(n2209), .B(n2208), .Z(n2211) );
  ANDN U2437 ( .B(n2211), .A(n2210), .Z(n2212) );
  OR U2438 ( .A(n2213), .B(n2212), .Z(n2214) );
  NANDN U2439 ( .A(n2215), .B(n2214), .Z(n2216) );
  NANDN U2440 ( .A(n2217), .B(n2216), .Z(n2218) );
  NANDN U2441 ( .A(n2219), .B(n2218), .Z(n2220) );
  NANDN U2442 ( .A(n2221), .B(n2220), .Z(n2223) );
  ANDN U2443 ( .B(n2223), .A(n2222), .Z(n2224) );
  OR U2444 ( .A(n2225), .B(n2224), .Z(n2226) );
  NANDN U2445 ( .A(n2227), .B(n2226), .Z(n2228) );
  NANDN U2446 ( .A(n2229), .B(n2228), .Z(n2230) );
  NANDN U2447 ( .A(n2231), .B(n2230), .Z(n2232) );
  NANDN U2448 ( .A(n2233), .B(n2232), .Z(n2235) );
  ANDN U2449 ( .B(n2235), .A(n2234), .Z(n2236) );
  OR U2450 ( .A(n2237), .B(n2236), .Z(n2238) );
  NANDN U2451 ( .A(n2239), .B(n2238), .Z(n2240) );
  NANDN U2452 ( .A(n2241), .B(n2240), .Z(n2242) );
  NANDN U2453 ( .A(n2243), .B(n2242), .Z(n2244) );
  NANDN U2454 ( .A(n2245), .B(n2244), .Z(n2246) );
  AND U2455 ( .A(n2247), .B(n2246), .Z(n2248) );
  OR U2456 ( .A(n2249), .B(n2248), .Z(n2250) );
  AND U2457 ( .A(n2251), .B(n2250), .Z(n2252) );
  OR U2458 ( .A(n2253), .B(n2252), .Z(n2255) );
  NAND U2459 ( .A(n2255), .B(n2254), .Z(n2256) );
  NANDN U2460 ( .A(n2257), .B(n2256), .Z(n2258) );
  NANDN U2461 ( .A(n2259), .B(n2258), .Z(n2260) );
  NANDN U2462 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U2463 ( .A(n2263), .B(n2262), .Z(n2264) );
  OR U2464 ( .A(n2265), .B(n2264), .Z(n2267) );
  NAND U2465 ( .A(n2267), .B(n2266), .Z(n2268) );
  NANDN U2466 ( .A(n2269), .B(n2268), .Z(n2270) );
  NANDN U2467 ( .A(n2271), .B(n2270), .Z(n2272) );
  NANDN U2468 ( .A(n2273), .B(n2272), .Z(n2275) );
  ANDN U2469 ( .B(n2275), .A(n2274), .Z(n2279) );
  NOR U2470 ( .A(n2277), .B(n2276), .Z(n2278) );
  NANDN U2471 ( .A(n2279), .B(n2278), .Z(n2281) );
  ANDN U2472 ( .B(n2281), .A(n2280), .Z(n2282) );
  OR U2473 ( .A(n2283), .B(n2282), .Z(n2287) );
  NANDN U2474 ( .A(x[339]), .B(y[339]), .Z(n2285) );
  AND U2475 ( .A(n2285), .B(n2284), .Z(n2286) );
  NAND U2476 ( .A(n2287), .B(n2286), .Z(n2288) );
  NANDN U2477 ( .A(n2289), .B(n2288), .Z(n2290) );
  NANDN U2478 ( .A(n2291), .B(n2290), .Z(n2292) );
  NANDN U2479 ( .A(n2293), .B(n2292), .Z(n2294) );
  AND U2480 ( .A(n2295), .B(n2294), .Z(n2296) );
  OR U2481 ( .A(n2297), .B(n2296), .Z(n2298) );
  NANDN U2482 ( .A(n2299), .B(n2298), .Z(n2300) );
  NANDN U2483 ( .A(n2301), .B(n2300), .Z(n2302) );
  NANDN U2484 ( .A(n2303), .B(n2302), .Z(n2304) );
  OR U2485 ( .A(n2319), .B(n2318), .Z(n2320) );
  NANDN U2486 ( .A(n2321), .B(n2320), .Z(n2322) );
  NANDN U2487 ( .A(n2323), .B(n2322), .Z(n2324) );
  NANDN U2488 ( .A(n2325), .B(n2324), .Z(n2326) );
  NANDN U2489 ( .A(n2327), .B(n2326), .Z(n2329) );
  ANDN U2490 ( .B(n2329), .A(n2328), .Z(n2330) );
  OR U2491 ( .A(n2331), .B(n2330), .Z(n2332) );
  NANDN U2492 ( .A(n2333), .B(n2332), .Z(n2334) );
  NANDN U2493 ( .A(n2335), .B(n2334), .Z(n2336) );
  NANDN U2494 ( .A(n2337), .B(n2336), .Z(n2338) );
  NANDN U2495 ( .A(n2339), .B(n2338), .Z(n2341) );
  ANDN U2496 ( .B(n2341), .A(n2340), .Z(n2342) );
  OR U2497 ( .A(n2343), .B(n2342), .Z(n2344) );
  NANDN U2498 ( .A(n2345), .B(n2344), .Z(n2346) );
  NANDN U2499 ( .A(n2347), .B(n2346), .Z(n2348) );
  NANDN U2500 ( .A(n2349), .B(n2348), .Z(n2350) );
  NANDN U2501 ( .A(n2351), .B(n2350), .Z(n2353) );
  ANDN U2502 ( .B(n2353), .A(n2352), .Z(n2354) );
  OR U2503 ( .A(n2355), .B(n2354), .Z(n2356) );
  NANDN U2504 ( .A(n2357), .B(n2356), .Z(n2358) );
  NANDN U2505 ( .A(n2359), .B(n2358), .Z(n2360) );
  NANDN U2506 ( .A(n2361), .B(n2360), .Z(n2362) );
  NANDN U2507 ( .A(n2363), .B(n2362), .Z(n2365) );
  ANDN U2508 ( .B(n2365), .A(n2364), .Z(n2366) );
  OR U2509 ( .A(n2367), .B(n2366), .Z(n2369) );
  NAND U2510 ( .A(n2369), .B(n2368), .Z(n2370) );
  NANDN U2511 ( .A(n2370), .B(x[384]), .Z(n2373) );
  XNOR U2512 ( .A(n2370), .B(x[384]), .Z(n2371) );
  NANDN U2513 ( .A(y[384]), .B(n2371), .Z(n2372) );
  AND U2514 ( .A(n2373), .B(n2372), .Z(n2376) );
  OR U2515 ( .A(n2376), .B(y[385]), .Z(n2375) );
  ANDN U2516 ( .B(n2375), .A(n2374), .Z(n2380) );
  XNOR U2517 ( .A(n2377), .B(n2376), .Z(n2378) );
  NAND U2518 ( .A(x[385]), .B(n2378), .Z(n2379) );
  NAND U2519 ( .A(n2380), .B(n2379), .Z(n2381) );
  NANDN U2520 ( .A(n2382), .B(n2381), .Z(n2383) );
  NANDN U2521 ( .A(n2384), .B(n2383), .Z(n2386) );
  ANDN U2522 ( .B(n2386), .A(n2385), .Z(n2387) );
  OR U2523 ( .A(n2388), .B(n2387), .Z(n2389) );
  NANDN U2524 ( .A(n2390), .B(n2389), .Z(n2391) );
  NANDN U2525 ( .A(n2392), .B(n2391), .Z(n2393) );
  NANDN U2526 ( .A(n2394), .B(n2393), .Z(n2395) );
  NANDN U2527 ( .A(n2396), .B(n2395), .Z(n2398) );
  ANDN U2528 ( .B(n2398), .A(n2397), .Z(n2399) );
  OR U2529 ( .A(n2400), .B(n2399), .Z(n2401) );
  NANDN U2530 ( .A(n2402), .B(n2401), .Z(n2403) );
  NANDN U2531 ( .A(n2404), .B(n2403), .Z(n2405) );
  NANDN U2532 ( .A(n2406), .B(n2405), .Z(n2407) );
  NANDN U2533 ( .A(n2408), .B(n2407), .Z(n2410) );
  ANDN U2534 ( .B(n2410), .A(n2409), .Z(n2411) );
  OR U2535 ( .A(n2412), .B(n2411), .Z(n2413) );
  NANDN U2536 ( .A(n2414), .B(n2413), .Z(n2415) );
  NANDN U2537 ( .A(n2416), .B(n2415), .Z(n2417) );
  NANDN U2538 ( .A(n2418), .B(n2417), .Z(n2419) );
  NANDN U2539 ( .A(n2420), .B(n2419), .Z(n2422) );
  ANDN U2540 ( .B(n2422), .A(n2421), .Z(n2423) );
  OR U2541 ( .A(n2424), .B(n2423), .Z(n2425) );
  NANDN U2542 ( .A(n2426), .B(n2425), .Z(n2427) );
  NANDN U2543 ( .A(n2428), .B(n2427), .Z(n2429) );
  NANDN U2544 ( .A(n2430), .B(n2429), .Z(n2431) );
  NANDN U2545 ( .A(n2432), .B(n2431), .Z(n2434) );
  ANDN U2546 ( .B(n2434), .A(n2433), .Z(n2435) );
  OR U2547 ( .A(n2436), .B(n2435), .Z(n2437) );
  NANDN U2548 ( .A(n2438), .B(n2437), .Z(n2439) );
  NANDN U2549 ( .A(n2440), .B(n2439), .Z(n2441) );
  NANDN U2550 ( .A(n2442), .B(n2441), .Z(n2443) );
  NANDN U2551 ( .A(n2444), .B(n2443), .Z(n2446) );
  ANDN U2552 ( .B(n2446), .A(n2445), .Z(n2447) );
  OR U2553 ( .A(n2448), .B(n2447), .Z(n2449) );
  NANDN U2554 ( .A(n2450), .B(n2449), .Z(n2451) );
  NANDN U2555 ( .A(n2452), .B(n2451), .Z(n2453) );
  NANDN U2556 ( .A(n2454), .B(n2453), .Z(n2455) );
  NANDN U2557 ( .A(n2456), .B(n2455), .Z(n2458) );
  ANDN U2558 ( .B(n2458), .A(n2457), .Z(n2459) );
  OR U2559 ( .A(n2460), .B(n2459), .Z(n2461) );
  NANDN U2560 ( .A(n2462), .B(n2461), .Z(n2463) );
  NANDN U2561 ( .A(n2464), .B(n2463), .Z(n2465) );
  NANDN U2562 ( .A(n2466), .B(n2465), .Z(n2467) );
  NANDN U2563 ( .A(n2468), .B(n2467), .Z(n2470) );
  ANDN U2564 ( .B(n2470), .A(n2469), .Z(n2471) );
  OR U2565 ( .A(n2472), .B(n2471), .Z(n2474) );
  ANDN U2566 ( .B(n2474), .A(n2473), .Z(n2475) );
  OR U2567 ( .A(n2476), .B(n2475), .Z(n2477) );
  NANDN U2568 ( .A(n2478), .B(n2477), .Z(n2480) );
  ANDN U2569 ( .B(n2480), .A(n2479), .Z(n2481) );
  OR U2570 ( .A(n2481), .B(y[436]), .Z(n2485) );
  XNOR U2571 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U2572 ( .A(n2483), .B(x[436]), .Z(n2484) );
  NAND U2573 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2574 ( .A(n2487), .B(n2486), .Z(n2488) );
  OR U2575 ( .A(n2489), .B(n2488), .Z(n2490) );
  NANDN U2576 ( .A(n2491), .B(n2490), .Z(n2492) );
  NANDN U2577 ( .A(n2493), .B(n2492), .Z(n2494) );
  NANDN U2578 ( .A(n2495), .B(n2494), .Z(n2496) );
  NANDN U2579 ( .A(n2497), .B(n2496), .Z(n2499) );
  ANDN U2580 ( .B(n2499), .A(n2498), .Z(n2500) );
  OR U2581 ( .A(n2501), .B(n2500), .Z(n2502) );
  NANDN U2582 ( .A(n2503), .B(n2502), .Z(n2504) );
  NANDN U2583 ( .A(n2505), .B(n2504), .Z(n2506) );
  NANDN U2584 ( .A(n2507), .B(n2506), .Z(n2508) );
  NANDN U2585 ( .A(n2509), .B(n2508), .Z(n2511) );
  ANDN U2586 ( .B(n2511), .A(n2510), .Z(n2512) );
  OR U2587 ( .A(n2513), .B(n2512), .Z(n2514) );
  NANDN U2588 ( .A(n2515), .B(n2514), .Z(n2516) );
  NANDN U2589 ( .A(n2517), .B(n2516), .Z(n2518) );
  NANDN U2590 ( .A(n2519), .B(n2518), .Z(n2520) );
  NANDN U2591 ( .A(n2521), .B(n2520), .Z(n2523) );
  ANDN U2592 ( .B(n2523), .A(n2522), .Z(n2524) );
  OR U2593 ( .A(n2525), .B(n2524), .Z(n2526) );
  NANDN U2594 ( .A(n2527), .B(n2526), .Z(n2528) );
  NANDN U2595 ( .A(n2529), .B(n2528), .Z(n2530) );
  NANDN U2596 ( .A(n2531), .B(n2530), .Z(n2532) );
  NANDN U2597 ( .A(n2533), .B(n2532), .Z(n2535) );
  ANDN U2598 ( .B(n2535), .A(n2534), .Z(n2539) );
  ANDN U2599 ( .B(n2537), .A(n2536), .Z(n2538) );
  NANDN U2600 ( .A(n2539), .B(n2538), .Z(n2541) );
  ANDN U2601 ( .B(n2541), .A(n2540), .Z(n2542) );
  OR U2602 ( .A(n2543), .B(n2542), .Z(n2545) );
  ANDN U2603 ( .B(n2545), .A(n2544), .Z(n2546) );
  OR U2604 ( .A(n2547), .B(n2546), .Z(n2548) );
  NAND U2605 ( .A(n2565), .B(n2564), .Z(n2566) );
  NANDN U2606 ( .A(n2567), .B(n2566), .Z(n2569) );
  ANDN U2607 ( .B(n2569), .A(n2568), .Z(n2570) );
  OR U2608 ( .A(n2571), .B(n2570), .Z(n2572) );
  AND U2609 ( .A(n2573), .B(n2572), .Z(n2574) );
  OR U2610 ( .A(n2575), .B(n2574), .Z(n2576) );
  NANDN U2611 ( .A(n2577), .B(n2576), .Z(n2578) );
  NANDN U2612 ( .A(n2579), .B(n2578), .Z(n2580) );
  NANDN U2613 ( .A(n2581), .B(n2580), .Z(n2582) );
  NANDN U2614 ( .A(n2583), .B(n2582), .Z(n2585) );
  ANDN U2615 ( .B(n2585), .A(n2584), .Z(n2586) );
  OR U2616 ( .A(n2587), .B(n2586), .Z(n2588) );
  NANDN U2617 ( .A(n2589), .B(n2588), .Z(n2590) );
  NANDN U2618 ( .A(n2591), .B(n2590), .Z(n2592) );
  OR U2619 ( .A(n2593), .B(n2592), .Z(n2594) );
  NANDN U2620 ( .A(n2595), .B(n2594), .Z(n2596) );
  NANDN U2621 ( .A(n2597), .B(n2596), .Z(n2598) );
  NANDN U2622 ( .A(n2599), .B(n2598), .Z(n2600) );
  NANDN U2623 ( .A(n2601), .B(n2600), .Z(n2603) );
  ANDN U2624 ( .B(n2603), .A(n2602), .Z(n2604) );
  OR U2625 ( .A(n2605), .B(n2604), .Z(n2606) );
  NANDN U2626 ( .A(n2607), .B(n2606), .Z(n2608) );
  NANDN U2627 ( .A(n2609), .B(n2608), .Z(n2610) );
  NANDN U2628 ( .A(n2611), .B(n2610), .Z(n2612) );
  NANDN U2629 ( .A(n2613), .B(n2612), .Z(n2615) );
  ANDN U2630 ( .B(n2615), .A(n2614), .Z(n2619) );
  ANDN U2631 ( .B(n2617), .A(n2616), .Z(n2618) );
  NANDN U2632 ( .A(n2619), .B(n2618), .Z(n2621) );
  ANDN U2633 ( .B(n2621), .A(n2620), .Z(n2622) );
  OR U2634 ( .A(n2623), .B(n2622), .Z(n2624) );
  NANDN U2635 ( .A(n2625), .B(n2624), .Z(n2626) );
  NANDN U2636 ( .A(n2627), .B(n2626), .Z(n2628) );
  OR U2637 ( .A(n2629), .B(n2628), .Z(n2630) );
  NANDN U2638 ( .A(n2631), .B(n2630), .Z(n2632) );
  NANDN U2639 ( .A(n2633), .B(n2632), .Z(n2634) );
  NANDN U2640 ( .A(n2635), .B(n2634), .Z(n2637) );
  NAND U2641 ( .A(n2635), .B(g), .Z(n2636) );
  NAND U2642 ( .A(n2637), .B(n2636), .Z(n4) );
endmodule

