
module k_nns_seq_W31_K4 ( clk, rst, q, DB, min_val_out );
  input [30:0] q;
  input [30:0] DB;
  output [123:0] min_val_out;
  input clk, rst;
  wire   \min_dist_reg[3][4] , \min_dist_reg[3][3] , \min_dist_reg[3][2] ,
         \min_dist_reg[3][1] , \min_dist_reg[3][0] , \min_dist_reg[2][4] ,
         \min_dist_reg[2][3] , \min_dist_reg[2][2] , \min_dist_reg[2][1] ,
         \min_dist_reg[2][0] , \min_dist_reg[1][4] , \min_dist_reg[1][3] ,
         \min_dist_reg[1][2] , \min_dist_reg[1][1] , \min_dist_reg[1][0] ,
         \min_dist_reg[0][4] , \min_dist_reg[0][3] , \min_dist_reg[0][2] ,
         \min_dist_reg[0][1] , \min_dist_reg[0][0] , \local_min_dist[0][4] ,
         \local_min_dist[0][3] , \local_min_dist[0][2] ,
         \local_min_dist[0][1] , \local_min_dist[0][0] , \min_dist[3][4] ,
         \min_dist[3][3] , \min_dist[3][2] , \min_dist[3][1] ,
         \min_dist[3][0] , \min_dist[2][4] , \min_dist[2][3] ,
         \min_dist[2][2] , \min_dist[2][1] , \min_dist[2][0] ,
         \min_dist[1][4] , \min_dist[1][3] , \min_dist[1][2] ,
         \min_dist[1][1] , \min_dist[1][0] , \min_val_reg[3][30] ,
         \min_val_reg[3][29] , \min_val_reg[3][28] , \min_val_reg[3][27] ,
         \min_val_reg[3][26] , \min_val_reg[3][25] , \min_val_reg[3][24] ,
         \min_val_reg[3][23] , \min_val_reg[3][22] , \min_val_reg[3][21] ,
         \min_val_reg[3][20] , \min_val_reg[3][19] , \min_val_reg[3][18] ,
         \min_val_reg[3][17] , \min_val_reg[3][16] , \min_val_reg[3][15] ,
         \min_val_reg[3][14] , \min_val_reg[3][13] , \min_val_reg[3][12] ,
         \min_val_reg[3][11] , \min_val_reg[3][10] , \min_val_reg[3][9] ,
         \min_val_reg[3][8] , \min_val_reg[3][7] , \min_val_reg[3][6] ,
         \min_val_reg[3][5] , \min_val_reg[3][4] , \min_val_reg[3][3] ,
         \min_val_reg[3][2] , \min_val_reg[3][1] , \min_val_reg[3][0] ,
         \min_val_reg[2][30] , \min_val_reg[2][29] , \min_val_reg[2][28] ,
         \min_val_reg[2][27] , \min_val_reg[2][26] , \min_val_reg[2][25] ,
         \min_val_reg[2][24] , \min_val_reg[2][23] , \min_val_reg[2][22] ,
         \min_val_reg[2][21] , \min_val_reg[2][20] , \min_val_reg[2][19] ,
         \min_val_reg[2][18] , \min_val_reg[2][17] , \min_val_reg[2][16] ,
         \min_val_reg[2][15] , \min_val_reg[2][14] , \min_val_reg[2][13] ,
         \min_val_reg[2][12] , \min_val_reg[2][11] , \min_val_reg[2][10] ,
         \min_val_reg[2][9] , \min_val_reg[2][8] , \min_val_reg[2][7] ,
         \min_val_reg[2][6] , \min_val_reg[2][5] , \min_val_reg[2][4] ,
         \min_val_reg[2][3] , \min_val_reg[2][2] , \min_val_reg[2][1] ,
         \min_val_reg[2][0] , \min_val_reg[1][30] , \min_val_reg[1][29] ,
         \min_val_reg[1][28] , \min_val_reg[1][27] , \min_val_reg[1][26] ,
         \min_val_reg[1][25] , \min_val_reg[1][24] , \min_val_reg[1][23] ,
         \min_val_reg[1][22] , \min_val_reg[1][21] , \min_val_reg[1][20] ,
         \min_val_reg[1][19] , \min_val_reg[1][18] , \min_val_reg[1][17] ,
         \min_val_reg[1][16] , \min_val_reg[1][15] , \min_val_reg[1][14] ,
         \min_val_reg[1][13] , \min_val_reg[1][12] , \min_val_reg[1][11] ,
         \min_val_reg[1][10] , \min_val_reg[1][9] , \min_val_reg[1][8] ,
         \min_val_reg[1][7] , \min_val_reg[1][6] , \min_val_reg[1][5] ,
         \min_val_reg[1][4] , \min_val_reg[1][3] , \min_val_reg[1][2] ,
         \min_val_reg[1][1] , \min_val_reg[1][0] , \min_val_reg[0][30] ,
         \min_val_reg[0][29] , \min_val_reg[0][28] , \min_val_reg[0][27] ,
         \min_val_reg[0][26] , \min_val_reg[0][25] , \min_val_reg[0][24] ,
         \min_val_reg[0][23] , \min_val_reg[0][22] , \min_val_reg[0][21] ,
         \min_val_reg[0][20] , \min_val_reg[0][19] , \min_val_reg[0][18] ,
         \min_val_reg[0][17] , \min_val_reg[0][16] , \min_val_reg[0][15] ,
         \min_val_reg[0][14] , \min_val_reg[0][13] , \min_val_reg[0][12] ,
         \min_val_reg[0][11] , \min_val_reg[0][10] , \min_val_reg[0][9] ,
         \min_val_reg[0][8] , \min_val_reg[0][7] , \min_val_reg[0][6] ,
         \min_val_reg[0][5] , \min_val_reg[0][4] , \min_val_reg[0][3] ,
         \min_val_reg[0][2] , \min_val_reg[0][1] , \min_val_reg[0][0] , n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968;

  DFF \min_dist_reg_reg[0][0]  ( .D(\local_min_dist[0][0] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][0] ) );
  DFF \min_dist_reg_reg[0][1]  ( .D(\local_min_dist[0][1] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][1] ) );
  DFF \min_dist_reg_reg[0][2]  ( .D(\local_min_dist[0][2] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][2] ) );
  DFF \min_dist_reg_reg[0][3]  ( .D(\local_min_dist[0][3] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][3] ) );
  DFF \min_dist_reg_reg[0][4]  ( .D(\local_min_dist[0][4] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][4] ) );
  DFF \min_dist_reg_reg[1][0]  ( .D(\min_dist[1][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][0] ) );
  DFF \min_dist_reg_reg[1][1]  ( .D(\min_dist[1][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][1] ) );
  DFF \min_dist_reg_reg[1][2]  ( .D(\min_dist[1][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][2] ) );
  DFF \min_dist_reg_reg[1][3]  ( .D(\min_dist[1][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][3] ) );
  DFF \min_dist_reg_reg[1][4]  ( .D(\min_dist[1][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][4] ) );
  DFF \min_dist_reg_reg[2][0]  ( .D(\min_dist[2][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][0] ) );
  DFF \min_dist_reg_reg[2][1]  ( .D(\min_dist[2][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][1] ) );
  DFF \min_dist_reg_reg[2][2]  ( .D(\min_dist[2][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][2] ) );
  DFF \min_dist_reg_reg[2][3]  ( .D(\min_dist[2][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][3] ) );
  DFF \min_dist_reg_reg[2][4]  ( .D(\min_dist[2][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][4] ) );
  DFF \min_dist_reg_reg[3][0]  ( .D(\min_dist[3][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][0] ) );
  DFF \min_dist_reg_reg[3][1]  ( .D(\min_dist[3][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][1] ) );
  DFF \min_dist_reg_reg[3][2]  ( .D(\min_dist[3][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][2] ) );
  DFF \min_dist_reg_reg[3][3]  ( .D(\min_dist[3][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][3] ) );
  DFF \min_dist_reg_reg[3][4]  ( .D(\min_dist[3][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][4] ) );
  DFF \min_val_reg_reg[0][0]  ( .D(min_val_out[0]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][0] ) );
  DFF \min_val_reg_reg[0][1]  ( .D(min_val_out[1]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][1] ) );
  DFF \min_val_reg_reg[0][2]  ( .D(min_val_out[2]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][2] ) );
  DFF \min_val_reg_reg[0][3]  ( .D(min_val_out[3]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][3] ) );
  DFF \min_val_reg_reg[0][4]  ( .D(min_val_out[4]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][4] ) );
  DFF \min_val_reg_reg[0][5]  ( .D(min_val_out[5]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][5] ) );
  DFF \min_val_reg_reg[0][6]  ( .D(min_val_out[6]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][6] ) );
  DFF \min_val_reg_reg[0][7]  ( .D(min_val_out[7]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][7] ) );
  DFF \min_val_reg_reg[0][8]  ( .D(min_val_out[8]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][8] ) );
  DFF \min_val_reg_reg[0][9]  ( .D(min_val_out[9]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][9] ) );
  DFF \min_val_reg_reg[0][10]  ( .D(min_val_out[10]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][10] ) );
  DFF \min_val_reg_reg[0][11]  ( .D(min_val_out[11]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][11] ) );
  DFF \min_val_reg_reg[0][12]  ( .D(min_val_out[12]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][12] ) );
  DFF \min_val_reg_reg[0][13]  ( .D(min_val_out[13]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][13] ) );
  DFF \min_val_reg_reg[0][14]  ( .D(min_val_out[14]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][14] ) );
  DFF \min_val_reg_reg[0][15]  ( .D(min_val_out[15]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][15] ) );
  DFF \min_val_reg_reg[0][16]  ( .D(min_val_out[16]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][16] ) );
  DFF \min_val_reg_reg[0][17]  ( .D(min_val_out[17]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][17] ) );
  DFF \min_val_reg_reg[0][18]  ( .D(min_val_out[18]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][18] ) );
  DFF \min_val_reg_reg[0][19]  ( .D(min_val_out[19]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][19] ) );
  DFF \min_val_reg_reg[0][20]  ( .D(min_val_out[20]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][20] ) );
  DFF \min_val_reg_reg[0][21]  ( .D(min_val_out[21]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][21] ) );
  DFF \min_val_reg_reg[0][22]  ( .D(min_val_out[22]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][22] ) );
  DFF \min_val_reg_reg[0][23]  ( .D(min_val_out[23]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][23] ) );
  DFF \min_val_reg_reg[0][24]  ( .D(min_val_out[24]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][24] ) );
  DFF \min_val_reg_reg[0][25]  ( .D(min_val_out[25]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][25] ) );
  DFF \min_val_reg_reg[0][26]  ( .D(min_val_out[26]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][26] ) );
  DFF \min_val_reg_reg[0][27]  ( .D(min_val_out[27]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][27] ) );
  DFF \min_val_reg_reg[0][28]  ( .D(min_val_out[28]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][28] ) );
  DFF \min_val_reg_reg[0][29]  ( .D(min_val_out[29]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][29] ) );
  DFF \min_val_reg_reg[0][30]  ( .D(min_val_out[30]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][30] ) );
  DFF \min_val_reg_reg[1][0]  ( .D(min_val_out[31]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][0] ) );
  DFF \min_val_reg_reg[1][1]  ( .D(min_val_out[32]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][1] ) );
  DFF \min_val_reg_reg[1][2]  ( .D(min_val_out[33]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][2] ) );
  DFF \min_val_reg_reg[1][3]  ( .D(min_val_out[34]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][3] ) );
  DFF \min_val_reg_reg[1][4]  ( .D(min_val_out[35]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][4] ) );
  DFF \min_val_reg_reg[1][5]  ( .D(min_val_out[36]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][5] ) );
  DFF \min_val_reg_reg[1][6]  ( .D(min_val_out[37]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][6] ) );
  DFF \min_val_reg_reg[1][7]  ( .D(min_val_out[38]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][7] ) );
  DFF \min_val_reg_reg[1][8]  ( .D(min_val_out[39]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][8] ) );
  DFF \min_val_reg_reg[1][9]  ( .D(min_val_out[40]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][9] ) );
  DFF \min_val_reg_reg[1][10]  ( .D(min_val_out[41]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][10] ) );
  DFF \min_val_reg_reg[1][11]  ( .D(min_val_out[42]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][11] ) );
  DFF \min_val_reg_reg[1][12]  ( .D(min_val_out[43]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][12] ) );
  DFF \min_val_reg_reg[1][13]  ( .D(min_val_out[44]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][13] ) );
  DFF \min_val_reg_reg[1][14]  ( .D(min_val_out[45]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][14] ) );
  DFF \min_val_reg_reg[1][15]  ( .D(min_val_out[46]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][15] ) );
  DFF \min_val_reg_reg[1][16]  ( .D(min_val_out[47]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][16] ) );
  DFF \min_val_reg_reg[1][17]  ( .D(min_val_out[48]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][17] ) );
  DFF \min_val_reg_reg[1][18]  ( .D(min_val_out[49]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][18] ) );
  DFF \min_val_reg_reg[1][19]  ( .D(min_val_out[50]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][19] ) );
  DFF \min_val_reg_reg[1][20]  ( .D(min_val_out[51]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][20] ) );
  DFF \min_val_reg_reg[1][21]  ( .D(min_val_out[52]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][21] ) );
  DFF \min_val_reg_reg[1][22]  ( .D(min_val_out[53]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][22] ) );
  DFF \min_val_reg_reg[1][23]  ( .D(min_val_out[54]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][23] ) );
  DFF \min_val_reg_reg[1][24]  ( .D(min_val_out[55]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][24] ) );
  DFF \min_val_reg_reg[1][25]  ( .D(min_val_out[56]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][25] ) );
  DFF \min_val_reg_reg[1][26]  ( .D(min_val_out[57]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][26] ) );
  DFF \min_val_reg_reg[1][27]  ( .D(min_val_out[58]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][27] ) );
  DFF \min_val_reg_reg[1][28]  ( .D(min_val_out[59]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][28] ) );
  DFF \min_val_reg_reg[1][29]  ( .D(min_val_out[60]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][29] ) );
  DFF \min_val_reg_reg[1][30]  ( .D(min_val_out[61]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][30] ) );
  DFF \min_val_reg_reg[2][0]  ( .D(min_val_out[62]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][0] ) );
  DFF \min_val_reg_reg[2][1]  ( .D(min_val_out[63]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][1] ) );
  DFF \min_val_reg_reg[2][2]  ( .D(min_val_out[64]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][2] ) );
  DFF \min_val_reg_reg[2][3]  ( .D(min_val_out[65]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][3] ) );
  DFF \min_val_reg_reg[2][4]  ( .D(min_val_out[66]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][4] ) );
  DFF \min_val_reg_reg[2][5]  ( .D(min_val_out[67]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][5] ) );
  DFF \min_val_reg_reg[2][6]  ( .D(min_val_out[68]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][6] ) );
  DFF \min_val_reg_reg[2][7]  ( .D(min_val_out[69]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][7] ) );
  DFF \min_val_reg_reg[2][8]  ( .D(min_val_out[70]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][8] ) );
  DFF \min_val_reg_reg[2][9]  ( .D(min_val_out[71]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][9] ) );
  DFF \min_val_reg_reg[2][10]  ( .D(min_val_out[72]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][10] ) );
  DFF \min_val_reg_reg[2][11]  ( .D(min_val_out[73]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][11] ) );
  DFF \min_val_reg_reg[2][12]  ( .D(min_val_out[74]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][12] ) );
  DFF \min_val_reg_reg[2][13]  ( .D(min_val_out[75]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][13] ) );
  DFF \min_val_reg_reg[2][14]  ( .D(min_val_out[76]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][14] ) );
  DFF \min_val_reg_reg[2][15]  ( .D(min_val_out[77]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][15] ) );
  DFF \min_val_reg_reg[2][16]  ( .D(min_val_out[78]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][16] ) );
  DFF \min_val_reg_reg[2][17]  ( .D(min_val_out[79]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][17] ) );
  DFF \min_val_reg_reg[2][18]  ( .D(min_val_out[80]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][18] ) );
  DFF \min_val_reg_reg[2][19]  ( .D(min_val_out[81]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][19] ) );
  DFF \min_val_reg_reg[2][20]  ( .D(min_val_out[82]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][20] ) );
  DFF \min_val_reg_reg[2][21]  ( .D(min_val_out[83]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][21] ) );
  DFF \min_val_reg_reg[2][22]  ( .D(min_val_out[84]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][22] ) );
  DFF \min_val_reg_reg[2][23]  ( .D(min_val_out[85]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][23] ) );
  DFF \min_val_reg_reg[2][24]  ( .D(min_val_out[86]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][24] ) );
  DFF \min_val_reg_reg[2][25]  ( .D(min_val_out[87]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][25] ) );
  DFF \min_val_reg_reg[2][26]  ( .D(min_val_out[88]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][26] ) );
  DFF \min_val_reg_reg[2][27]  ( .D(min_val_out[89]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][27] ) );
  DFF \min_val_reg_reg[2][28]  ( .D(min_val_out[90]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][28] ) );
  DFF \min_val_reg_reg[2][29]  ( .D(min_val_out[91]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][29] ) );
  DFF \min_val_reg_reg[2][30]  ( .D(min_val_out[92]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][30] ) );
  DFF \min_val_reg_reg[3][0]  ( .D(min_val_out[93]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][0] ) );
  DFF \min_val_reg_reg[3][1]  ( .D(min_val_out[94]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][1] ) );
  DFF \min_val_reg_reg[3][2]  ( .D(min_val_out[95]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][2] ) );
  DFF \min_val_reg_reg[3][3]  ( .D(min_val_out[96]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][3] ) );
  DFF \min_val_reg_reg[3][4]  ( .D(min_val_out[97]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][4] ) );
  DFF \min_val_reg_reg[3][5]  ( .D(min_val_out[98]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][5] ) );
  DFF \min_val_reg_reg[3][6]  ( .D(min_val_out[99]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][6] ) );
  DFF \min_val_reg_reg[3][7]  ( .D(min_val_out[100]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][7] ) );
  DFF \min_val_reg_reg[3][8]  ( .D(min_val_out[101]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][8] ) );
  DFF \min_val_reg_reg[3][9]  ( .D(min_val_out[102]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][9] ) );
  DFF \min_val_reg_reg[3][10]  ( .D(min_val_out[103]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][10] ) );
  DFF \min_val_reg_reg[3][11]  ( .D(min_val_out[104]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][11] ) );
  DFF \min_val_reg_reg[3][12]  ( .D(min_val_out[105]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][12] ) );
  DFF \min_val_reg_reg[3][13]  ( .D(min_val_out[106]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][13] ) );
  DFF \min_val_reg_reg[3][14]  ( .D(min_val_out[107]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][14] ) );
  DFF \min_val_reg_reg[3][15]  ( .D(min_val_out[108]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][15] ) );
  DFF \min_val_reg_reg[3][16]  ( .D(min_val_out[109]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][16] ) );
  DFF \min_val_reg_reg[3][17]  ( .D(min_val_out[110]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][17] ) );
  DFF \min_val_reg_reg[3][18]  ( .D(min_val_out[111]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][18] ) );
  DFF \min_val_reg_reg[3][19]  ( .D(min_val_out[112]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][19] ) );
  DFF \min_val_reg_reg[3][20]  ( .D(min_val_out[113]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][20] ) );
  DFF \min_val_reg_reg[3][21]  ( .D(min_val_out[114]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][21] ) );
  DFF \min_val_reg_reg[3][22]  ( .D(min_val_out[115]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][22] ) );
  DFF \min_val_reg_reg[3][23]  ( .D(min_val_out[116]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][23] ) );
  DFF \min_val_reg_reg[3][24]  ( .D(min_val_out[117]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][24] ) );
  DFF \min_val_reg_reg[3][25]  ( .D(min_val_out[118]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][25] ) );
  DFF \min_val_reg_reg[3][26]  ( .D(min_val_out[119]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][26] ) );
  DFF \min_val_reg_reg[3][27]  ( .D(min_val_out[120]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][27] ) );
  DFF \min_val_reg_reg[3][28]  ( .D(min_val_out[121]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][28] ) );
  DFF \min_val_reg_reg[3][29]  ( .D(min_val_out[122]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][29] ) );
  DFF \min_val_reg_reg[3][30]  ( .D(min_val_out[123]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][30] ) );
  XOR U178 ( .A(\min_val_reg[0][9] ), .B(n145), .Z(min_val_out[9]) );
  AND U179 ( .A(n146), .B(n147), .Z(n145) );
  XNOR U180 ( .A(n148), .B(n149), .Z(min_val_out[99]) );
  AND U181 ( .A(n150), .B(n151), .Z(n148) );
  XNOR U182 ( .A(n152), .B(n153), .Z(min_val_out[98]) );
  AND U183 ( .A(n150), .B(n154), .Z(n152) );
  XNOR U184 ( .A(n155), .B(n156), .Z(min_val_out[97]) );
  AND U185 ( .A(n150), .B(n157), .Z(n155) );
  XNOR U186 ( .A(n158), .B(n159), .Z(min_val_out[96]) );
  AND U187 ( .A(n150), .B(n160), .Z(n158) );
  XNOR U188 ( .A(n161), .B(n162), .Z(min_val_out[95]) );
  AND U189 ( .A(n150), .B(n163), .Z(n161) );
  XNOR U190 ( .A(n164), .B(n165), .Z(min_val_out[94]) );
  AND U191 ( .A(n150), .B(n166), .Z(n164) );
  XNOR U192 ( .A(n167), .B(n168), .Z(min_val_out[93]) );
  AND U193 ( .A(n150), .B(n169), .Z(n167) );
  XOR U194 ( .A(n170), .B(n171), .Z(min_val_out[92]) );
  AND U195 ( .A(n172), .B(n173), .Z(n170) );
  XOR U196 ( .A(n174), .B(n175), .Z(min_val_out[91]) );
  AND U197 ( .A(n172), .B(n176), .Z(n174) );
  XOR U198 ( .A(n177), .B(n178), .Z(min_val_out[90]) );
  AND U199 ( .A(n172), .B(n179), .Z(n177) );
  XOR U200 ( .A(\min_val_reg[0][8] ), .B(n180), .Z(min_val_out[8]) );
  AND U201 ( .A(n146), .B(n181), .Z(n180) );
  XOR U202 ( .A(n182), .B(n183), .Z(min_val_out[89]) );
  AND U203 ( .A(n172), .B(n184), .Z(n182) );
  XOR U204 ( .A(n185), .B(n186), .Z(min_val_out[88]) );
  AND U205 ( .A(n172), .B(n187), .Z(n185) );
  XOR U206 ( .A(n188), .B(n189), .Z(min_val_out[87]) );
  AND U207 ( .A(n172), .B(n190), .Z(n188) );
  XOR U208 ( .A(n191), .B(n192), .Z(min_val_out[86]) );
  AND U209 ( .A(n172), .B(n193), .Z(n191) );
  XOR U210 ( .A(n194), .B(n195), .Z(min_val_out[85]) );
  AND U211 ( .A(n172), .B(n196), .Z(n194) );
  XOR U212 ( .A(n197), .B(n198), .Z(min_val_out[84]) );
  AND U213 ( .A(n172), .B(n199), .Z(n197) );
  XOR U214 ( .A(n200), .B(n201), .Z(min_val_out[83]) );
  AND U215 ( .A(n172), .B(n202), .Z(n200) );
  XOR U216 ( .A(n203), .B(n204), .Z(min_val_out[82]) );
  AND U217 ( .A(n172), .B(n205), .Z(n203) );
  XOR U218 ( .A(n206), .B(n207), .Z(min_val_out[81]) );
  AND U219 ( .A(n172), .B(n208), .Z(n206) );
  XOR U220 ( .A(n209), .B(n210), .Z(min_val_out[80]) );
  AND U221 ( .A(n172), .B(n211), .Z(n209) );
  XOR U222 ( .A(\min_val_reg[0][7] ), .B(n212), .Z(min_val_out[7]) );
  AND U223 ( .A(n146), .B(n213), .Z(n212) );
  XOR U224 ( .A(n214), .B(n215), .Z(min_val_out[79]) );
  AND U225 ( .A(n172), .B(n216), .Z(n214) );
  XOR U226 ( .A(n217), .B(n218), .Z(min_val_out[78]) );
  AND U227 ( .A(n172), .B(n219), .Z(n217) );
  XOR U228 ( .A(n220), .B(n221), .Z(min_val_out[77]) );
  AND U229 ( .A(n172), .B(n222), .Z(n220) );
  XOR U230 ( .A(n223), .B(n224), .Z(min_val_out[76]) );
  AND U231 ( .A(n172), .B(n225), .Z(n223) );
  XOR U232 ( .A(n226), .B(n227), .Z(min_val_out[75]) );
  AND U233 ( .A(n172), .B(n228), .Z(n226) );
  XOR U234 ( .A(n229), .B(n230), .Z(min_val_out[74]) );
  AND U235 ( .A(n172), .B(n231), .Z(n229) );
  XOR U236 ( .A(n232), .B(n233), .Z(min_val_out[73]) );
  AND U237 ( .A(n172), .B(n234), .Z(n232) );
  XOR U238 ( .A(n235), .B(n236), .Z(min_val_out[72]) );
  AND U239 ( .A(n172), .B(n237), .Z(n235) );
  XOR U240 ( .A(n238), .B(n239), .Z(min_val_out[71]) );
  AND U241 ( .A(n172), .B(n240), .Z(n238) );
  XOR U242 ( .A(n241), .B(n242), .Z(min_val_out[70]) );
  AND U243 ( .A(n172), .B(n243), .Z(n241) );
  XOR U244 ( .A(\min_val_reg[0][6] ), .B(n244), .Z(min_val_out[6]) );
  AND U245 ( .A(n146), .B(n245), .Z(n244) );
  XOR U246 ( .A(n246), .B(n247), .Z(min_val_out[69]) );
  AND U247 ( .A(n172), .B(n248), .Z(n246) );
  XNOR U248 ( .A(n249), .B(n250), .Z(min_val_out[68]) );
  AND U249 ( .A(n172), .B(n251), .Z(n249) );
  XNOR U250 ( .A(n252), .B(n253), .Z(min_val_out[67]) );
  AND U251 ( .A(n172), .B(n254), .Z(n252) );
  XNOR U252 ( .A(n255), .B(n256), .Z(min_val_out[66]) );
  AND U253 ( .A(n172), .B(n257), .Z(n255) );
  XNOR U254 ( .A(n258), .B(n259), .Z(min_val_out[65]) );
  AND U255 ( .A(n172), .B(n260), .Z(n258) );
  XNOR U256 ( .A(n261), .B(n262), .Z(min_val_out[64]) );
  AND U257 ( .A(n172), .B(n263), .Z(n261) );
  XNOR U258 ( .A(n264), .B(n265), .Z(min_val_out[63]) );
  AND U259 ( .A(n172), .B(n266), .Z(n264) );
  XNOR U260 ( .A(n267), .B(n268), .Z(min_val_out[62]) );
  AND U261 ( .A(n172), .B(n269), .Z(n267) );
  XNOR U262 ( .A(n270), .B(n271), .Z(min_val_out[61]) );
  AND U263 ( .A(n272), .B(n273), .Z(n270) );
  XNOR U264 ( .A(n274), .B(n275), .Z(min_val_out[60]) );
  AND U265 ( .A(n272), .B(n276), .Z(n274) );
  XOR U266 ( .A(\min_val_reg[0][5] ), .B(n277), .Z(min_val_out[5]) );
  AND U267 ( .A(n146), .B(n278), .Z(n277) );
  XNOR U268 ( .A(n279), .B(n280), .Z(min_val_out[59]) );
  AND U269 ( .A(n272), .B(n281), .Z(n279) );
  XNOR U270 ( .A(n282), .B(n283), .Z(min_val_out[58]) );
  AND U271 ( .A(n272), .B(n284), .Z(n282) );
  XNOR U272 ( .A(n285), .B(n286), .Z(min_val_out[57]) );
  AND U273 ( .A(n272), .B(n287), .Z(n285) );
  XNOR U274 ( .A(n288), .B(n289), .Z(min_val_out[56]) );
  AND U275 ( .A(n272), .B(n290), .Z(n288) );
  XNOR U276 ( .A(n291), .B(n292), .Z(min_val_out[55]) );
  AND U277 ( .A(n272), .B(n293), .Z(n291) );
  XNOR U278 ( .A(n294), .B(n295), .Z(min_val_out[54]) );
  AND U279 ( .A(n272), .B(n296), .Z(n294) );
  XNOR U280 ( .A(n297), .B(n298), .Z(min_val_out[53]) );
  AND U281 ( .A(n272), .B(n299), .Z(n297) );
  XNOR U282 ( .A(n300), .B(n301), .Z(min_val_out[52]) );
  AND U283 ( .A(n272), .B(n302), .Z(n300) );
  XNOR U284 ( .A(n303), .B(n304), .Z(min_val_out[51]) );
  AND U285 ( .A(n272), .B(n305), .Z(n303) );
  XNOR U286 ( .A(n306), .B(n307), .Z(min_val_out[50]) );
  AND U287 ( .A(n272), .B(n308), .Z(n306) );
  XOR U288 ( .A(\min_val_reg[0][4] ), .B(n309), .Z(min_val_out[4]) );
  AND U289 ( .A(n146), .B(n310), .Z(n309) );
  XNOR U290 ( .A(n311), .B(n312), .Z(min_val_out[49]) );
  AND U291 ( .A(n272), .B(n313), .Z(n311) );
  XNOR U292 ( .A(n314), .B(n315), .Z(min_val_out[48]) );
  AND U293 ( .A(n272), .B(n316), .Z(n314) );
  XNOR U294 ( .A(n317), .B(n318), .Z(min_val_out[47]) );
  AND U295 ( .A(n272), .B(n319), .Z(n317) );
  XNOR U296 ( .A(n320), .B(n321), .Z(min_val_out[46]) );
  AND U297 ( .A(n272), .B(n322), .Z(n320) );
  XNOR U298 ( .A(n323), .B(n324), .Z(min_val_out[45]) );
  AND U299 ( .A(n272), .B(n325), .Z(n323) );
  XNOR U300 ( .A(n326), .B(n327), .Z(min_val_out[44]) );
  AND U301 ( .A(n272), .B(n328), .Z(n326) );
  XNOR U302 ( .A(n329), .B(n330), .Z(min_val_out[43]) );
  AND U303 ( .A(n272), .B(n331), .Z(n329) );
  XNOR U304 ( .A(n332), .B(n333), .Z(min_val_out[42]) );
  AND U305 ( .A(n272), .B(n334), .Z(n332) );
  XNOR U306 ( .A(n335), .B(n336), .Z(min_val_out[41]) );
  AND U307 ( .A(n272), .B(n337), .Z(n335) );
  XOR U308 ( .A(n338), .B(n339), .Z(min_val_out[40]) );
  AND U309 ( .A(n272), .B(n147), .Z(n338) );
  XOR U310 ( .A(\min_val_reg[0][9] ), .B(n339), .Z(n147) );
  XNOR U311 ( .A(\min_val_reg[1][9] ), .B(n340), .Z(n339) );
  NAND U312 ( .A(n240), .B(n172), .Z(n340) );
  XOR U313 ( .A(\min_val_reg[1][9] ), .B(n239), .Z(n240) );
  XNOR U314 ( .A(\min_val_reg[2][9] ), .B(n341), .Z(n239) );
  NAND U315 ( .A(n342), .B(n343), .Z(n341) );
  XOR U316 ( .A(\min_val_reg[0][3] ), .B(n344), .Z(min_val_out[3]) );
  AND U317 ( .A(n146), .B(n345), .Z(n344) );
  XOR U318 ( .A(n346), .B(n347), .Z(min_val_out[39]) );
  AND U319 ( .A(n272), .B(n181), .Z(n346) );
  XOR U320 ( .A(\min_val_reg[0][8] ), .B(n347), .Z(n181) );
  XNOR U321 ( .A(\min_val_reg[1][8] ), .B(n348), .Z(n347) );
  NAND U322 ( .A(n243), .B(n172), .Z(n348) );
  XOR U323 ( .A(\min_val_reg[1][8] ), .B(n242), .Z(n243) );
  XNOR U324 ( .A(\min_val_reg[2][8] ), .B(n349), .Z(n242) );
  NAND U325 ( .A(n350), .B(n343), .Z(n349) );
  XOR U326 ( .A(n351), .B(n352), .Z(min_val_out[38]) );
  AND U327 ( .A(n272), .B(n213), .Z(n351) );
  XOR U328 ( .A(\min_val_reg[0][7] ), .B(n352), .Z(n213) );
  XNOR U329 ( .A(\min_val_reg[1][7] ), .B(n353), .Z(n352) );
  NAND U330 ( .A(n248), .B(n172), .Z(n353) );
  XOR U331 ( .A(\min_val_reg[1][7] ), .B(n247), .Z(n248) );
  XNOR U332 ( .A(\min_val_reg[2][7] ), .B(n354), .Z(n247) );
  NAND U333 ( .A(n355), .B(n343), .Z(n354) );
  XOR U334 ( .A(n356), .B(n357), .Z(min_val_out[37]) );
  AND U335 ( .A(n272), .B(n245), .Z(n356) );
  XOR U336 ( .A(\min_val_reg[0][6] ), .B(n357), .Z(n245) );
  XNOR U337 ( .A(\min_val_reg[1][6] ), .B(n358), .Z(n357) );
  NAND U338 ( .A(n251), .B(n172), .Z(n358) );
  XNOR U339 ( .A(\min_val_reg[1][6] ), .B(n250), .Z(n251) );
  XOR U340 ( .A(\min_val_reg[2][6] ), .B(n359), .Z(n250) );
  NAND U341 ( .A(n151), .B(n343), .Z(n359) );
  XNOR U342 ( .A(\min_val_reg[2][6] ), .B(n149), .Z(n151) );
  XOR U343 ( .A(\min_val_reg[3][6] ), .B(n360), .Z(n149) );
  NAND U344 ( .A(n361), .B(n362), .Z(n360) );
  XOR U345 ( .A(\min_val_reg[3][6] ), .B(DB[6]), .Z(n361) );
  XNOR U346 ( .A(n363), .B(n364), .Z(min_val_out[36]) );
  AND U347 ( .A(n272), .B(n278), .Z(n363) );
  XNOR U348 ( .A(\min_val_reg[0][5] ), .B(n364), .Z(n278) );
  XOR U349 ( .A(\min_val_reg[1][5] ), .B(n365), .Z(n364) );
  NAND U350 ( .A(n254), .B(n172), .Z(n365) );
  XNOR U351 ( .A(\min_val_reg[1][5] ), .B(n253), .Z(n254) );
  XOR U352 ( .A(\min_val_reg[2][5] ), .B(n366), .Z(n253) );
  NAND U353 ( .A(n154), .B(n343), .Z(n366) );
  XNOR U354 ( .A(\min_val_reg[2][5] ), .B(n153), .Z(n154) );
  XOR U355 ( .A(\min_val_reg[3][5] ), .B(n367), .Z(n153) );
  NAND U356 ( .A(n368), .B(n362), .Z(n367) );
  XOR U357 ( .A(\min_val_reg[3][5] ), .B(DB[5]), .Z(n368) );
  XNOR U358 ( .A(n369), .B(n370), .Z(min_val_out[35]) );
  AND U359 ( .A(n272), .B(n310), .Z(n369) );
  XNOR U360 ( .A(\min_val_reg[0][4] ), .B(n370), .Z(n310) );
  XOR U361 ( .A(\min_val_reg[1][4] ), .B(n371), .Z(n370) );
  NAND U362 ( .A(n257), .B(n172), .Z(n371) );
  XNOR U363 ( .A(\min_val_reg[1][4] ), .B(n256), .Z(n257) );
  XOR U364 ( .A(\min_val_reg[2][4] ), .B(n372), .Z(n256) );
  NAND U365 ( .A(n157), .B(n343), .Z(n372) );
  XNOR U366 ( .A(\min_val_reg[2][4] ), .B(n156), .Z(n157) );
  XOR U367 ( .A(\min_val_reg[3][4] ), .B(n373), .Z(n156) );
  NAND U368 ( .A(n374), .B(n362), .Z(n373) );
  XOR U369 ( .A(\min_val_reg[3][4] ), .B(DB[4]), .Z(n374) );
  XNOR U370 ( .A(n375), .B(n376), .Z(min_val_out[34]) );
  AND U371 ( .A(n272), .B(n345), .Z(n375) );
  XNOR U372 ( .A(\min_val_reg[0][3] ), .B(n376), .Z(n345) );
  XOR U373 ( .A(\min_val_reg[1][3] ), .B(n377), .Z(n376) );
  NAND U374 ( .A(n260), .B(n172), .Z(n377) );
  XNOR U375 ( .A(\min_val_reg[1][3] ), .B(n259), .Z(n260) );
  XOR U376 ( .A(\min_val_reg[2][3] ), .B(n378), .Z(n259) );
  NAND U377 ( .A(n160), .B(n343), .Z(n378) );
  XNOR U378 ( .A(\min_val_reg[2][3] ), .B(n159), .Z(n160) );
  XOR U379 ( .A(\min_val_reg[3][3] ), .B(n379), .Z(n159) );
  NAND U380 ( .A(n380), .B(n362), .Z(n379) );
  XOR U381 ( .A(\min_val_reg[3][3] ), .B(DB[3]), .Z(n380) );
  XNOR U382 ( .A(n381), .B(n382), .Z(min_val_out[33]) );
  AND U383 ( .A(n272), .B(n383), .Z(n381) );
  XNOR U384 ( .A(n384), .B(n385), .Z(min_val_out[32]) );
  AND U385 ( .A(n272), .B(n386), .Z(n384) );
  XNOR U386 ( .A(n387), .B(n388), .Z(min_val_out[31]) );
  AND U387 ( .A(n272), .B(n389), .Z(n387) );
  XOR U388 ( .A(\min_val_reg[0][30] ), .B(n390), .Z(min_val_out[30]) );
  AND U389 ( .A(n146), .B(n273), .Z(n390) );
  XNOR U390 ( .A(\min_val_reg[0][30] ), .B(n271), .Z(n273) );
  XOR U391 ( .A(\min_val_reg[1][30] ), .B(n391), .Z(n271) );
  NAND U392 ( .A(n173), .B(n172), .Z(n391) );
  XOR U393 ( .A(\min_val_reg[1][30] ), .B(n171), .Z(n173) );
  XNOR U394 ( .A(\min_val_reg[2][30] ), .B(n392), .Z(n171) );
  NAND U395 ( .A(n393), .B(n343), .Z(n392) );
  XOR U396 ( .A(\min_val_reg[0][2] ), .B(n394), .Z(min_val_out[2]) );
  AND U397 ( .A(n146), .B(n383), .Z(n394) );
  XNOR U398 ( .A(\min_val_reg[0][2] ), .B(n382), .Z(n383) );
  XOR U399 ( .A(\min_val_reg[1][2] ), .B(n395), .Z(n382) );
  NAND U400 ( .A(n263), .B(n172), .Z(n395) );
  XNOR U401 ( .A(\min_val_reg[1][2] ), .B(n262), .Z(n263) );
  XOR U402 ( .A(\min_val_reg[2][2] ), .B(n396), .Z(n262) );
  NAND U403 ( .A(n163), .B(n343), .Z(n396) );
  XNOR U404 ( .A(\min_val_reg[2][2] ), .B(n162), .Z(n163) );
  XOR U405 ( .A(\min_val_reg[3][2] ), .B(n397), .Z(n162) );
  NAND U406 ( .A(n398), .B(n362), .Z(n397) );
  XOR U407 ( .A(\min_val_reg[3][2] ), .B(DB[2]), .Z(n398) );
  XOR U408 ( .A(\min_val_reg[0][29] ), .B(n399), .Z(min_val_out[29]) );
  AND U409 ( .A(n146), .B(n276), .Z(n399) );
  XNOR U410 ( .A(\min_val_reg[0][29] ), .B(n275), .Z(n276) );
  XOR U411 ( .A(\min_val_reg[1][29] ), .B(n400), .Z(n275) );
  NAND U412 ( .A(n176), .B(n172), .Z(n400) );
  XOR U413 ( .A(\min_val_reg[1][29] ), .B(n175), .Z(n176) );
  XNOR U414 ( .A(\min_val_reg[2][29] ), .B(n401), .Z(n175) );
  NAND U415 ( .A(n402), .B(n343), .Z(n401) );
  XOR U416 ( .A(\min_val_reg[0][28] ), .B(n403), .Z(min_val_out[28]) );
  AND U417 ( .A(n146), .B(n281), .Z(n403) );
  XNOR U418 ( .A(\min_val_reg[0][28] ), .B(n280), .Z(n281) );
  XOR U419 ( .A(\min_val_reg[1][28] ), .B(n404), .Z(n280) );
  NAND U420 ( .A(n179), .B(n172), .Z(n404) );
  XOR U421 ( .A(\min_val_reg[1][28] ), .B(n178), .Z(n179) );
  XNOR U422 ( .A(\min_val_reg[2][28] ), .B(n405), .Z(n178) );
  NAND U423 ( .A(n406), .B(n343), .Z(n405) );
  XOR U424 ( .A(\min_val_reg[0][27] ), .B(n407), .Z(min_val_out[27]) );
  AND U425 ( .A(n146), .B(n284), .Z(n407) );
  XNOR U426 ( .A(\min_val_reg[0][27] ), .B(n283), .Z(n284) );
  XOR U427 ( .A(\min_val_reg[1][27] ), .B(n408), .Z(n283) );
  NAND U428 ( .A(n184), .B(n172), .Z(n408) );
  XOR U429 ( .A(\min_val_reg[1][27] ), .B(n183), .Z(n184) );
  XNOR U430 ( .A(\min_val_reg[2][27] ), .B(n409), .Z(n183) );
  NAND U431 ( .A(n410), .B(n343), .Z(n409) );
  XOR U432 ( .A(\min_val_reg[0][26] ), .B(n411), .Z(min_val_out[26]) );
  AND U433 ( .A(n146), .B(n287), .Z(n411) );
  XNOR U434 ( .A(\min_val_reg[0][26] ), .B(n286), .Z(n287) );
  XOR U435 ( .A(\min_val_reg[1][26] ), .B(n412), .Z(n286) );
  NAND U436 ( .A(n187), .B(n172), .Z(n412) );
  XOR U437 ( .A(\min_val_reg[1][26] ), .B(n186), .Z(n187) );
  XNOR U438 ( .A(\min_val_reg[2][26] ), .B(n413), .Z(n186) );
  NAND U439 ( .A(n414), .B(n343), .Z(n413) );
  XOR U440 ( .A(\min_val_reg[0][25] ), .B(n415), .Z(min_val_out[25]) );
  AND U441 ( .A(n146), .B(n290), .Z(n415) );
  XNOR U442 ( .A(\min_val_reg[0][25] ), .B(n289), .Z(n290) );
  XOR U443 ( .A(\min_val_reg[1][25] ), .B(n416), .Z(n289) );
  NAND U444 ( .A(n190), .B(n172), .Z(n416) );
  XOR U445 ( .A(\min_val_reg[1][25] ), .B(n189), .Z(n190) );
  XNOR U446 ( .A(\min_val_reg[2][25] ), .B(n417), .Z(n189) );
  NAND U447 ( .A(n418), .B(n343), .Z(n417) );
  XOR U448 ( .A(\min_val_reg[0][24] ), .B(n419), .Z(min_val_out[24]) );
  AND U449 ( .A(n146), .B(n293), .Z(n419) );
  XNOR U450 ( .A(\min_val_reg[0][24] ), .B(n292), .Z(n293) );
  XOR U451 ( .A(\min_val_reg[1][24] ), .B(n420), .Z(n292) );
  NAND U452 ( .A(n193), .B(n172), .Z(n420) );
  XOR U453 ( .A(\min_val_reg[1][24] ), .B(n192), .Z(n193) );
  XNOR U454 ( .A(\min_val_reg[2][24] ), .B(n421), .Z(n192) );
  NAND U455 ( .A(n422), .B(n343), .Z(n421) );
  XOR U456 ( .A(\min_val_reg[0][23] ), .B(n423), .Z(min_val_out[23]) );
  AND U457 ( .A(n146), .B(n296), .Z(n423) );
  XNOR U458 ( .A(\min_val_reg[0][23] ), .B(n295), .Z(n296) );
  XOR U459 ( .A(\min_val_reg[1][23] ), .B(n424), .Z(n295) );
  NAND U460 ( .A(n196), .B(n172), .Z(n424) );
  XOR U461 ( .A(\min_val_reg[1][23] ), .B(n195), .Z(n196) );
  XNOR U462 ( .A(\min_val_reg[2][23] ), .B(n425), .Z(n195) );
  NAND U463 ( .A(n426), .B(n343), .Z(n425) );
  XOR U464 ( .A(\min_val_reg[0][22] ), .B(n427), .Z(min_val_out[22]) );
  AND U465 ( .A(n146), .B(n299), .Z(n427) );
  XNOR U466 ( .A(\min_val_reg[0][22] ), .B(n298), .Z(n299) );
  XOR U467 ( .A(\min_val_reg[1][22] ), .B(n428), .Z(n298) );
  NAND U468 ( .A(n199), .B(n172), .Z(n428) );
  XOR U469 ( .A(\min_val_reg[1][22] ), .B(n198), .Z(n199) );
  XNOR U470 ( .A(\min_val_reg[2][22] ), .B(n429), .Z(n198) );
  NAND U471 ( .A(n430), .B(n343), .Z(n429) );
  XOR U472 ( .A(\min_val_reg[0][21] ), .B(n431), .Z(min_val_out[21]) );
  AND U473 ( .A(n146), .B(n302), .Z(n431) );
  XNOR U474 ( .A(\min_val_reg[0][21] ), .B(n301), .Z(n302) );
  XOR U475 ( .A(\min_val_reg[1][21] ), .B(n432), .Z(n301) );
  NAND U476 ( .A(n202), .B(n172), .Z(n432) );
  XOR U477 ( .A(\min_val_reg[1][21] ), .B(n201), .Z(n202) );
  XNOR U478 ( .A(\min_val_reg[2][21] ), .B(n433), .Z(n201) );
  NAND U479 ( .A(n434), .B(n343), .Z(n433) );
  XOR U480 ( .A(\min_val_reg[0][20] ), .B(n435), .Z(min_val_out[20]) );
  AND U481 ( .A(n146), .B(n305), .Z(n435) );
  XNOR U482 ( .A(\min_val_reg[0][20] ), .B(n304), .Z(n305) );
  XOR U483 ( .A(\min_val_reg[1][20] ), .B(n436), .Z(n304) );
  NAND U484 ( .A(n205), .B(n172), .Z(n436) );
  XOR U485 ( .A(\min_val_reg[1][20] ), .B(n204), .Z(n205) );
  XNOR U486 ( .A(\min_val_reg[2][20] ), .B(n437), .Z(n204) );
  NAND U487 ( .A(n438), .B(n343), .Z(n437) );
  XOR U488 ( .A(\min_val_reg[0][1] ), .B(n439), .Z(min_val_out[1]) );
  AND U489 ( .A(n146), .B(n386), .Z(n439) );
  XNOR U490 ( .A(\min_val_reg[0][1] ), .B(n385), .Z(n386) );
  XOR U491 ( .A(\min_val_reg[1][1] ), .B(n440), .Z(n385) );
  NAND U492 ( .A(n266), .B(n172), .Z(n440) );
  XNOR U493 ( .A(\min_val_reg[1][1] ), .B(n265), .Z(n266) );
  XOR U494 ( .A(\min_val_reg[2][1] ), .B(n441), .Z(n265) );
  NAND U495 ( .A(n166), .B(n343), .Z(n441) );
  XNOR U496 ( .A(\min_val_reg[2][1] ), .B(n165), .Z(n166) );
  XOR U497 ( .A(\min_val_reg[3][1] ), .B(n442), .Z(n165) );
  NAND U498 ( .A(n443), .B(n362), .Z(n442) );
  XOR U499 ( .A(\min_val_reg[3][1] ), .B(DB[1]), .Z(n443) );
  XOR U500 ( .A(\min_val_reg[0][19] ), .B(n444), .Z(min_val_out[19]) );
  AND U501 ( .A(n146), .B(n308), .Z(n444) );
  XNOR U502 ( .A(\min_val_reg[0][19] ), .B(n307), .Z(n308) );
  XOR U503 ( .A(\min_val_reg[1][19] ), .B(n445), .Z(n307) );
  NAND U504 ( .A(n208), .B(n172), .Z(n445) );
  XOR U505 ( .A(\min_val_reg[1][19] ), .B(n207), .Z(n208) );
  XNOR U506 ( .A(\min_val_reg[2][19] ), .B(n446), .Z(n207) );
  NAND U507 ( .A(n447), .B(n343), .Z(n446) );
  XOR U508 ( .A(\min_val_reg[0][18] ), .B(n448), .Z(min_val_out[18]) );
  AND U509 ( .A(n146), .B(n313), .Z(n448) );
  XNOR U510 ( .A(\min_val_reg[0][18] ), .B(n312), .Z(n313) );
  XOR U511 ( .A(\min_val_reg[1][18] ), .B(n449), .Z(n312) );
  NAND U512 ( .A(n211), .B(n172), .Z(n449) );
  XOR U513 ( .A(\min_val_reg[1][18] ), .B(n210), .Z(n211) );
  XNOR U514 ( .A(\min_val_reg[2][18] ), .B(n450), .Z(n210) );
  NAND U515 ( .A(n451), .B(n343), .Z(n450) );
  XOR U516 ( .A(\min_val_reg[0][17] ), .B(n452), .Z(min_val_out[17]) );
  AND U517 ( .A(n146), .B(n316), .Z(n452) );
  XNOR U518 ( .A(\min_val_reg[0][17] ), .B(n315), .Z(n316) );
  XOR U519 ( .A(\min_val_reg[1][17] ), .B(n453), .Z(n315) );
  NAND U520 ( .A(n216), .B(n172), .Z(n453) );
  XOR U521 ( .A(\min_val_reg[1][17] ), .B(n215), .Z(n216) );
  XNOR U522 ( .A(\min_val_reg[2][17] ), .B(n454), .Z(n215) );
  NAND U523 ( .A(n455), .B(n343), .Z(n454) );
  XOR U524 ( .A(\min_val_reg[0][16] ), .B(n456), .Z(min_val_out[16]) );
  AND U525 ( .A(n146), .B(n319), .Z(n456) );
  XNOR U526 ( .A(\min_val_reg[0][16] ), .B(n318), .Z(n319) );
  XOR U527 ( .A(\min_val_reg[1][16] ), .B(n457), .Z(n318) );
  NAND U528 ( .A(n219), .B(n172), .Z(n457) );
  XOR U529 ( .A(\min_val_reg[1][16] ), .B(n218), .Z(n219) );
  XNOR U530 ( .A(\min_val_reg[2][16] ), .B(n458), .Z(n218) );
  NAND U531 ( .A(n459), .B(n343), .Z(n458) );
  XOR U532 ( .A(\min_val_reg[0][15] ), .B(n460), .Z(min_val_out[15]) );
  AND U533 ( .A(n146), .B(n322), .Z(n460) );
  XNOR U534 ( .A(\min_val_reg[0][15] ), .B(n321), .Z(n322) );
  XOR U535 ( .A(\min_val_reg[1][15] ), .B(n461), .Z(n321) );
  NAND U536 ( .A(n222), .B(n172), .Z(n461) );
  XOR U537 ( .A(\min_val_reg[1][15] ), .B(n221), .Z(n222) );
  XNOR U538 ( .A(\min_val_reg[2][15] ), .B(n462), .Z(n221) );
  NAND U539 ( .A(n463), .B(n343), .Z(n462) );
  XOR U540 ( .A(\min_val_reg[0][14] ), .B(n464), .Z(min_val_out[14]) );
  AND U541 ( .A(n146), .B(n325), .Z(n464) );
  XNOR U542 ( .A(\min_val_reg[0][14] ), .B(n324), .Z(n325) );
  XOR U543 ( .A(\min_val_reg[1][14] ), .B(n465), .Z(n324) );
  NAND U544 ( .A(n225), .B(n172), .Z(n465) );
  XOR U545 ( .A(\min_val_reg[1][14] ), .B(n224), .Z(n225) );
  XNOR U546 ( .A(\min_val_reg[2][14] ), .B(n466), .Z(n224) );
  NAND U547 ( .A(n467), .B(n343), .Z(n466) );
  XOR U548 ( .A(\min_val_reg[0][13] ), .B(n468), .Z(min_val_out[13]) );
  AND U549 ( .A(n146), .B(n328), .Z(n468) );
  XNOR U550 ( .A(\min_val_reg[0][13] ), .B(n327), .Z(n328) );
  XOR U551 ( .A(\min_val_reg[1][13] ), .B(n469), .Z(n327) );
  NAND U552 ( .A(n228), .B(n172), .Z(n469) );
  XOR U553 ( .A(\min_val_reg[1][13] ), .B(n227), .Z(n228) );
  XNOR U554 ( .A(\min_val_reg[2][13] ), .B(n470), .Z(n227) );
  NAND U555 ( .A(n471), .B(n343), .Z(n470) );
  XOR U556 ( .A(\min_val_reg[0][12] ), .B(n472), .Z(min_val_out[12]) );
  AND U557 ( .A(n146), .B(n331), .Z(n472) );
  XNOR U558 ( .A(\min_val_reg[0][12] ), .B(n330), .Z(n331) );
  XOR U559 ( .A(\min_val_reg[1][12] ), .B(n473), .Z(n330) );
  NAND U560 ( .A(n231), .B(n172), .Z(n473) );
  XOR U561 ( .A(\min_val_reg[1][12] ), .B(n230), .Z(n231) );
  XNOR U562 ( .A(\min_val_reg[2][12] ), .B(n474), .Z(n230) );
  NAND U563 ( .A(n475), .B(n343), .Z(n474) );
  XNOR U564 ( .A(n476), .B(n477), .Z(min_val_out[123]) );
  AND U565 ( .A(n150), .B(n393), .Z(n476) );
  XNOR U566 ( .A(\min_val_reg[2][30] ), .B(n477), .Z(n393) );
  XOR U567 ( .A(\min_val_reg[3][30] ), .B(n478), .Z(n477) );
  NAND U568 ( .A(n479), .B(n362), .Z(n478) );
  XOR U569 ( .A(\min_val_reg[3][30] ), .B(DB[30]), .Z(n479) );
  XNOR U570 ( .A(n480), .B(n481), .Z(min_val_out[122]) );
  AND U571 ( .A(n150), .B(n402), .Z(n480) );
  XNOR U572 ( .A(\min_val_reg[2][29] ), .B(n481), .Z(n402) );
  XOR U573 ( .A(\min_val_reg[3][29] ), .B(n482), .Z(n481) );
  NAND U574 ( .A(n483), .B(n362), .Z(n482) );
  XOR U575 ( .A(\min_val_reg[3][29] ), .B(DB[29]), .Z(n483) );
  XNOR U576 ( .A(n484), .B(n485), .Z(min_val_out[121]) );
  AND U577 ( .A(n150), .B(n406), .Z(n484) );
  XNOR U578 ( .A(\min_val_reg[2][28] ), .B(n485), .Z(n406) );
  XOR U579 ( .A(\min_val_reg[3][28] ), .B(n486), .Z(n485) );
  NAND U580 ( .A(n487), .B(n362), .Z(n486) );
  XOR U581 ( .A(\min_val_reg[3][28] ), .B(DB[28]), .Z(n487) );
  XNOR U582 ( .A(n488), .B(n489), .Z(min_val_out[120]) );
  AND U583 ( .A(n150), .B(n410), .Z(n488) );
  XNOR U584 ( .A(\min_val_reg[2][27] ), .B(n489), .Z(n410) );
  XOR U585 ( .A(\min_val_reg[3][27] ), .B(n490), .Z(n489) );
  NAND U586 ( .A(n491), .B(n362), .Z(n490) );
  XOR U587 ( .A(\min_val_reg[3][27] ), .B(DB[27]), .Z(n491) );
  XOR U588 ( .A(\min_val_reg[0][11] ), .B(n492), .Z(min_val_out[11]) );
  AND U589 ( .A(n146), .B(n334), .Z(n492) );
  XNOR U590 ( .A(\min_val_reg[0][11] ), .B(n333), .Z(n334) );
  XOR U591 ( .A(\min_val_reg[1][11] ), .B(n493), .Z(n333) );
  NAND U592 ( .A(n234), .B(n172), .Z(n493) );
  XOR U593 ( .A(\min_val_reg[1][11] ), .B(n233), .Z(n234) );
  XNOR U594 ( .A(\min_val_reg[2][11] ), .B(n494), .Z(n233) );
  NAND U595 ( .A(n495), .B(n343), .Z(n494) );
  XNOR U596 ( .A(n496), .B(n497), .Z(min_val_out[119]) );
  AND U597 ( .A(n150), .B(n414), .Z(n496) );
  XNOR U598 ( .A(\min_val_reg[2][26] ), .B(n497), .Z(n414) );
  XOR U599 ( .A(\min_val_reg[3][26] ), .B(n498), .Z(n497) );
  NAND U600 ( .A(n499), .B(n362), .Z(n498) );
  XOR U601 ( .A(\min_val_reg[3][26] ), .B(DB[26]), .Z(n499) );
  XNOR U602 ( .A(n500), .B(n501), .Z(min_val_out[118]) );
  AND U603 ( .A(n150), .B(n418), .Z(n500) );
  XNOR U604 ( .A(\min_val_reg[2][25] ), .B(n501), .Z(n418) );
  XOR U605 ( .A(\min_val_reg[3][25] ), .B(n502), .Z(n501) );
  NAND U606 ( .A(n503), .B(n362), .Z(n502) );
  XOR U607 ( .A(\min_val_reg[3][25] ), .B(DB[25]), .Z(n503) );
  XNOR U608 ( .A(n504), .B(n505), .Z(min_val_out[117]) );
  AND U609 ( .A(n150), .B(n422), .Z(n504) );
  XNOR U610 ( .A(\min_val_reg[2][24] ), .B(n505), .Z(n422) );
  XOR U611 ( .A(\min_val_reg[3][24] ), .B(n506), .Z(n505) );
  NAND U612 ( .A(n507), .B(n362), .Z(n506) );
  XOR U613 ( .A(\min_val_reg[3][24] ), .B(DB[24]), .Z(n507) );
  XNOR U614 ( .A(n508), .B(n509), .Z(min_val_out[116]) );
  AND U615 ( .A(n150), .B(n426), .Z(n508) );
  XNOR U616 ( .A(\min_val_reg[2][23] ), .B(n509), .Z(n426) );
  XOR U617 ( .A(\min_val_reg[3][23] ), .B(n510), .Z(n509) );
  NAND U618 ( .A(n511), .B(n362), .Z(n510) );
  XOR U619 ( .A(\min_val_reg[3][23] ), .B(DB[23]), .Z(n511) );
  XNOR U620 ( .A(n512), .B(n513), .Z(min_val_out[115]) );
  AND U621 ( .A(n150), .B(n430), .Z(n512) );
  XNOR U622 ( .A(\min_val_reg[2][22] ), .B(n513), .Z(n430) );
  XOR U623 ( .A(\min_val_reg[3][22] ), .B(n514), .Z(n513) );
  NAND U624 ( .A(n515), .B(n362), .Z(n514) );
  XOR U625 ( .A(\min_val_reg[3][22] ), .B(DB[22]), .Z(n515) );
  XNOR U626 ( .A(n516), .B(n517), .Z(min_val_out[114]) );
  AND U627 ( .A(n150), .B(n434), .Z(n516) );
  XNOR U628 ( .A(\min_val_reg[2][21] ), .B(n517), .Z(n434) );
  XOR U629 ( .A(\min_val_reg[3][21] ), .B(n518), .Z(n517) );
  NAND U630 ( .A(n519), .B(n362), .Z(n518) );
  XOR U631 ( .A(\min_val_reg[3][21] ), .B(DB[21]), .Z(n519) );
  XNOR U632 ( .A(n520), .B(n521), .Z(min_val_out[113]) );
  AND U633 ( .A(n150), .B(n438), .Z(n520) );
  XNOR U634 ( .A(\min_val_reg[2][20] ), .B(n521), .Z(n438) );
  XOR U635 ( .A(\min_val_reg[3][20] ), .B(n522), .Z(n521) );
  NAND U636 ( .A(n523), .B(n362), .Z(n522) );
  XOR U637 ( .A(\min_val_reg[3][20] ), .B(DB[20]), .Z(n523) );
  XNOR U638 ( .A(n524), .B(n525), .Z(min_val_out[112]) );
  AND U639 ( .A(n150), .B(n447), .Z(n524) );
  XNOR U640 ( .A(\min_val_reg[2][19] ), .B(n525), .Z(n447) );
  XOR U641 ( .A(\min_val_reg[3][19] ), .B(n526), .Z(n525) );
  NAND U642 ( .A(n527), .B(n362), .Z(n526) );
  XOR U643 ( .A(\min_val_reg[3][19] ), .B(DB[19]), .Z(n527) );
  XNOR U644 ( .A(n528), .B(n529), .Z(min_val_out[111]) );
  AND U645 ( .A(n150), .B(n451), .Z(n528) );
  XNOR U646 ( .A(\min_val_reg[2][18] ), .B(n529), .Z(n451) );
  XOR U647 ( .A(\min_val_reg[3][18] ), .B(n530), .Z(n529) );
  NAND U648 ( .A(n531), .B(n362), .Z(n530) );
  XOR U649 ( .A(\min_val_reg[3][18] ), .B(DB[18]), .Z(n531) );
  XNOR U650 ( .A(n532), .B(n533), .Z(min_val_out[110]) );
  AND U651 ( .A(n150), .B(n455), .Z(n532) );
  XNOR U652 ( .A(\min_val_reg[2][17] ), .B(n533), .Z(n455) );
  XOR U653 ( .A(\min_val_reg[3][17] ), .B(n534), .Z(n533) );
  NAND U654 ( .A(n535), .B(n362), .Z(n534) );
  XOR U655 ( .A(\min_val_reg[3][17] ), .B(DB[17]), .Z(n535) );
  XOR U656 ( .A(\min_val_reg[0][10] ), .B(n536), .Z(min_val_out[10]) );
  AND U657 ( .A(n146), .B(n337), .Z(n536) );
  XNOR U658 ( .A(\min_val_reg[0][10] ), .B(n336), .Z(n337) );
  XOR U659 ( .A(\min_val_reg[1][10] ), .B(n537), .Z(n336) );
  NAND U660 ( .A(n237), .B(n172), .Z(n537) );
  XOR U661 ( .A(\min_val_reg[1][10] ), .B(n236), .Z(n237) );
  XNOR U662 ( .A(\min_val_reg[2][10] ), .B(n538), .Z(n236) );
  NAND U663 ( .A(n539), .B(n343), .Z(n538) );
  XNOR U664 ( .A(n540), .B(n541), .Z(min_val_out[109]) );
  AND U665 ( .A(n150), .B(n459), .Z(n540) );
  XNOR U666 ( .A(\min_val_reg[2][16] ), .B(n541), .Z(n459) );
  XOR U667 ( .A(\min_val_reg[3][16] ), .B(n542), .Z(n541) );
  NAND U668 ( .A(n543), .B(n362), .Z(n542) );
  XOR U669 ( .A(\min_val_reg[3][16] ), .B(DB[16]), .Z(n543) );
  XNOR U670 ( .A(n544), .B(n545), .Z(min_val_out[108]) );
  AND U671 ( .A(n150), .B(n463), .Z(n544) );
  XNOR U672 ( .A(\min_val_reg[2][15] ), .B(n545), .Z(n463) );
  XOR U673 ( .A(\min_val_reg[3][15] ), .B(n546), .Z(n545) );
  NAND U674 ( .A(n547), .B(n362), .Z(n546) );
  XOR U675 ( .A(\min_val_reg[3][15] ), .B(DB[15]), .Z(n547) );
  XNOR U676 ( .A(n548), .B(n549), .Z(min_val_out[107]) );
  AND U677 ( .A(n150), .B(n467), .Z(n548) );
  XNOR U678 ( .A(\min_val_reg[2][14] ), .B(n549), .Z(n467) );
  XOR U679 ( .A(\min_val_reg[3][14] ), .B(n550), .Z(n549) );
  NAND U680 ( .A(n551), .B(n362), .Z(n550) );
  XOR U681 ( .A(\min_val_reg[3][14] ), .B(DB[14]), .Z(n551) );
  XNOR U682 ( .A(n552), .B(n553), .Z(min_val_out[106]) );
  AND U683 ( .A(n150), .B(n471), .Z(n552) );
  XNOR U684 ( .A(\min_val_reg[2][13] ), .B(n553), .Z(n471) );
  XOR U685 ( .A(\min_val_reg[3][13] ), .B(n554), .Z(n553) );
  NAND U686 ( .A(n555), .B(n362), .Z(n554) );
  XOR U687 ( .A(\min_val_reg[3][13] ), .B(DB[13]), .Z(n555) );
  XNOR U688 ( .A(n556), .B(n557), .Z(min_val_out[105]) );
  AND U689 ( .A(n150), .B(n475), .Z(n556) );
  XNOR U690 ( .A(\min_val_reg[2][12] ), .B(n557), .Z(n475) );
  XOR U691 ( .A(\min_val_reg[3][12] ), .B(n558), .Z(n557) );
  NAND U692 ( .A(n559), .B(n362), .Z(n558) );
  XOR U693 ( .A(\min_val_reg[3][12] ), .B(DB[12]), .Z(n559) );
  XNOR U694 ( .A(n560), .B(n561), .Z(min_val_out[104]) );
  AND U695 ( .A(n150), .B(n495), .Z(n560) );
  XNOR U696 ( .A(\min_val_reg[2][11] ), .B(n561), .Z(n495) );
  XOR U697 ( .A(\min_val_reg[3][11] ), .B(n562), .Z(n561) );
  NAND U698 ( .A(n563), .B(n362), .Z(n562) );
  XOR U699 ( .A(\min_val_reg[3][11] ), .B(DB[11]), .Z(n563) );
  XNOR U700 ( .A(n564), .B(n565), .Z(min_val_out[103]) );
  AND U701 ( .A(n150), .B(n539), .Z(n564) );
  XNOR U702 ( .A(\min_val_reg[2][10] ), .B(n565), .Z(n539) );
  XOR U703 ( .A(\min_val_reg[3][10] ), .B(n566), .Z(n565) );
  NAND U704 ( .A(n567), .B(n362), .Z(n566) );
  XOR U705 ( .A(\min_val_reg[3][10] ), .B(DB[10]), .Z(n567) );
  XNOR U706 ( .A(n568), .B(n569), .Z(min_val_out[102]) );
  AND U707 ( .A(n150), .B(n342), .Z(n568) );
  XNOR U708 ( .A(\min_val_reg[2][9] ), .B(n569), .Z(n342) );
  XOR U709 ( .A(\min_val_reg[3][9] ), .B(n570), .Z(n569) );
  NAND U710 ( .A(n571), .B(n362), .Z(n570) );
  XOR U711 ( .A(\min_val_reg[3][9] ), .B(DB[9]), .Z(n571) );
  XNOR U712 ( .A(n572), .B(n573), .Z(min_val_out[101]) );
  AND U713 ( .A(n150), .B(n350), .Z(n572) );
  XNOR U714 ( .A(\min_val_reg[2][8] ), .B(n573), .Z(n350) );
  XOR U715 ( .A(\min_val_reg[3][8] ), .B(n574), .Z(n573) );
  NAND U716 ( .A(n575), .B(n362), .Z(n574) );
  XOR U717 ( .A(\min_val_reg[3][8] ), .B(DB[8]), .Z(n575) );
  XNOR U718 ( .A(n576), .B(n577), .Z(min_val_out[100]) );
  AND U719 ( .A(n150), .B(n355), .Z(n576) );
  XNOR U720 ( .A(\min_val_reg[2][7] ), .B(n577), .Z(n355) );
  XOR U721 ( .A(\min_val_reg[3][7] ), .B(n578), .Z(n577) );
  NAND U722 ( .A(n579), .B(n362), .Z(n578) );
  XOR U723 ( .A(\min_val_reg[3][7] ), .B(DB[7]), .Z(n579) );
  XOR U724 ( .A(\min_val_reg[0][0] ), .B(n580), .Z(min_val_out[0]) );
  AND U725 ( .A(n146), .B(n389), .Z(n580) );
  XNOR U726 ( .A(\min_val_reg[0][0] ), .B(n388), .Z(n389) );
  XOR U727 ( .A(\min_val_reg[1][0] ), .B(n581), .Z(n388) );
  NAND U728 ( .A(n269), .B(n172), .Z(n581) );
  XNOR U729 ( .A(\min_val_reg[1][0] ), .B(n268), .Z(n269) );
  XOR U730 ( .A(\min_val_reg[2][0] ), .B(n582), .Z(n268) );
  NAND U731 ( .A(n169), .B(n343), .Z(n582) );
  XNOR U732 ( .A(\min_val_reg[2][0] ), .B(n168), .Z(n169) );
  XOR U733 ( .A(\min_val_reg[3][0] ), .B(n583), .Z(n168) );
  NAND U734 ( .A(n584), .B(n362), .Z(n583) );
  XOR U735 ( .A(\min_val_reg[3][0] ), .B(DB[0]), .Z(n584) );
  XOR U736 ( .A(n585), .B(n586), .Z(\min_dist[3][4] ) );
  AND U737 ( .A(n150), .B(n587), .Z(n585) );
  XOR U738 ( .A(\min_dist_reg[2][4] ), .B(n586), .Z(n587) );
  XOR U739 ( .A(n588), .B(n589), .Z(\min_dist[3][3] ) );
  AND U740 ( .A(n150), .B(n590), .Z(n588) );
  XNOR U741 ( .A(\min_dist_reg[2][3] ), .B(n591), .Z(n590) );
  XOR U742 ( .A(n592), .B(n593), .Z(\min_dist[3][2] ) );
  AND U743 ( .A(n150), .B(n594), .Z(n592) );
  XNOR U744 ( .A(\min_dist_reg[2][2] ), .B(n595), .Z(n594) );
  XOR U745 ( .A(n596), .B(n597), .Z(\min_dist[3][1] ) );
  AND U746 ( .A(n150), .B(n598), .Z(n596) );
  XNOR U747 ( .A(\min_dist_reg[2][1] ), .B(n599), .Z(n598) );
  XOR U748 ( .A(n600), .B(n601), .Z(\min_dist[3][0] ) );
  AND U749 ( .A(n150), .B(n602), .Z(n600) );
  XOR U750 ( .A(n603), .B(n604), .Z(n150) );
  AND U751 ( .A(n605), .B(n606), .Z(n603) );
  XNOR U752 ( .A(n586), .B(n604), .Z(n606) );
  XNOR U753 ( .A(n607), .B(n604), .Z(n605) );
  XOR U754 ( .A(n608), .B(n609), .Z(n604) );
  AND U755 ( .A(n610), .B(n611), .Z(n608) );
  XNOR U756 ( .A(n591), .B(n612), .Z(n611) );
  IV U757 ( .A(n609), .Z(n612) );
  IV U758 ( .A(n589), .Z(n591) );
  XOR U759 ( .A(n613), .B(n614), .Z(\min_dist[2][4] ) );
  AND U760 ( .A(n172), .B(n615), .Z(n613) );
  XOR U761 ( .A(\min_dist_reg[1][4] ), .B(n614), .Z(n615) );
  XOR U762 ( .A(n616), .B(n617), .Z(\min_dist[2][3] ) );
  AND U763 ( .A(n172), .B(n618), .Z(n616) );
  XOR U764 ( .A(\min_dist_reg[1][3] ), .B(n617), .Z(n618) );
  XOR U765 ( .A(n619), .B(n620), .Z(\min_dist[2][2] ) );
  AND U766 ( .A(n172), .B(n621), .Z(n619) );
  XOR U767 ( .A(\min_dist_reg[1][2] ), .B(n620), .Z(n621) );
  XOR U768 ( .A(n622), .B(n623), .Z(\min_dist[2][1] ) );
  AND U769 ( .A(n172), .B(n624), .Z(n622) );
  XOR U770 ( .A(\min_dist_reg[1][1] ), .B(n623), .Z(n624) );
  XOR U771 ( .A(n625), .B(n626), .Z(\min_dist[2][0] ) );
  AND U772 ( .A(n172), .B(n627), .Z(n625) );
  XOR U773 ( .A(n628), .B(n629), .Z(\min_dist[1][4] ) );
  AND U774 ( .A(n272), .B(n630), .Z(n628) );
  XOR U775 ( .A(\min_dist_reg[0][4] ), .B(n629), .Z(n630) );
  XOR U776 ( .A(n631), .B(n632), .Z(\min_dist[1][3] ) );
  AND U777 ( .A(n272), .B(n633), .Z(n631) );
  XOR U778 ( .A(n634), .B(n635), .Z(\min_dist[1][2] ) );
  AND U779 ( .A(n272), .B(n636), .Z(n634) );
  XOR U780 ( .A(n637), .B(n638), .Z(\min_dist[1][1] ) );
  AND U781 ( .A(n272), .B(n639), .Z(n637) );
  XNOR U782 ( .A(n640), .B(n641), .Z(\min_dist[1][0] ) );
  AND U783 ( .A(n272), .B(n642), .Z(n640) );
  XNOR U784 ( .A(\min_dist_reg[0][0] ), .B(n641), .Z(n642) );
  XNOR U785 ( .A(n643), .B(n644), .Z(n272) );
  AND U786 ( .A(n645), .B(n646), .Z(n643) );
  XOR U787 ( .A(n629), .B(n644), .Z(n646) );
  XNOR U788 ( .A(\min_dist_reg[0][4] ), .B(n644), .Z(n645) );
  XOR U789 ( .A(n647), .B(n648), .Z(n644) );
  AND U790 ( .A(n649), .B(n650), .Z(n647) );
  XNOR U791 ( .A(n632), .B(n651), .Z(n650) );
  XNOR U792 ( .A(\min_dist_reg[0][3] ), .B(n648), .Z(n649) );
  IV U793 ( .A(n651), .Z(n648) );
  XOR U794 ( .A(n652), .B(n653), .Z(n651) );
  AND U795 ( .A(n654), .B(n655), .Z(n652) );
  XNOR U796 ( .A(n635), .B(n653), .Z(n655) );
  XOR U797 ( .A(\min_dist_reg[0][2] ), .B(n653), .Z(n654) );
  XOR U798 ( .A(n656), .B(n657), .Z(n653) );
  NAND U799 ( .A(n658), .B(n659), .Z(n657) );
  XOR U800 ( .A(n656), .B(n638), .Z(n659) );
  XNOR U801 ( .A(\min_dist_reg[0][1] ), .B(n656), .Z(n658) );
  NOR U802 ( .A(n641), .B(\min_dist_reg[0][0] ), .Z(n656) );
  AND U803 ( .A(\min_dist_reg[0][4] ), .B(n660), .Z(\local_min_dist[0][4] ) );
  NANDN U804 ( .A(n629), .B(n146), .Z(n660) );
  XOR U805 ( .A(\min_dist_reg[0][3] ), .B(n661), .Z(\local_min_dist[0][3] ) );
  AND U806 ( .A(n146), .B(n633), .Z(n661) );
  XOR U807 ( .A(\min_dist_reg[0][3] ), .B(n632), .Z(n633) );
  XOR U808 ( .A(\min_dist_reg[0][2] ), .B(n662), .Z(\local_min_dist[0][2] ) );
  AND U809 ( .A(n146), .B(n636), .Z(n662) );
  XOR U810 ( .A(\min_dist_reg[0][2] ), .B(n635), .Z(n636) );
  XOR U811 ( .A(\min_dist_reg[0][1] ), .B(n663), .Z(\local_min_dist[0][1] ) );
  AND U812 ( .A(n146), .B(n639), .Z(n663) );
  XOR U813 ( .A(\min_dist_reg[0][1] ), .B(n638), .Z(n639) );
  XOR U814 ( .A(\min_dist_reg[0][0] ), .B(n664), .Z(\local_min_dist[0][0] ) );
  AND U815 ( .A(n146), .B(n665), .Z(n664) );
  XOR U816 ( .A(\min_dist_reg[0][0] ), .B(n666), .Z(n665) );
  XNOR U817 ( .A(n667), .B(n668), .Z(n146) );
  AND U818 ( .A(n669), .B(n670), .Z(n667) );
  XOR U819 ( .A(n629), .B(n668), .Z(n670) );
  AND U820 ( .A(n671), .B(\min_dist_reg[1][4] ), .Z(n629) );
  NANDN U821 ( .A(n614), .B(n172), .Z(n671) );
  XNOR U822 ( .A(\min_dist_reg[0][4] ), .B(n668), .Z(n669) );
  XOR U823 ( .A(n672), .B(n673), .Z(n668) );
  AND U824 ( .A(n674), .B(n675), .Z(n672) );
  XNOR U825 ( .A(n676), .B(n632), .Z(n675) );
  XNOR U826 ( .A(\min_dist_reg[1][3] ), .B(n677), .Z(n632) );
  NAND U827 ( .A(n678), .B(n172), .Z(n677) );
  XNOR U828 ( .A(n679), .B(n617), .Z(n678) );
  XNOR U829 ( .A(\min_dist_reg[0][3] ), .B(n673), .Z(n674) );
  IV U830 ( .A(n676), .Z(n673) );
  XOR U831 ( .A(n680), .B(n681), .Z(n676) );
  AND U832 ( .A(n682), .B(n683), .Z(n680) );
  XNOR U833 ( .A(n681), .B(n635), .Z(n683) );
  XNOR U834 ( .A(\min_dist_reg[1][2] ), .B(n684), .Z(n635) );
  NAND U835 ( .A(n685), .B(n172), .Z(n684) );
  XNOR U836 ( .A(n686), .B(n620), .Z(n685) );
  XOR U837 ( .A(\min_dist_reg[0][2] ), .B(n681), .Z(n682) );
  XOR U838 ( .A(n687), .B(n688), .Z(n681) );
  NAND U839 ( .A(n689), .B(n690), .Z(n688) );
  XOR U840 ( .A(n687), .B(n638), .Z(n690) );
  XNOR U841 ( .A(\min_dist_reg[1][1] ), .B(n691), .Z(n638) );
  NAND U842 ( .A(n692), .B(n172), .Z(n691) );
  XNOR U843 ( .A(n693), .B(n623), .Z(n692) );
  XNOR U844 ( .A(\min_dist_reg[0][1] ), .B(n687), .Z(n689) );
  ANDN U845 ( .B(n666), .A(\min_dist_reg[0][0] ), .Z(n687) );
  IV U846 ( .A(n641), .Z(n666) );
  XOR U847 ( .A(\min_dist_reg[1][0] ), .B(n694), .Z(n641) );
  NAND U848 ( .A(n627), .B(n172), .Z(n694) );
  XOR U849 ( .A(n695), .B(n696), .Z(n172) );
  AND U850 ( .A(n697), .B(n698), .Z(n695) );
  XNOR U851 ( .A(n614), .B(n696), .Z(n698) );
  AND U852 ( .A(n699), .B(\min_dist_reg[2][4] ), .Z(n614) );
  NANDN U853 ( .A(n586), .B(n343), .Z(n699) );
  XNOR U854 ( .A(n700), .B(n696), .Z(n697) );
  XOR U855 ( .A(n701), .B(n702), .Z(n696) );
  AND U856 ( .A(n703), .B(n704), .Z(n701) );
  XNOR U857 ( .A(n617), .B(n702), .Z(n704) );
  XNOR U858 ( .A(\min_dist_reg[2][3] ), .B(n705), .Z(n617) );
  NAND U859 ( .A(n706), .B(n343), .Z(n705) );
  XNOR U860 ( .A(n707), .B(n589), .Z(n706) );
  XNOR U861 ( .A(n679), .B(n702), .Z(n703) );
  XOR U862 ( .A(n708), .B(n709), .Z(n702) );
  AND U863 ( .A(n710), .B(n711), .Z(n708) );
  XNOR U864 ( .A(n620), .B(n709), .Z(n711) );
  XNOR U865 ( .A(\min_dist_reg[2][2] ), .B(n712), .Z(n620) );
  NAND U866 ( .A(n713), .B(n343), .Z(n712) );
  XNOR U867 ( .A(n714), .B(n593), .Z(n713) );
  XNOR U868 ( .A(n686), .B(n709), .Z(n710) );
  XOR U869 ( .A(n715), .B(n716), .Z(n709) );
  NAND U870 ( .A(n717), .B(n718), .Z(n716) );
  XOR U871 ( .A(n715), .B(n623), .Z(n718) );
  XNOR U872 ( .A(\min_dist_reg[2][1] ), .B(n719), .Z(n623) );
  NAND U873 ( .A(n720), .B(n343), .Z(n719) );
  XNOR U874 ( .A(n721), .B(n597), .Z(n720) );
  XOR U875 ( .A(n693), .B(n715), .Z(n717) );
  IV U876 ( .A(\min_dist_reg[1][1] ), .Z(n693) );
  AND U877 ( .A(n626), .B(n722), .Z(n715) );
  IV U878 ( .A(\min_dist_reg[1][2] ), .Z(n686) );
  IV U879 ( .A(\min_dist_reg[1][3] ), .Z(n679) );
  IV U880 ( .A(\min_dist_reg[1][4] ), .Z(n700) );
  XNOR U881 ( .A(n722), .B(n626), .Z(n627) );
  XNOR U882 ( .A(\min_dist_reg[2][0] ), .B(n723), .Z(n626) );
  NAND U883 ( .A(n602), .B(n343), .Z(n723) );
  XOR U884 ( .A(n724), .B(n725), .Z(n343) );
  AND U885 ( .A(n726), .B(n727), .Z(n724) );
  XNOR U886 ( .A(n725), .B(n586), .Z(n727) );
  XNOR U887 ( .A(\min_dist_reg[3][4] ), .B(n728), .Z(n586) );
  NAND U888 ( .A(n729), .B(n362), .Z(n728) );
  XOR U889 ( .A(\min_dist_reg[3][4] ), .B(n730), .Z(n729) );
  XNOR U890 ( .A(n607), .B(n725), .Z(n726) );
  XOR U891 ( .A(n731), .B(n609), .Z(n725) );
  AND U892 ( .A(n610), .B(n732), .Z(n731) );
  XNOR U893 ( .A(n609), .B(n589), .Z(n732) );
  XNOR U894 ( .A(\min_dist_reg[3][3] ), .B(n733), .Z(n589) );
  NAND U895 ( .A(n734), .B(n362), .Z(n733) );
  XNOR U896 ( .A(\min_dist_reg[3][3] ), .B(n735), .Z(n734) );
  XNOR U897 ( .A(n707), .B(n609), .Z(n610) );
  XOR U898 ( .A(n736), .B(n737), .Z(n609) );
  AND U899 ( .A(n738), .B(n739), .Z(n736) );
  XOR U900 ( .A(n595), .B(n737), .Z(n739) );
  IV U901 ( .A(n593), .Z(n595) );
  XNOR U902 ( .A(\min_dist_reg[3][2] ), .B(n740), .Z(n593) );
  NAND U903 ( .A(n741), .B(n362), .Z(n740) );
  XNOR U904 ( .A(\min_dist_reg[3][2] ), .B(n742), .Z(n741) );
  XNOR U905 ( .A(n714), .B(n737), .Z(n738) );
  XOR U906 ( .A(n743), .B(n744), .Z(n737) );
  NAND U907 ( .A(n745), .B(n746), .Z(n744) );
  XNOR U908 ( .A(n743), .B(n599), .Z(n746) );
  IV U909 ( .A(n597), .Z(n599) );
  XNOR U910 ( .A(\min_dist_reg[3][1] ), .B(n747), .Z(n597) );
  NAND U911 ( .A(n748), .B(n362), .Z(n747) );
  XNOR U912 ( .A(\min_dist_reg[3][1] ), .B(n749), .Z(n748) );
  XOR U913 ( .A(n721), .B(n743), .Z(n745) );
  IV U914 ( .A(\min_dist_reg[2][1] ), .Z(n721) );
  ANDN U915 ( .B(n601), .A(\min_dist_reg[2][0] ), .Z(n743) );
  IV U916 ( .A(\min_dist_reg[2][2] ), .Z(n714) );
  IV U917 ( .A(\min_dist_reg[2][3] ), .Z(n707) );
  IV U918 ( .A(\min_dist_reg[2][4] ), .Z(n607) );
  XOR U919 ( .A(\min_dist_reg[2][0] ), .B(n601), .Z(n602) );
  XOR U920 ( .A(n750), .B(n751), .Z(n601) );
  NAND U921 ( .A(n752), .B(n362), .Z(n751) );
  XNOR U922 ( .A(n753), .B(n754), .Z(n362) );
  AND U923 ( .A(n755), .B(n756), .Z(n753) );
  XNOR U924 ( .A(n757), .B(n730), .Z(n756) );
  XNOR U925 ( .A(n758), .B(n759), .Z(n730) );
  ANDN U926 ( .B(n760), .A(n761), .Z(n758) );
  XOR U927 ( .A(n759), .B(n762), .Z(n760) );
  XNOR U928 ( .A(\min_dist_reg[3][4] ), .B(n754), .Z(n755) );
  IV U929 ( .A(n757), .Z(n754) );
  XOR U930 ( .A(n763), .B(n764), .Z(n757) );
  AND U931 ( .A(n765), .B(n766), .Z(n763) );
  XOR U932 ( .A(n764), .B(n735), .Z(n766) );
  XOR U933 ( .A(n767), .B(n762), .Z(n735) );
  XNOR U934 ( .A(n768), .B(n769), .Z(n762) );
  ANDN U935 ( .B(n770), .A(n771), .Z(n768) );
  XOR U936 ( .A(n772), .B(n773), .Z(n770) );
  IV U937 ( .A(n761), .Z(n767) );
  XOR U938 ( .A(n774), .B(n775), .Z(n761) );
  XNOR U939 ( .A(n776), .B(n777), .Z(n775) );
  ANDN U940 ( .B(n778), .A(n779), .Z(n776) );
  XNOR U941 ( .A(n780), .B(n781), .Z(n778) );
  IV U942 ( .A(n759), .Z(n774) );
  XOR U943 ( .A(n782), .B(n783), .Z(n759) );
  ANDN U944 ( .B(n784), .A(n785), .Z(n782) );
  XOR U945 ( .A(n783), .B(n786), .Z(n784) );
  XNOR U946 ( .A(\min_dist_reg[3][3] ), .B(n787), .Z(n765) );
  IV U947 ( .A(n764), .Z(n787) );
  XOR U948 ( .A(n788), .B(n789), .Z(n764) );
  AND U949 ( .A(n790), .B(n791), .Z(n788) );
  XOR U950 ( .A(n789), .B(n742), .Z(n791) );
  XOR U951 ( .A(n792), .B(n786), .Z(n742) );
  XOR U952 ( .A(n793), .B(n773), .Z(n786) );
  XNOR U953 ( .A(n794), .B(n795), .Z(n773) );
  ANDN U954 ( .B(n796), .A(n797), .Z(n794) );
  XOR U955 ( .A(n798), .B(n799), .Z(n796) );
  IV U956 ( .A(n771), .Z(n793) );
  XOR U957 ( .A(n769), .B(n800), .Z(n771) );
  XNOR U958 ( .A(n801), .B(n802), .Z(n800) );
  ANDN U959 ( .B(n803), .A(n804), .Z(n801) );
  XNOR U960 ( .A(n805), .B(n806), .Z(n803) );
  IV U961 ( .A(n772), .Z(n769) );
  XOR U962 ( .A(n807), .B(n808), .Z(n772) );
  ANDN U963 ( .B(n809), .A(n810), .Z(n807) );
  XOR U964 ( .A(n808), .B(n811), .Z(n809) );
  IV U965 ( .A(n785), .Z(n792) );
  XOR U966 ( .A(n812), .B(n813), .Z(n785) );
  XNOR U967 ( .A(n780), .B(n814), .Z(n813) );
  IV U968 ( .A(n783), .Z(n814) );
  XOR U969 ( .A(n815), .B(n816), .Z(n783) );
  ANDN U970 ( .B(n817), .A(n818), .Z(n815) );
  XOR U971 ( .A(n816), .B(n819), .Z(n817) );
  XNOR U972 ( .A(n820), .B(n821), .Z(n780) );
  ANDN U973 ( .B(n822), .A(n823), .Z(n820) );
  XOR U974 ( .A(n821), .B(n824), .Z(n822) );
  IV U975 ( .A(n779), .Z(n812) );
  XOR U976 ( .A(n777), .B(n825), .Z(n779) );
  XNOR U977 ( .A(n826), .B(n827), .Z(n825) );
  ANDN U978 ( .B(n828), .A(n829), .Z(n826) );
  XNOR U979 ( .A(n830), .B(n831), .Z(n828) );
  IV U980 ( .A(n781), .Z(n777) );
  XOR U981 ( .A(n832), .B(n833), .Z(n781) );
  ANDN U982 ( .B(n834), .A(n835), .Z(n832) );
  XOR U983 ( .A(n836), .B(n833), .Z(n834) );
  XOR U984 ( .A(\min_dist_reg[3][2] ), .B(n789), .Z(n790) );
  XOR U985 ( .A(n837), .B(n838), .Z(n789) );
  NAND U986 ( .A(n839), .B(n840), .Z(n838) );
  XNOR U987 ( .A(n837), .B(n749), .Z(n840) );
  XOR U988 ( .A(n841), .B(n819), .Z(n749) );
  XOR U989 ( .A(n842), .B(n811), .Z(n819) );
  XOR U990 ( .A(n843), .B(n799), .Z(n811) );
  XNOR U991 ( .A(n844), .B(n845), .Z(n799) );
  ANDN U992 ( .B(n846), .A(n847), .Z(n844) );
  XNOR U993 ( .A(n845), .B(n848), .Z(n846) );
  IV U994 ( .A(n797), .Z(n843) );
  XOR U995 ( .A(n795), .B(n849), .Z(n797) );
  XNOR U996 ( .A(n850), .B(n851), .Z(n849) );
  ANDN U997 ( .B(n852), .A(n853), .Z(n850) );
  XNOR U998 ( .A(n854), .B(n855), .Z(n852) );
  IV U999 ( .A(n851), .Z(n855) );
  IV U1000 ( .A(n798), .Z(n795) );
  XNOR U1001 ( .A(n856), .B(n857), .Z(n798) );
  ANDN U1002 ( .B(n858), .A(n859), .Z(n856) );
  XNOR U1003 ( .A(n857), .B(n860), .Z(n858) );
  IV U1004 ( .A(n810), .Z(n842) );
  XOR U1005 ( .A(n861), .B(n862), .Z(n810) );
  XNOR U1006 ( .A(n805), .B(n863), .Z(n862) );
  IV U1007 ( .A(n808), .Z(n863) );
  XNOR U1008 ( .A(n864), .B(n865), .Z(n808) );
  ANDN U1009 ( .B(n866), .A(n867), .Z(n864) );
  XNOR U1010 ( .A(n865), .B(n868), .Z(n866) );
  XOR U1011 ( .A(n869), .B(n870), .Z(n805) );
  ANDN U1012 ( .B(n871), .A(n872), .Z(n869) );
  XNOR U1013 ( .A(n870), .B(n873), .Z(n871) );
  IV U1014 ( .A(n804), .Z(n861) );
  XOR U1015 ( .A(n802), .B(n874), .Z(n804) );
  XNOR U1016 ( .A(n875), .B(n876), .Z(n874) );
  ANDN U1017 ( .B(n877), .A(n878), .Z(n875) );
  XNOR U1018 ( .A(n879), .B(n880), .Z(n877) );
  IV U1019 ( .A(n876), .Z(n880) );
  IV U1020 ( .A(n806), .Z(n802) );
  XNOR U1021 ( .A(n881), .B(n882), .Z(n806) );
  ANDN U1022 ( .B(n883), .A(n884), .Z(n881) );
  XNOR U1023 ( .A(n885), .B(n882), .Z(n883) );
  IV U1024 ( .A(n818), .Z(n841) );
  XOR U1025 ( .A(n886), .B(n887), .Z(n818) );
  XOR U1026 ( .A(n836), .B(n888), .Z(n887) );
  IV U1027 ( .A(n816), .Z(n888) );
  XNOR U1028 ( .A(n889), .B(n890), .Z(n816) );
  ANDN U1029 ( .B(n891), .A(n892), .Z(n889) );
  XNOR U1030 ( .A(n890), .B(n893), .Z(n891) );
  XOR U1031 ( .A(n894), .B(n824), .Z(n836) );
  XNOR U1032 ( .A(n895), .B(n896), .Z(n824) );
  ANDN U1033 ( .B(n897), .A(n898), .Z(n895) );
  XNOR U1034 ( .A(n896), .B(n899), .Z(n897) );
  IV U1035 ( .A(n823), .Z(n894) );
  XOR U1036 ( .A(n900), .B(n901), .Z(n823) );
  XNOR U1037 ( .A(n902), .B(n903), .Z(n901) );
  ANDN U1038 ( .B(n904), .A(n905), .Z(n902) );
  XNOR U1039 ( .A(n906), .B(n907), .Z(n904) );
  IV U1040 ( .A(n903), .Z(n907) );
  IV U1041 ( .A(n821), .Z(n900) );
  XNOR U1042 ( .A(n908), .B(n909), .Z(n821) );
  ANDN U1043 ( .B(n910), .A(n911), .Z(n908) );
  XNOR U1044 ( .A(n909), .B(n912), .Z(n910) );
  IV U1045 ( .A(n835), .Z(n886) );
  XOR U1046 ( .A(n913), .B(n914), .Z(n835) );
  XNOR U1047 ( .A(n830), .B(n915), .Z(n914) );
  IV U1048 ( .A(n833), .Z(n915) );
  XNOR U1049 ( .A(n916), .B(n917), .Z(n833) );
  ANDN U1050 ( .B(n918), .A(n919), .Z(n916) );
  XNOR U1051 ( .A(n920), .B(n917), .Z(n918) );
  XOR U1052 ( .A(n921), .B(n922), .Z(n830) );
  ANDN U1053 ( .B(n923), .A(n924), .Z(n921) );
  XNOR U1054 ( .A(n922), .B(n925), .Z(n923) );
  IV U1055 ( .A(n829), .Z(n913) );
  XOR U1056 ( .A(n827), .B(n926), .Z(n829) );
  XNOR U1057 ( .A(n927), .B(n928), .Z(n926) );
  ANDN U1058 ( .B(n929), .A(n930), .Z(n927) );
  XNOR U1059 ( .A(n931), .B(n932), .Z(n929) );
  IV U1060 ( .A(n928), .Z(n932) );
  IV U1061 ( .A(n831), .Z(n827) );
  XNOR U1062 ( .A(n933), .B(n934), .Z(n831) );
  ANDN U1063 ( .B(n935), .A(n936), .Z(n933) );
  XNOR U1064 ( .A(n937), .B(n934), .Z(n935) );
  XNOR U1065 ( .A(\min_dist_reg[3][1] ), .B(n837), .Z(n839) );
  NOR U1066 ( .A(\min_dist_reg[3][0] ), .B(n938), .Z(n837) );
  XOR U1067 ( .A(n750), .B(n938), .Z(n752) );
  XOR U1068 ( .A(n939), .B(n893), .Z(n938) );
  XOR U1069 ( .A(n940), .B(n868), .Z(n893) );
  XOR U1070 ( .A(n941), .B(n860), .Z(n868) );
  XOR U1071 ( .A(n942), .B(n848), .Z(n860) );
  XNOR U1072 ( .A(q[30]), .B(DB[30]), .Z(n848) );
  IV U1073 ( .A(n847), .Z(n942) );
  XOR U1074 ( .A(n845), .B(n943), .Z(n847) );
  XNOR U1075 ( .A(q[29]), .B(DB[29]), .Z(n943) );
  XOR U1076 ( .A(q[28]), .B(DB[28]), .Z(n845) );
  IV U1077 ( .A(n859), .Z(n941) );
  XOR U1078 ( .A(n944), .B(n945), .Z(n859) );
  XNOR U1079 ( .A(n854), .B(n857), .Z(n945) );
  XOR U1080 ( .A(q[24]), .B(DB[24]), .Z(n857) );
  XOR U1081 ( .A(q[27]), .B(DB[27]), .Z(n854) );
  IV U1082 ( .A(n853), .Z(n944) );
  XOR U1083 ( .A(n851), .B(n946), .Z(n853) );
  XNOR U1084 ( .A(q[26]), .B(DB[26]), .Z(n946) );
  XOR U1085 ( .A(q[25]), .B(DB[25]), .Z(n851) );
  IV U1086 ( .A(n867), .Z(n940) );
  XOR U1087 ( .A(n947), .B(n948), .Z(n867) );
  XOR U1088 ( .A(n885), .B(n865), .Z(n948) );
  XOR U1089 ( .A(q[16]), .B(DB[16]), .Z(n865) );
  XOR U1090 ( .A(n949), .B(n873), .Z(n885) );
  XNOR U1091 ( .A(q[23]), .B(DB[23]), .Z(n873) );
  IV U1092 ( .A(n872), .Z(n949) );
  XOR U1093 ( .A(n870), .B(n950), .Z(n872) );
  XNOR U1094 ( .A(q[22]), .B(DB[22]), .Z(n950) );
  XOR U1095 ( .A(q[21]), .B(DB[21]), .Z(n870) );
  IV U1096 ( .A(n884), .Z(n947) );
  XOR U1097 ( .A(n951), .B(n952), .Z(n884) );
  XNOR U1098 ( .A(n879), .B(n882), .Z(n952) );
  XOR U1099 ( .A(q[17]), .B(DB[17]), .Z(n882) );
  XOR U1100 ( .A(q[20]), .B(DB[20]), .Z(n879) );
  IV U1101 ( .A(n878), .Z(n951) );
  XOR U1102 ( .A(n876), .B(n953), .Z(n878) );
  XNOR U1103 ( .A(q[19]), .B(DB[19]), .Z(n953) );
  XOR U1104 ( .A(q[18]), .B(DB[18]), .Z(n876) );
  IV U1105 ( .A(n892), .Z(n939) );
  XOR U1106 ( .A(n954), .B(n955), .Z(n892) );
  XOR U1107 ( .A(n920), .B(n890), .Z(n955) );
  XOR U1108 ( .A(q[0]), .B(DB[0]), .Z(n890) );
  XOR U1109 ( .A(n956), .B(n912), .Z(n920) );
  XOR U1110 ( .A(n957), .B(n899), .Z(n912) );
  XNOR U1111 ( .A(q[15]), .B(DB[15]), .Z(n899) );
  IV U1112 ( .A(n898), .Z(n957) );
  XOR U1113 ( .A(n896), .B(n958), .Z(n898) );
  XNOR U1114 ( .A(q[14]), .B(DB[14]), .Z(n958) );
  XOR U1115 ( .A(q[13]), .B(DB[13]), .Z(n896) );
  IV U1116 ( .A(n911), .Z(n956) );
  XOR U1117 ( .A(n959), .B(n960), .Z(n911) );
  XNOR U1118 ( .A(n906), .B(n909), .Z(n960) );
  XOR U1119 ( .A(q[9]), .B(DB[9]), .Z(n909) );
  XOR U1120 ( .A(q[12]), .B(DB[12]), .Z(n906) );
  IV U1121 ( .A(n905), .Z(n959) );
  XOR U1122 ( .A(n903), .B(n961), .Z(n905) );
  XNOR U1123 ( .A(q[11]), .B(DB[11]), .Z(n961) );
  XOR U1124 ( .A(q[10]), .B(DB[10]), .Z(n903) );
  IV U1125 ( .A(n919), .Z(n954) );
  XOR U1126 ( .A(n962), .B(n963), .Z(n919) );
  XOR U1127 ( .A(n937), .B(n917), .Z(n963) );
  XOR U1128 ( .A(q[1]), .B(DB[1]), .Z(n917) );
  XOR U1129 ( .A(n964), .B(n925), .Z(n937) );
  XNOR U1130 ( .A(q[8]), .B(DB[8]), .Z(n925) );
  IV U1131 ( .A(n924), .Z(n964) );
  XOR U1132 ( .A(n922), .B(n965), .Z(n924) );
  XNOR U1133 ( .A(q[7]), .B(DB[7]), .Z(n965) );
  XOR U1134 ( .A(q[6]), .B(DB[6]), .Z(n922) );
  IV U1135 ( .A(n936), .Z(n962) );
  XOR U1136 ( .A(n966), .B(n967), .Z(n936) );
  XNOR U1137 ( .A(n931), .B(n934), .Z(n967) );
  XOR U1138 ( .A(q[2]), .B(DB[2]), .Z(n934) );
  XOR U1139 ( .A(q[5]), .B(DB[5]), .Z(n931) );
  IV U1140 ( .A(n930), .Z(n966) );
  XOR U1141 ( .A(n928), .B(n968), .Z(n930) );
  XNOR U1142 ( .A(q[4]), .B(DB[4]), .Z(n968) );
  XOR U1143 ( .A(q[3]), .B(DB[3]), .Z(n928) );
  IV U1144 ( .A(\min_dist_reg[3][0] ), .Z(n750) );
  IV U1145 ( .A(\min_dist_reg[1][0] ), .Z(n722) );
endmodule

